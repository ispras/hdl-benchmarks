module test ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , 
 n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , 
 n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , 
 n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , 
 n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , 
 n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , 
 n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , 
 n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , 
 n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , 
 n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , 
 n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , 
 n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , 
 n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , 
 n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , 
 n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , 
 n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , 
 n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , 
 n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , 
 n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , 
 n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , 
 n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , 
 n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , 
 n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , 
 n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , 
 n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , 
 n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , 
 n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , 
 n271 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , 
 n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , 
 n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , 
 n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , 
 n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , 
 n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , 
 n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , 
 n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 ;
output n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , 
 n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , 
 n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , 
 n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , 
 n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , 
 n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , 
 n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , 
 n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , 
 n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , 
 n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , 
 n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , 
 n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , 
 n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , 
 n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , 
 n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , 
 n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , 
 n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , 
 n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , 
 n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , 
 n271 ;
wire n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , 
 n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , 
 n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , 
 n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , 
 n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , 
 n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , 
 n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , 
 n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , 
 n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , 
 n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , 
 n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , 
 n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , 
 n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , 
 n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , 
 n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , 
 n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , 
 n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , 
 n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , 
 n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , 
 n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , 
 n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , 
 n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , 
 n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , 
 n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , 
 n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , 
 n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , 
 n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , 
 n815 , n347310 , n347311 , n347312 , n347313 , n347314 , n347315 , n347316 , n347317 , n347318 , 
 n347319 , n347320 , n347321 , n347322 , n347323 , n347324 , n347325 , n347326 , n347327 , n347328 , 
 n347329 , n347330 , n347331 , n347332 , n347333 , n347334 , n347335 , n347336 , n347337 , n347338 , 
 n347339 , n347340 , n347341 , n347342 , n347343 , n347344 , n347345 , n347346 , n347347 , n347348 , 
 n347349 , n347350 , n347351 , n347352 , n347353 , n347354 , n347355 , n347356 , n347357 , n347358 , 
 n347359 , n347360 , n347361 , n347362 , n347363 , n347364 , n347365 , n347366 , n347367 , n347368 , 
 n347369 , n347370 , n347371 , n347372 , n347373 , n347374 , n347375 , n347376 , n347377 , n347378 , 
 n347379 , n347380 , n347381 , n347382 , n347383 , n347384 , n347385 , n347386 , n347387 , n347388 , 
 n347389 , n347390 , n347391 , n347392 , n347393 , n347394 , n347395 , n347396 , n347397 , n347398 , 
 n347399 , n347400 , n347401 , n347402 , n347403 , n347404 , n347405 , n347406 , n347407 , n347408 , 
 n347409 , n347410 , n347411 , n347412 , n347413 , n347414 , n347415 , n347416 , n347417 , n347418 , 
 n347419 , n347420 , n347421 , n347422 , n347423 , n347424 , n347425 , n347426 , n347427 , n347428 , 
 n347429 , n347430 , n347431 , n347432 , n347433 , n347434 , n347435 , n347436 , n347437 , n347438 , 
 n347439 , n347440 , n347441 , n347442 , n347443 , n347444 , n347445 , n347446 , n347447 , n347448 , 
 n347449 , n347450 , n347451 , n347452 , n347453 , n347454 , n347455 , n347456 , n347457 , n347458 , 
 n347459 , n347460 , n347461 , n347462 , n347463 , n347464 , n347465 , n347466 , n347467 , n347468 , 
 n347469 , n347470 , n347471 , n347472 , n347473 , n347474 , n347475 , n347476 , n347477 , n347478 , 
 n347479 , n347480 , n347481 , n347482 , n347483 , n347484 , n347485 , n347486 , n347487 , n347488 , 
 n347489 , n347490 , n347491 , n347492 , n347493 , n347494 , n347495 , n347496 , n347497 , n347498 , 
 n347499 , n347500 , n347501 , n347502 , n347503 , n347504 , n347505 , n347506 , n347507 , n347508 , 
 n347509 , n347510 , n347511 , n347512 , n347513 , n347514 , n347515 , n347516 , n347517 , n347518 , 
 n347519 , n347520 , n347521 , n347522 , n347523 , n347524 , n347525 , n347526 , n347527 , n347528 , 
 n347529 , n347530 , n347531 , n347532 , n347533 , n347534 , n347535 , n347536 , n347537 , n347538 , 
 n347539 , n347540 , n347541 , n347542 , n347543 , n347544 , n347545 , n347546 , n347547 , n347548 , 
 n347549 , n347550 , n347551 , n347552 , n347553 , n347554 , n347555 , n347556 , n347557 , n347558 , 
 n347559 , n347560 , n347561 , n347562 , n347563 , n347564 , n347565 , n347566 , n347567 , n347568 , 
 n347569 , n347570 , n347571 , n347572 , n347573 , n347574 , n347575 , n347576 , n347577 , n347578 , 
 n347579 , n347580 , n347581 , n347582 , n347583 , n347584 , n347585 , n347586 , n347587 , n347588 , 
 n347589 , n347590 , n347591 , n347592 , n347593 , n347594 , n347595 , n347596 , n347597 , n347598 , 
 n347599 , n347600 , n347601 , n347602 , n347603 , n347604 , n347605 , n347606 , n347607 , n347608 , 
 n347609 , n347610 , n347611 , n347612 , n347613 , n347614 , n347615 , n347616 , n347617 , n347618 , 
 n347619 , n347620 , n347621 , n347622 , n347623 , n347624 , n347625 , n347626 , n347627 , n347628 , 
 n347629 , n347630 , n347631 , n347632 , n347633 , n347634 , n347635 , n347636 , n347637 , n347638 , 
 n347639 , n347640 , n347641 , n347642 , n347643 , n347644 , n347645 , n347646 , n347647 , n347648 , 
 n347649 , n347650 , n347651 , n347652 , n347653 , n347654 , n347655 , n347656 , n347657 , n347658 , 
 n347659 , n347660 , n347661 , n347662 , n347663 , n347664 , n347665 , n347666 , n347667 , n347668 , 
 n347669 , n347670 , n347671 , n347672 , n347673 , n347674 , n347675 , n347676 , n347677 , n347678 , 
 n347679 , n347680 , n347681 , n347682 , n347683 , n347684 , n347685 , n347686 , n347687 , n347688 , 
 n347689 , n347690 , n347691 , n347692 , n347693 , n347694 , n347695 , n347696 , n347697 , n347698 , 
 n347699 , n347700 , n347701 , n347702 , n347703 , n347704 , n347705 , n347706 , n347707 , n347708 , 
 n347709 , n347710 , n347711 , n347712 , n347713 , n347714 , n347715 , n347716 , n347717 , n347718 , 
 n347719 , n347720 , n347721 , n347722 , n347723 , n347724 , n347725 , n347726 , n347727 , n347728 , 
 n347729 , n347730 , n347731 , n347732 , n347733 , n347734 , n347735 , n347736 , n347737 , n347738 , 
 n347739 , n347740 , n347741 , n347742 , n347743 , n347744 , n347745 , n347746 , n347747 , n347748 , 
 n347749 , n347750 , n347751 , n347752 , n347753 , n347754 , n347755 , n347756 , n347757 , n347758 , 
 n347759 , n347760 , n347761 , n347762 , n347763 , n347764 , n347765 , n347766 , n347767 , n347768 , 
 n347769 , n347770 , n347771 , n347772 , n347773 , n347774 , n347775 , n347776 , n347777 , n347778 , 
 n347779 , n347780 , n347781 , n347782 , n347783 , n347784 , n347785 , n347786 , n347787 , n347788 , 
 n347789 , n347790 , n347791 , n347792 , n347793 , n347794 , n347795 , n347796 , n347797 , n347798 , 
 n347799 , n347800 , n347801 , n347802 , n347803 , n347804 , n347805 , n347806 , n347807 , n347808 , 
 n347809 , n347810 , n347811 , n347812 , n347813 , n347814 , n347815 , n347816 , n347817 , n347818 , 
 n347819 , n347820 , n347821 , n347822 , n347823 , n347824 , n347825 , n347826 , n347827 , n347828 , 
 n347829 , n347830 , n347831 , n347832 , n347833 , n347834 , n347835 , n347836 , n347837 , n347838 , 
 n347839 , n347840 , n347841 , n347842 , n347843 , n347844 , n347845 , n347846 , n347847 , n347848 , 
 n347849 , n347850 , n347851 , n347852 , n347853 , n347854 , n347855 , n347856 , n347857 , n347858 , 
 n347859 , n347860 , n347861 , n347862 , n347863 , n347864 , n347865 , n347866 , n347867 , n347868 , 
 n347869 , n347870 , n347871 , n347872 , n347873 , n347874 , n347875 , n347876 , n347877 , n347878 , 
 n347879 , n347880 , n347881 , n347882 , n347883 , n347884 , n347885 , n347886 , n347887 , n347888 , 
 n347889 , n347890 , n347891 , n347892 , n347893 , n347894 , n347895 , n347896 , n347897 , n347898 , 
 n347899 , n347900 , n347901 , n347902 , n347903 , n347904 , n347905 , n347906 , n347907 , n347908 , 
 n347909 , n347910 , n347911 , n347912 , n347913 , n347914 , n347915 , n347916 , n347917 , n347918 , 
 n347919 , n347920 , n347921 , n347922 , n347923 , n347924 , n347925 , n347926 , n347927 , n347928 , 
 n347929 , n347930 , n347931 , n347932 , n347933 , n347934 , n347935 , n347936 , n347937 , n347938 , 
 n347939 , n347940 , n347941 , n347942 , n347943 , n347944 , n347945 , n347946 , n347947 , n347948 , 
 n347949 , n347950 , n347951 , n347952 , n347953 , n347954 , n347955 , n347956 , n347957 , n347958 , 
 n347959 , n347960 , n347961 , n347962 , n347963 , n347964 , n347965 , n347966 , n347967 , n347968 , 
 n347969 , n347970 , n347971 , n347972 , n347973 , n347974 , n347975 , n347976 , n347977 , n347978 , 
 n347979 , n347980 , n347981 , n347982 , n347983 , n347984 , n347985 , n347986 , n347987 , n347988 , 
 n347989 , n347990 , n347991 , n347992 , n347993 , n347994 , n347995 , n347996 , n347997 , n347998 , 
 n347999 , n348000 , n348001 , n348002 , n348003 , n348004 , n348005 , n348006 , n348007 , n348008 , 
 n348009 , n348010 , n348011 , n348012 , n348013 , n348014 , n348015 , n348016 , n348017 , n348018 , 
 n348019 , n348020 , n348021 , n348022 , n348023 , n348024 , n348025 , n348026 , n348027 , n348028 , 
 n348029 , n348030 , n348031 , n348032 , n348033 , n348034 , n348035 , n348036 , n348037 , n348038 , 
 n348039 , n348040 , n348041 , n348042 , n348043 , n348044 , n348045 , n348046 , n348047 , n348048 , 
 n348049 , n348050 , n348051 , n348052 , n348053 , n348054 , n348055 , n348056 , n348057 , n348058 , 
 n348059 , n348060 , n348061 , n348062 , n348063 , n348064 , n348065 , n348066 , n348067 , n348068 , 
 n348069 , n348070 , n348071 , n348072 , n348073 , n348074 , n348075 , n348076 , n348077 , n348078 , 
 n348079 , n348080 , n348081 , n348082 , n348083 , n348084 , n348085 , n348086 , n348087 , n348088 , 
 n348089 , n348090 , n348091 , n348092 , n348093 , n348094 , n348095 , n348096 , n348097 , n348098 , 
 n348099 , n348100 , n348101 , n348102 , n348103 , n348104 , n348105 , n348106 , n348107 , n348108 , 
 n348109 , n348110 , n348111 , n348112 , n348113 , n348114 , n348115 , n348116 , n348117 , n348118 , 
 n348119 , n348120 , n348121 , n348122 , n348123 , n348124 , n348125 , n348126 , n348127 , n348128 , 
 n348129 , n348130 , n348131 , n348132 , n348133 , n348134 , n348135 , n348136 , n348137 , n348138 , 
 n348139 , n348140 , n348141 , n348142 , n348143 , n348144 , n348145 , n348146 , n348147 , n348148 , 
 n348149 , n348150 , n348151 , n348152 , n348153 , n348154 , n348155 , n348156 , n348157 , n348158 , 
 n348159 , n348160 , n348161 , n348162 , n348163 , n348164 , n348165 , n348166 , n348167 , n348168 , 
 n348169 , n348170 , n348171 , n348172 , n348173 , n348174 , n348175 , n348176 , n348177 , n348178 , 
 n348179 , n348180 , n348181 , n348182 , n348183 , n348184 , n348185 , n348186 , n348187 , n348188 , 
 n348189 , n348190 , n348191 , n348192 , n348193 , n348194 , n348195 , n348196 , n348197 , n348198 , 
 n348199 , n348200 , n348201 , n348202 , n348203 , n348204 , n348205 , n348206 , n348207 , n348208 , 
 n348209 , n348210 , n348211 , n348212 , n348213 , n348214 , n348215 , n348216 , n348217 , n348218 , 
 n348219 , n348220 , n348221 , n348222 , n348223 , n348224 , n348225 , n348226 , n348227 , n348228 , 
 n348229 , n348230 , n348231 , n348232 , n348233 , n348234 , n348235 , n348236 , n348237 , n348238 , 
 n348239 , n348240 , n348241 , n348242 , n348243 , n348244 , n348245 , n348246 , n348247 , n348248 , 
 n348249 , n348250 , n348251 , n348252 , n348253 , n348254 , n348255 , n348256 , n348257 , n348258 , 
 n348259 , n348260 , n348261 , n348262 , n348263 , n348264 , n348265 , n348266 , n348267 , n348268 , 
 n348269 , n348270 , n348271 , n348272 , n348273 , n348274 , n348275 , n348276 , n348277 , n348278 , 
 n348279 , n348280 , n348281 , n348282 , n348283 , n348284 , n348285 , n348286 , n348287 , n348288 , 
 n348289 , n348290 , n348291 , n348292 , n348293 , n348294 , n348295 , n348296 , n348297 , n348298 , 
 n348299 , n348300 , n348301 , n348302 , n348303 , n348304 , n348305 , n348306 , n348307 , n348308 , 
 n348309 , n348310 , n348311 , n348312 , n348313 , n348314 , n348315 , n348316 , n348317 , n348318 , 
 n348319 , n348320 , n348321 , n348322 , n348323 , n348324 , n348325 , n348326 , n348327 , n348328 , 
 n348329 , n348330 , n348331 , n348332 , n348333 , n348334 , n348335 , n348336 , n348337 , n348338 , 
 n348339 , n348340 , n348341 , n348342 , n348343 , n348344 , n348345 , n348346 , n348347 , n348348 , 
 n348349 , n348350 , n348351 , n348352 , n348353 , n348354 , n348355 , n348356 , n348357 , n348358 , 
 n348359 , n348360 , n348361 , n348362 , n348363 , n348364 , n348365 , n348366 , n348367 , n348368 , 
 n348369 , n348370 , n348371 , n348372 , n348373 , n348374 , n348375 , n348376 , n348377 , n348378 , 
 n348379 , n348380 , n348381 , n348382 , n348383 , n348384 , n348385 , n348386 , n348387 , n348388 , 
 n348389 , n348390 , n348391 , n348392 , n348393 , n348394 , n348395 , n348396 , n348397 , n348398 , 
 n348399 , n348400 , n348401 , n348402 , n348403 , n348404 , n348405 , n348406 , n348407 , n348408 , 
 n348409 , n348410 , n348411 , n348412 , n348413 , n348414 , n348415 , n348416 , n348417 , n348418 , 
 n348419 , n348420 , n348421 , n348422 , n348423 , n348424 , n348425 , n348426 , n348427 , n348428 , 
 n348429 , n348430 , n348431 , n348432 , n348433 , n348434 , n348435 , n348436 , n348437 , n348438 , 
 n348439 , n348440 , n348441 , n348442 , n348443 , n348444 , n348445 , n348446 , n348447 , n348448 , 
 n348449 , n348450 , n348451 , n348452 , n348453 , n348454 , n348455 , n348456 , n348457 , n348458 , 
 n348459 , n348460 , n348461 , n348462 , n348463 , n348464 , n348465 , n348466 , n348467 , n348468 , 
 n348469 , n348470 , n348471 , n348472 , n348473 , n348474 , n348475 , n348476 , n348477 , n348478 , 
 n348479 , n348480 , n348481 , n348482 , n348483 , n348484 , n348485 , n348486 , n348487 , n348488 , 
 n348489 , n348490 , n348491 , n348492 , n348493 , n348494 , n348495 , n348496 , n348497 , n348498 , 
 n348499 , n348500 , n348501 , n348502 , n348503 , n348504 , n348505 , n348506 , n348507 , n348508 , 
 n348509 , n348510 , n348511 , n348512 , n348513 , n348514 , n348515 , n348516 , n348517 , n348518 , 
 n348519 , n348520 , n348521 , n348522 , n348523 , n348524 , n348525 , n348526 , n348527 , n348528 , 
 n348529 , n348530 , n348531 , n348532 , n348533 , n348534 , n348535 , n348536 , n348537 , n348538 , 
 n348539 , n348540 , n348541 , n348542 , n348543 , n348544 , n348545 , n348546 , n348547 , n348548 , 
 n348549 , n348550 , n348551 , n348552 , n348553 , n348554 , n348555 , n348556 , n348557 , n348558 , 
 n348559 , n348560 , n348561 , n348562 , n348563 , n348564 , n348565 , n348566 , n348567 , n348568 , 
 n348569 , n348570 , n348571 , n348572 , n348573 , n348574 , n348575 , n348576 , n348577 , n348578 , 
 n348579 , n348580 , n348581 , n348582 , n835 , n348584 , n837 , n348586 , n839 , n348588 , 
 n841 , n348590 , n843 , n348592 , n845 , n348594 , n348595 , n848 , n348597 , n850 , 
 n851 , n852 , n348601 , n854 , n348603 , n348604 , n857 , n348606 , n859 , n348608 , 
 n348609 , n348610 , n348611 , n348612 , n865 , n348614 , n348615 , n868 , n348617 , n348618 , 
 n871 , n348620 , n348621 , n874 , n875 , n348624 , n348625 , n348626 , n348627 , n880 , 
 n348629 , n348630 , n348631 , n348632 , n348633 , n348634 , n348635 , n888 , n889 , n348638 , 
 n348639 , n348640 , n893 , n348642 , n895 , n348644 , n348645 , n348646 , n348647 , n348648 , 
 n348649 , n348650 , n903 , n348652 , n348653 , n906 , n348655 , n348656 , n909 , n348658 , 
 n348659 , n912 , n348661 , n914 , n915 , n348664 , n348665 , n918 , n348667 , n920 , 
 n921 , n922 , n923 , n924 , n925 , n926 , n348675 , n928 , n929 , n930 , 
 n931 , n348680 , n348681 , n934 , n348683 , n348684 , n937 , n348686 , n939 , n348688 , 
 n941 , n348690 , n943 , n944 , n945 , n348694 , n348695 , n948 , n348697 , n950 , 
 n951 , n952 , n348701 , n954 , n348703 , n348704 , n957 , n348706 , n959 , n960 , 
 n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , 
 n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , 
 n981 , n982 , n348731 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , 
 n991 , n992 , n993 , n994 , n995 , n348744 , n997 , n348746 , n999 , n1000 , 
 n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n348757 , n1010 , 
 n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , 
 n1021 , n1022 , n1023 , n348772 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , 
 n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , 
 n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , 
 n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , 
 n1061 , n1062 , n1063 , n1064 , n1065 , n1086 , n1091 , n1092 , n1093 , n1094 , 
 n1095 , n1096 , n1110 , n1111 , n1112 , n1114 , n1115 , n1116 , n1117 , n1118 , 
 n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n348835 , n1128 , n1129 , n1130 , 
 n1131 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , 
 n1142 , n1143 , n1144 , n1145 , n348853 , n1147 , n348855 , n348856 , n1150 , n348858 , 
 n348859 , n1153 , n1154 , n348862 , n348863 , n1157 , n348865 , n348866 , n1160 , n348868 , 
 n348869 , n1163 , n348871 , n348872 , n1166 , n1167 , n1171 , n1172 , n1173 , n1174 , 
 n1175 , n1176 , n1177 , n348882 , n1179 , n348884 , n1181 , n1182 , n1183 , n1184 , 
 n348889 , n348890 , n348891 , n1188 , n348893 , n348894 , n1191 , n348896 , n1193 , n348898 , 
 n348899 , n1196 , n348901 , n348902 , n1199 , n348904 , n348905 , n1202 , n348907 , n348908 , 
 n1205 , n348910 , n348911 , n1208 , n348913 , n348914 , n348915 , n1212 , n1213 , n1214 , 
 n1215 , n348920 , n1217 , n348922 , n348923 , n1220 , n348925 , n348926 , n348927 , n1224 , 
 n348929 , n1226 , n348931 , n348932 , n1229 , n348934 , n348935 , n348936 , n1233 , n348938 , 
 n348939 , n1236 , n348941 , n348942 , n348943 , n348944 , n348945 , n348946 , n348947 , n1244 , 
 n348949 , n1246 , n348951 , n1248 , n1249 , n1250 , n348955 , n1252 , n348957 , n348958 , 
 n1255 , n1256 , n348961 , n348962 , n1259 , n1260 , n348965 , n348966 , n1263 , n348968 , 
 n348969 , n1266 , n348971 , n348972 , n348973 , n1270 , n348975 , n348976 , n348977 , n1274 , 
 n348979 , n348980 , n1277 , n348982 , n1279 , n348984 , n348985 , n348986 , n1283 , n348988 , 
 n348989 , n1286 , n348991 , n348992 , n348993 , n348994 , n1291 , n1292 , n1296 , n1297 , 
 n1300 , n1301 , n349001 , n1303 , n1304 , n1305 , n349005 , n349006 , n1308 , n1309 , 
 n349009 , n349010 , n349011 , n1313 , n349013 , n349014 , n1316 , n349016 , n349017 , n1319 , 
 n349019 , n349020 , n1322 , n349022 , n349023 , n1325 , n349025 , n349026 , n1328 , n349028 , 
 n1330 , n349030 , n1332 , n1333 , n1334 , n1335 , n349035 , n349036 , n1338 , n1340 , 
 n1341 , n1342 , n1343 , n1344 , n1349 , n349044 , n349045 , n349046 , n349047 , n1354 , 
 n349049 , n349050 , n1357 , n349052 , n1359 , n1360 , n1361 , n1362 , n349057 , n1364 , 
 n1365 , n349060 , n1367 , n1368 , n1372 , n1375 , n349065 , n1377 , n349067 , n349068 , 
 n1380 , n349070 , n349071 , n1383 , n1384 , n349074 , n349075 , n1387 , n349077 , n349078 , 
 n1390 , n349080 , n349081 , n1393 , n1394 , n1395 , n1396 , n1397 , n349087 , n1399 , 
 n349089 , n349090 , n1402 , n349092 , n349093 , n1405 , n1406 , n349096 , n349097 , n1409 , 
 n349099 , n1411 , n349101 , n349102 , n1414 , n349104 , n1416 , n349106 , n349107 , n1419 , 
 n1420 , n349110 , n349111 , n1423 , n349113 , n349114 , n1426 , n349116 , n349117 , n349118 , 
 n1430 , n349120 , n349121 , n1433 , n349123 , n349124 , n1436 , n349126 , n349127 , n1439 , 
 n349129 , n349130 , n349131 , n1443 , n349133 , n1445 , n349135 , n1447 , n1448 , n349138 , 
 n349139 , n1451 , n349141 , n349142 , n1454 , n349144 , n349145 , n1457 , n1458 , n349148 , 
 n349149 , n349150 , n1462 , n1463 , n349153 , n349154 , n1466 , n349156 , n349157 , n349158 , 
 n1470 , n349160 , n349161 , n1473 , n349163 , n349164 , n1476 , n1477 , n349167 , n349168 , 
 n1480 , n349170 , n349171 , n1483 , n349173 , n349174 , n1486 , n349176 , n349177 , n1489 , 
 n349179 , n1491 , n349181 , n349182 , n349183 , n1495 , n349185 , n349186 , n1498 , n349188 , 
 n349189 , n1501 , n349191 , n1503 , n349193 , n1505 , n1506 , n349196 , n349197 , n1509 , 
 n349199 , n349200 , n1512 , n349202 , n349203 , n1515 , n1517 , n349206 , n349207 , n1520 , 
 n1521 , n1522 , n349211 , n349212 , n1525 , n349214 , n349215 , n1528 , n349217 , n1530 , 
 n349219 , n1532 , n1533 , n349222 , n1535 , n349224 , n1537 , n1538 , n349227 , n1540 , 
 n349229 , n349230 , n1543 , n349232 , n349233 , n1546 , n349235 , n1548 , n349237 , n349238 , 
 n1551 , n349240 , n349241 , n349242 , n1555 , n349244 , n349245 , n1558 , n349247 , n349248 , 
 n1561 , n1562 , n349251 , n349252 , n1565 , n1566 , n1567 , n349256 , n349257 , n349258 , 
 n349259 , n349260 , n1573 , n1574 , n349263 , n1576 , n349265 , n1578 , n1579 , n349268 , 
 n349269 , n1582 , n349271 , n349272 , n1585 , n349274 , n349275 , n349276 , n1589 , n349278 , 
 n349279 , n1592 , n349281 , n349282 , n1595 , n349284 , n1597 , n349286 , n1599 , n1600 , 
 n349289 , n349290 , n1603 , n1604 , n349293 , n349294 , n349295 , n1608 , n349297 , n1610 , 
 n1611 , n349300 , n1613 , n349302 , n1615 , n1616 , n349305 , n349306 , n1619 , n349308 , 
 n349309 , n1622 , n349311 , n349312 , n349313 , n1626 , n349315 , n349316 , n1629 , n349318 , 
 n349319 , n1632 , n349321 , n349322 , n1635 , n349324 , n349325 , n1638 , n1639 , n1640 , 
 n1641 , n349330 , n349331 , n1644 , n349333 , n1646 , n1647 , n1648 , n1649 , n1650 , 
 n1651 , n1652 , n1653 , n1654 , n349343 , n1656 , n349345 , n349346 , n1659 , n349348 , 
 n1661 , n349350 , n349351 , n349352 , n349353 , n1666 , n349355 , n349356 , n349357 , n1670 , 
 n349359 , n349360 , n349361 , n349362 , n349363 , n1676 , n349365 , n1678 , n349367 , n1680 , 
 n1681 , n349370 , n349371 , n1684 , n349373 , n349374 , n1687 , n349376 , n349377 , n1690 , 
 n1692 , n349380 , n349381 , n1695 , n1696 , n1697 , n349385 , n349386 , n1700 , n349388 , 
 n1702 , n349390 , n349391 , n1705 , n1706 , n1707 , n349395 , n349396 , n1710 , n1711 , 
 n1712 , n349400 , n349401 , n1715 , n1716 , n349404 , n1718 , n349406 , n1720 , n1721 , 
 n1722 , n349410 , n1724 , n349412 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , 
 n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , 
 n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , 
 n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , 
 n1762 , n1763 , n1764 , n1765 , n349453 , n1767 , n1768 , n1769 , n1770 , n1771 , 
 n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n349468 , 
 n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , 
 n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , 
 n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , 
 n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , 
 n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , 
 n349519 , n1833 , n1834 , n1835 , n1836 , n1837 , n349525 , n1839 , n349527 , n1841 , 
 n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , 
 n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , 
 n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , 
 n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , 
 n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , 
 n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , 
 n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , 
 n1912 , n1913 , n349601 , n1915 , n1916 , n1917 , n1918 , n1919 , n349607 , n1921 , 
 n349609 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , 
 n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , 
 n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , 
 n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , 
 n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , 
 n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , 
 n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , 
 n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , 
 n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , 
 n2012 , n2013 , n349701 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , 
 n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , 
 n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , 
 n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , 
 n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , 
 n2062 , n2063 , n2064 , n2065 , n2066 , n349754 , n2068 , n2069 , n2070 , n2071 , 
 n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , 
 n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , 
 n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , 
 n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , 
 n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , 
 n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , 
 n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , 
 n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , 
 n2152 , n2153 , n2154 , n2155 , n2156 , n349844 , n2158 , n2159 , n2160 , n2161 , 
 n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , 
 n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n349868 , 
 n2182 , n349870 , n2184 , n349872 , n349873 , n349874 , n2188 , n349876 , n349877 , n349878 , 
 n2192 , n349880 , n349881 , n2195 , n349883 , n349884 , n349885 , n349886 , n2200 , n349888 , 
 n2202 , n349890 , n349891 , n349892 , n349893 , n2207 , n349895 , n349896 , n349897 , n2211 , 
 n349899 , n349900 , n2214 , n2215 , n349903 , n2217 , n349905 , n349906 , n2220 , n2221 , 
 n349909 , n2223 , n349911 , n349912 , n2226 , n349914 , n349915 , n2229 , n2230 , n2231 , 
 n2232 , n2233 , n2234 , n2235 , n2236 , n349924 , n2238 , n2239 , n2240 , n2241 , 
 n2242 , n2243 , n349931 , n2245 , n349933 , n349934 , n349935 , n349936 , n2250 , n349938 , 
 n349939 , n2253 , n349941 , n349942 , n2256 , n349944 , n349945 , n2259 , n349947 , n2261 , 
 n349949 , n2263 , n2264 , n349952 , n349953 , n349954 , n2268 , n349956 , n349957 , n2271 , 
 n349959 , n349960 , n2274 , n349962 , n349963 , n2277 , n349965 , n349966 , n2280 , n2281 , 
 n349969 , n349970 , n2284 , n349972 , n349973 , n2287 , n349975 , n349976 , n2290 , n349978 , 
 n349979 , n349980 , n2294 , n349982 , n2296 , n2297 , n349985 , n349986 , n349987 , n2301 , 
 n349989 , n349990 , n2304 , n349992 , n349993 , n2307 , n349995 , n349996 , n2310 , n2311 , 
 n349999 , n2313 , n350001 , n350002 , n2316 , n2317 , n350005 , n2319 , n2320 , n2321 , 
 n2322 , n2323 , n350011 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , 
 n350019 , n2333 , n2334 , n350022 , n2336 , n2337 , n2338 , n2339 , n2340 , n350028 , 
 n350029 , n2343 , n2344 , n350032 , n350033 , n2347 , n350035 , n2349 , n2350 , n350038 , 
 n350039 , n2353 , n350041 , n350042 , n2356 , n350044 , n350045 , n2359 , n350047 , n350048 , 
 n2362 , n350050 , n2364 , n350052 , n350053 , n350054 , n350055 , n2369 , n350057 , n350058 , 
 n350059 , n2373 , n350061 , n350062 , n2376 , n350064 , n2378 , n350066 , n2380 , n2381 , 
 n350069 , n350070 , n2384 , n350072 , n350073 , n350074 , n2388 , n350076 , n350077 , n2391 , 
 n350079 , n350080 , n2394 , n2395 , n350083 , n350084 , n2398 , n2399 , n350087 , n350088 , 
 n350089 , n2403 , n350091 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , 
 n350099 , n2413 , n350101 , n2415 , n350103 , n350104 , n2418 , n350106 , n350107 , n350108 , 
 n2422 , n350110 , n350111 , n2425 , n2426 , n350114 , n350115 , n350116 , n2430 , n350118 , 
 n350119 , n2433 , n350121 , n350122 , n2436 , n350124 , n350125 , n350126 , n2440 , n350128 , 
 n2442 , n350130 , n350131 , n2445 , n350133 , n350134 , n2448 , n2449 , n350137 , n350138 , 
 n350139 , n2453 , n350141 , n350142 , n2456 , n350144 , n350145 , n2459 , n350147 , n350148 , 
 n2462 , n350150 , n350151 , n2465 , n350153 , n350154 , n2468 , n2469 , n2470 , n2471 , 
 n350159 , n2473 , n2474 , n350162 , n350163 , n350164 , n2478 , n350166 , n350167 , n2481 , 
 n350169 , n350170 , n2484 , n350172 , n350173 , n2487 , n350175 , n350176 , n2490 , n350178 , 
 n350179 , n2493 , n350181 , n350182 , n2496 , n350184 , n350185 , n2499 , n2500 , n2501 , 
 n2502 , n2503 , n2504 , n2505 , n2506 , n350194 , n2508 , n350196 , n350197 , n2511 , 
 n350199 , n350200 , n350201 , n350202 , n350203 , n2517 , n350205 , n350206 , n350207 , n2521 , 
 n350209 , n350210 , n2524 , n350212 , n350213 , n350214 , n2528 , n350216 , n2530 , n350218 , 
 n350219 , n2533 , n350221 , n350222 , n2536 , n350224 , n350225 , n2539 , n350227 , n350228 , 
 n2542 , n350230 , n350231 , n2545 , n350233 , n2547 , n2548 , n2549 , n2550 , n350238 , 
 n350239 , n2553 , n350241 , n350242 , n350243 , n2557 , n350245 , n2559 , n2560 , n350248 , 
 n350249 , n2563 , n350251 , n350252 , n350253 , n2567 , n350255 , n350256 , n2570 , n350258 , 
 n350259 , n2573 , n350261 , n2575 , n350263 , n2577 , n2578 , n2579 , n350267 , n350268 , 
 n350269 , n2583 , n350271 , n350272 , n2586 , n350274 , n350275 , n2589 , n350277 , n350278 , 
 n2592 , n350280 , n350281 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , 
 n2602 , n350290 , n2604 , n350292 , n2606 , n350294 , n2608 , n2609 , n350297 , n350298 , 
 n350299 , n2613 , n350301 , n350302 , n2616 , n350304 , n350305 , n2619 , n350307 , n350308 , 
 n350309 , n2623 , n350311 , n2625 , n2626 , n350314 , n350315 , n350316 , n2630 , n350318 , 
 n350319 , n2633 , n350321 , n350322 , n2636 , n350324 , n350325 , n2639 , n350327 , n350328 , 
 n2642 , n350330 , n350331 , n2645 , n350333 , n350334 , n2648 , n350336 , n2650 , n2651 , 
 n2652 , n2653 , n2654 , n350342 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , 
 n2662 , n2663 , n2664 , n2665 , n2666 , n350354 , n2668 , n350356 , n2670 , n350358 , 
 n2672 , n350360 , n2674 , n2675 , n2676 , n2677 , n350365 , n350366 , n2680 , n350368 , 
 n350369 , n2683 , n350371 , n350372 , n2686 , n350374 , n350375 , n2689 , n350377 , n350378 , 
 n350379 , n2693 , n350381 , n350382 , n350383 , n2697 , n350385 , n2699 , n2700 , n350388 , 
 n350389 , n2703 , n350391 , n350392 , n350393 , n2707 , n350395 , n350396 , n2710 , n350398 , 
 n350399 , n2713 , n350401 , n2715 , n350403 , n2717 , n2718 , n350406 , n350407 , n350408 , 
 n2722 , n350410 , n350411 , n2725 , n350413 , n350414 , n2728 , n350416 , n350417 , n2731 , 
 n350419 , n350420 , n2734 , n2735 , n2736 , n2737 , n350425 , n350426 , n2740 , n350428 , 
 n2742 , n350430 , n2744 , n2745 , n350433 , n350434 , n350435 , n2749 , n350437 , n350438 , 
 n2752 , n350440 , n350441 , n2755 , n350443 , n350444 , n2758 , n350446 , n350447 , n2761 , 
 n350449 , n2763 , n350451 , n2765 , n2766 , n350454 , n350455 , n350456 , n2770 , n350458 , 
 n350459 , n2773 , n350461 , n350462 , n2776 , n350464 , n350465 , n2779 , n2780 , n350468 , 
 n2782 , n350470 , n2784 , n2785 , n350473 , n2787 , n350475 , n350476 , n350477 , n2791 , 
 n2792 , n350480 , n350481 , n350482 , n2796 , n350484 , n2798 , n350486 , n350487 , n2801 , 
 n350489 , n350490 , n2804 , n350492 , n350493 , n2807 , n350495 , n350496 , n2810 , n350498 , 
 n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , 
 n350509 , n2823 , n2824 , n350512 , n2826 , n2827 , n2828 , n350516 , n2830 , n2831 , 
 n350519 , n2833 , n2834 , n2835 , n2836 , n350524 , n2838 , n350526 , n350527 , n2841 , 
 n350529 , n350530 , n350531 , n2845 , n350533 , n350534 , n2848 , n2849 , n2850 , n2851 , 
 n350539 , n2853 , n2854 , n350542 , n350543 , n350544 , n2858 , n350546 , n350547 , n2861 , 
 n350549 , n350550 , n2864 , n350552 , n2866 , n350554 , n2868 , n350556 , n2870 , n2871 , 
 n350559 , n350560 , n2874 , n350562 , n350563 , n350564 , n2878 , n350566 , n350567 , n2881 , 
 n350569 , n2883 , n350571 , n2885 , n2886 , n2887 , n2888 , n350576 , n350577 , n2891 , 
 n350579 , n2893 , n350581 , n2895 , n2896 , n350584 , n350585 , n350586 , n2900 , n350588 , 
 n350589 , n2903 , n350591 , n350592 , n2906 , n350594 , n350595 , n2909 , n2910 , n2911 , 
 n350599 , n350600 , n350601 , n2915 , n350603 , n350604 , n2918 , n350606 , n2920 , n350608 , 
 n350609 , n2923 , n350611 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , 
 n2932 , n350620 , n2934 , n2935 , n2936 , n2937 , n2938 , n350626 , n350627 , n2941 , 
 n350629 , n350630 , n2944 , n350632 , n350633 , n2947 , n2948 , n2949 , n2950 , n350638 , 
 n350639 , n2953 , n2954 , n2955 , n2956 , n2957 , n350645 , n350646 , n2960 , n2961 , 
 n2962 , n2963 , n350651 , n350652 , n2966 , n350654 , n2968 , n350656 , n2970 , n2971 , 
 n350659 , n2973 , n350661 , n350662 , n350663 , n350664 , n2978 , n350666 , n350667 , n2981 , 
 n350669 , n350670 , n350671 , n2985 , n350673 , n2987 , n2988 , n350676 , n350677 , n2991 , 
 n350679 , n350680 , n350681 , n2995 , n350683 , n350684 , n2998 , n350686 , n350687 , n350688 , 
 n350689 , n3003 , n350691 , n350692 , n3006 , n3007 , n3008 , n3009 , n350697 , n3011 , 
 n350699 , n350700 , n3014 , n3015 , n350703 , n3017 , n350705 , n350706 , n350707 , n350708 , 
 n3022 , n350710 , n350711 , n3025 , n350713 , n350714 , n3028 , n350716 , n350717 , n3031 , 
 n350719 , n3033 , n350721 , n3035 , n3036 , n350724 , n3038 , n350726 , n350727 , n350728 , 
 n350729 , n3043 , n350731 , n350732 , n3046 , n350734 , n350735 , n3049 , n350737 , n350738 , 
 n3052 , n350740 , n350741 , n3055 , n350743 , n3057 , n350745 , n3059 , n3060 , n350748 , 
 n3062 , n3063 , n3064 , n3065 , n3066 , n350754 , n3068 , n350756 , n350757 , n3071 , 
 n350759 , n350760 , n350761 , n350762 , n3076 , n350764 , n3078 , n350766 , n350767 , n350768 , 
 n350769 , n3083 , n350771 , n350772 , n350773 , n3087 , n350775 , n350776 , n3090 , n3091 , 
 n3092 , n3093 , n350781 , n3095 , n3096 , n350784 , n350785 , n350786 , n3100 , n350788 , 
 n350789 , n3103 , n350791 , n350792 , n3106 , n350794 , n3108 , n350796 , n3110 , n3111 , 
 n3112 , n3113 , n3114 , n350802 , n350803 , n3117 , n350805 , n350806 , n3120 , n350808 , 
 n350809 , n3123 , n350811 , n350812 , n3126 , n350814 , n350815 , n3129 , n3130 , n3131 , 
 n3132 , n3133 , n3134 , n350822 , n3136 , n350824 , n3138 , n3139 , n3140 , n350828 , 
 n350829 , n3143 , n350831 , n350832 , n350833 , n3147 , n350835 , n350836 , n3150 , n350838 , 
 n350839 , n3153 , n350841 , n350842 , n3156 , n350844 , n3158 , n3159 , n3160 , n3161 , 
 n3162 , n350850 , n3164 , n350852 , n3166 , n350854 , n3168 , n3169 , n3170 , n3171 , 
 n3172 , n3173 , n3174 , n350862 , n350863 , n3177 , n350865 , n350866 , n3180 , n350868 , 
 n350869 , n3183 , n3184 , n350872 , n3186 , n350874 , n350875 , n3189 , n3190 , n3191 , 
 n3192 , n3193 , n350881 , n3195 , n350883 , n3197 , n350885 , n3199 , n350887 , n3201 , 
 n3202 , n350890 , n350891 , n350892 , n3206 , n350894 , n350895 , n3209 , n350897 , n350898 , 
 n3212 , n350900 , n3214 , n350902 , n3216 , n3217 , n3218 , n3219 , n350907 , n350908 , 
 n3222 , n3223 , n3224 , n3225 , n3226 , n350914 , n350915 , n3229 , n350917 , n3231 , 
 n350919 , n3233 , n3234 , n3235 , n350923 , n350924 , n3238 , n350926 , n3240 , n3241 , 
 n3242 , n3243 , n3244 , n350932 , n350933 , n3247 , n350935 , n3249 , n3250 , n3251 , 
 n3252 , n3253 , n3254 , n350942 , n350943 , n350944 , n3258 , n350946 , n350947 , n3261 , 
 n350949 , n3263 , n3264 , n350952 , n3266 , n350954 , n3268 , n350956 , n3270 , n350958 , 
 n350959 , n3273 , n3274 , n3275 , n3276 , n350964 , n350965 , n3279 , n3280 , n3281 , 
 n3282 , n3283 , n350971 , n350972 , n3286 , n3287 , n3288 , n3289 , n350977 , n350978 , 
 n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , 
 n3302 , n3303 , n3304 , n3305 , n350993 , n350994 , n3308 , n350996 , n3310 , n3311 , 
 n3312 , n3313 , n3314 , n351002 , n351003 , n351004 , n3318 , n351006 , n351007 , n3321 , 
 n351009 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , 
 n351019 , n3333 , n3334 , n3335 , n3336 , n351024 , n351025 , n3339 , n351027 , n351028 , 
 n3342 , n351030 , n351031 , n3345 , n351033 , n3347 , n351035 , n351036 , n3350 , n351038 , 
 n351039 , n351040 , n3354 , n351042 , n351043 , n3357 , n351045 , n3359 , n3360 , n3361 , 
 n3362 , n3363 , n351051 , n351052 , n3366 , n351054 , n3368 , n351056 , n3370 , n351058 , 
 n3372 , n351060 , n3374 , n351062 , n3376 , n3377 , n351065 , n351066 , n351067 , n3381 , 
 n351069 , n351070 , n3384 , n351072 , n351073 , n3387 , n351075 , n3389 , n351077 , n3391 , 
 n3392 , n3393 , n3394 , n3395 , n351083 , n351084 , n3398 , n351086 , n351087 , n3401 , 
 n351089 , n351090 , n3404 , n351092 , n351093 , n3407 , n351095 , n3409 , n3410 , n351098 , 
 n3412 , n351100 , n351101 , n3415 , n351103 , n3417 , n3418 , n3419 , n3420 , n3421 , 
 n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n351116 , n3430 , n351118 , 
 n3432 , n351120 , n3434 , n351122 , n3436 , n351124 , n3438 , n351126 , n351127 , n351128 , 
 n3442 , n351130 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , 
 n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , 
 n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , 
 n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , 
 n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , 
 n351179 , n3493 , n351181 , n3495 , n351183 , n351184 , n3498 , n351186 , n3500 , n3501 , 
 n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , 
 n3512 , n3513 , n351201 , n351202 , n351203 , n3517 , n351205 , n351206 , n3520 , n351208 , 
 n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , 
 n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , 
 n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3551 , n3552 , n3553 , n3554 , 
 n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , 
 n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , 
 n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , 
 n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n351275 , n3592 , n351277 , n3594 , 
 n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , 
 n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n351295 , n351296 , n3613 , n351298 , 
 n351299 , n351300 , n351301 , n3618 , n351303 , n351304 , n3621 , n351306 , n3623 , n3624 , 
 n3625 , n3626 , n3627 , n3628 , n3629 , n351314 , n351315 , n3632 , n351317 , n351318 , 
 n3635 , n351320 , n3637 , n351322 , n351323 , n3640 , n351325 , n3642 , n351327 , n351328 , 
 n3645 , n351330 , n351331 , n3648 , n3649 , n3650 , n351335 , n351336 , n351337 , n3654 , 
 n351339 , n351340 , n3657 , n351342 , n351343 , n3660 , n351345 , n351346 , n351347 , n3664 , 
 n351349 , n3666 , n3667 , n351352 , n351353 , n351354 , n3671 , n351356 , n351357 , n3674 , 
 n351359 , n351360 , n3677 , n351362 , n351363 , n3680 , n351365 , n351366 , n3683 , n351368 , 
 n3685 , n351370 , n351371 , n351372 , n351373 , n3690 , n351375 , n351376 , n351377 , n3694 , 
 n351379 , n351380 , n351381 , n3698 , n351383 , n3700 , n3701 , n351386 , n3703 , n351388 , 
 n3705 , n351390 , n351391 , n3708 , n351393 , n351394 , n3711 , n351396 , n351397 , n3714 , 
 n351399 , n351400 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , 
 n3725 , n351410 , n3727 , n351412 , n3729 , n351414 , n3731 , n3732 , n351417 , n351418 , 
 n3735 , n351420 , n3737 , n351422 , n351423 , n3740 , n351425 , n351426 , n351427 , n3744 , 
 n351429 , n3746 , n3747 , n3748 , n3749 , n351434 , n3751 , n351436 , n351437 , n3754 , 
 n3755 , n351440 , n351441 , n3758 , n351443 , n3760 , n3761 , n3762 , n3763 , n3764 , 
 n3765 , n351450 , n3767 , n3768 , n3769 , n3770 , n351455 , n351456 , n351457 , n3774 , 
 n351459 , n351460 , n3777 , n351462 , n3779 , n351464 , n3781 , n351466 , n3783 , n351468 , 
 n3785 , n3786 , n351471 , n3788 , n351473 , n3790 , n351475 , n351476 , n3793 , n351478 , 
 n351479 , n3796 , n351481 , n351482 , n3799 , n351484 , n351485 , n3802 , n351487 , n351488 , 
 n3805 , n3806 , n3807 , n3808 , n351493 , n351494 , n3811 , n3812 , n3813 , n3814 , 
 n3815 , n351500 , n351501 , n3818 , n3819 , n3820 , n3821 , n351506 , n351507 , n3824 , 
 n351509 , n351510 , n3827 , n351512 , n3829 , n351514 , n351515 , n351516 , n351517 , n3834 , 
 n351519 , n351520 , n351521 , n3838 , n351523 , n351524 , n3841 , n351526 , n3843 , n3844 , 
 n351529 , n351530 , n351531 , n3848 , n351533 , n351534 , n3851 , n351536 , n351537 , n3854 , 
 n351539 , n3856 , n3857 , n351542 , n351543 , n3860 , n351545 , n3862 , n3863 , n3864 , 
 n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n351557 , n3874 , 
 n351559 , n351560 , n351561 , n351562 , n3879 , n351564 , n351565 , n3882 , n351567 , n3884 , 
 n3885 , n3886 , n3887 , n351572 , n351573 , n351574 , n3891 , n351576 , n351577 , n3894 , 
 n351579 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , 
 n3905 , n351590 , n3907 , n3908 , n3909 , n3910 , n351595 , n351596 , n3913 , n3914 , 
 n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , 
 n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n351618 , 
 n351619 , n351620 , n3937 , n351622 , n351623 , n3940 , n351625 , n3942 , n3943 , n351628 , 
 n351629 , n3946 , n351631 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n351638 , 
 n3955 , n351640 , n351641 , n3958 , n351643 , n351644 , n3961 , n351646 , n351647 , n3964 , 
 n351649 , n3966 , n3967 , n3968 , n3969 , n351654 , n351655 , n3972 , n351657 , n3974 , 
 n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n351666 , n3983 , n351668 , 
 n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , 
 n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , 
 n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , 
 n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , 
 n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , 
 n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n351725 , n351726 , n351727 , n351728 , 
 n4045 , n351730 , n351731 , n4048 , n351733 , n351734 , n4051 , n351736 , n351737 , n4054 , 
 n351739 , n351740 , n4057 , n351742 , n351743 , n4060 , n351745 , n351746 , n4063 , n351748 , 
 n351749 , n4066 , n351751 , n351752 , n4069 , n351754 , n351755 , n4072 , n351757 , n351758 , 
 n4075 , n351760 , n351761 , n4078 , n351763 , n351764 , n4081 , n351766 , n351767 , n4084 , 
 n351769 , n351770 , n4087 , n351772 , n351773 , n4090 , n4091 , n4092 , n4093 , n4094 , 
 n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , 
 n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , 
 n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , 
 n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , 
 n4135 , n351820 , n351821 , n4138 , n351823 , n4140 , n351825 , n4142 , n4143 , n351828 , 
 n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , 
 n4155 , n4156 , n4157 , n4158 , n4159 , n351844 , n351845 , n4162 , n351847 , n4164 , 
 n351849 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , 
 n4175 , n4176 , n4177 , n4178 , n4179 , n351864 , n4181 , n4182 , n4183 , n351868 , 
 n4185 , n351870 , n351871 , n4188 , n351873 , n351874 , n351875 , n4192 , n4193 , n351878 , 
 n4195 , n351880 , n351881 , n4198 , n351883 , n351884 , n351885 , n4202 , n351887 , n4204 , 
 n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , 
 n4215 , n4216 , n351901 , n351902 , n351903 , n4220 , n4221 , n351906 , n351907 , n4224 , 
 n351909 , n351910 , n4227 , n351912 , n351913 , n351914 , n351915 , n351916 , n351917 , n351918 , 
 n351919 , n4236 , n351921 , n351922 , n4239 , n351924 , n351925 , n4242 , n351927 , n351928 , 
 n4245 , n351930 , n351931 , n4248 , n351933 , n4250 , n351935 , n4252 , n4253 , n351938 , 
 n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , 
 n4266 , n351950 , n4268 , n351952 , n351953 , n4271 , n4272 , n351956 , n4274 , n351958 , 
 n351959 , n351960 , n4278 , n351962 , n351963 , n351964 , n351965 , n351966 , n4284 , n4285 , 
 n351969 , n351970 , n4288 , n351972 , n351973 , n4291 , n351975 , n351976 , n351977 , n4295 , 
 n351979 , n4297 , n4298 , n351982 , n4300 , n4301 , n351985 , n351986 , n4304 , n351988 , 
 n351989 , n4307 , n351991 , n351992 , n4310 , n4311 , n351995 , n351996 , n351997 , n351998 , 
 n351999 , n4317 , n352001 , n352002 , n352003 , n352004 , n4322 , n352006 , n352007 , n4325 , 
 n4326 , n4328 , n352011 , n352012 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , 
 n352019 , n4338 , n352021 , n4340 , n352023 , n4342 , n352025 , n4344 , n352027 , n352028 , 
 n4347 , n4348 , n4349 , n4350 , n4351 , n352034 , n352035 , n4354 , n352037 , n352038 , 
 n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n352045 , n4364 , n352047 , n4366 , 
 n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , 
 n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n352065 , n352066 , n352067 , n4386 , 
 n4387 , n4388 , n352071 , n352072 , n4391 , n352074 , n352075 , n4394 , n352077 , n352078 , 
 n4397 , n4398 , n352081 , n4400 , n4401 , n352084 , n4403 , n352086 , n4405 , n4406 , 
 n4407 , n4408 , n4409 , n4410 , n352093 , n4412 , n352095 , n352096 , n4415 , n4416 , 
 n352099 , n352100 , n352101 , n352102 , n352103 , n4422 , n352105 , n352106 , n4425 , n352108 , 
 n352109 , n352110 , n4429 , n352112 , n352113 , n352114 , n352115 , n4434 , n352117 , n352118 , 
 n4437 , n4438 , n352121 , n352122 , n4441 , n352124 , n4443 , n352126 , n4445 , n352128 , 
 n352129 , n4448 , n352131 , n352132 , n4451 , n352134 , n352135 , n4454 , n4455 , n4456 , 
 n352139 , n352140 , n4459 , n352142 , n352143 , n4462 , n352145 , n4464 , n352147 , n4466 , 
 n352149 , n352150 , n4469 , n352152 , n4471 , n4472 , n4473 , n4474 , n4475 , n352158 , 
 n4477 , n352160 , n352161 , n4480 , n352163 , n4482 , n4483 , n4484 , n4485 , n4486 , 
 n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n352175 , n352176 , n352177 , n4496 , 
 n352179 , n352180 , n4499 , n352182 , n4501 , n4502 , n4503 , n4504 , n4505 , n352188 , 
 n352189 , n352190 , n4509 , n352192 , n352193 , n352194 , n352195 , n4514 , n4515 , n4516 , 
 n352199 , n352200 , n4519 , n352202 , n352203 , n352204 , n352205 , n4524 , n352207 , n352208 , 
 n352209 , n4528 , n352211 , n4530 , n4531 , n352214 , n4533 , n352216 , n4535 , n352218 , 
 n352219 , n4538 , n352221 , n352222 , n4541 , n352224 , n4543 , n352226 , n4545 , n352228 , 
 n352229 , n352230 , n352231 , n4550 , n352233 , n352234 , n4553 , n352236 , n352237 , n4556 , 
 n352239 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , 
 n4567 , n4568 , n352251 , n352252 , n4571 , n352254 , n4573 , n4574 , n4575 , n4576 , 
 n352259 , n4578 , n352261 , n352262 , n352263 , n352264 , n4583 , n352266 , n4585 , n4586 , 
 n4587 , n4588 , n352271 , n4590 , n4591 , n352274 , n4593 , n4594 , n352277 , n4596 , 
 n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , 
 n4607 , n4608 , n4609 , n4610 , n352293 , n4612 , n352295 , n4614 , n352297 , n352298 , 
 n4617 , n352300 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , 
 n352309 , n352310 , n4629 , n352312 , n4631 , n4632 , n4633 , n4634 , n352317 , n352318 , 
 n352319 , n4638 , n352321 , n352322 , n4641 , n352324 , n4643 , n4644 , n352327 , n352328 , 
 n352329 , n4648 , n352331 , n352332 , n4651 , n352334 , n352335 , n4654 , n352337 , n352338 , 
 n4657 , n352340 , n4659 , n352342 , n352343 , n4662 , n352345 , n352346 , n352347 , n4666 , 
 n352349 , n352350 , n4669 , n352352 , n352353 , n4672 , n352355 , n352356 , n4675 , n352358 , 
 n352359 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n352366 , n4685 , n4686 , 
 n4687 , n352370 , n352371 , n4690 , n352373 , n4692 , n4693 , n352376 , n4695 , n352378 , 
 n4697 , n352380 , n4699 , n4700 , n352383 , n352384 , n352385 , n4704 , n352387 , n352388 , 
 n4707 , n352390 , n352391 , n4710 , n352393 , n352394 , n4713 , n352396 , n352397 , n4716 , 
 n352399 , n4718 , n352401 , n4720 , n4721 , n352404 , n352405 , n4724 , n352407 , n352408 , 
 n4727 , n352410 , n352411 , n4730 , n4731 , n4732 , n4733 , n352416 , n352417 , n4736 , 
 n4737 , n352420 , n352421 , n4740 , n4741 , n4742 , n352425 , n352426 , n4745 , n352428 , 
 n4747 , n4748 , n4749 , n4750 , n4751 , n352434 , n4753 , n4754 , n4755 , n4756 , 
 n352439 , n352440 , n4759 , n4760 , n4761 , n4762 , n352445 , n352446 , n4765 , n352448 , 
 n4767 , n352450 , n4769 , n4770 , n352453 , n352454 , n352455 , n4774 , n352457 , n352458 , 
 n4777 , n352460 , n352461 , n4780 , n352463 , n352464 , n352465 , n352466 , n352467 , n352468 , 
 n352469 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n352478 , 
 n4797 , n352480 , n352481 , n4800 , n4801 , n4802 , n4803 , n352486 , n4805 , n352488 , 
 n352489 , n4808 , n352491 , n352492 , n352493 , n4812 , n352495 , n352496 , n4815 , n352498 , 
 n4817 , n352500 , n4819 , n4820 , n352503 , n352504 , n4823 , n352506 , n4825 , n352508 , 
 n4827 , n352510 , n352511 , n4830 , n352513 , n352514 , n4833 , n4834 , n352517 , n352518 , 
 n352519 , n4838 , n352521 , n352522 , n4841 , n352524 , n352525 , n4844 , n352527 , n352528 , 
 n352529 , n4848 , n352531 , n4850 , n4851 , n352534 , n4853 , n4854 , n4855 , n4856 , 
 n352539 , n4858 , n352541 , n352542 , n4861 , n352544 , n352545 , n4864 , n352547 , n352548 , 
 n4867 , n4868 , n352551 , n4870 , n4871 , n352554 , n4873 , n4874 , n352557 , n4876 , 
 n352559 , n4878 , n4879 , n352562 , n352563 , n4882 , n352565 , n352566 , n352567 , n4886 , 
 n352569 , n352570 , n4889 , n352572 , n352573 , n352574 , n4893 , n352576 , n4895 , n4896 , 
 n352579 , n352580 , n352581 , n4900 , n352583 , n352584 , n4903 , n352586 , n352587 , n4906 , 
 n352589 , n352590 , n4909 , n352592 , n4911 , n352594 , n4913 , n352596 , n352597 , n352598 , 
 n352599 , n4918 , n352601 , n352602 , n4921 , n352604 , n352605 , n352606 , n352607 , n352608 , 
 n4927 , n352610 , n4929 , n4930 , n4931 , n4932 , n4933 , n352616 , n4935 , n352618 , 
 n4937 , n352620 , n352621 , n4940 , n352623 , n4942 , n4943 , n352626 , n352627 , n4946 , 
 n352629 , n352630 , n352631 , n352632 , n4951 , n4952 , n4953 , n4954 , n4955 , n352638 , 
 n4957 , n352640 , n352641 , n4960 , n4961 , n4962 , n352645 , n352646 , n4965 , n4966 , 
 n4967 , n4968 , n4969 , n352652 , n4971 , n4972 , n4973 , n352656 , n4975 , n4976 , 
 n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , 
 n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n352675 , n4994 , n4995 , n4996 , 
 n4997 , n352680 , n352681 , n5000 , n352683 , n5002 , n352685 , n5004 , n5005 , n352688 , 
 n5007 , n352690 , n352691 , n352692 , n5011 , n352694 , n5013 , n352696 , n352697 , n5016 , 
 n352699 , n352700 , n352701 , n5020 , n352703 , n5022 , n5023 , n352706 , n5025 , n352708 , 
 n352709 , n352710 , n5029 , n352712 , n5031 , n352714 , n352715 , n5034 , n352717 , n352718 , 
 n352719 , n5038 , n352721 , n5040 , n352723 , n352724 , n352725 , n5044 , n352727 , n5046 , 
 n352729 , n5048 , n352731 , n5050 , n5051 , n352734 , n352735 , n5054 , n352737 , n352738 , 
 n352739 , n5058 , n352741 , n352742 , n5061 , n352744 , n5063 , n5064 , n5065 , n5066 , 
 n5067 , n5068 , n352751 , n5070 , n352753 , n352754 , n5073 , n352756 , n5075 , n5076 , 
 n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n352765 , n5084 , n5085 , n5086 , 
 n5087 , n352770 , n352771 , n5090 , n352773 , n5092 , n5093 , n5094 , n352777 , n352778 , 
 n5097 , n352780 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , 
 n5107 , n352790 , n352791 , n352792 , n5111 , n352794 , n352795 , n5114 , n352797 , n5116 , 
 n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , 
 n5127 , n352810 , n352811 , n5130 , n352813 , n5132 , n5133 , n352816 , n352817 , n352818 , 
 n5137 , n352820 , n352821 , n5140 , n352823 , n352824 , n5143 , n352826 , n352827 , n5146 , 
 n352829 , n352830 , n5149 , n352832 , n352833 , n5152 , n5153 , n5154 , n5155 , n5156 , 
 n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n352845 , n5164 , n5165 , n352848 , 
 n352849 , n352850 , n5169 , n352852 , n352853 , n5172 , n352855 , n352856 , n5175 , n352858 , 
 n352859 , n5178 , n352861 , n5180 , n352863 , n5182 , n352865 , n5184 , n352867 , n352868 , 
 n5187 , n5188 , n352871 , n5190 , n352873 , n352874 , n5193 , n352876 , n5195 , n5196 , 
 n352879 , n5198 , n352881 , n352882 , n5201 , n352884 , n5203 , n352886 , n5205 , n352888 , 
 n352889 , n5208 , n352891 , n352892 , n5211 , n352894 , n5213 , n5214 , n5215 , n5216 , 
 n5217 , n5218 , n5219 , n5220 , n352903 , n5222 , n5223 , n5224 , n5225 , n352908 , 
 n352909 , n5228 , n5229 , n5230 , n352913 , n352914 , n5233 , n5234 , n5235 , n352918 , 
 n5237 , n5238 , n5239 , n352922 , n5241 , n5242 , n5243 , n5244 , n352927 , n5246 , 
 n5247 , n5248 , n5249 , n352932 , n5251 , n5252 , n5253 , n352936 , n5255 , n5256 , 
 n5257 , n5258 , n5259 , n5260 , n5261 , n352944 , n5263 , n352946 , n352947 , n5266 , 
 n352949 , n5268 , n352951 , n352952 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , 
 n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n352967 , n5286 , 
 n352969 , n352970 , n352971 , n5290 , n5291 , n352974 , n5293 , n5294 , n352977 , n352978 , 
 n352979 , n5298 , n352981 , n352982 , n5301 , n352984 , n352985 , n5304 , n352987 , n352988 , 
 n352989 , n5308 , n352991 , n5310 , n5311 , n352994 , n352995 , n352996 , n5315 , n352998 , 
 n352999 , n5318 , n353001 , n353002 , n5321 , n353004 , n353005 , n5324 , n353007 , n353008 , 
 n5327 , n353010 , n353011 , n5330 , n353013 , n5332 , n5333 , n5334 , n5335 , n5336 , 
 n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n353025 , n353026 , n353027 , n5346 , 
 n353029 , n353030 , n5349 , n353032 , n5351 , n5352 , n5353 , n5354 , n5355 , n353038 , 
 n353039 , n353040 , n5359 , n353042 , n353043 , n5362 , n353045 , n5364 , n5365 , n5366 , 
 n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n353057 , n353058 , 
 n5377 , n353060 , n5379 , n353062 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , 
 n353069 , n5388 , n5389 , n5390 , n5391 , n353074 , n353075 , n5394 , n353077 , n353078 , 
 n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , 
 n5407 , n353090 , n353091 , n5410 , n353093 , n5412 , n353095 , n5414 , n353097 , n5416 , 
 n5417 , n353100 , n353101 , n353102 , n5421 , n353104 , n353105 , n5424 , n353107 , n353108 , 
 n5427 , n353110 , n5429 , n353112 , n5431 , n5432 , n353115 , n5434 , n353117 , n353118 , 
 n5437 , n5438 , n353121 , n353122 , n5441 , n5442 , n5443 , n5444 , n353127 , n353128 , 
 n5447 , n5448 , n353131 , n5450 , n353133 , n353134 , n5453 , n5454 , n353137 , n353138 , 
 n5457 , n5458 , n353141 , n5460 , n353143 , n353144 , n5463 , n5464 , n353147 , n5466 , 
 n5467 , n5468 , n5469 , n353152 , n5471 , n353154 , n5473 , n5474 , n5475 , n5476 , 
 n353159 , n353160 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , 
 n5487 , n5488 , n5489 , n5490 , n353173 , n5492 , n353175 , n5494 , n353177 , n5496 , 
 n5497 , n353180 , n353181 , n5500 , n353183 , n5502 , n353185 , n353186 , n5505 , n353188 , 
 n353189 , n353190 , n353191 , n5510 , n353193 , n353194 , n353195 , n5514 , n353197 , n353198 , 
 n5517 , n353200 , n353201 , n5520 , n353203 , n5522 , n5523 , n5524 , n5525 , n353208 , 
 n5527 , n353210 , n5529 , n353212 , n5531 , n5532 , n353215 , n353216 , n5535 , n353218 , 
 n5537 , n353220 , n5539 , n353222 , n353223 , n5542 , n353225 , n353226 , n5545 , n5546 , 
 n5547 , n5548 , n353231 , n5550 , n5551 , n5552 , n5553 , n5554 , n353237 , n353238 , 
 n5557 , n353240 , n353241 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , 
 n5567 , n353250 , n5569 , n5570 , n353253 , n5572 , n5573 , n353256 , n353257 , n353258 , 
 n5577 , n353260 , n353261 , n5580 , n353263 , n353264 , n5583 , n353266 , n353267 , n5586 , 
 n353269 , n5588 , n5589 , n353272 , n353273 , n353274 , n5593 , n353276 , n353277 , n5596 , 
 n353279 , n353280 , n5599 , n353282 , n353283 , n5602 , n353285 , n5604 , n5605 , n5606 , 
 n5607 , n5608 , n353291 , n353292 , n5611 , n353294 , n5613 , n5614 , n5615 , n5616 , 
 n5617 , n5618 , n5619 , n5620 , n5621 , n353304 , n5623 , n353306 , n5625 , n5626 , 
 n353309 , n353310 , n353311 , n5630 , n353313 , n353314 , n5633 , n353316 , n353317 , n5636 , 
 n353319 , n353320 , n353321 , n5640 , n353323 , n5642 , n5643 , n5644 , n5645 , n5646 , 
 n353329 , n5648 , n353331 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , 
 n5657 , n5658 , n353341 , n5660 , n353343 , n5662 , n5663 , n5664 , n5665 , n5666 , 
 n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n353358 , 
 n5677 , n353360 , n5679 , n353362 , n5681 , n353364 , n353365 , n5684 , n5685 , n5686 , 
 n5687 , n353370 , n353371 , n5690 , n353373 , n353374 , n5693 , n353376 , n353377 , n353378 , 
 n353379 , n5698 , n353381 , n353382 , n5701 , n353384 , n353385 , n5704 , n353387 , n353388 , 
 n5707 , n353390 , n353391 , n5710 , n5711 , n353394 , n5713 , n5714 , n353397 , n5716 , 
 n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , 
 n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , 
 n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , 
 n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , 
 n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , 
 n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , 
 n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n353465 , n353466 , n5785 , n5786 , 
 n5787 , n353470 , n353471 , n5790 , n353473 , n353474 , n5793 , n5794 , n5795 , n353478 , 
 n353479 , n5798 , n353481 , n353482 , n5801 , n5802 , n5803 , n353486 , n353487 , n5806 , 
 n353489 , n353490 , n5809 , n5810 , n5811 , n353494 , n353495 , n5814 , n353497 , n353498 , 
 n5817 , n5818 , n5819 , n353502 , n353503 , n5822 , n353505 , n353506 , n5825 , n5826 , 
 n5827 , n353510 , n353511 , n5830 , n353513 , n353514 , n5833 , n5834 , n5835 , n353518 , 
 n353519 , n5838 , n353521 , n353522 , n5841 , n5842 , n5843 , n353526 , n353527 , n5846 , 
 n353529 , n353530 , n5849 , n5850 , n5851 , n353534 , n353535 , n5854 , n353537 , n353538 , 
 n5857 , n5858 , n5859 , n353542 , n353543 , n5862 , n353545 , n353546 , n5865 , n5866 , 
 n5867 , n353550 , n353551 , n5870 , n353553 , n353554 , n5873 , n5874 , n5875 , n353558 , 
 n353559 , n5878 , n353561 , n353562 , n5881 , n5882 , n5883 , n353566 , n353567 , n5886 , 
 n353569 , n353570 , n5889 , n5890 , n5891 , n353574 , n353575 , n5894 , n353577 , n353578 , 
 n5897 , n5898 , n5899 , n353582 , n353583 , n5902 , n353585 , n353586 , n5905 , n5906 , 
 n5907 , n353590 , n353591 , n5910 , n353593 , n353594 , n5913 , n5914 , n5915 , n353598 , 
 n353599 , n5918 , n353601 , n353602 , n5921 , n5922 , n5923 , n353606 , n353607 , n5926 , 
 n353609 , n353610 , n5929 , n5930 , n5931 , n353614 , n353615 , n5934 , n353617 , n353618 , 
 n5937 , n5938 , n5939 , n353622 , n353623 , n5942 , n353625 , n353626 , n5945 , n5946 , 
 n5947 , n353630 , n353631 , n5950 , n353633 , n353634 , n5953 , n5954 , n5955 , n353638 , 
 n353639 , n5958 , n353641 , n353642 , n5961 , n5962 , n5963 , n353646 , n353647 , n5966 , 
 n353649 , n353650 , n5969 , n5970 , n5971 , n353654 , n353655 , n5974 , n353657 , n353658 , 
 n5977 , n5978 , n5979 , n353662 , n353663 , n5982 , n353665 , n353666 , n5985 , n5986 , 
 n5987 , n353670 , n353671 , n5990 , n353673 , n353674 , n5993 , n5994 , n5995 , n353678 , 
 n353679 , n5998 , n353681 , n353682 , n6001 , n6002 , n6003 , n353686 , n353687 , n6006 , 
 n353689 , n353690 , n6009 , n6010 , n6011 , n353694 , n353695 , n6014 , n353697 , n353698 , 
 n6017 , n6018 , n6019 , n353702 , n353703 , n6022 , n353705 , n353706 , n6025 , n6026 , 
 n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , 
 n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , 
 n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , 
 n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , 
 n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , 
 n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , 
 n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , 
 n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , 
 n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , 
 n6117 , n6118 , n6119 , n6120 , n353803 , n353804 , n353805 , n353806 , n353807 , n353808 , 
 n353809 , n353810 , n353811 , n353812 , n353813 , n353814 , n353815 , n353816 , n353817 , n353818 , 
 n353819 , n353820 , n353821 , n353822 , n353823 , n353824 , n353825 , n353826 , n353827 , n353828 , 
 n353829 , n353830 , n353831 , n353832 , n353833 , n353834 , n353835 , n353836 , n353837 , n353838 , 
 n353839 , n353840 , n353841 , n353842 , n353843 , n353844 , n353845 , n353846 , n353847 , n353848 , 
 n353849 , n353850 , n353851 , n353852 , n353853 , n353854 , n353855 , n353856 , n353857 , n353858 , 
 n353859 , n353860 , n353861 , n353862 , n353863 , n353864 , n353865 , n353866 , n353867 , n353868 , 
 n353869 , n353870 , n353871 , n353872 , n353873 , n353874 , n353875 , n353876 , n353877 , n353878 , 
 n353879 , n353880 , n353881 , n353882 , n353883 , n353884 , n353885 , n353886 , n353887 , n353888 , 
 n353889 , n353890 , n353891 , n353892 , n353893 , n353894 , n353895 , n353896 , n353897 , n353898 , 
 n353899 , n353900 , n353901 , n353902 , n353903 , n353904 , n353905 , n353906 , n353907 , n353908 , 
 n353909 , n353910 , n353911 , n353912 , n353913 , n353914 , n353915 , n353916 , n353917 , n353918 , 
 n353919 , n353920 , n353921 , n353922 , n353923 , n353924 , n353925 , n353926 , n353927 , n353928 , 
 n353929 , n353930 , n353931 , n353932 , n353933 , n353934 , n353935 , n353936 , n353937 , n353938 , 
 n353939 , n353940 , n353941 , n353942 , n353943 , n353944 , n353945 , n353946 , n353947 , n353948 , 
 n353949 , n353950 , n353951 , n353952 , n353953 , n353954 , n353955 , n353956 , n353957 , n353958 , 
 n353959 , n353960 , n353961 , n353962 , n353963 , n353964 , n353965 , n353966 , n353967 , n353968 , 
 n353969 , n353970 , n353971 , n353972 , n353973 , n353974 , n353975 , n353976 , n353977 , n353978 , 
 n353979 , n353980 , n353981 , n353982 , n353983 , n353984 , n353985 , n353986 , n353987 , n353988 , 
 n353989 , n353990 , n353991 , n353992 , n353993 , n353994 , n6311 , n6312 , n353997 , n353998 , 
 n6315 , n6316 , n354001 , n354002 , n6319 , n6320 , n354005 , n354006 , n6323 , n6324 , 
 n354009 , n354010 , n6327 , n6328 , n354013 , n354014 , n6331 , n6332 , n354017 , n354018 , 
 n6335 , n6336 , n354021 , n354022 , n6339 , n6340 , n354025 , n354026 , n6343 , n6344 , 
 n354029 , n354030 , n6347 , n6348 , n354033 , n354034 , n6351 , n6352 , n354037 , n354038 , 
 n6355 , n6356 , n354041 , n354042 , n6359 , n6360 , n354045 , n354046 , n6363 , n6364 , 
 n354049 , n354050 , n354051 , n6368 , n354053 , n354054 , n6371 , n354056 , n354057 , n354058 , 
 n6375 , n354060 , n354061 , n354062 , n354063 , n354064 , n6381 , n354066 , n354067 , n354068 , 
 n354069 , n354070 , n6387 , n6388 , n354073 , n354074 , n354075 , n6392 , n6393 , n6394 , 
 n354079 , n354080 , n354081 , n6398 , n6399 , n6400 , n354085 , n354086 , n354087 , n354088 , 
 n6405 , n6406 , n354091 , n354092 , n354093 , n354094 , n354095 , n6412 , n354097 , n354098 , 
 n354099 , n354100 , n354101 , n354102 , n354103 , n354104 , n354105 , n6422 , n354107 , n6424 , 
 n354109 , n354110 , n354111 , n6428 , n354113 , n354114 , n354115 , n354116 , n354117 , n6434 , 
 n354119 , n354120 , n354121 , n354122 , n354123 , n6440 , n6441 , n354126 , n354127 , n354128 , 
 n354129 , n6446 , n6447 , n6448 , n354133 , n354134 , n354135 , n6452 , n6453 , n6454 , 
 n354139 , n354140 , n354141 , n6458 , n6459 , n6460 , n354145 , n354146 , n354147 , n6464 , 
 n354149 , n6466 , n6467 , n6468 , n6469 , n6470 , n354155 , n354156 , n354157 , n6474 , 
 n354159 , n6476 , n354161 , n6478 , n6479 , n354164 , n354165 , n6482 , n354167 , n354168 , 
 n6485 , n354170 , n354171 , n6488 , n6489 , n354174 , n354175 , n6492 , n354177 , n354178 , 
 n6495 , n354180 , n354181 , n6498 , n354183 , n6500 , n6501 , n6502 , n6503 , n6504 , 
 n354189 , n6506 , n6507 , n354192 , n354193 , n6510 , n354195 , n354196 , n6513 , n354198 , 
 n354199 , n354200 , n354201 , n6518 , n354203 , n354204 , n6521 , n354206 , n6523 , n354208 , 
 n6525 , n6526 , n354211 , n6528 , n354213 , n354214 , n354215 , n6532 , n354217 , n354218 , 
 n6535 , n354220 , n6537 , n6538 , n6539 , n6540 , n6541 , n354226 , n6543 , n6544 , 
 n6545 , n6546 , n6547 , n354232 , n354233 , n6550 , n354235 , n354236 , n6553 , n354238 , 
 n6555 , n354240 , n6557 , n354242 , n6559 , n6560 , n6561 , n354246 , n6563 , n354248 , 
 n354249 , n6566 , n354251 , n354252 , n354253 , n6570 , n354255 , n354256 , n6573 , n354258 , 
 n354259 , n6576 , n6577 , n354262 , n354263 , n6580 , n354265 , n354266 , n6583 , n354268 , 
 n354269 , n6586 , n354271 , n354272 , n6589 , n354274 , n354275 , n6592 , n354277 , n354278 , 
 n6595 , n354280 , n354281 , n6598 , n6599 , n6600 , n354285 , n6602 , n6603 , n6604 , 
 n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , 
 n6615 , n6616 , n354301 , n354302 , n354303 , n354304 , n354305 , n6618 , n354307 , n354308 , 
 n6621 , n354310 , n354311 , n354312 , n354313 , n354314 , n354315 , n354316 , n354317 , n6630 , 
 n354319 , n354320 , n6633 , n354322 , n354323 , n6636 , n354325 , n354326 , n6639 , n354328 , 
 n354329 , n6642 , n354331 , n354332 , n6645 , n354334 , n354335 , n354336 , n354337 , n354338 , 
 n6651 , n354340 , n354341 , n354342 , n354343 , n354344 , n354345 , n354346 , n354347 , n6660 , 
 n354349 , n354350 , n6663 , n354352 , n354353 , n6666 , n354355 , n354356 , n6669 , n354358 , 
 n354359 , n6672 , n354361 , n354362 , n354363 , n354364 , n354365 , n354366 , n354367 , n354368 , 
 n6681 , n354370 , n354371 , n354372 , n354373 , n354374 , n354375 , n354376 , n354377 , n354378 , 
 n354379 , n354380 , n354381 , n354382 , n354383 , n354384 , n354385 , n354386 , n6699 , n354388 , 
 n354389 , n6702 , n354391 , n354392 , n6705 , n354394 , n354395 , n354396 , n354397 , n354398 , 
 n354399 , n354400 , n354401 , n6714 , n354403 , n354404 , n6717 , n354406 , n354407 , n6720 , 
 n354409 , n354410 , n6723 , n354412 , n354413 , n354414 , n354415 , n354416 , n6729 , n354418 , 
 n354419 , n6732 , n354421 , n354422 , n354423 , n354424 , n354425 , n354426 , n354427 , n354428 , 
 n354429 , n354430 , n354431 , n354432 , n354433 , n354434 , n6747 , n354436 , n354437 , n6750 , 
 n354439 , n354440 , n6753 , n354442 , n354443 , n354444 , n354445 , n354446 , n354447 , n354448 , 
 n354449 , n6762 , n354451 , n354452 , n6765 , n354454 , n354455 , n6768 , n354457 , n354458 , 
 n6771 , n354460 , n354461 , n354462 , n354463 , n354464 , n6777 , n354466 , n354467 , n6780 , 
 n354469 , n354470 , n354471 , n354472 , n354473 , n6786 , n354475 , n354476 , n6789 , n354478 , 
 n354479 , n6792 , n354481 , n354482 , n354483 , n354484 , n354485 , n354486 , n354487 , n354488 , 
 n354489 , n354490 , n354491 , n354492 , n354493 , n354494 , n354495 , n354496 , n354497 , n6810 , 
 n354499 , n354500 , n354501 , n354502 , n354503 , n354504 , n354505 , n354506 , n6819 , n354508 , 
 n354509 , n6822 , n354511 , n354512 , n354513 , n354514 , n354515 , n354516 , n354517 , n354518 , 
 n354519 , n354520 , n354521 , n6834 , n354523 , n354524 , n6837 , n354526 , n354527 , n6840 , 
 n354529 , n354530 , n354531 , n354532 , n354533 , n354534 , n354535 , n354536 , n354537 , n354538 , 
 n354539 , n6852 , n354541 , n354542 , n6855 , n354544 , n354545 , n6858 , n354547 , n354548 , 
 n354549 , n354550 , n354551 , n6864 , n354553 , n354554 , n6867 , n354556 , n354557 , n6870 , 
 n354559 , n354560 , n6873 , n354562 , n354563 , n354564 , n354565 , n354566 , n354567 , n354568 , 
 n354569 , n354570 , n354571 , n354572 , n6885 , n354574 , n354575 , n6888 , n354577 , n354578 , 
 n6891 , n354580 , n354581 , n354582 , n354583 , n354584 , n6897 , n354586 , n354587 , n6900 , 
 n354589 , n354590 , n354591 , n354592 , n354593 , n354594 , n354595 , n354596 , n354597 , n354598 , 
 n354599 , n354600 , n354601 , n354602 , n354603 , n354604 , n354605 , n6918 , n354607 , n354608 , 
 n354609 , n354610 , n354611 , n6924 , n354613 , n354614 , n6927 , n354616 , n354617 , n6930 , 
 n354619 , n354620 , n6933 , n354622 , n354623 , n6936 , n354625 , n354626 , n6939 , n354628 , 
 n354629 , n354630 , n354631 , n354632 , n6945 , n354634 , n354635 , n354636 , n354637 , n354638 , 
 n354639 , n354640 , n354641 , n354642 , n354643 , n354644 , n354645 , n354646 , n354647 , n6960 , 
 n354649 , n354650 , n6963 , n6964 , n354653 , n354654 , n6967 , n6968 , n354657 , n354658 , 
 n6971 , n6972 , n354661 , n354662 , n6975 , n6976 , n354665 , n354666 , n6979 , n6980 , 
 n354669 , n354670 , n6983 , n354672 , n354673 , n354674 , n354675 , n6988 , n354677 , n354678 , 
 n354679 , n6992 , n354681 , n354682 , n354683 , n354684 , n354685 , n354686 , n354687 , n354688 , 
 n354689 , n354690 , n7003 , n7004 , n354693 , n354694 , n354695 , n7008 , n354697 , n354698 , 
 n354699 , n354700 , n354701 , n354702 , n7015 , n7016 , n7017 , n354706 , n354707 , n354708 , 
 n7021 , n354710 , n354711 , n7024 , n354713 , n7026 , n7027 , n354716 , n7029 , n354718 , 
 n354719 , n7032 , n354721 , n354722 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , 
 n7041 , n7042 , n7043 , n7044 , n7045 , n354734 , n7047 , n7048 , n7049 , n7050 , 
 n7051 , n7052 , n7053 , n7054 , n7055 , n354744 , n354745 , n354746 , n7059 , n354748 , 
 n7061 , n354750 , n354751 , n354752 , n354753 , n7066 , n354755 , n354756 , n354757 , n7070 , 
 n354759 , n354760 , n354761 , n7074 , n354763 , n7076 , n7077 , n354766 , n354767 , n7080 , 
 n354769 , n354770 , n354771 , n7084 , n354773 , n354774 , n7087 , n354776 , n354777 , n7090 , 
 n354779 , n354780 , n354781 , n7094 , n354783 , n7096 , n7097 , n354786 , n7099 , n354788 , 
 n354789 , n7102 , n354791 , n7104 , n354793 , n354794 , n7107 , n354796 , n354797 , n7110 , 
 n7111 , n7112 , n7113 , n7114 , n354803 , n354804 , n7117 , n354806 , n354807 , n7120 , 
 n7121 , n7122 , n7123 , n7124 , n354813 , n354814 , n7127 , n354816 , n354817 , n7130 , 
 n354819 , n354820 , n7133 , n354822 , n354823 , n7136 , n354825 , n354826 , n7139 , n7140 , 
 n7141 , n7142 , n354831 , n354832 , n7145 , n354834 , n7147 , n354836 , n7149 , n354838 , 
 n354839 , n354840 , n7153 , n354842 , n354843 , n7156 , n354845 , n7158 , n7159 , n7160 , 
 n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , 
 n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , 
 n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , 
 n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , 
 n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , 
 n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , 
 n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , 
 n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , 
 n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , 
 n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , 
 n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , 
 n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , 
 n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , 
 n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , 
 n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , 
 n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , 
 n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , 
 n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , 
 n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , 
 n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , 
 n7361 , n7362 , n7363 , n7364 , n7365 , n355054 , n7367 , n7368 , n7369 , n7370 , 
 n7371 , n7372 , n355061 , n355062 , n355063 , n7376 , n355065 , n355066 , n355067 , n7380 , 
 n355069 , n355070 , n7383 , n355072 , n355073 , n7386 , n355075 , n355076 , n7389 , n355078 , 
 n355079 , n7392 , n355081 , n355082 , n355083 , n7396 , n355085 , n7398 , n355087 , n7400 , 
 n355089 , n355090 , n7403 , n7404 , n355093 , n7406 , n355095 , n7408 , n355097 , n355098 , 
 n7411 , n355100 , n355101 , n7414 , n7415 , n355104 , n7417 , n355106 , n7419 , n7420 , 
 n355109 , n355110 , n7423 , n355112 , n355113 , n7426 , n355115 , n355116 , n355117 , n7430 , 
 n355119 , n355120 , n7433 , n355122 , n355123 , n7436 , n7437 , n355126 , n355127 , n7440 , 
 n355129 , n7442 , n355131 , n7444 , n7445 , n355134 , n7447 , n7448 , n355137 , n355138 , 
 n7451 , n355140 , n355141 , n7454 , n355143 , n355144 , n7457 , n7458 , n355147 , n7460 , 
 n355149 , n7462 , n7463 , n355152 , n355153 , n7466 , n355155 , n355156 , n7469 , n355158 , 
 n355159 , n355160 , n7473 , n355162 , n355163 , n7476 , n355165 , n355166 , n7479 , n7480 , 
 n7481 , n355170 , n355171 , n355172 , n7485 , n355174 , n7487 , n355176 , n7489 , n355178 , 
 n355179 , n7492 , n7493 , n355182 , n355183 , n7496 , n355185 , n355186 , n7499 , n355188 , 
 n355189 , n7502 , n7503 , n355192 , n7505 , n355194 , n7507 , n7508 , n355197 , n355198 , 
 n7511 , n355200 , n355201 , n7514 , n355203 , n355204 , n355205 , n7518 , n355207 , n355208 , 
 n7521 , n355210 , n355211 , n7524 , n355213 , n7526 , n355215 , n7528 , n7529 , n355218 , 
 n355219 , n7532 , n355221 , n355222 , n7535 , n355224 , n355225 , n355226 , n7539 , n355228 , 
 n7541 , n7542 , n355231 , n355232 , n7545 , n355234 , n355235 , n7548 , n355237 , n355238 , 
 n7551 , n7552 , n7553 , n355242 , n355243 , n7556 , n355245 , n355246 , n7559 , n7560 , 
 n7561 , n355250 , n355251 , n7564 , n7565 , n7566 , n7567 , n7568 , n355257 , n355258 , 
 n7571 , n7572 , n355261 , n355262 , n7575 , n355264 , n7577 , n355266 , n7579 , n7580 , 
 n355269 , n355270 , n7583 , n355272 , n355273 , n7586 , n355275 , n355276 , n7589 , n355278 , 
 n355279 , n7592 , n7593 , n7594 , n355283 , n355284 , n7597 , n7598 , n7599 , n7600 , 
 n7601 , n355290 , n355291 , n355292 , n7605 , n7606 , n7607 , n7608 , n7609 , n355298 , 
 n355299 , n355300 , n7613 , n355302 , n7615 , n355304 , n355305 , n7618 , n355307 , n7620 , 
 n7621 , n355310 , n355311 , n7624 , n355313 , n7626 , n355315 , n355316 , n7629 , n355318 , 
 n7631 , n7632 , n355321 , n7634 , n355323 , n7636 , n7637 , n355326 , n7639 , n355328 , 
 n7641 , n7642 , n355331 , n355332 , n7645 , n355334 , n7647 , n7648 , n7649 , n355338 , 
 n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n355348 , 
 n7661 , n355350 , n7663 , n7664 , n7665 , n7666 , n355355 , n7668 , n355357 , n355358 , 
 n7671 , n355360 , n355361 , n7674 , n7675 , n355364 , n355365 , n7678 , n355367 , n355368 , 
 n355369 , n7682 , n355371 , n7684 , n7685 , n355374 , n7687 , n355376 , n7689 , n7690 , 
 n355379 , n7692 , n355381 , n7694 , n7695 , n355384 , n355385 , n355386 , n7699 , n355388 , 
 n355389 , n7702 , n355391 , n355392 , n7705 , n355394 , n7707 , n7708 , n7709 , n7710 , 
 n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n355405 , n355406 , n355407 , n7720 , 
 n355409 , n355410 , n7723 , n355412 , n7725 , n355414 , n7727 , n355416 , n7729 , n7730 , 
 n355419 , n355420 , n355421 , n7734 , n355423 , n355424 , n7737 , n355426 , n355427 , n7740 , 
 n355429 , n7742 , n355431 , n7744 , n355433 , n7746 , n7747 , n355436 , n355437 , n355438 , 
 n7751 , n355440 , n355441 , n7754 , n355443 , n355444 , n7757 , n355446 , n7759 , n355448 , 
 n7761 , n355450 , n7763 , n7764 , n355453 , n355454 , n7767 , n355456 , n7769 , n355458 , 
 n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n355468 , 
 n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n355478 , 
 n7791 , n355480 , n7793 , n355482 , n7795 , n7796 , n355485 , n355486 , n355487 , n7800 , 
 n355489 , n355490 , n7803 , n355492 , n355493 , n7806 , n355495 , n355496 , n7809 , n355498 , 
 n355499 , n7812 , n355501 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , 
 n355509 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , 
 n355519 , n355520 , n7833 , n355522 , n355523 , n7836 , n355525 , n7838 , n7839 , n355528 , 
 n355529 , n7842 , n355531 , n7844 , n355533 , n355534 , n7847 , n355536 , n7849 , n355538 , 
 n7851 , n355540 , n355541 , n7854 , n355543 , n355544 , n7857 , n7858 , n355547 , n7860 , 
 n355549 , n7862 , n355551 , n355552 , n7865 , n355554 , n7867 , n7868 , n7869 , n355558 , 
 n355559 , n355560 , n7873 , n355562 , n355563 , n7876 , n355565 , n7878 , n7879 , n7880 , 
 n7881 , n7882 , n355571 , n7884 , n355573 , n7886 , n355575 , n7888 , n7889 , n355578 , 
 n7891 , n355580 , n7893 , n7894 , n355583 , n355584 , n7897 , n355586 , n355587 , n7900 , 
 n355589 , n355590 , n355591 , n7904 , n355593 , n7906 , n355595 , n7908 , n355597 , n7910 , 
 n7911 , n355600 , n355601 , n7914 , n355603 , n355604 , n355605 , n7918 , n355607 , n355608 , 
 n7921 , n355610 , n7923 , n7924 , n7925 , n355614 , n7927 , n355616 , n7929 , n7930 , 
 n355619 , n355620 , n355621 , n7934 , n355623 , n355624 , n7937 , n355626 , n355627 , n7940 , 
 n355629 , n355630 , n355631 , n7944 , n355633 , n7946 , n7947 , n355636 , n355637 , n355638 , 
 n7951 , n355640 , n355641 , n7954 , n355643 , n355644 , n7957 , n355646 , n355647 , n7960 , 
 n355649 , n7962 , n355651 , n7964 , n7965 , n355654 , n355655 , n355656 , n7969 , n355658 , 
 n355659 , n7972 , n355661 , n355662 , n7975 , n355664 , n355665 , n7978 , n355667 , n355668 , 
 n7981 , n355670 , n7983 , n355672 , n7985 , n7986 , n7987 , n7988 , n355677 , n355678 , 
 n7991 , n7992 , n7993 , n7994 , n7995 , n355684 , n355685 , n355686 , n7999 , n355688 , 
 n8001 , n8002 , n355691 , n8004 , n355693 , n355694 , n355695 , n8008 , n355697 , n8010 , 
 n355699 , n355700 , n8013 , n355702 , n355703 , n8016 , n8017 , n355706 , n355707 , n8020 , 
 n8021 , n8022 , n8023 , n355712 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , 
 n8031 , n355720 , n8033 , n355722 , n355723 , n8036 , n355725 , n355726 , n8039 , n355728 , 
 n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , 
 n355739 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n355746 , n8059 , n355748 , 
 n355749 , n8062 , n355751 , n355752 , n355753 , n8066 , n355755 , n355756 , n8069 , n8070 , 
 n355759 , n355760 , n8073 , n355762 , n355763 , n8076 , n355765 , n8078 , n355767 , n355768 , 
 n8081 , n355770 , n355771 , n8084 , n355773 , n355774 , n355775 , n355776 , n8089 , n355778 , 
 n8091 , n355780 , n355781 , n355782 , n355783 , n355784 , n8097 , n355786 , n355787 , n8100 , 
 n355789 , n355790 , n8103 , n355792 , n355793 , n8106 , n355795 , n8108 , n8109 , n8110 , 
 n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , 
 n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , 
 n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , 
 n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , 
 n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , 
 n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , 
 n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , 
 n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , 
 n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , 
 n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , 
 n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , 
 n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , 
 n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , 
 n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , 
 n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , 
 n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , 
 n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , 
 n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , 
 n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , 
 n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , 
 n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , 
 n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , 
 n8331 , n8332 , n8333 , n8334 , n8335 , n356024 , n8337 , n8338 , n356027 , n356028 , 
 n8341 , n356030 , n356031 , n8344 , n356033 , n356034 , n8347 , n356036 , n8349 , n356038 , 
 n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , 
 n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , 
 n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , 
 n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , 
 n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , 
 n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , 
 n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , 
 n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , 
 n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , 
 n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , 
 n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , 
 n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , 
 n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , 
 n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , 
 n8491 , n8492 , n8493 , n8494 , n356183 , n356184 , n356185 , n356186 , n8499 , n356188 , 
 n356189 , n8502 , n8503 , n356192 , n356193 , n8506 , n356195 , n8508 , n8509 , n8510 , 
 n8511 , n356200 , n8513 , n356202 , n356203 , n8516 , n356205 , n356206 , n8519 , n356208 , 
 n8521 , n356210 , n8523 , n8524 , n356213 , n356214 , n356215 , n8528 , n356217 , n356218 , 
 n8531 , n356220 , n356221 , n8534 , n356223 , n356224 , n8537 , n356226 , n8539 , n8540 , 
 n356229 , n356230 , n356231 , n8544 , n356233 , n356234 , n8547 , n356236 , n356237 , n8550 , 
 n356239 , n8552 , n356241 , n8554 , n356243 , n8556 , n8557 , n356246 , n8559 , n356248 , 
 n8561 , n356250 , n356251 , n8564 , n356253 , n8566 , n8567 , n8568 , n8569 , n8570 , 
 n356259 , n8572 , n8573 , n8574 , n8575 , n356264 , n8577 , n356266 , n356267 , n8580 , 
 n8581 , n8582 , n8583 , n356272 , n8585 , n356274 , n356275 , n8588 , n8589 , n356278 , 
 n8591 , n8592 , n356281 , n8594 , n8595 , n356284 , n8597 , n356286 , n8599 , n8600 , 
 n356289 , n8602 , n8603 , n8604 , n356293 , n8606 , n8607 , n356296 , n356297 , n356298 , 
 n8611 , n356300 , n356301 , n8614 , n356303 , n356304 , n8617 , n356306 , n356307 , n8620 , 
 n356309 , n8622 , n8623 , n356312 , n356313 , n356314 , n8627 , n356316 , n356317 , n8630 , 
 n356319 , n356320 , n8633 , n356322 , n8635 , n356324 , n8637 , n356326 , n8639 , n8640 , 
 n356329 , n356330 , n356331 , n8644 , n356333 , n356334 , n8647 , n356336 , n356337 , n8650 , 
 n356339 , n8652 , n356341 , n8654 , n356343 , n356344 , n8657 , n356346 , n356347 , n8660 , 
 n8661 , n356350 , n356351 , n8664 , n356353 , n356354 , n8667 , n356356 , n356357 , n8670 , 
 n8671 , n356360 , n8673 , n356362 , n8675 , n356364 , n356365 , n8678 , n8679 , n8680 , 
 n8681 , n8682 , n356371 , n356372 , n8685 , n356374 , n8687 , n8688 , n8689 , n8690 , 
 n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n356385 , n8698 , n356387 , n8700 , 
 n356389 , n356390 , n8703 , n356392 , n8705 , n8706 , n356395 , n356396 , n8709 , n356398 , 
 n8711 , n356400 , n356401 , n8714 , n356403 , n356404 , n8717 , n356406 , n8719 , n356408 , 
 n8721 , n8722 , n356411 , n356412 , n8725 , n356414 , n8727 , n356416 , n356417 , n8730 , 
 n356419 , n356420 , n8733 , n8734 , n8735 , n8736 , n356425 , n356426 , n8739 , n356428 , 
 n356429 , n8742 , n356431 , n356432 , n356433 , n8746 , n356435 , n8748 , n356437 , n356438 , 
 n8751 , n356440 , n356441 , n8754 , n8755 , n356444 , n8757 , n356446 , n356447 , n8760 , 
 n356449 , n8762 , n356451 , n356452 , n8765 , n356454 , n356455 , n8768 , n356457 , n356458 , 
 n356459 , n8772 , n356461 , n8774 , n8775 , n356464 , n8777 , n356466 , n8779 , n356468 , 
 n356469 , n8782 , n356471 , n356472 , n8785 , n356474 , n356475 , n8788 , n356477 , n8790 , 
 n8791 , n356480 , n356481 , n356482 , n8795 , n356484 , n356485 , n8798 , n356487 , n356488 , 
 n8801 , n356490 , n8803 , n8804 , n8805 , n8806 , n356495 , n356496 , n8809 , n356498 , 
 n356499 , n356500 , n8813 , n356502 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , 
 n8821 , n356510 , n8823 , n8824 , n8825 , n8826 , n8827 , n356516 , n356517 , n8830 , 
 n356519 , n356520 , n8833 , n8834 , n8835 , n8836 , n356525 , n356526 , n8839 , n356528 , 
 n8841 , n356530 , n8843 , n8844 , n356533 , n8846 , n356535 , n8848 , n356537 , n356538 , 
 n8851 , n356540 , n356541 , n356542 , n8855 , n356544 , n8857 , n8858 , n356547 , n8860 , 
 n356549 , n8862 , n356551 , n356552 , n8865 , n356554 , n356555 , n8868 , n356557 , n8870 , 
 n356559 , n8872 , n8873 , n356562 , n8875 , n356564 , n8877 , n356566 , n356567 , n8880 , 
 n356569 , n356570 , n8883 , n356572 , n356573 , n8886 , n356575 , n356576 , n356577 , n8890 , 
 n356579 , n8892 , n356581 , n356582 , n8895 , n8896 , n8897 , n8898 , n356587 , n8900 , 
 n356589 , n356590 , n8903 , n356592 , n8905 , n356594 , n8907 , n356596 , n8909 , n356598 , 
 n356599 , n8912 , n8913 , n356602 , n8915 , n356604 , n8917 , n356606 , n356607 , n8920 , 
 n356609 , n356610 , n356611 , n356612 , n8925 , n356614 , n8927 , n356616 , n356617 , n356618 , 
 n356619 , n8932 , n356621 , n356622 , n8935 , n356624 , n356625 , n8938 , n8939 , n8940 , 
 n8941 , n356630 , n356631 , n8944 , n356633 , n356634 , n8947 , n356636 , n8949 , n8950 , 
 n356639 , n8952 , n356641 , n356642 , n8955 , n356644 , n356645 , n8958 , n356647 , n356648 , 
 n8961 , n356650 , n356651 , n8964 , n356653 , n8966 , n8967 , n8968 , n8969 , n8970 , 
 n8971 , n8972 , n8973 , n8974 , n356663 , n356664 , n8977 , n356666 , n8979 , n8980 , 
 n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , 
 n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , 
 n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , 
 n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , 
 n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , 
 n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , 
 n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , 
 n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , 
 n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , 
 n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , 
 n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , 
 n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , 
 n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , 
 n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , 
 n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , 
 n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n356828 , 
 n9141 , n356830 , n9143 , n356832 , n356833 , n9146 , n356835 , n356836 , n356837 , n9150 , 
 n356839 , n9152 , n9153 , n356842 , n9155 , n356844 , n9157 , n356846 , n356847 , n9160 , 
 n356849 , n356850 , n9163 , n356852 , n9165 , n356854 , n9167 , n9168 , n356857 , n356858 , 
 n356859 , n9172 , n356861 , n356862 , n9175 , n356864 , n356865 , n9178 , n356867 , n356868 , 
 n9181 , n356870 , n356871 , n356872 , n9185 , n9186 , n356875 , n9188 , n9189 , n356878 , 
 n356879 , n356880 , n9193 , n356882 , n356883 , n9196 , n356885 , n356886 , n9199 , n356888 , 
 n356889 , n356890 , n9203 , n356892 , n9205 , n356894 , n9207 , n9208 , n356897 , n356898 , 
 n9211 , n356900 , n356901 , n9214 , n356903 , n356904 , n9217 , n356906 , n356907 , n9220 , 
 n356909 , n356910 , n9223 , n9224 , n9225 , n9226 , n9227 , n356916 , n356917 , n9230 , 
 n356919 , n356920 , n356921 , n9234 , n356923 , n9236 , n356925 , n356926 , n9239 , n9240 , 
 n356929 , n9242 , n356931 , n356932 , n356933 , n9246 , n356935 , n9248 , n356937 , n356938 , 
 n9251 , n356940 , n356941 , n9254 , n356943 , n356944 , n9257 , n356946 , n356947 , n356948 , 
 n9261 , n356950 , n356951 , n9264 , n356953 , n356954 , n9267 , n356956 , n356957 , n356958 , 
 n356959 , n9272 , n356961 , n9274 , n9275 , n9276 , n9277 , n9278 , n356967 , n356968 , 
 n9281 , n356970 , n9283 , n9284 , n9285 , n9286 , n356975 , n9288 , n356977 , n356978 , 
 n9291 , n356980 , n9293 , n356982 , n9295 , n9296 , n9297 , n9298 , n356987 , n9300 , 
 n356989 , n356990 , n356991 , n9304 , n356993 , n9306 , n9307 , n356996 , n356997 , n356998 , 
 n9311 , n357000 , n357001 , n9314 , n357003 , n357004 , n9317 , n357006 , n357007 , n9320 , 
 n357009 , n9322 , n357011 , n9324 , n9325 , n357014 , n357015 , n357016 , n9329 , n357018 , 
 n357019 , n9332 , n357021 , n357022 , n9335 , n357024 , n357025 , n9338 , n357027 , n357028 , 
 n9341 , n357030 , n357031 , n9344 , n9345 , n9346 , n357035 , n357036 , n357037 , n9350 , 
 n357039 , n357040 , n9353 , n357042 , n357043 , n9356 , n357045 , n357046 , n9359 , n357048 , 
 n357049 , n9362 , n9363 , n9364 , n9365 , n357054 , n357055 , n9368 , n9369 , n357058 , 
 n9371 , n357060 , n9373 , n9374 , n9375 , n9376 , n9377 , n357066 , n9379 , n9380 , 
 n9381 , n9382 , n357071 , n357072 , n9385 , n357074 , n9387 , n357076 , n9389 , n9390 , 
 n357079 , n357080 , n357081 , n9394 , n357083 , n357084 , n9397 , n357086 , n357087 , n9400 , 
 n357089 , n357090 , n357091 , n357092 , n9405 , n357094 , n357095 , n9408 , n357097 , n357098 , 
 n9411 , n9412 , n357101 , n9414 , n9415 , n357104 , n357105 , n9418 , n357107 , n9420 , 
 n9421 , n357110 , n9423 , n357112 , n9425 , n357114 , n357115 , n9428 , n357117 , n9430 , 
 n357119 , n357120 , n9433 , n357122 , n9435 , n9436 , n357125 , n357126 , n357127 , n9440 , 
 n357129 , n357130 , n9443 , n357132 , n357133 , n9446 , n357135 , n357136 , n357137 , n9450 , 
 n357139 , n9452 , n9453 , n357142 , n357143 , n9456 , n357145 , n357146 , n9459 , n357148 , 
 n357149 , n9462 , n357151 , n357152 , n9465 , n357154 , n9467 , n357156 , n357157 , n9470 , 
 n9471 , n9472 , n9473 , n9474 , n357163 , n357164 , n9477 , n357166 , n357167 , n9480 , 
 n9481 , n9482 , n9483 , n357172 , n357173 , n9486 , n9487 , n9488 , n9489 , n9490 , 
 n357179 , n357180 , n9493 , n9494 , n9495 , n9496 , n357185 , n357186 , n357187 , n9500 , 
 n357189 , n9502 , n9503 , n357192 , n9505 , n357194 , n9507 , n9508 , n357197 , n9510 , 
 n357199 , n357200 , n9513 , n357202 , n357203 , n9516 , n357205 , n357206 , n9519 , n357208 , 
 n9521 , n9522 , n9523 , n9524 , n9525 , n357214 , n357215 , n9528 , n357217 , n9530 , 
 n9531 , n357220 , n357221 , n357222 , n9535 , n357224 , n357225 , n9538 , n357227 , n357228 , 
 n9541 , n357230 , n357231 , n9544 , n357233 , n9546 , n357235 , n9548 , n9549 , n357238 , 
 n9551 , n357240 , n9553 , n357242 , n357243 , n9556 , n357245 , n357246 , n9559 , n357248 , 
 n357249 , n9562 , n357251 , n357252 , n9565 , n9566 , n9567 , n9568 , n9569 , n357258 , 
 n357259 , n9572 , n357261 , n357262 , n9575 , n357264 , n357265 , n9578 , n357267 , n357268 , 
 n9581 , n357270 , n9583 , n9584 , n9585 , n9586 , n357275 , n9588 , n357277 , n357278 , 
 n9591 , n357280 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , 
 n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , 
 n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , 
 n9621 , n9622 , n9623 , n9624 , n9625 , n357314 , n9627 , n357316 , n9629 , n9630 , 
 n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n357326 , n9639 , n9640 , 
 n357329 , n9642 , n357331 , n9644 , n357333 , n357334 , n9647 , n357336 , n357337 , n9650 , 
 n9651 , n357340 , n9653 , n9654 , n9655 , n9656 , n9657 , n357346 , n9659 , n357348 , 
 n9661 , n9662 , n9663 , n9664 , n357353 , n9666 , n357355 , n357356 , n9669 , n9670 , 
 n357359 , n357360 , n9673 , n357362 , n357363 , n9676 , n357365 , n357366 , n357367 , n357368 , 
 n9681 , n357370 , n357371 , n9684 , n357373 , n357374 , n9687 , n357376 , n357377 , n9690 , 
 n357379 , n357380 , n9693 , n357382 , n357383 , n9696 , n357385 , n357386 , n9699 , n357388 , 
 n357389 , n9702 , n357391 , n9704 , n357393 , n9706 , n9707 , n9708 , n9709 , n9710 , 
 n9711 , n9712 , n357401 , n357402 , n9715 , n357404 , n357405 , n9718 , n357407 , n357408 , 
 n357409 , n9722 , n357411 , n9724 , n9725 , n357414 , n357415 , n9728 , n357417 , n9730 , 
 n9731 , n357420 , n357421 , n9734 , n357423 , n357424 , n9737 , n357426 , n357427 , n9740 , 
 n357429 , n357430 , n9743 , n357432 , n357433 , n9746 , n9747 , n357436 , n357437 , n9750 , 
 n9751 , n357440 , n9753 , n357442 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , 
 n357449 , n357450 , n9763 , n357452 , n357453 , n9766 , n357455 , n357456 , n9769 , n9770 , 
 n9771 , n357460 , n357461 , n9774 , n9775 , n9776 , n357465 , n9778 , n357467 , n9780 , 
 n9781 , n357470 , n357471 , n9784 , n357473 , n357474 , n9787 , n357476 , n357477 , n357478 , 
 n9791 , n357480 , n9793 , n357482 , n9795 , n9796 , n9797 , n357486 , n357487 , n9800 , 
 n9801 , n9802 , n357491 , n357492 , n357493 , n9806 , n357495 , n9808 , n9809 , n9810 , 
 n9811 , n9812 , n9813 , n9814 , n357503 , n9816 , n357505 , n9818 , n9819 , n9820 , 
 n9821 , n357510 , n357511 , n9824 , n357513 , n357514 , n9827 , n357516 , n357517 , n9830 , 
 n9831 , n9832 , n357521 , n357522 , n9835 , n9836 , n9837 , n357526 , n357527 , n9840 , 
 n9841 , n9842 , n357531 , n357532 , n9845 , n9846 , n9847 , n357536 , n357537 , n9850 , 
 n357539 , n357540 , n9853 , n357542 , n9855 , n357544 , n9857 , n357546 , n9859 , n357548 , 
 n9861 , n9862 , n357551 , n357552 , n9865 , n357554 , n357555 , n9868 , n357557 , n357558 , 
 n9871 , n9872 , n357561 , n9874 , n357563 , n9876 , n9877 , n357566 , n357567 , n9880 , 
 n357569 , n357570 , n9883 , n357572 , n357573 , n357574 , n9887 , n357576 , n357577 , n9890 , 
 n357579 , n357580 , n357581 , n9894 , n357583 , n9896 , n9897 , n357586 , n9899 , n357588 , 
 n9901 , n357590 , n357591 , n9904 , n9905 , n357594 , n9907 , n357596 , n357597 , n357598 , 
 n9911 , n357600 , n357601 , n9914 , n357603 , n357604 , n357605 , n9918 , n357607 , n357608 , 
 n9921 , n357610 , n357611 , n357612 , n9925 , n357614 , n9927 , n9928 , n357617 , n9930 , 
 n357619 , n9932 , n9933 , n357622 , n357623 , n9936 , n357625 , n357626 , n9939 , n357628 , 
 n357629 , n357630 , n9943 , n357632 , n357633 , n9946 , n357635 , n357636 , n9949 , n9950 , 
 n357639 , n357640 , n9953 , n9954 , n9955 , n357644 , n357645 , n357646 , n9959 , n357648 , 
 n9961 , n9962 , n357651 , n9964 , n357653 , n9966 , n9967 , n357656 , n357657 , n9970 , 
 n357659 , n357660 , n9973 , n357662 , n357663 , n357664 , n9977 , n357666 , n357667 , n9980 , 
 n357669 , n357670 , n9983 , n357672 , n9985 , n357674 , n9987 , n9988 , n357677 , n357678 , 
 n9991 , n9992 , n357681 , n357682 , n357683 , n9996 , n357685 , n9998 , n9999 , n357688 , 
 n10001 , n357690 , n10003 , n10004 , n357693 , n357694 , n10007 , n357696 , n357697 , n10010 , 
 n357699 , n357700 , n357701 , n10014 , n357703 , n357704 , n10017 , n357706 , n357707 , n10020 , 
 n357709 , n357710 , n10023 , n357712 , n357713 , n10026 , n357715 , n357716 , n10029 , n10030 , 
 n10031 , n10032 , n357721 , n357722 , n10035 , n357724 , n10037 , n10038 , n10039 , n357728 , 
 n357729 , n10042 , n357731 , n357732 , n10045 , n357734 , n10047 , n10048 , n357737 , n357738 , 
 n357739 , n10052 , n10053 , n357742 , n357743 , n10056 , n10057 , n357746 , n10059 , n357748 , 
 n357749 , n357750 , n10063 , n357752 , n10065 , n357754 , n357755 , n357756 , n357757 , n10070 , 
 n357759 , n10072 , n357761 , n357762 , n10075 , n357764 , n357765 , n10078 , n10079 , n357768 , 
 n357769 , n10082 , n357771 , n10084 , n357773 , n10086 , n10087 , n10088 , n357777 , n10090 , 
 n357779 , n357780 , n10093 , n10095 , n357783 , n357784 , n10098 , n10099 , n10100 , n357788 , 
 n357789 , n10103 , n10104 , n10105 , n357793 , n357794 , n10108 , n357796 , n357797 , n10111 , 
 n357799 , n10113 , n357801 , n10115 , n357803 , n10117 , n10118 , n357806 , n357807 , n10121 , 
 n357809 , n357810 , n10124 , n357812 , n357813 , n10127 , n10128 , n357816 , n10130 , n357818 , 
 n10132 , n10133 , n357821 , n357822 , n10136 , n357824 , n357825 , n10139 , n357827 , n357828 , 
 n357829 , n10143 , n357831 , n357832 , n10146 , n357834 , n357835 , n10149 , n10150 , n10151 , 
 n357839 , n357840 , n357841 , n10155 , n357843 , n357844 , n10158 , n10159 , n357847 , n10161 , 
 n10162 , n357850 , n357851 , n10165 , n10166 , n10167 , n10168 , n357856 , n10170 , n357858 , 
 n10172 , n10173 , n357861 , n357862 , n10176 , n357864 , n357865 , n10179 , n357867 , n357868 , 
 n10182 , n10183 , n10184 , n10185 , n10186 , n357874 , n357875 , n357876 , n10190 , n357878 , 
 n10192 , n10193 , n357881 , n357882 , n10196 , n357884 , n357885 , n10199 , n357887 , n357888 , 
 n10202 , n10203 , n10204 , n357892 , n357893 , n10207 , n357895 , n357896 , n10210 , n10211 , 
 n10212 , n357900 , n357901 , n10215 , n10216 , n10217 , n10218 , n10219 , n357907 , n357908 , 
 n10222 , n10223 , n357911 , n357912 , n10226 , n357914 , n10228 , n357916 , n10230 , n10231 , 
 n357919 , n357920 , n10234 , n357922 , n357923 , n10237 , n357925 , n357926 , n10240 , n357928 , 
 n357929 , n10243 , n357931 , n357932 , n357933 , n10247 , n357935 , n10249 , n10250 , n357938 , 
 n10252 , n357940 , n10254 , n10255 , n357943 , n357944 , n10258 , n357946 , n357947 , n10261 , 
 n357949 , n357950 , n357951 , n10265 , n357953 , n357954 , n10268 , n357956 , n357957 , n10271 , 
 n10272 , n357960 , n357961 , n10275 , n357963 , n10277 , n357965 , n10279 , n10280 , n357968 , 
 n10282 , n357970 , n10284 , n10285 , n357973 , n357974 , n10288 , n357976 , n357977 , n10291 , 
 n357979 , n357980 , n357981 , n10295 , n357983 , n357984 , n10298 , n357986 , n357987 , n10301 , 
 n10302 , n357990 , n357991 , n10305 , n10306 , n10307 , n357995 , n357996 , n357997 , n10311 , 
 n357999 , n10313 , n10314 , n358002 , n10316 , n358004 , n10318 , n10319 , n358007 , n358008 , 
 n10322 , n358010 , n358011 , n10325 , n358013 , n358014 , n358015 , n10329 , n358017 , n358018 , 
 n10332 , n358020 , n358021 , n10335 , n358023 , n10337 , n358025 , n10339 , n10340 , n358028 , 
 n358029 , n10343 , n10344 , n358032 , n358033 , n358034 , n358035 , n10349 , n358037 , n358038 , 
 n358039 , n10353 , n358041 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , 
 n10362 , n358050 , n358051 , n358052 , n10366 , n10367 , n358055 , n358056 , n10370 , n358058 , 
 n358059 , n358060 , n10374 , n358062 , n358063 , n10377 , n358065 , n358066 , n10380 , n10381 , 
 n358069 , n10383 , n10384 , n10385 , n358073 , n10387 , n358075 , n358076 , n10390 , n358078 , 
 n10392 , n358080 , n358081 , n358082 , n358083 , n10397 , n358085 , n358086 , n358087 , n10401 , 
 n358089 , n358090 , n10404 , n358092 , n358093 , n10407 , n10408 , n10409 , n10413 , n10414 , 
 n10415 , n10416 , n10417 , n10419 , n10420 , n10424 , n10425 , n10426 , n10427 , n10428 , 
 n10429 , n10430 , n10431 , n10432 , n358113 , n10434 , n10436 , n358116 , n358117 , n10439 , 
 n358119 , n10441 , n358121 , n10443 , n10444 , n10445 , n358125 , n10447 , n358127 , n358128 , 
 n10450 , n10451 , n10452 , n358132 , n358133 , n10455 , n10456 , n10457 , n358137 , n358138 , 
 n10460 , n10461 , n10462 , n358142 , n358143 , n10465 , n10466 , n10467 , n358147 , n358148 , 
 n358149 , n10471 , n358151 , n10473 , n10474 , n358154 , n10476 , n10477 , n10478 , n10479 , 
 n358159 , n10481 , n358161 , n358162 , n10484 , n358164 , n358165 , n10487 , n10488 , n10489 , 
 n358169 , n358170 , n10492 , n10493 , n10494 , n358174 , n358175 , n358176 , n10498 , n358178 , 
 n10500 , n10501 , n358181 , n10503 , n358183 , n10505 , n10506 , n358186 , n358187 , n10509 , 
 n358189 , n358190 , n10512 , n358192 , n358193 , n358194 , n10516 , n358196 , n358197 , n10519 , 
 n358199 , n358200 , n10522 , n10523 , n10524 , n358204 , n358205 , n10527 , n10528 , n10529 , 
 n358209 , n358210 , n10532 , n358212 , n358213 , n10535 , n358215 , n10537 , n10538 , n10539 , 
 n358219 , n358220 , n358221 , n10543 , n358223 , n10545 , n10546 , n358226 , n10548 , n358228 , 
 n10550 , n10551 , n358231 , n358232 , n10554 , n358234 , n358235 , n10557 , n358237 , n358238 , 
 n358239 , n10561 , n358241 , n358242 , n10564 , n358244 , n358245 , n358246 , n10568 , n358248 , 
 n10570 , n10571 , n358251 , n10573 , n10574 , n358254 , n10576 , n10577 , n358257 , n10579 , 
 n358259 , n10581 , n358261 , n358262 , n10584 , n358264 , n358265 , n358266 , n10588 , n358268 , 
 n358269 , n10591 , n358271 , n358272 , n10594 , n10595 , n10596 , n358276 , n358277 , n10599 , 
 n10600 , n10601 , n358281 , n358282 , n10604 , n10605 , n358285 , n358286 , n10608 , n358288 , 
 n10610 , n358290 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , 
 n358299 , n358300 , n10622 , n358302 , n358303 , n10625 , n358305 , n358306 , n10628 , n10629 , 
 n10630 , n358310 , n358311 , n10633 , n358313 , n10635 , n10636 , n358316 , n10638 , n358318 , 
 n10640 , n358320 , n10642 , n10643 , n358323 , n358324 , n10646 , n358326 , n358327 , n10649 , 
 n358329 , n358330 , n10652 , n10653 , n358333 , n10655 , n358335 , n10657 , n10658 , n358338 , 
 n358339 , n10661 , n358341 , n358342 , n10664 , n358344 , n358345 , n358346 , n10668 , n358348 , 
 n358349 , n10671 , n358351 , n358352 , n10674 , n10675 , n358355 , n358356 , n10678 , n10679 , 
 n10680 , n358360 , n358361 , n358362 , n10684 , n358364 , n10686 , n10687 , n358367 , n10689 , 
 n358369 , n10691 , n10692 , n10693 , n10694 , n358374 , n10696 , n358376 , n358377 , n358378 , 
 n10700 , n358380 , n358381 , n10703 , n358383 , n358384 , n10706 , n358386 , n10708 , n358388 , 
 n10710 , n10711 , n358391 , n358392 , n10714 , n10715 , n358395 , n358396 , n358397 , n358398 , 
 n10720 , n358400 , n358401 , n358402 , n358403 , n10725 , n10726 , n358406 , n10728 , n10729 , 
 n358409 , n358410 , n358411 , n10733 , n358413 , n358414 , n358415 , n10737 , n358417 , n358418 , 
 n10740 , n358420 , n358421 , n358422 , n10744 , n358424 , n358425 , n10747 , n10748 , n358428 , 
 n358429 , n10751 , n358431 , n358432 , n10754 , n358434 , n358435 , n10757 , n358437 , n10759 , 
 n358439 , n358440 , n358441 , n358442 , n10764 , n358444 , n358445 , n10767 , n358447 , n358448 , 
 n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n358458 , 
 n10780 , n10782 , n358461 , n358462 , n10785 , n358464 , n10787 , n358466 , n10789 , n10790 , 
 n10791 , n10792 , n358471 , n10794 , n358473 , n358474 , n10797 , n10798 , n10799 , n358478 , 
 n358479 , n10802 , n10803 , n10804 , n358483 , n358484 , n10807 , n10808 , n10809 , n358488 , 
 n358489 , n358490 , n10813 , n358492 , n358493 , n10816 , n10817 , n358496 , n10819 , n10820 , 
 n358499 , n358500 , n10823 , n10824 , n358503 , n10826 , n358505 , n10828 , n10829 , n358508 , 
 n358509 , n10832 , n358511 , n358512 , n10835 , n358514 , n358515 , n358516 , n10839 , n358518 , 
 n358519 , n10842 , n358521 , n358522 , n10845 , n358524 , n10847 , n358526 , n10849 , n358528 , 
 n10851 , n10852 , n358531 , n358532 , n10855 , n358534 , n358535 , n10858 , n358537 , n358538 , 
 n10861 , n10862 , n358541 , n358542 , n10865 , n358544 , n358545 , n10868 , n358547 , n358548 , 
 n10871 , n10872 , n358551 , n358552 , n10875 , n358554 , n10877 , n358556 , n10879 , n358558 , 
 n10881 , n10882 , n358561 , n10884 , n358563 , n10886 , n358565 , n358566 , n10889 , n358568 , 
 n358569 , n10892 , n10893 , n10894 , n10895 , n10896 , n358575 , n10898 , n358577 , n10900 , 
 n358579 , n10902 , n358581 , n358582 , n10905 , n358584 , n358585 , n10908 , n358587 , n358588 , 
 n10911 , n358590 , n358591 , n10914 , n358593 , n358594 , n10917 , n10918 , n10919 , n10920 , 
 n10921 , n10922 , n10923 , n358602 , n10925 , n10926 , n358605 , n358606 , n10929 , n358608 , 
 n10931 , n358610 , n10933 , n10934 , n358613 , n10936 , n358615 , n10938 , n10939 , n10940 , 
 n10941 , n358620 , n10943 , n358622 , n358623 , n358624 , n10947 , n358626 , n358627 , n10950 , 
 n358629 , n358630 , n10953 , n10954 , n10955 , n358634 , n358635 , n10958 , n358637 , n358638 , 
 n10961 , n358640 , n10963 , n358642 , n10965 , n358644 , n10967 , n10968 , n10969 , n10970 , 
 n10971 , n10972 , n10973 , n358652 , n358653 , n10976 , n358655 , n358656 , n10979 , n358658 , 
 n358659 , n10982 , n10983 , n358662 , n358663 , n10986 , n358665 , n10988 , n358667 , n10990 , 
 n10991 , n358670 , n358671 , n10994 , n358673 , n358674 , n358675 , n10998 , n358677 , n358678 , 
 n11001 , n358680 , n358681 , n11004 , n11005 , n11006 , n358685 , n11008 , n11009 , n358688 , 
 n11011 , n358690 , n11013 , n358692 , n11015 , n11016 , n358695 , n11018 , n358697 , n11020 , 
 n11021 , n358700 , n11023 , n358702 , n11025 , n358704 , n358705 , n11028 , n358707 , n358708 , 
 n358709 , n11032 , n358711 , n358712 , n11035 , n358714 , n358715 , n11038 , n11039 , n358718 , 
 n358719 , n11042 , n11043 , n11044 , n358723 , n358724 , n358725 , n11048 , n358727 , n11050 , 
 n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n358735 , n358736 , n11059 , n358738 , 
 n358739 , n11062 , n358741 , n358742 , n11065 , n358744 , n11067 , n358746 , n11069 , n11070 , 
 n358749 , n358750 , n11073 , n11074 , n358753 , n358754 , n358755 , n11078 , n358757 , n11080 , 
 n11081 , n11082 , n11083 , n11084 , n11085 , n358764 , n358765 , n11088 , n358767 , n358768 , 
 n11091 , n358770 , n358771 , n11094 , n358773 , n358774 , n11097 , n358776 , n358777 , n358778 , 
 n11101 , n358780 , n11103 , n358782 , n11105 , n11106 , n358785 , n11108 , n358787 , n11110 , 
 n358789 , n358790 , n11113 , n358792 , n358793 , n11116 , n11117 , n358796 , n358797 , n11120 , 
 n11121 , n358800 , n11123 , n11124 , n358803 , n358804 , n358805 , n11128 , n358807 , n358808 , 
 n11131 , n358810 , n358811 , n11134 , n358813 , n358814 , n11137 , n358816 , n11139 , n358818 , 
 n358819 , n358820 , n358821 , n11144 , n11145 , n358824 , n11147 , n358826 , n358827 , n11150 , 
 n358829 , n358830 , n11153 , n358832 , n358833 , n11156 , n358835 , n11158 , n358837 , n11160 , 
 n11161 , n358840 , n358841 , n11164 , n358843 , n358844 , n11167 , n358846 , n358847 , n11170 , 
 n11172 , n358850 , n358851 , n11175 , n11176 , n11177 , n358855 , n358856 , n11180 , n11181 , 
 n11182 , n358860 , n358861 , n11185 , n11186 , n11187 , n358865 , n11189 , n11190 , n358868 , 
 n11192 , n11193 , n11194 , n358872 , n11196 , n358874 , n11198 , n358876 , n358877 , n11201 , 
 n11202 , n358880 , n11204 , n11205 , n358883 , n358884 , n11208 , n11209 , n11210 , n11211 , 
 n11212 , n358890 , n358891 , n11215 , n358893 , n11217 , n358895 , n358896 , n11220 , n358898 , 
 n358899 , n11223 , n358901 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , 
 n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n358917 , n11241 , 
 n11242 , n358920 , n358921 , n11245 , n358923 , n11247 , n358925 , n11249 , n11250 , n358928 , 
 n358929 , n11253 , n11254 , n358932 , n358933 , n358934 , n358935 , n11259 , n358937 , n358938 , 
 n11262 , n358940 , n358941 , n358942 , n11266 , n358944 , n11268 , n11269 , n358947 , n358948 , 
 n11272 , n358950 , n358951 , n11275 , n358953 , n358954 , n358955 , n11279 , n358957 , n11281 , 
 n358959 , n11283 , n358961 , n358962 , n11286 , n358964 , n358965 , n358966 , n358967 , n11291 , 
 n358969 , n358970 , n11294 , n358972 , n358973 , n11297 , n358975 , n358976 , n358977 , n11301 , 
 n358979 , n358980 , n11304 , n358982 , n358983 , n11307 , n11308 , n358986 , n358987 , n11311 , 
 n358989 , n358990 , n11314 , n358992 , n358993 , n11317 , n358995 , n358996 , n11320 , n11322 , 
 n358999 , n359000 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n359007 , n359008 , 
 n11333 , n359010 , n11335 , n359012 , n11337 , n359014 , n359015 , n11340 , n359017 , n359018 , 
 n11343 , n11344 , n11345 , n359022 , n11347 , n359024 , n11349 , n359026 , n11351 , n11352 , 
 n359029 , n11354 , n359031 , n11356 , n359033 , n359034 , n11359 , n359036 , n11361 , n11362 , 
 n359039 , n11364 , n11365 , n11366 , n11367 , n359044 , n11369 , n11370 , n11371 , n359048 , 
 n11373 , n11374 , n11375 , n359052 , n11377 , n11378 , n359055 , n359056 , n11381 , n11382 , 
 n11383 , n359060 , n11385 , n359062 , n11387 , n11388 , n359065 , n11390 , n359067 , n359068 , 
 n11393 , n359070 , n359071 , n11396 , n359073 , n359074 , n11399 , n359076 , n11401 , n11402 , 
 n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n359085 , n359086 , n11411 , n359088 , 
 n11413 , n359090 , n11415 , n11416 , n11417 , n11418 , n11419 , n359096 , n11421 , n359098 , 
 n11423 , n11424 , n11425 , n11426 , n11427 , n359104 , n11429 , n11430 , n359107 , n359108 , 
 n11433 , n359110 , n359111 , n11436 , n359113 , n359114 , n11439 , n11440 , n11441 , n11442 , 
 n359119 , n359120 , n11445 , n359122 , n11447 , n359124 , n11449 , n11450 , n359127 , n359128 , 
 n11453 , n359130 , n359131 , n11456 , n359133 , n359134 , n11459 , n11460 , n359137 , n359138 , 
 n11463 , n359140 , n11465 , n359142 , n11467 , n11468 , n359145 , n11470 , n359147 , n359148 , 
 n359149 , n11474 , n359151 , n359152 , n11477 , n359154 , n359155 , n11480 , n359157 , n359158 , 
 n11483 , n359160 , n359161 , n11486 , n359163 , n11488 , n359165 , n11490 , n11491 , n359168 , 
 n11493 , n359170 , n11495 , n359172 , n359173 , n11498 , n359175 , n359176 , n11501 , n11502 , 
 n11503 , n11504 , n11505 , n359182 , n359183 , n11508 , n11509 , n359186 , n359187 , n11512 , 
 n359189 , n11514 , n359191 , n11516 , n11517 , n359194 , n359195 , n11520 , n359197 , n359198 , 
 n11523 , n359200 , n359201 , n11526 , n359203 , n359204 , n11529 , n11530 , n11531 , n11532 , 
 n359209 , n359210 , n11535 , n359212 , n359213 , n11538 , n359215 , n359216 , n11541 , n11542 , 
 n359219 , n359220 , n11545 , n359222 , n359223 , n11548 , n359225 , n11550 , n11551 , n11552 , 
 n359229 , n359230 , n11555 , n11556 , n11557 , n11558 , n11559 , n359236 , n359237 , n11562 , 
 n359239 , n359240 , n11565 , n359242 , n11567 , n11568 , n359245 , n359246 , n11571 , n359248 , 
 n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n359256 , n359257 , n11582 , 
 n359259 , n11584 , n359261 , n11586 , n359263 , n11588 , n11589 , n11590 , n11591 , n359268 , 
 n359269 , n11594 , n11595 , n11596 , n11597 , n11598 , n359275 , n11600 , n11601 , n11602 , 
 n359279 , n359280 , n11605 , n359282 , n359283 , n11608 , n11609 , n11610 , n11611 , n359288 , 
 n359289 , n11614 , n359291 , n11616 , n359293 , n359294 , n11619 , n359296 , n11621 , n11622 , 
 n11623 , n11624 , n359301 , n359302 , n11627 , n11628 , n11629 , n11630 , n11631 , n359308 , 
 n359309 , n11634 , n359311 , n359312 , n11637 , n359314 , n11639 , n11640 , n359317 , n359318 , 
 n11643 , n359320 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , 
 n11653 , n11654 , n359331 , n359332 , n359333 , n11658 , n359335 , n11660 , n359337 , n11662 , 
 n11663 , n359340 , n359341 , n11666 , n359343 , n359344 , n11669 , n359346 , n359347 , n11672 , 
 n11673 , n359350 , n359351 , n11676 , n359353 , n359354 , n11679 , n359356 , n359357 , n11682 , 
 n11683 , n11684 , n11685 , n11686 , n359363 , n359364 , n359365 , n11690 , n359367 , n11692 , 
 n359369 , n11694 , n11695 , n359372 , n359373 , n11698 , n359375 , n359376 , n11701 , n359378 , 
 n359379 , n11704 , n11705 , n11706 , n359383 , n11708 , n359385 , n359386 , n11711 , n11712 , 
 n11713 , n11714 , n11715 , n359392 , n359393 , n11718 , n11719 , n11720 , n11721 , n359398 , 
 n359399 , n11724 , n359401 , n11726 , n11727 , n11728 , n11729 , n11730 , n359407 , n11732 , 
 n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n359417 , n359418 , 
 n11743 , n359420 , n11745 , n359422 , n359423 , n359424 , n11749 , n359426 , n359427 , n359428 , 
 n11753 , n359430 , n11755 , n359432 , n11757 , n359434 , n359435 , n11760 , n11761 , n359438 , 
 n359439 , n11764 , n359441 , n359442 , n11767 , n359444 , n359445 , n11770 , n11771 , n11772 , 
 n11773 , n11774 , n359451 , n359452 , n11777 , n359454 , n359455 , n11780 , n359457 , n11782 , 
 n359459 , n11784 , n359461 , n11786 , n11787 , n359464 , n359465 , n11790 , n359467 , n359468 , 
 n11793 , n359470 , n359471 , n11796 , n11797 , n359474 , n359475 , n11800 , n359477 , n359478 , 
 n11803 , n359480 , n359481 , n11806 , n359483 , n359484 , n11809 , n359486 , n359487 , n11812 , 
 n359489 , n359490 , n11815 , n359492 , n359493 , n11818 , n11819 , n11820 , n11821 , n359498 , 
 n359499 , n11824 , n11825 , n11826 , n11827 , n11828 , n359505 , n359506 , n359507 , n11832 , 
 n11833 , n11834 , n11835 , n11836 , n359513 , n11838 , n11839 , n359516 , n359517 , n11842 , 
 n359519 , n359520 , n11845 , n359522 , n359523 , n11848 , n359525 , n11850 , n359527 , n11852 , 
 n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , 
 n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n359545 , n359546 , n359547 , n359548 , 
 n11873 , n359550 , n359551 , n359552 , n11877 , n359554 , n11879 , n11880 , n359557 , n359558 , 
 n359559 , n11884 , n359561 , n359562 , n11887 , n359564 , n359565 , n11890 , n359567 , n359568 , 
 n11893 , n359570 , n11895 , n359572 , n11897 , n11898 , n359575 , n11900 , n359577 , n11902 , 
 n359579 , n359580 , n11905 , n359582 , n359583 , n11908 , n359585 , n359586 , n11911 , n11912 , 
 n11913 , n11914 , n359591 , n359592 , n359593 , n11918 , n359595 , n359596 , n11921 , n359598 , 
 n11923 , n11924 , n359601 , n11926 , n359603 , n11928 , n11929 , n359606 , n359607 , n359608 , 
 n11933 , n359610 , n359611 , n11936 , n359613 , n359614 , n11939 , n359616 , n11941 , n11942 , 
 n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n359626 , n11951 , n359628 , 
 n359629 , n11954 , n11955 , n11956 , n11957 , n359634 , n359635 , n11960 , n11961 , n11962 , 
 n11963 , n11964 , n359641 , n359642 , n11967 , n11968 , n11969 , n11970 , n359647 , n359648 , 
 n11973 , n11974 , n11975 , n11976 , n359653 , n359654 , n11979 , n359656 , n11981 , n359658 , 
 n11983 , n11984 , n359661 , n359662 , n359663 , n11988 , n359665 , n359666 , n11991 , n359668 , 
 n359669 , n11994 , n359671 , n359672 , n11997 , n11998 , n359675 , n12000 , n359677 , n12002 , 
 n359679 , n12004 , n12005 , n359682 , n359683 , n359684 , n12009 , n359686 , n359687 , n12012 , 
 n359689 , n359690 , n12015 , n359692 , n359693 , n12018 , n359695 , n359696 , n12021 , n359698 , 
 n359699 , n12024 , n12025 , n12026 , n12027 , n12028 , n359705 , n359706 , n12031 , n359708 , 
 n359709 , n12034 , n359711 , n359712 , n12037 , n12038 , n12039 , n12040 , n359717 , n359718 , 
 n12043 , n12044 , n12045 , n12046 , n12047 , n359724 , n359725 , n12050 , n12051 , n12052 , 
 n12053 , n359730 , n359731 , n12056 , n12057 , n12058 , n12059 , n12060 , n359737 , n359738 , 
 n359739 , n359740 , n12065 , n359742 , n359743 , n12068 , n12069 , n12070 , n12071 , n12072 , 
 n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n359755 , n12080 , n359757 , n12082 , 
 n359759 , n12084 , n12085 , n359762 , n12087 , n359764 , n12089 , n359766 , n359767 , n12092 , 
 n359769 , n359770 , n12095 , n359772 , n359773 , n12098 , n359775 , n12100 , n359777 , n12102 , 
 n12103 , n359780 , n359781 , n359782 , n12107 , n359784 , n359785 , n12110 , n359787 , n359788 , 
 n12113 , n359790 , n359791 , n359792 , n12117 , n359794 , n12119 , n12120 , n359797 , n12122 , 
 n359799 , n12124 , n359801 , n359802 , n12127 , n359804 , n359805 , n12130 , n359807 , n359808 , 
 n359809 , n12134 , n359811 , n359812 , n12137 , n359814 , n359815 , n12140 , n12141 , n12142 , 
 n12143 , n359820 , n359821 , n12146 , n12147 , n12148 , n12149 , n12150 , n359827 , n359828 , 
 n359829 , n359830 , n12155 , n359832 , n12157 , n359834 , n359835 , n359836 , n359837 , n12162 , 
 n359839 , n359840 , n12165 , n359842 , n359843 , n12168 , n12169 , n12170 , n12171 , n359848 , 
 n359849 , n12174 , n359851 , n12176 , n359853 , n12178 , n12179 , n359856 , n359857 , n359858 , 
 n12183 , n359860 , n359861 , n12186 , n359863 , n359864 , n12189 , n359866 , n359867 , n12192 , 
 n359869 , n12194 , n12195 , n359872 , n359873 , n359874 , n12199 , n359876 , n359877 , n12202 , 
 n359879 , n359880 , n12205 , n359882 , n12207 , n12208 , n359885 , n12210 , n359887 , n12212 , 
 n12213 , n359890 , n12215 , n359892 , n12217 , n359894 , n12219 , n359896 , n359897 , n12222 , 
 n12223 , n12224 , n12225 , n12226 , n359903 , n359904 , n12229 , n359906 , n359907 , n12232 , 
 n359909 , n359910 , n12235 , n359912 , n359913 , n12238 , n359915 , n12240 , n12241 , n12242 , 
 n12243 , n359920 , n12245 , n12246 , n359923 , n359924 , n12249 , n359926 , n12251 , n12252 , 
 n12253 , n359930 , n12255 , n359932 , n12257 , n12258 , n359935 , n12260 , n359937 , n359938 , 
 n12263 , n359940 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , 
 n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , 
 n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , 
 n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , 
 n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , 
 n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , 
 n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , 
 n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , 
 n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , 
 n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , 
 n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , 
 n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , 
 n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , 
 n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , 
 n12403 , n12404 , n12405 , n12406 , n12407 , n360084 , n12409 , n360086 , n12411 , n12412 , 
 n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n360097 , n12422 , 
 n360099 , n360100 , n12425 , n12426 , n360103 , n12428 , n360105 , n360106 , n360107 , n12432 , 
 n360109 , n360110 , n12435 , n360112 , n360113 , n12438 , n12439 , n360116 , n360117 , n12442 , 
 n360119 , n360120 , n12445 , n360122 , n360123 , n12448 , n360125 , n360126 , n12451 , n360128 , 
 n12453 , n12454 , n12455 , n12456 , n360133 , n12458 , n360135 , n360136 , n360137 , n12462 , 
 n360139 , n360140 , n12465 , n360142 , n360143 , n12468 , n360145 , n12470 , n12471 , n12472 , 
 n12473 , n12474 , n12475 , n360152 , n12477 , n360154 , n12479 , n12480 , n12481 , n12482 , 
 n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , 
 n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , 
 n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , 
 n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , 
 n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , 
 n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , 
 n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , 
 n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , 
 n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , 
 n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , 
 n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , 
 n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , 
 n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , 
 n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , 
 n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , 
 n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , 
 n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n360328 , 
 n360329 , n12654 , n12655 , n12656 , n12657 , n360334 , n360335 , n12660 , n12661 , n12662 , 
 n12663 , n12664 , n360341 , n360342 , n360343 , n12668 , n360345 , n12670 , n12671 , n360348 , 
 n360349 , n12674 , n360351 , n360352 , n12677 , n360354 , n360355 , n12680 , n360357 , n360358 , 
 n12683 , n12684 , n12685 , n12686 , n360363 , n360364 , n12689 , n12690 , n12691 , n12692 , 
 n12693 , n360370 , n360371 , n12696 , n360373 , n360374 , n12699 , n360376 , n12701 , n360378 , 
 n12703 , n12704 , n360381 , n12706 , n360383 , n360384 , n360385 , n360386 , n12711 , n360388 , 
 n360389 , n12714 , n360391 , n360392 , n360393 , n360394 , n12719 , n360396 , n360397 , n360398 , 
 n12723 , n360400 , n12725 , n12726 , n360403 , n360404 , n360405 , n12730 , n360407 , n360408 , 
 n12733 , n360410 , n360411 , n12736 , n360413 , n360414 , n12739 , n360416 , n12741 , n360418 , 
 n12743 , n360420 , n360421 , n12746 , n12747 , n360424 , n360425 , n360426 , n12751 , n360428 , 
 n360429 , n12754 , n360431 , n360432 , n12757 , n360434 , n360435 , n12760 , n360437 , n360438 , 
 n12763 , n360440 , n12765 , n360442 , n12767 , n12768 , n360445 , n360446 , n360447 , n12772 , 
 n360449 , n360450 , n12775 , n360452 , n360453 , n12778 , n360455 , n360456 , n360457 , n12782 , 
 n360459 , n12784 , n12785 , n360462 , n360463 , n360464 , n12789 , n360466 , n360467 , n12792 , 
 n360469 , n360470 , n12795 , n360472 , n360473 , n12798 , n360475 , n12800 , n360477 , n12802 , 
 n12803 , n360480 , n360481 , n360482 , n12807 , n360484 , n360485 , n12810 , n360487 , n360488 , 
 n12813 , n360490 , n360491 , n12816 , n360493 , n360494 , n12819 , n360496 , n360497 , n12822 , 
 n360499 , n360500 , n12825 , n360502 , n360503 , n12828 , n12829 , n12830 , n12831 , n360508 , 
 n360509 , n12834 , n12835 , n12836 , n12837 , n12838 , n360515 , n360516 , n12841 , n12842 , 
 n12843 , n12844 , n360521 , n360522 , n12847 , n12848 , n12849 , n12850 , n12851 , n360528 , 
 n360529 , n360530 , n12855 , n360532 , n12857 , n12858 , n360535 , n360536 , n12861 , n360538 , 
 n360539 , n12864 , n360541 , n360542 , n12867 , n360544 , n360545 , n12870 , n12871 , n12872 , 
 n12873 , n360550 , n360551 , n12876 , n360553 , n360554 , n12879 , n360556 , n12881 , n360558 , 
 n360559 , n360560 , n360561 , n12886 , n360563 , n360564 , n12889 , n360566 , n360567 , n12892 , 
 n360569 , n360570 , n12895 , n12896 , n12897 , n12898 , n360575 , n360576 , n12901 , n360578 , 
 n12903 , n360580 , n12905 , n12906 , n360583 , n360584 , n12909 , n360586 , n12911 , n360588 , 
 n360589 , n12914 , n360591 , n360592 , n12917 , n12918 , n12919 , n12920 , n360597 , n360598 , 
 n360599 , n12924 , n360601 , n360602 , n12927 , n360604 , n12929 , n12930 , n12931 , n12932 , 
 n12933 , n360610 , n360611 , n360612 , n12937 , n360614 , n360615 , n12940 , n360617 , n12942 , 
 n12943 , n360620 , n12945 , n12946 , n12947 , n12948 , n360625 , n360626 , n360627 , n12952 , 
 n360629 , n360630 , n12955 , n360632 , n12957 , n360634 , n12959 , n360636 , n12961 , n12962 , 
 n360639 , n12964 , n360641 , n12966 , n360643 , n360644 , n12969 , n360646 , n12971 , n360648 , 
 n360649 , n12974 , n360651 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n360658 , 
 n12983 , n360660 , n360661 , n12986 , n360663 , n360664 , n12989 , n12990 , n12991 , n12992 , 
 n12993 , n360670 , n360671 , n12996 , n360673 , n360674 , n12999 , n360676 , n360677 , n13002 , 
 n360679 , n360680 , n13005 , n360682 , n360683 , n13008 , n13009 , n13010 , n13011 , n360688 , 
 n360689 , n13014 , n360691 , n360692 , n13017 , n360694 , n360695 , n13020 , n360697 , n13022 , 
 n13023 , n13024 , n13025 , n13026 , n13027 , n360704 , n13029 , n360706 , n13031 , n13032 , 
 n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n360717 , n13042 , 
 n360719 , n13044 , n13045 , n360722 , n13047 , n360724 , n13049 , n360726 , n13051 , n360728 , 
 n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , 
 n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , 
 n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , 
 n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , 
 n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , 
 n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , 
 n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , 
 n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , 
 n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , 
 n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , 
 n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , 
 n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , 
 n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , 
 n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n360866 , n13191 , n360868 , 
 n13193 , n360870 , n13195 , n360872 , n360873 , n13198 , n13199 , n13200 , n13201 , n13202 , 
 n13203 , n360880 , n13205 , n360882 , n360883 , n13208 , n360885 , n13210 , n13211 , n13212 , 
 n13213 , n360890 , n360891 , n360892 , n13217 , n360894 , n13219 , n13220 , n360897 , n360898 , 
 n360899 , n13224 , n360901 , n360902 , n13227 , n360904 , n360905 , n13230 , n360907 , n360908 , 
 n360909 , n13234 , n360911 , n13236 , n360913 , n360914 , n13239 , n13240 , n360917 , n360918 , 
 n360919 , n13244 , n360921 , n360922 , n13247 , n360924 , n360925 , n13250 , n360927 , n360928 , 
 n13253 , n360930 , n360931 , n13256 , n360933 , n13258 , n360935 , n360936 , n13261 , n360938 , 
 n360939 , n13264 , n360941 , n13266 , n360943 , n13268 , n13269 , n360946 , n360947 , n360948 , 
 n13273 , n360950 , n360951 , n13276 , n360953 , n360954 , n13279 , n360956 , n360957 , n360958 , 
 n13283 , n360960 , n13285 , n13286 , n360963 , n360964 , n360965 , n13290 , n360967 , n360968 , 
 n13293 , n360970 , n360971 , n13296 , n360973 , n360974 , n13299 , n360976 , n13301 , n360978 , 
 n13303 , n13304 , n360981 , n360982 , n360983 , n13308 , n360985 , n360986 , n13311 , n360988 , 
 n360989 , n13314 , n360991 , n360992 , n13317 , n360994 , n360995 , n13320 , n360997 , n360998 , 
 n13323 , n13324 , n13325 , n13326 , n361003 , n361004 , n13329 , n361006 , n361007 , n13332 , 
 n361009 , n361010 , n361011 , n13336 , n13337 , n13338 , n13339 , n13340 , n361017 , n361018 , 
 n13343 , n361020 , n361021 , n13346 , n13347 , n13348 , n13349 , n361026 , n361027 , n13352 , 
 n13353 , n13354 , n13355 , n13356 , n361033 , n361034 , n13359 , n361036 , n361037 , n13362 , 
 n361039 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n361048 , 
 n361049 , n361050 , n13375 , n361052 , n13377 , n361054 , n361055 , n361056 , n13381 , n361058 , 
 n13383 , n13384 , n13385 , n13386 , n361063 , n13388 , n361065 , n361066 , n13391 , n361068 , 
 n13393 , n361070 , n13395 , n13396 , n361073 , n361074 , n361075 , n13400 , n361077 , n361078 , 
 n13403 , n361080 , n361081 , n13406 , n361083 , n361084 , n13409 , n361086 , n361087 , n13412 , 
 n361089 , n13414 , n361091 , n13416 , n13417 , n361094 , n361095 , n361096 , n13421 , n361098 , 
 n361099 , n13424 , n361101 , n361102 , n13427 , n361104 , n361105 , n361106 , n13431 , n361108 , 
 n13433 , n361110 , n361111 , n13436 , n13437 , n361114 , n361115 , n361116 , n13441 , n361118 , 
 n361119 , n13444 , n361121 , n361122 , n13447 , n361124 , n361125 , n13450 , n361127 , n13452 , 
 n361129 , n13454 , n361131 , n361132 , n13457 , n13458 , n361135 , n361136 , n361137 , n13462 , 
 n361139 , n361140 , n13465 , n361142 , n361143 , n13468 , n361145 , n361146 , n13471 , n361148 , 
 n361149 , n13474 , n361151 , n361152 , n361153 , n361154 , n13479 , n361156 , n13481 , n13482 , 
 n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n361165 , n13490 , n13491 , n13492 , 
 n13493 , n361170 , n361171 , n13496 , n13497 , n13498 , n13499 , n13500 , n361177 , n361178 , 
 n13503 , n361180 , n361181 , n13506 , n13507 , n13508 , n13509 , n13510 , n361187 , n361188 , 
 n13513 , n361190 , n13515 , n13516 , n13517 , n13518 , n361195 , n13520 , n13521 , n13522 , 
 n13523 , n13524 , n361201 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n361208 , 
 n13533 , n361210 , n13535 , n361212 , n361213 , n13538 , n13539 , n13540 , n13541 , n361218 , 
 n361219 , n13544 , n361221 , n361222 , n13547 , n361224 , n361225 , n13550 , n361227 , n13552 , 
 n13553 , n361230 , n13555 , n361232 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , 
 n13563 , n13564 , n13565 , n13566 , n13567 , n361244 , n13569 , n361246 , n13571 , n361248 , 
 n361249 , n13574 , n361251 , n361252 , n13577 , n361254 , n13579 , n13580 , n361257 , n13582 , 
 n361259 , n13584 , n13585 , n13586 , n361263 , n361264 , n13589 , n361266 , n361267 , n13592 , 
 n361269 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n361277 , n361278 , 
 n13603 , n361280 , n361281 , n361282 , n13607 , n361284 , n13609 , n13610 , n361287 , n361288 , 
 n361289 , n13614 , n361291 , n361292 , n13617 , n361294 , n361295 , n13620 , n361297 , n361298 , 
 n13623 , n361300 , n361301 , n13626 , n361303 , n361304 , n361305 , n13630 , n361307 , n361308 , 
 n13633 , n13634 , n361311 , n361312 , n13637 , n361314 , n361315 , n13640 , n13641 , n13642 , 
 n13643 , n361320 , n361321 , n13646 , n13647 , n13648 , n13649 , n13650 , n361327 , n361328 , 
 n13653 , n361330 , n13655 , n13656 , n13657 , n13658 , n361335 , n361336 , n361337 , n13662 , 
 n361339 , n13664 , n13665 , n361342 , n361343 , n13668 , n361345 , n361346 , n13671 , n361348 , 
 n361349 , n13674 , n361351 , n13676 , n13677 , n361354 , n13679 , n361356 , n13681 , n361358 , 
 n361359 , n13684 , n361361 , n13686 , n361363 , n13688 , n361365 , n13690 , n13691 , n361368 , 
 n361369 , n361370 , n13695 , n361372 , n361373 , n13698 , n361375 , n361376 , n13701 , n361378 , 
 n13703 , n361380 , n13705 , n13706 , n13707 , n13708 , n13709 , n361386 , n361387 , n13712 , 
 n361389 , n13714 , n13715 , n13716 , n13717 , n13718 , n361395 , n13720 , n13721 , n13722 , 
 n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , 
 n13733 , n13734 , n13735 , n13736 , n13737 , n361414 , n13739 , n13740 , n13741 , n13742 , 
 n361419 , n361420 , n13745 , n13746 , n13747 , n13748 , n361425 , n361426 , n13751 , n13752 , 
 n13753 , n13754 , n13755 , n13756 , n13757 , n361434 , n13759 , n361436 , n13761 , n13762 , 
 n361439 , n361440 , n361441 , n13766 , n361443 , n361444 , n13769 , n361446 , n361447 , n13772 , 
 n361449 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n361456 , n13781 , n361458 , 
 n13783 , n13784 , n361461 , n361462 , n361463 , n13788 , n361465 , n361466 , n13791 , n361468 , 
 n361469 , n13794 , n361471 , n13796 , n13797 , n13798 , n13799 , n13800 , n361477 , n13802 , 
 n361479 , n361480 , n361481 , n361482 , n13807 , n361484 , n361485 , n361486 , n13811 , n361488 , 
 n13813 , n13814 , n361491 , n361492 , n361493 , n13818 , n361495 , n361496 , n13821 , n361498 , 
 n361499 , n13824 , n361501 , n361502 , n13827 , n13828 , n13829 , n13830 , n361507 , n361508 , 
 n361509 , n13834 , n361511 , n361512 , n13837 , n361514 , n13839 , n361516 , n13841 , n361518 , 
 n361519 , n13844 , n361521 , n361522 , n361523 , n361524 , n13849 , n361526 , n361527 , n13852 , 
 n361529 , n13854 , n13855 , n361532 , n13857 , n361534 , n13859 , n361536 , n361537 , n13862 , 
 n361539 , n361540 , n13865 , n13866 , n13867 , n13868 , n13869 , n361546 , n361547 , n13872 , 
 n361549 , n361550 , n13875 , n13876 , n13877 , n13878 , n13879 , n361556 , n361557 , n13882 , 
 n361559 , n13884 , n13885 , n13886 , n13887 , n13888 , n361565 , n13890 , n13891 , n13892 , 
 n361569 , n13894 , n361571 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , 
 n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , 
 n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , 
 n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , 
 n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , 
 n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , 
 n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , 
 n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , 
 n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , 
 n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , 
 n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , 
 n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , 
 n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , 
 n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , 
 n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , 
 n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , 
 n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , 
 n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , 
 n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , 
 n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , 
 n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , 
 n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , 
 n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , 
 n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , 
 n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n361815 , n361816 , n14141 , n361818 , 
 n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , 
 n14153 , n14154 , n14155 , n361832 , n14157 , n14158 , n14159 , n14160 , n361837 , n361838 , 
 n361839 , n14164 , n361841 , n361842 , n361843 , n14168 , n361845 , n14170 , n14171 , n361848 , 
 n361849 , n14174 , n361851 , n14176 , n361853 , n361854 , n14179 , n361856 , n361857 , n14182 , 
 n361859 , n361860 , n14185 , n361862 , n361863 , n361864 , n14189 , n361866 , n14191 , n14192 , 
 n361869 , n361870 , n361871 , n14196 , n361873 , n361874 , n14199 , n361876 , n361877 , n14202 , 
 n361879 , n361880 , n14205 , n361882 , n14207 , n361884 , n14209 , n14210 , n361887 , n361888 , 
 n361889 , n14214 , n361891 , n361892 , n14217 , n361894 , n361895 , n14220 , n361897 , n361898 , 
 n14223 , n361900 , n361901 , n14226 , n361903 , n361904 , n14229 , n361906 , n14231 , n14232 , 
 n361909 , n361910 , n361911 , n14236 , n361913 , n361914 , n14239 , n361916 , n361917 , n14242 , 
 n361919 , n361920 , n14245 , n361922 , n361923 , n14248 , n361925 , n14250 , n361927 , n361928 , 
 n14253 , n361930 , n361931 , n14256 , n14257 , n361934 , n361935 , n14260 , n14261 , n361938 , 
 n361939 , n361940 , n361941 , n14266 , n361943 , n14268 , n14269 , n14270 , n14271 , n361948 , 
 n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n361955 , n14280 , n14281 , n361958 , 
 n361959 , n14284 , n361961 , n14286 , n14287 , n14288 , n14289 , n361966 , n361967 , n14292 , 
 n361969 , n14294 , n14295 , n361972 , n14297 , n14298 , n14299 , n14300 , n14301 , n361978 , 
 n361979 , n14304 , n361981 , n361982 , n14307 , n14308 , n14309 , n14310 , n361987 , n14312 , 
 n14313 , n14314 , n14315 , n14316 , n361993 , n361994 , n14319 , n14320 , n14321 , n14322 , 
 n361999 , n362000 , n14325 , n14326 , n14327 , n14328 , n362005 , n362006 , n14331 , n14332 , 
 n14333 , n14334 , n14335 , n362012 , n362013 , n362014 , n14339 , n362016 , n14341 , n14342 , 
 n362019 , n362020 , n362021 , n14346 , n362023 , n362024 , n14349 , n362026 , n362027 , n14352 , 
 n362029 , n362030 , n14355 , n14356 , n14357 , n14358 , n362035 , n14360 , n362037 , n14362 , 
 n362039 , n14364 , n14365 , n362042 , n362043 , n362044 , n14369 , n362046 , n362047 , n14372 , 
 n362049 , n362050 , n14375 , n362052 , n362053 , n14378 , n362055 , n362056 , n14381 , n14382 , 
 n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n362065 , n362066 , n14391 , n362068 , 
 n362069 , n14394 , n362071 , n14396 , n14397 , n362074 , n362075 , n362076 , n14401 , n362078 , 
 n362079 , n14404 , n362081 , n362082 , n14407 , n362084 , n14409 , n362086 , n14411 , n362088 , 
 n14413 , n14414 , n362091 , n362092 , n362093 , n14418 , n362095 , n362096 , n14421 , n362098 , 
 n362099 , n14424 , n362101 , n14426 , n14427 , n362104 , n14429 , n362106 , n362107 , n14432 , 
 n362109 , n362110 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n362118 , 
 n14443 , n362120 , n362121 , n14446 , n362123 , n362124 , n14449 , n362126 , n362127 , n14452 , 
 n362129 , n14454 , n362131 , n362132 , n14457 , n362134 , n14459 , n14460 , n14461 , n14462 , 
 n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , 
 n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , 
 n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , 
 n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , 
 n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , 
 n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , 
 n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , 
 n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , 
 n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , 
 n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , 
 n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , 
 n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , 
 n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , 
 n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , 
 n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , 
 n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , 
 n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , 
 n362309 , n362310 , n14635 , n14636 , n14637 , n14638 , n362315 , n362316 , n362317 , n14642 , 
 n362319 , n14644 , n14645 , n14646 , n362323 , n362324 , n14649 , n362326 , n14651 , n14652 , 
 n362329 , n14654 , n362331 , n14656 , n14657 , n362334 , n362335 , n362336 , n14661 , n362338 , 
 n362339 , n14664 , n362341 , n362342 , n14667 , n362344 , n14669 , n362346 , n14671 , n14672 , 
 n14673 , n14674 , n362351 , n362352 , n14677 , n362354 , n14679 , n362356 , n14681 , n14682 , 
 n362359 , n362360 , n362361 , n14686 , n362363 , n362364 , n14689 , n362366 , n362367 , n14692 , 
 n362369 , n362370 , n362371 , n14696 , n362373 , n14698 , n362375 , n362376 , n14701 , n14702 , 
 n362379 , n362380 , n362381 , n14706 , n362383 , n362384 , n14709 , n362386 , n362387 , n14712 , 
 n362389 , n362390 , n14715 , n362392 , n362393 , n14718 , n14719 , n14720 , n14721 , n14722 , 
 n14723 , n14724 , n362401 , n14726 , n362403 , n362404 , n14729 , n362406 , n362407 , n14732 , 
 n14733 , n14734 , n14735 , n14736 , n362413 , n362414 , n14739 , n362416 , n362417 , n14742 , 
 n362419 , n362420 , n14745 , n14746 , n362423 , n14748 , n14749 , n362426 , n14751 , n14752 , 
 n14753 , n14754 , n362431 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , 
 n14763 , n14764 , n14765 , n14766 , n362443 , n14768 , n14769 , n14770 , n14771 , n362448 , 
 n362449 , n362450 , n362451 , n14776 , n362453 , n362454 , n362455 , n14780 , n362457 , n14782 , 
 n14783 , n362460 , n362461 , n362462 , n14787 , n362464 , n362465 , n14790 , n362467 , n362468 , 
 n14793 , n362470 , n362471 , n14796 , n362473 , n14798 , n362475 , n14800 , n14801 , n362478 , 
 n362479 , n14804 , n362481 , n362482 , n14807 , n362484 , n362485 , n14810 , n362487 , n362488 , 
 n362489 , n14814 , n362491 , n14816 , n14817 , n362494 , n14819 , n362496 , n362497 , n362498 , 
 n362499 , n14824 , n362501 , n362502 , n14827 , n362504 , n362505 , n14830 , n362507 , n14832 , 
 n362509 , n14834 , n14835 , n362512 , n362513 , n362514 , n14839 , n362516 , n362517 , n14842 , 
 n362519 , n362520 , n14845 , n362522 , n362523 , n362524 , n14849 , n362526 , n14851 , n14852 , 
 n362529 , n362530 , n362531 , n14856 , n362533 , n362534 , n14859 , n362536 , n362537 , n14862 , 
 n362539 , n362540 , n14865 , n362542 , n362543 , n14868 , n14869 , n14870 , n14871 , n14872 , 
 n362549 , n362550 , n14875 , n362552 , n362553 , n14878 , n362555 , n362556 , n14881 , n362558 , 
 n362559 , n14884 , n362561 , n362562 , n14887 , n362564 , n14889 , n14890 , n362567 , n362568 , 
 n14893 , n362570 , n362571 , n14896 , n362573 , n362574 , n14899 , n362576 , n362577 , n14902 , 
 n362579 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , 
 n362589 , n14914 , n14915 , n14916 , n14917 , n362594 , n362595 , n14920 , n362597 , n362598 , 
 n14923 , n362600 , n362601 , n362602 , n362603 , n14928 , n362605 , n362606 , n14931 , n362608 , 
 n14933 , n362610 , n14935 , n362612 , n14937 , n362614 , n362615 , n362616 , n14941 , n362618 , 
 n362619 , n14944 , n362621 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , 
 n14953 , n14954 , n14955 , n14956 , n362633 , n14958 , n362635 , n14960 , n14961 , n14962 , 
 n14963 , n14964 , n14965 , n14966 , n362643 , n14968 , n362645 , n14970 , n14971 , n14972 , 
 n14973 , n14974 , n14975 , n362652 , n362653 , n14978 , n362655 , n14980 , n14981 , n14982 , 
 n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n362665 , n362666 , n14991 , n362668 , 
 n14993 , n362670 , n14995 , n14996 , n362673 , n362674 , n14999 , n362676 , n362677 , n15002 , 
 n362679 , n15004 , n362681 , n362682 , n15007 , n362684 , n362685 , n15010 , n362687 , n362688 , 
 n15013 , n362690 , n362691 , n15016 , n15017 , n15018 , n15019 , n362696 , n362697 , n15022 , 
 n15023 , n15024 , n15025 , n362702 , n362703 , n15028 , n15029 , n15030 , n15031 , n15032 , 
 n362709 , n362710 , n15035 , n362712 , n362713 , n362714 , n15039 , n362716 , n15041 , n362718 , 
 n15043 , n15044 , n362721 , n362722 , n362723 , n15048 , n362725 , n362726 , n15051 , n362728 , 
 n362729 , n15054 , n362731 , n362732 , n15057 , n362734 , n15059 , n15060 , n15061 , n15062 , 
 n15063 , n15064 , n362741 , n15066 , n362743 , n362744 , n15069 , n362746 , n15071 , n15072 , 
 n362749 , n15074 , n362751 , n362752 , n15077 , n362754 , n15079 , n15080 , n362757 , n362758 , 
 n362759 , n15084 , n362761 , n362762 , n15087 , n362764 , n362765 , n15090 , n362767 , n15092 , 
 n15093 , n15094 , n15095 , n15096 , n15097 , n362774 , n15099 , n362776 , n15101 , n15102 , 
 n362779 , n362780 , n362781 , n15106 , n362783 , n362784 , n15109 , n362786 , n362787 , n15112 , 
 n362789 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n362798 , 
 n15123 , n15124 , n15125 , n15126 , n15127 , n362804 , n362805 , n15130 , n362807 , n362808 , 
 n15133 , n15134 , n15135 , n15136 , n362813 , n362814 , n15139 , n15140 , n15141 , n15142 , 
 n15143 , n362820 , n362821 , n15146 , n15147 , n15148 , n15149 , n362826 , n362827 , n362828 , 
 n362829 , n15154 , n362831 , n362832 , n362833 , n15158 , n362835 , n15160 , n362837 , n15162 , 
 n15163 , n362840 , n362841 , n362842 , n15167 , n362844 , n362845 , n15170 , n362847 , n362848 , 
 n15173 , n362850 , n362851 , n15176 , n362853 , n362854 , n15179 , n362856 , n15181 , n362858 , 
 n15183 , n15184 , n362861 , n362862 , n362863 , n15188 , n362865 , n362866 , n15191 , n362868 , 
 n362869 , n15194 , n362871 , n362872 , n362873 , n15198 , n362875 , n15200 , n15201 , n362878 , 
 n15203 , n362880 , n15205 , n362882 , n362883 , n15208 , n362885 , n362886 , n15211 , n362888 , 
 n362889 , n15214 , n362891 , n15216 , n362893 , n362894 , n15219 , n362896 , n362897 , n15222 , 
 n362899 , n362900 , n15225 , n15226 , n15227 , n15228 , n15229 , n362906 , n362907 , n15232 , 
 n362909 , n362910 , n15235 , n362912 , n362913 , n15238 , n362915 , n15240 , n362917 , n15242 , 
 n15243 , n362920 , n362921 , n15246 , n362923 , n15248 , n362925 , n362926 , n15251 , n362928 , 
 n362929 , n15254 , n362931 , n362932 , n15257 , n362934 , n15259 , n362936 , n362937 , n15262 , 
 n362939 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , 
 n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , 
 n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , 
 n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , 
 n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , 
 n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , 
 n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , 
 n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , 
 n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , 
 n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n363037 , n363038 , 
 n15363 , n15364 , n15365 , n15366 , n363043 , n363044 , n15369 , n15370 , n15371 , n15372 , 
 n15373 , n363050 , n363051 , n363052 , n15377 , n363054 , n15379 , n15380 , n363057 , n363058 , 
 n15383 , n363060 , n363061 , n15386 , n363063 , n363064 , n15389 , n363066 , n363067 , n15392 , 
 n15393 , n15394 , n15395 , n363072 , n363073 , n15398 , n363075 , n363076 , n15401 , n363078 , 
 n363079 , n363080 , n15405 , n363082 , n15407 , n15408 , n363085 , n15410 , n363087 , n15412 , 
 n363089 , n363090 , n15415 , n363092 , n363093 , n15418 , n363095 , n15420 , n363097 , n15422 , 
 n15423 , n363100 , n363101 , n363102 , n15427 , n363104 , n363105 , n15430 , n363107 , n363108 , 
 n15433 , n363110 , n363111 , n15436 , n363113 , n363114 , n15439 , n363116 , n363117 , n15442 , 
 n15443 , n15444 , n15445 , n15446 , n363123 , n363124 , n15449 , n363126 , n363127 , n15452 , 
 n15453 , n15454 , n15455 , n363132 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , 
 n15463 , n15464 , n15465 , n15466 , n15467 , n363144 , n363145 , n15470 , n363147 , n15472 , 
 n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n363158 , 
 n363159 , n15484 , n363161 , n363162 , n15487 , n363164 , n15489 , n15490 , n363167 , n363168 , 
 n363169 , n15494 , n363171 , n363172 , n15497 , n363174 , n363175 , n15500 , n363177 , n15502 , 
 n363179 , n15504 , n363181 , n15506 , n15507 , n363184 , n363185 , n363186 , n15511 , n363188 , 
 n363189 , n15514 , n363191 , n363192 , n15517 , n363194 , n15519 , n15520 , n15521 , n363198 , 
 n15523 , n15524 , n15525 , n15526 , n15527 , n363204 , n363205 , n15530 , n363207 , n363208 , 
 n15533 , n363210 , n363211 , n15536 , n15537 , n15538 , n15539 , n363216 , n363217 , n15542 , 
 n363219 , n363220 , n15545 , n363222 , n363223 , n363224 , n15549 , n363226 , n363227 , n15552 , 
 n363229 , n15554 , n15555 , n15556 , n363233 , n363234 , n15559 , n363236 , n363237 , n15562 , 
 n363239 , n15564 , n15565 , n363242 , n363243 , n15568 , n363245 , n15570 , n363247 , n15572 , 
 n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , 
 n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , 
 n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , 
 n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , 
 n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , 
 n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , 
 n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , 
 n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , 
 n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , 
 n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , 
 n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , 
 n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , 
 n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , 
 n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , 
 n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , 
 n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n363405 , n363406 , n15731 , n15732 , 
 n15733 , n15734 , n363411 , n363412 , n363413 , n363414 , n15739 , n363416 , n363417 , n363418 , 
 n15743 , n363420 , n15745 , n15746 , n363423 , n15748 , n15749 , n15750 , n15751 , n363428 , 
 n15753 , n363430 , n363431 , n15756 , n363433 , n363434 , n15759 , n363436 , n363437 , n15762 , 
 n363439 , n15764 , n363441 , n363442 , n15767 , n363444 , n363445 , n363446 , n363447 , n15772 , 
 n363449 , n15774 , n15775 , n363452 , n363453 , n363454 , n15779 , n363456 , n363457 , n15782 , 
 n363459 , n363460 , n15785 , n363462 , n363463 , n15788 , n15789 , n15790 , n15791 , n15792 , 
 n363469 , n363470 , n15795 , n363472 , n363473 , n15798 , n15799 , n15800 , n15801 , n15802 , 
 n363479 , n363480 , n15805 , n363482 , n363483 , n15808 , n15809 , n15810 , n15811 , n363488 , 
 n15813 , n363490 , n15815 , n15816 , n363493 , n363494 , n363495 , n15820 , n363497 , n363498 , 
 n15823 , n363500 , n363501 , n15826 , n363503 , n15828 , n15829 , n15830 , n15831 , n15832 , 
 n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n363515 , n363516 , n15841 , n363518 , 
 n363519 , n363520 , n15845 , n363522 , n15847 , n15848 , n363525 , n363526 , n363527 , n15852 , 
 n363529 , n363530 , n15855 , n363532 , n363533 , n15858 , n363535 , n363536 , n15861 , n363538 , 
 n363539 , n15864 , n363541 , n15866 , n363543 , n363544 , n15869 , n363546 , n15871 , n363548 , 
 n15873 , n15874 , n15875 , n15876 , n15877 , n363554 , n15879 , n363556 , n363557 , n15882 , 
 n15883 , n15884 , n15885 , n15886 , n363563 , n363564 , n15889 , n363566 , n363567 , n15892 , 
 n363569 , n363570 , n363571 , n15896 , n363573 , n15898 , n15899 , n15900 , n15901 , n15902 , 
 n363579 , n15904 , n363581 , n15906 , n15907 , n363584 , n15909 , n363586 , n15911 , n15912 , 
 n15913 , n15914 , n15915 , n363592 , n15917 , n363594 , n15919 , n15920 , n15921 , n15922 , 
 n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , 
 n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , 
 n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , 
 n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , 
 n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , 
 n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , 
 n15983 , n15984 , n15985 , n363662 , n363663 , n15988 , n363665 , n363666 , n15991 , n363668 , 
 n15993 , n15994 , n363671 , n363672 , n15997 , n363674 , n15999 , n363676 , n363677 , n16002 , 
 n363679 , n16004 , n363681 , n363682 , n16007 , n363684 , n16009 , n363686 , n363687 , n16012 , 
 n363689 , n363690 , n363691 , n16016 , n363693 , n16018 , n16019 , n16020 , n16021 , n16022 , 
 n363699 , n363700 , n16025 , n16026 , n16027 , n16028 , n16029 , n363706 , n363707 , n16032 , 
 n16033 , n16034 , n16035 , n363712 , n363713 , n16038 , n363715 , n363716 , n363717 , n16042 , 
 n363719 , n16044 , n16045 , n363722 , n363723 , n363724 , n16049 , n363726 , n363727 , n16052 , 
 n363729 , n363730 , n16055 , n363732 , n363733 , n16058 , n363735 , n16060 , n363737 , n16062 , 
 n16063 , n363740 , n363741 , n16066 , n363743 , n363744 , n16069 , n363746 , n363747 , n16072 , 
 n363749 , n363750 , n16075 , n363752 , n363753 , n16078 , n16079 , n16080 , n16081 , n16082 , 
 n16083 , n16084 , n363761 , n16086 , n363763 , n363764 , n16089 , n16090 , n16091 , n16092 , 
 n363769 , n363770 , n16095 , n16096 , n16097 , n363774 , n363775 , n363776 , n16101 , n363778 , 
 n363779 , n16104 , n363781 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , 
 n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , 
 n363799 , n16124 , n16125 , n16126 , n16127 , n16128 , n363805 , n363806 , n16131 , n363808 , 
 n363809 , n16134 , n16135 , n16136 , n16137 , n16138 , n363815 , n16140 , n363817 , n363818 , 
 n16143 , n16144 , n16145 , n16146 , n16147 , n363824 , n363825 , n16150 , n363827 , n363828 , 
 n16153 , n363830 , n363831 , n16156 , n363833 , n363834 , n16159 , n363836 , n16161 , n363838 , 
 n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , 
 n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , 
 n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , 
 n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , 
 n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , 
 n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , 
 n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , 
 n16233 , n16234 , n363911 , n363912 , n16237 , n16238 , n16239 , n16240 , n16241 , n363918 , 
 n363919 , n363920 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n363928 , 
 n16253 , n16254 , n363931 , n363932 , n16257 , n16258 , n363935 , n16260 , n363937 , n16262 , 
 n363939 , n16264 , n16265 , n363942 , n363943 , n16268 , n363945 , n363946 , n16271 , n363948 , 
 n16273 , n363950 , n363951 , n16276 , n363953 , n363954 , n16279 , n363956 , n363957 , n16282 , 
 n363959 , n363960 , n363961 , n16286 , n16287 , n16288 , n16289 , n363966 , n363967 , n16292 , 
 n16293 , n363970 , n363971 , n363972 , n16297 , n363974 , n16299 , n16300 , n363977 , n363978 , 
 n16303 , n363980 , n363981 , n16306 , n363983 , n16308 , n363985 , n363986 , n16311 , n363988 , 
 n363989 , n16314 , n363991 , n363992 , n16317 , n363994 , n16319 , n363996 , n363997 , n16322 , 
 n363999 , n364000 , n16325 , n364002 , n364003 , n16328 , n16329 , n16330 , n16331 , n16332 , 
 n364009 , n364010 , n16335 , n364012 , n364013 , n16338 , n16339 , n16340 , n16341 , n16342 , 
 n364019 , n364020 , n16345 , n364022 , n364023 , n16348 , n364025 , n364026 , n16351 , n364028 , 
 n364029 , n364030 , n16355 , n364032 , n16357 , n364034 , n364035 , n16360 , n364037 , n16362 , 
 n16363 , n16364 , n16365 , n364042 , n364043 , n16368 , n364045 , n364046 , n16371 , n364048 , 
 n16373 , n16374 , n364051 , n16376 , n364053 , n16378 , n364055 , n364056 , n16381 , n16382 , 
 n364059 , n16384 , n364061 , n364062 , n16387 , n364064 , n364065 , n16390 , n364067 , n364068 , 
 n16393 , n364070 , n364071 , n364072 , n16397 , n364074 , n364075 , n16400 , n364077 , n364078 , 
 n364079 , n364080 , n364081 , n16406 , n364083 , n364084 , n16409 , n364086 , n16411 , n16412 , 
 n16413 , n16414 , n364091 , n364092 , n16417 , n16418 , n16419 , n16420 , n364097 , n364098 , 
 n364099 , n364100 , n16425 , n364102 , n364103 , n364104 , n16429 , n364106 , n364107 , n364108 , 
 n16433 , n364110 , n16435 , n364112 , n364113 , n364114 , n16439 , n16440 , n364117 , n364118 , 
 n16443 , n16444 , n16445 , n16446 , n16447 , n364124 , n364125 , n16450 , n364127 , n364128 , 
 n364129 , n364130 , n16455 , n364132 , n364133 , n364134 , n16459 , n364136 , n364137 , n364138 , 
 n16463 , n364140 , n16465 , n364142 , n364143 , n364144 , n16469 , n16470 , n364147 , n364148 , 
 n16473 , n16474 , n16475 , n16476 , n16477 , n364154 , n364155 , n16480 , n364157 , n364158 , 
 n16483 , n16484 , n16485 , n16486 , n16487 , n364164 , n364165 , n16490 , n364167 , n364168 , 
 n16493 , n16494 , n16495 , n16496 , n16497 , n364174 , n364175 , n16500 , n364177 , n364178 , 
 n16503 , n364180 , n364181 , n364182 , n364183 , n16508 , n364185 , n364186 , n16511 , n364188 , 
 n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , 
 n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , 
 n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , 
 n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , 
 n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , 
 n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , 
 n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , 
 n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , 
 n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , 
 n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , 
 n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , 
 n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , 
 n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , 
 n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n364327 , n16652 , 
 n364329 , n16654 , n364331 , n364332 , n16657 , n364334 , n16659 , n16660 , n364337 , n16662 , 
 n364339 , n16664 , n16665 , n364342 , n16667 , n364344 , n364345 , n16670 , n364347 , n364348 , 
 n16673 , n364350 , n364351 , n364352 , n16677 , n364354 , n364355 , n16680 , n364357 , n364358 , 
 n364359 , n364360 , n364361 , n16686 , n364363 , n364364 , n16689 , n364366 , n364367 , n364368 , 
 n16693 , n364370 , n364371 , n16696 , n364373 , n364374 , n16699 , n364376 , n16701 , n364378 , 
 n364379 , n16704 , n16705 , n364382 , n364383 , n16708 , n16709 , n364386 , n364387 , n364388 , 
 n16713 , n364390 , n364391 , n16716 , n16717 , n16718 , n16719 , n16720 , n364397 , n364398 , 
 n364399 , n364400 , n16725 , n364402 , n364403 , n16728 , n364405 , n364406 , n16731 , n364408 , 
 n16733 , n364410 , n364411 , n16736 , n16737 , n364414 , n364415 , n16740 , n16741 , n364418 , 
 n364419 , n364420 , n16745 , n364422 , n364423 , n16748 , n364425 , n364426 , n16751 , n16752 , 
 n364429 , n364430 , n16755 , n16756 , n364433 , n364434 , n16759 , n16760 , n16761 , n16762 , 
 n364439 , n364440 , n16765 , n16766 , n16767 , n16768 , n364445 , n364446 , n16771 , n364448 , 
 n364449 , n16774 , n364451 , n364452 , n16777 , n16778 , n16779 , n16780 , n16781 , n364458 , 
 n364459 , n16784 , n16785 , n364462 , n364463 , n16788 , n16789 , n364466 , n16791 , n16792 , 
 n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , 
 n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , 
 n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , 
 n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , 
 n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , 
 n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , 
 n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , 
 n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , 
 n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , 
 n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , 
 n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , 
 n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , 
 n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , 
 n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , 
 n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , 
 n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , 
 n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , 
 n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , 
 n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , 
 n364659 , n16984 , n364661 , n364662 , n16987 , n364664 , n16989 , n16990 , n16991 , n16992 , 
 n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , 
 n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , 
 n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , 
 n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n364708 , 
 n364709 , n17034 , n17035 , n17036 , n17037 , n364714 , n17039 , n364716 , n17041 , n364718 , 
 n17043 , n364720 , n364721 , n17046 , n17047 , n364724 , n364725 , n17050 , n364727 , n364728 , 
 n17053 , n364730 , n364731 , n17056 , n364733 , n364734 , n17059 , n17060 , n364737 , n17062 , 
 n364739 , n17064 , n17065 , n364742 , n364743 , n17068 , n364745 , n364746 , n17071 , n364748 , 
 n364749 , n364750 , n364751 , n17076 , n364753 , n17078 , n17079 , n17080 , n17081 , n17082 , 
 n364759 , n17084 , n364761 , n364762 , n17087 , n364764 , n364765 , n364766 , n364767 , n17092 , 
 n364769 , n17094 , n364771 , n364772 , n364773 , n17098 , n17099 , n364776 , n364777 , n17102 , 
 n364779 , n364780 , n17105 , n17106 , n364783 , n17108 , n17109 , n364786 , n17111 , n364788 , 
 n17113 , n364790 , n364791 , n17116 , n17117 , n364794 , n364795 , n17120 , n364797 , n364798 , 
 n17123 , n364800 , n364801 , n17126 , n364803 , n364804 , n17129 , n17130 , n17131 , n17132 , 
 n364809 , n17133 , n364811 , n17135 , n364813 , n364814 , n17138 , n364816 , n364817 , n17141 , 
 n364819 , n17143 , n364821 , n17145 , n364823 , n364824 , n17148 , n364826 , n364827 , n17151 , 
 n364829 , n364830 , n364831 , n364832 , n17156 , n364834 , n364835 , n17159 , n364837 , n17161 , 
 n364839 , n17163 , n364841 , n364842 , n17166 , n17167 , n364845 , n17169 , n17170 , n17171 , 
 n17172 , n17173 , n17174 , n364852 , n17176 , n364854 , n364855 , n17179 , n17180 , n17181 , 
 n17182 , n364860 , n17184 , n364862 , n364863 , n17187 , n364865 , n364866 , n17190 , n364868 , 
 n364869 , n17193 , n17194 , n17195 , n17196 , n17197 , n364875 , n364876 , n364877 , n17201 , 
 n364879 , n364880 , n17204 , n364882 , n364883 , n17207 , n364885 , n17209 , n17210 , n17211 , 
 n364889 , n17213 , n364891 , n17215 , n17216 , n364894 , n17218 , n364896 , n17220 , n364898 , 
 n364899 , n364900 , n364901 , n17221 , n364903 , n364904 , n17223 , n364906 , n364907 , n17226 , 
 n364909 , n17228 , n17229 , n17230 , n17231 , n17232 , n364915 , n17234 , n364917 , n364918 , 
 n17237 , n364920 , n364921 , n364922 , n364923 , n17242 , n364925 , n364926 , n17245 , n364928 , 
 n17247 , n17248 , n17249 , n17250 , n17251 , n364934 , n17253 , n364936 , n364937 , n17256 , 
 n17257 , n17258 , n364941 , n17260 , n364943 , n364944 , n17263 , n17264 , n364947 , n17266 , 
 n364949 , n17268 , n364951 , n364952 , n17271 , n17272 , n364955 , n364956 , n17275 , n364958 , 
 n364959 , n17278 , n364961 , n364962 , n364963 , n364964 , n17283 , n364966 , n364967 , n364968 , 
 n17287 , n364970 , n364971 , n17290 , n364973 , n364974 , n17293 , n364976 , n364977 , n17296 , 
 n364979 , n364980 , n364981 , n17300 , n17301 , n364984 , n17303 , n364986 , n364987 , n364988 , 
 n364989 , n364990 , n364991 , n364992 , n17306 , n364994 , n17307 , n17308 , n17309 , n364998 , 
 n364999 , n365000 , n17313 , n365002 , n365003 , n17316 , n365005 , n365006 , n17319 , n365008 , 
 n17321 , n17322 , n17323 , n17324 , n17325 , n365014 , n17327 , n17328 , n365017 , n17330 , 
 n365019 , n17332 , n17333 , n365022 , n17335 , n365024 , n365025 , n17338 , n365027 , n365028 , 
 n17341 , n365030 , n17343 , n365032 , n365033 , n17346 , n365035 , n365036 , n365037 , n17350 , 
 n365039 , n365040 , n365041 , n17354 , n365043 , n17356 , n365045 , n17358 , n17359 , n365048 , 
 n365049 , n17362 , n365051 , n365052 , n17365 , n365054 , n365055 , n17368 , n17369 , n365058 , 
 n17371 , n17372 , n365061 , n17374 , n365063 , n365064 , n17377 , n17378 , n365067 , n365068 , 
 n17381 , n365070 , n365071 , n365072 , n365073 , n365074 , n365075 , n17383 , n365077 , n365078 , 
 n17385 , n365080 , n365081 , n17388 , n365083 , n17390 , n17391 , n365086 , n17393 , n17394 , 
 n365089 , n17396 , n365091 , n17398 , n365093 , n365094 , n17401 , n17402 , n365097 , n17404 , 
 n365099 , n365100 , n365101 , n17408 , n365103 , n365104 , n17411 , n365106 , n365107 , n365108 , 
 n17415 , n365110 , n365111 , n17418 , n365113 , n365114 , n17421 , n17422 , n17423 , n365118 , 
 n365119 , n365120 , n17427 , n365122 , n17429 , n17430 , n365125 , n17432 , n365127 , n17434 , 
 n365129 , n365130 , n17437 , n17438 , n365133 , n365134 , n17441 , n365136 , n365137 , n17444 , 
 n365139 , n365140 , n365141 , n17448 , n365143 , n365144 , n17451 , n365146 , n365147 , n17454 , 
 n365149 , n365150 , n365151 , n365152 , n365153 , n365154 , n17456 , n365156 , n17457 , n17458 , 
 n365159 , n17460 , n365161 , n365162 , n365163 , n17464 , n365165 , n365166 , n17467 , n365168 , 
 n365169 , n17470 , n17471 , n365172 , n17473 , n365174 , n17475 , n365176 , n365177 , n17478 , 
 n17479 , n17480 , n365181 , n17482 , n365183 , n365184 , n365185 , n17486 , n365187 , n365188 , 
 n17489 , n365190 , n365191 , n17492 , n17493 , n17494 , n365195 , n365196 , n17497 , n17498 , 
 n17499 , n365200 , n365201 , n17502 , n17503 , n17504 , n17505 , n17506 , n365207 , n365208 , 
 n365209 , n17510 , n365211 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , 
 n17519 , n17520 , n365221 , n365222 , n365223 , n365224 , n365225 , n17521 , n365227 , n365228 , 
 n17523 , n365230 , n365231 , n17526 , n17527 , n365234 , n365235 , n17530 , n365237 , n365238 , 
 n17533 , n365240 , n365241 , n17536 , n365243 , n17538 , n365245 , n17540 , n17541 , n365248 , 
 n17543 , n365250 , n17545 , n17546 , n17547 , n365254 , n365255 , n17550 , n365257 , n365258 , 
 n17553 , n365260 , n365261 , n365262 , n17557 , n365264 , n365265 , n17560 , n365267 , n365268 , 
 n365269 , n17564 , n365271 , n17566 , n17567 , n365274 , n365275 , n17570 , n365277 , n365278 , 
 n17573 , n365280 , n365281 , n17576 , n365283 , n365284 , n17579 , n365286 , n365287 , n365288 , 
 n365289 , n365290 , n365291 , n17581 , n365293 , n365294 , n17583 , n365296 , n365297 , n17586 , 
 n365299 , n365300 , n17589 , n365302 , n17591 , n365304 , n17593 , n17594 , n365307 , n365308 , 
 n17597 , n365310 , n365311 , n17600 , n365313 , n365314 , n17603 , n17604 , n17605 , n365318 , 
 n365319 , n17608 , n17609 , n17610 , n365323 , n365324 , n17613 , n365326 , n365327 , n17616 , 
 n365329 , n365330 , n365331 , n365332 , n17621 , n365334 , n365335 , n17624 , n365337 , n17626 , 
 n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n365347 , n365348 , 
 n365349 , n365350 , n365351 , n17635 , n365353 , n365354 , n365355 , n365356 , n365357 , n17640 , 
 n365359 , n365360 , n17643 , n365362 , n17645 , n17646 , n365365 , n365366 , n17649 , n365368 , 
 n365369 , n365370 , n17653 , n365372 , n365373 , n17656 , n365375 , n17658 , n17659 , n17660 , 
 n365379 , n365380 , n17663 , n365382 , n17665 , n17666 , n17667 , n365386 , n17669 , n365388 , 
 n17671 , n17672 , n365391 , n365392 , n17675 , n365394 , n17677 , n17678 , n365397 , n17680 , 
 n365399 , n365400 , n365401 , n365402 , n365403 , n365404 , n365405 , n365406 , n365407 , n365408 , 
 n17685 , n365410 , n17687 , n17688 , n17689 , n365414 , n17691 , n365416 , n17693 , n17694 , 
 n365419 , n365420 , n17697 , n365422 , n365423 , n17700 , n365425 , n17702 , n365427 , n365428 , 
 n17705 , n365430 , n17707 , n17708 , n365433 , n17710 , n365435 , n17712 , n365437 , n17714 , 
 n365439 , n17716 , n17717 , n365442 , n365443 , n17720 , n365445 , n365446 , n17723 , n365448 , 
 n365449 , n365450 , n365451 , n365452 , n365453 , n17725 , n365455 , n365456 , n17727 , n365458 , 
 n365459 , n17730 , n365461 , n365462 , n17733 , n365464 , n365465 , n365466 , n17737 , n365468 , 
 n365469 , n17740 , n365471 , n365472 , n365473 , n17744 , n365475 , n365476 , n365477 , n17748 , 
 n365479 , n365480 , n365481 , n17752 , n17753 , n17754 , n17755 , n17756 , n365487 , n17758 , 
 n17759 , n365490 , n365491 , n365492 , n365493 , n365494 , n365495 , n17761 , n365497 , n365498 , 
 n17763 , n365500 , n365501 , n365502 , n17767 , n365504 , n365505 , n17770 , n365507 , n365508 , 
 n17773 , n365510 , n17775 , n365512 , n17777 , n365514 , n17779 , n365516 , n365517 , n17782 , 
 n17783 , n365520 , n17785 , n365522 , n17787 , n365524 , n365525 , n17790 , n365527 , n365528 , 
 n365529 , n365530 , n365531 , n17791 , n365533 , n365534 , n17793 , n365536 , n365537 , n17796 , 
 n365539 , n365540 , n17799 , n365542 , n365543 , n365544 , n17803 , n365546 , n365547 , n17806 , 
 n365549 , n365550 , n17809 , n17810 , n17811 , n365554 , n365555 , n17814 , n365557 , n365558 , 
 n365559 , n365560 , n365561 , n365562 , n17816 , n365564 , n365565 , n365566 , n17819 , n365568 , 
 n365569 , n17822 , n365571 , n365572 , n17825 , n365574 , n17827 , n365576 , n17829 , n17830 , 
 n365579 , n365580 , n365581 , n365582 , n365583 , n365584 , n365585 , n365586 , n17834 , n365588 , 
 n365589 , n17836 , n17837 , n17838 , n365593 , n365594 , n17841 , n17842 , n17843 , n365598 , 
 n365599 , n365600 , n365601 , n365602 , n365603 , n365604 , n17846 , n365606 , n17847 , n365608 , 
 n365609 , n17850 , n365611 , n365612 , n365613 , n365614 , n365615 , n365616 , n365617 , n365618 , 
 n365619 , n365620 , n365621 , n365622 , n365623 , n365624 , n365625 , n365626 , n365627 , n365628 , 
 n17859 , n365630 , n17861 , n365632 , n17863 , n365634 , n17865 , n365636 , n17867 , n365638 , 
 n17869 , n365640 , n365641 , n365642 , n365643 , n365644 , n17875 , n365646 , n365647 , n365648 , 
 n365649 , n365650 , n365651 , n365652 , n365653 , n365654 , n17885 , n365656 , n365657 , n365658 , 
 n365659 , n365660 , n365661 , n365662 , n17893 , n365664 , n365665 , n365666 , n365667 , n365668 , 
 n17899 , n365670 , n17901 , n365672 , n17903 , n365674 , n17905 , n365676 , n17907 , n365678 , 
 n17909 , n365680 , n365681 , n365682 , n365683 , n365684 , n17915 , n365686 , n365687 , n365688 , 
 n17919 , n365690 , n365691 , n365692 , n17923 , n365694 , n365695 , n365696 , n365697 , n365698 , 
 n17929 , n365700 , n17931 , n365702 , n17933 , n365704 , n365705 , n365706 , n17937 , n365708 , 
 n17939 , n365710 , n17941 , n365712 , n365713 , n365714 , n17945 , n365716 , n17947 , n365718 , 
 n17949 , n365720 , n365721 , n365722 , n365723 , n365724 , n365725 , n365726 , n365727 , n365728 , 
 n365729 , n365730 , n17961 , n365732 , n365733 , n365734 , n365735 , n365736 , n17967 , n365738 , 
 n365739 , n365740 , n365741 , n365742 , n17973 , n365744 , n365745 , n365746 , n17977 , n365748 , 
 n17979 , n365750 , n17981 , n365752 , n365753 , n365754 , n17985 , n365756 , n365757 , n365758 , 
 n365759 , n365760 , n17991 , n365762 , n365763 , n365764 , n17995 , n365766 , n365767 , n365768 , 
 n365769 , n365770 , n365771 , n365772 , n18003 , n365774 , n18005 , n365776 , n365777 , n365778 , 
 n18009 , n365780 , n365781 , n365782 , n365783 , n365784 , n18015 , n365786 , n365787 , n365788 , 
 n18019 , n365790 , n18021 , n365792 , n365793 , n365794 , n365795 , n365796 , n18027 , n365798 , 
 n18029 , n365800 , n18031 , n365802 , n365803 , n365804 , n18035 , n365806 , n365807 , n365808 , 
 n365809 , n365810 , n365811 , n365812 , n18043 , n365814 , n365815 , n365816 , n365817 , n365818 , 
 n18049 , n365820 , n365821 , n365822 , n18053 , n365824 , n365825 , n365826 , n18057 , n365828 , 
 n365829 , n365830 , n18061 , n365832 , n365833 , n365834 , n18065 , n365836 , n18067 , n365838 , 
 n365839 , n365840 , n18071 , n365842 , n18073 , n365844 , n365845 , n365846 , n365847 , n365848 , 
 n18079 , n365850 , n18081 , n365852 , n365853 , n365854 , n18085 , n365856 , n18087 , n365858 , 
 n18089 , n365860 , n365861 , n365862 , n18093 , n365864 , n365865 , n365866 , n365867 , n365868 , 
 n365869 , n365870 , n365871 , n365872 , n18103 , n365874 , n365875 , n365876 , n365877 , n365878 , 
 n365879 , n365880 , n365881 , n365882 , n365883 , n365884 , n365885 , n365886 , n365887 , n365888 , 
 n365889 , n365890 , n365891 , n365892 , n365893 , n365894 , n365895 , n365896 , n365897 , n365898 , 
 n365899 , n365900 , n365901 , n365902 , n365903 , n365904 , n365905 , n365906 , n18130 , n365908 , 
 n365909 , n18133 , n365911 , n365912 , n365913 , n18137 , n18138 , n365916 , n365917 , n365918 , 
 n18142 , n365920 , n365921 , n365922 , n18146 , n365924 , n365925 , n18149 , n365927 , n365928 , 
 n365929 , n18153 , n18154 , n365932 , n365933 , n18157 , n18158 , n365936 , n365937 , n365938 , 
 n18162 , n365940 , n365941 , n18165 , n365943 , n365944 , n365945 , n365946 , n18170 , n365948 , 
 n365949 , n365950 , n365951 , n365952 , n365953 , n18177 , n365955 , n365956 , n365957 , n365958 , 
 n365959 , n365960 , n365961 , n365962 , n18186 , n365964 , n365965 , n18189 , n18190 , n365968 , 
 n365969 , n18193 , n18194 , n365972 , n365973 , n18197 , n365975 , n365976 , n365977 , n365978 , 
 n18202 , n365980 , n365981 , n365982 , n18206 , n365984 , n365985 , n365986 , n18210 , n365988 , 
 n365989 , n18213 , n365991 , n365992 , n365993 , n18217 , n365995 , n365996 , n365997 , n365998 , 
 n365999 , n366000 , n366001 , n366002 , n18226 , n366004 , n366005 , n366006 , n18230 , n366008 , 
 n366009 , n18233 , n366011 , n366012 , n366013 , n366014 , n366015 , n366016 , n366017 , n366018 , 
 n366019 , n366020 , n366021 , n18245 , n366023 , n18247 , n18248 , n366026 , n18250 , n366028 , 
 n366029 , n366030 , n18254 , n366032 , n366033 , n366034 , n18258 , n366036 , n18260 , n18261 , 
 n366039 , n18263 , n366041 , n18265 , n366043 , n366044 , n18268 , n18269 , n366047 , n18271 , 
 n366049 , n366050 , n366051 , n18275 , n366053 , n366054 , n18278 , n366056 , n366057 , n366058 , 
 n18282 , n366060 , n366061 , n18285 , n366063 , n366064 , n18288 , n366066 , n18290 , n366068 , 
 n18292 , n18293 , n366071 , n18295 , n366073 , n18297 , n18298 , n366076 , n366077 , n18301 , 
 n366079 , n366080 , n18304 , n366082 , n366083 , n366084 , n18308 , n366086 , n366087 , n18311 , 
 n366089 , n366090 , n18314 , n18315 , n18316 , n366094 , n366095 , n366096 , n18320 , n366098 , 
 n18322 , n18323 , n366101 , n18325 , n366103 , n18327 , n18328 , n366106 , n366107 , n18331 , 
 n366109 , n366110 , n18334 , n366112 , n366113 , n366114 , n18338 , n366116 , n366117 , n366118 , 
 n366119 , n366120 , n366121 , n366122 , n366123 , n366124 , n366125 , n366126 , n366127 , n366128 , 
 n366129 , n366130 , n366131 , n366132 , n366133 , n366134 , n366135 , n366136 , n366137 , n366138 , 
 n366139 , n366140 , n366141 , n366142 , n366143 , n366144 , n366145 , n366146 , n366147 , n366148 , 
 n366149 , n366150 , n366151 , n366152 , n366153 , n366154 , n366155 , n366156 , n366157 , n366158 , 
 n366159 , n366160 , n366161 , n366162 , n366163 , n366164 , n366165 , n366166 , n366167 , n366168 , 
 n366169 , n366170 , n366171 , n366172 , n366173 , n366174 , n366175 , n366176 , n366177 , n366178 , 
 n366179 , n366180 , n366181 , n366182 , n366183 , n366184 , n366185 , n366186 , n366187 , n366188 , 
 n366189 , n366190 , n366191 , n366192 , n366193 , n366194 , n366195 , n366196 , n366197 , n366198 , 
 n366199 , n366200 , n366201 , n366202 , n366203 , n366204 , n366205 , n366206 , n366207 , n366208 , 
 n366209 , n366210 , n366211 , n366212 , n366213 , n366214 , n366215 , n366216 , n366217 , n366218 , 
 n366219 , n366220 , n366221 , n366222 , n366223 , n366224 , n366225 , n366226 , n366227 , n366228 , 
 n366229 , n366230 , n366231 , n366232 , n366233 , n366234 , n366235 , n366236 , n366237 , n366238 , 
 n366239 , n366240 , n366241 , n366242 , n366243 , n366244 , n366245 , n366246 , n366247 , n366248 , 
 n366249 , n366250 , n366251 , n366252 , n366253 , n366254 , n366255 , n366256 , n366257 , n366258 , 
 n366259 , n366260 , n366261 , n366262 , n366263 , n366264 , n366265 , n366266 , n366267 , n366268 , 
 n366269 , n366270 , n366271 , n366272 , n366273 , n366274 , n366275 , n366276 , n366277 , n366278 , 
 n366279 , n366280 , n366281 , n366282 , n366283 , n366284 , n366285 , n366286 , n366287 , n366288 , 
 n366289 , n366290 , n366291 , n366292 , n366293 , n366294 , n366295 , n366296 , n366297 , n366298 , 
 n366299 , n366300 , n366301 , n366302 , n366303 , n366304 , n366305 , n366306 , n366307 , n366308 , 
 n366309 , n18533 , n366311 , n366312 , n366313 , n366314 , n18538 , n366316 , n366317 , n18541 , 
 n18542 , n366320 , n366321 , n18545 , n366323 , n366324 , n366325 , n18549 , n366327 , n366328 , 
 n366329 , n18553 , n18554 , n366332 , n366333 , n366334 , n366335 , n366336 , n366337 , n366338 , 
 n18562 , n366340 , n366341 , n18565 , n18566 , n366344 , n366345 , n18569 , n18570 , n366348 , 
 n366349 , n366350 , n366351 , n366352 , n366353 , n18577 , n18578 , n366356 , n366357 , n366358 , 
 n18582 , n366360 , n366361 , n366362 , n18586 , n366364 , n366365 , n18589 , n366367 , n366368 , 
 n366369 , n18593 , n366371 , n366372 , n366373 , n366374 , n366375 , n366376 , n366377 , n18601 , 
 n18602 , n366380 , n366381 , n18605 , n366383 , n366384 , n366385 , n366386 , n366387 , n366388 , 
 n366389 , n366390 , n18614 , n366392 , n366393 , n18617 , n18618 , n366396 , n366397 , n366398 , 
 n18622 , n366400 , n366401 , n366402 , n366403 , n366404 , n366405 , n366406 , n366407 , n366408 , 
 n366409 , n18633 , n366411 , n366412 , n366413 , n18637 , n18638 , n366416 , n366417 , n366418 , 
 n366419 , n366420 , n366421 , n366422 , n18646 , n366424 , n366425 , n18649 , n18650 , n366428 , 
 n366429 , n18653 , n366431 , n366432 , n366433 , n18657 , n18658 , n366436 , n18660 , n366438 , 
 n18662 , n366440 , n366441 , n18665 , n18666 , n366444 , n366445 , n18669 , n366447 , n366448 , 
 n18672 , n366450 , n366451 , n366452 , n18676 , n366454 , n366455 , n18679 , n366457 , n366458 , 
 n18682 , n18683 , n366461 , n366462 , n18686 , n366464 , n18688 , n366466 , n366467 , n18691 , 
 n366469 , n366470 , n366471 , n18695 , n366473 , n366474 , n366475 , n18699 , n366477 , n18701 , 
 n18702 , n366480 , n18704 , n366482 , n18706 , n18707 , n366485 , n366486 , n18710 , n366488 , 
 n366489 , n18713 , n366491 , n366492 , n366493 , n18717 , n366495 , n366496 , n18720 , n366498 , 
 n366499 , n18723 , n366501 , n18725 , n366503 , n18727 , n18728 , n366506 , n18730 , n366508 , 
 n18732 , n18733 , n366511 , n366512 , n18736 , n366514 , n366515 , n18739 , n366517 , n366518 , 
 n366519 , n18743 , n366521 , n366522 , n18746 , n366524 , n366525 , n18749 , n18750 , n18751 , 
 n366529 , n366530 , n18754 , n18755 , n366533 , n366534 , n18758 , n366536 , n18760 , n366538 , 
 n18762 , n18763 , n18764 , n18765 , n18766 , n366544 , n366545 , n18769 , n366547 , n18771 , 
 n18772 , n366550 , n18774 , n366552 , n366553 , n18777 , n18778 , n18779 , n366557 , n366558 , 
 n366559 , n18783 , n366561 , n18785 , n18786 , n366564 , n18788 , n366566 , n18790 , n18791 , 
 n366569 , n366570 , n18794 , n366572 , n366573 , n18797 , n366575 , n366576 , n366577 , n18801 , 
 n366579 , n366580 , n18804 , n366582 , n366583 , n18807 , n18808 , n18809 , n366587 , n366588 , 
 n18812 , n18813 , n18814 , n366592 , n366593 , n18817 , n18818 , n18819 , n366597 , n366598 , 
 n18822 , n18823 , n18824 , n366602 , n366603 , n18827 , n18828 , n18829 , n366607 , n366608 , 
 n18832 , n18833 , n18834 , n366612 , n366613 , n18837 , n18838 , n18839 , n366617 , n18841 , 
 n18842 , n18843 , n366621 , n366622 , n18846 , n18847 , n366625 , n366626 , n366627 , n18851 , 
 n18852 , n18853 , n18854 , n18855 , n18856 , n366634 , n18858 , n18859 , n366637 , n366638 , 
 n18862 , n366640 , n366641 , n18865 , n366643 , n366644 , n18868 , n18869 , n366647 , n366648 , 
 n18872 , n366650 , n18874 , n366652 , n18876 , n366654 , n366655 , n18879 , n366657 , n18881 , 
 n18882 , n18883 , n18884 , n366662 , n18886 , n18887 , n366665 , n366666 , n18890 , n366668 , 
 n366669 , n18893 , n366671 , n366672 , n18896 , n18897 , n366675 , n366676 , n18900 , n366678 , 
 n18902 , n366680 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n366687 , n366688 , 
 n18912 , n366690 , n366691 , n18915 , n366693 , n366694 , n366695 , n18919 , n366697 , n18921 , 
 n18922 , n366700 , n18924 , n366702 , n18926 , n18927 , n366705 , n366706 , n18930 , n366708 , 
 n366709 , n18933 , n366711 , n366712 , n366713 , n18937 , n366715 , n366716 , n18940 , n366718 , 
 n366719 , n18943 , n366721 , n18945 , n366723 , n18947 , n18948 , n366726 , n18950 , n366728 , 
 n18952 , n18953 , n366731 , n366732 , n18956 , n366734 , n366735 , n18959 , n366737 , n366738 , 
 n366739 , n18963 , n366741 , n366742 , n18966 , n366744 , n366745 , n18969 , n18970 , n18971 , 
 n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n366755 , n366756 , n366757 , n18981 , 
 n366759 , n366760 , n366761 , n18985 , n366763 , n18987 , n18988 , n366766 , n18990 , n366768 , 
 n18992 , n18993 , n366771 , n366772 , n18996 , n366774 , n366775 , n18999 , n366777 , n366778 , 
 n366779 , n19003 , n366781 , n366782 , n19006 , n366784 , n366785 , n19009 , n366787 , n19011 , 
 n366789 , n19013 , n19014 , n366792 , n19016 , n366794 , n19018 , n19019 , n366797 , n366798 , 
 n19022 , n366800 , n366801 , n19025 , n366803 , n366804 , n366805 , n19029 , n366807 , n366808 , 
 n19032 , n366810 , n366811 , n19035 , n19036 , n19037 , n366815 , n366816 , n19040 , n19041 , 
 n19042 , n366820 , n366821 , n19045 , n19046 , n19047 , n366825 , n366826 , n19050 , n19051 , 
 n19052 , n366830 , n366831 , n19055 , n19056 , n19057 , n366835 , n366836 , n19060 , n19061 , 
 n19062 , n366840 , n366841 , n19065 , n19066 , n19067 , n366845 , n366846 , n19070 , n19071 , 
 n19072 , n366850 , n366851 , n19075 , n19076 , n19077 , n366855 , n366856 , n19080 , n19081 , 
 n19082 , n366860 , n366861 , n19085 , n366863 , n19087 , n366865 , n19089 , n19090 , n19091 , 
 n366869 , n19093 , n19094 , n366872 , n366873 , n19097 , n19098 , n366876 , n366877 , n366878 , 
 n19102 , n366880 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n366888 , 
 n366889 , n19113 , n366891 , n366892 , n19116 , n366894 , n366895 , n19119 , n19120 , n19121 , 
 n366899 , n366900 , n366901 , n19125 , n366903 , n19127 , n19128 , n19129 , n366907 , n366908 , 
 n19132 , n366910 , n366911 , n19135 , n366913 , n366914 , n19138 , n366916 , n19140 , n366918 , 
 n19142 , n19143 , n366921 , n19145 , n19146 , n366924 , n19148 , n19149 , n366927 , n366928 , 
 n19152 , n366930 , n366931 , n19155 , n366933 , n366934 , n366935 , n19159 , n366937 , n366938 , 
 n19162 , n366940 , n366941 , n366942 , n19166 , n366944 , n19168 , n366946 , n366947 , n19171 , 
 n366949 , n366950 , n19174 , n366952 , n366953 , n366954 , n19178 , n366956 , n19180 , n19181 , 
 n19182 , n366960 , n366961 , n366962 , n19186 , n366964 , n366965 , n19189 , n366967 , n366968 , 
 n19192 , n366970 , n19194 , n366972 , n19196 , n19197 , n366975 , n19199 , n366977 , n19201 , 
 n19202 , n366980 , n19204 , n366982 , n366983 , n366984 , n19208 , n366986 , n19210 , n19211 , 
 n19212 , n366990 , n19214 , n366992 , n366993 , n19217 , n19218 , n19219 , n366997 , n366998 , 
 n366999 , n19223 , n367001 , n19225 , n19226 , n367004 , n19228 , n367006 , n19230 , n19231 , 
 n367009 , n367010 , n19234 , n367012 , n367013 , n19237 , n367015 , n367016 , n367017 , n19241 , 
 n367019 , n367020 , n19244 , n367022 , n367023 , n19247 , n19248 , n19249 , n367027 , n367028 , 
 n19252 , n19253 , n19254 , n367032 , n367033 , n367034 , n19258 , n367036 , n19260 , n19261 , 
 n367039 , n19263 , n367041 , n19265 , n19266 , n367044 , n367045 , n19269 , n367047 , n367048 , 
 n19272 , n367050 , n367051 , n367052 , n19276 , n367054 , n367055 , n19279 , n367057 , n367058 , 
 n19282 , n19283 , n19284 , n367062 , n367063 , n19287 , n19288 , n19289 , n367067 , n367068 , 
 n19292 , n367070 , n19294 , n367072 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , 
 n19302 , n367080 , n19304 , n367082 , n367083 , n19307 , n19308 , n19309 , n367087 , n367088 , 
 n19312 , n19313 , n19314 , n367092 , n367093 , n19317 , n19318 , n19319 , n367097 , n367098 , 
 n19322 , n19323 , n19324 , n367102 , n367103 , n19327 , n19328 , n19329 , n367107 , n19331 , 
 n367109 , n19333 , n367111 , n19335 , n19336 , n367114 , n19338 , n367116 , n367117 , n19341 , 
 n19342 , n19343 , n367121 , n19345 , n367123 , n19347 , n19348 , n367126 , n19350 , n367128 , 
 n367129 , n19353 , n367131 , n367132 , n19356 , n19357 , n367135 , n367136 , n19360 , n19361 , 
 n19362 , n367140 , n367141 , n367142 , n19366 , n367144 , n19368 , n19369 , n19370 , n19371 , 
 n19372 , n19373 , n367151 , n367152 , n19376 , n367154 , n367155 , n19379 , n367157 , n367158 , 
 n19382 , n367160 , n19384 , n19385 , n19386 , n19387 , n19388 , n367166 , n19390 , n19391 , 
 n367169 , n367170 , n19394 , n367172 , n367173 , n19397 , n367175 , n367176 , n19400 , n19401 , 
 n19402 , n367180 , n367181 , n19405 , n19406 , n19407 , n367185 , n367186 , n19410 , n19411 , 
 n367189 , n367190 , n19414 , n19415 , n19416 , n367194 , n367195 , n19419 , n367197 , n19421 , 
 n19422 , n367200 , n367201 , n19425 , n19426 , n367204 , n367205 , n19429 , n367207 , n19431 , 
 n367209 , n19433 , n19434 , n367212 , n19436 , n367214 , n19438 , n19439 , n367217 , n367218 , 
 n19442 , n367220 , n367221 , n19445 , n367223 , n367224 , n367225 , n19449 , n367227 , n367228 , 
 n19452 , n367230 , n367231 , n367232 , n367233 , n367234 , n19461 , n367236 , n19463 , n19464 , 
 n19465 , n367240 , n367241 , n367242 , n19469 , n367244 , n367245 , n19472 , n367247 , n367248 , 
 n19475 , n367250 , n367251 , n367252 , n367253 , n367254 , n19487 , n367256 , n19493 , n367258 , 
 n367259 , n19499 , n367261 , n19501 , n19502 , n19503 , n367265 , n19505 , n367267 , n19511 , 
 n367269 , n367270 , n19520 , n367272 , n367273 , n367274 , n19524 , n367276 , n19526 , n367278 , 
 n19528 , n367280 , n367281 , n367282 , n367283 , n19533 , n367285 , n19535 , n367287 , n367288 , 
 n19538 , n367290 , n367291 , n19541 , n19542 , n19543 , n367295 , n367296 , n19546 , n367298 , 
 n367299 , n367300 , n19550 , n367302 , n19552 , n367304 , n19554 , n367306 , n367307 , n19557 , 
 n19558 , n367310 , n367311 , n19561 , n367313 , n19563 , n367315 , n19565 , n19566 , n367318 , 
 n367319 , n19569 , n367321 , n367322 , n19572 , n367324 , n367325 , n19575 , n19577 , n367328 , 
 n367329 , n19580 , n19582 , n367332 , n367333 , n19585 , n19586 , n367336 , n367337 , n19589 , 
 n367339 , n19591 , n367341 , n19593 , n19594 , n19595 , n19596 , n19597 , n367347 , n367348 , 
 n19600 , n367350 , n19602 , n19603 , n367353 , n19605 , n367355 , n367356 , n19608 , n19609 , 
 n19610 , n367360 , n367361 , n367362 , n19614 , n367364 , n19616 , n19617 , n367367 , n19619 , 
 n367369 , n19621 , n19622 , n367372 , n367373 , n19625 , n367375 , n367376 , n19628 , n367378 , 
 n367379 , n367380 , n19632 , n367382 , n367383 , n19635 , n367385 , n367386 , n19638 , n19639 , 
 n19640 , n367390 , n367391 , n19643 , n19644 , n19645 , n367395 , n367396 , n19648 , n19649 , 
 n19650 , n367400 , n367401 , n19653 , n19654 , n19655 , n367405 , n367406 , n19658 , n19659 , 
 n367409 , n367410 , n19662 , n367412 , n19664 , n367414 , n19666 , n19667 , n367417 , n19669 , 
 n367419 , n19671 , n19672 , n367422 , n367423 , n19675 , n367425 , n367426 , n19678 , n367428 , 
 n367429 , n367430 , n19682 , n367432 , n367433 , n19685 , n367435 , n367436 , n367437 , n19689 , 
 n19690 , n367440 , n19692 , n19693 , n367443 , n367444 , n19696 , n367446 , n367447 , n19699 , 
 n367449 , n367450 , n19702 , n367452 , n19704 , n367454 , n19706 , n19707 , n367457 , n19709 , 
 n367459 , n19711 , n19712 , n367462 , n19714 , n367464 , n19716 , n367466 , n367467 , n19719 , 
 n367469 , n367470 , n367471 , n19723 , n367473 , n367474 , n19726 , n367476 , n367477 , n367478 , 
 n19730 , n19731 , n367481 , n19733 , n19734 , n367484 , n19736 , n367486 , n19738 , n19739 , 
 n367489 , n367490 , n19742 , n367492 , n367493 , n19745 , n367495 , n367496 , n19748 , n367498 , 
 n367499 , n367500 , n19752 , n367502 , n367503 , n19755 , n367505 , n367506 , n19758 , n19759 , 
 n367509 , n367510 , n19762 , n19763 , n19764 , n19765 , n367515 , n19767 , n367517 , n19769 , 
 n19770 , n367520 , n367521 , n19773 , n367523 , n367524 , n19776 , n367526 , n367527 , n367528 , 
 n19780 , n367530 , n19782 , n367532 , n19784 , n19785 , n19786 , n367536 , n367537 , n367538 , 
 n19790 , n367540 , n19792 , n19793 , n367543 , n19795 , n367545 , n19797 , n19798 , n367548 , 
 n367549 , n19801 , n367551 , n367552 , n19804 , n367554 , n367555 , n367556 , n19808 , n367558 , 
 n367559 , n19811 , n367561 , n367562 , n19814 , n19815 , n19816 , n367566 , n367567 , n19819 , 
 n19820 , n19821 , n367571 , n367572 , n19824 , n19825 , n19826 , n367576 , n367577 , n19829 , 
 n19830 , n19831 , n367581 , n367582 , n19834 , n19835 , n19836 , n367586 , n367587 , n19839 , 
 n19840 , n19841 , n367591 , n367592 , n19844 , n19845 , n19846 , n367596 , n19848 , n19849 , 
 n19850 , n367600 , n19852 , n19853 , n19854 , n19855 , n367605 , n19857 , n19858 , n19859 , 
 n19860 , n19861 , n367611 , n367612 , n19864 , n367614 , n367615 , n19867 , n19868 , n367618 , 
 n367619 , n367620 , n19872 , n367622 , n19874 , n19875 , n367625 , n19877 , n367627 , n19879 , 
 n19880 , n367630 , n19882 , n367632 , n19884 , n367634 , n367635 , n19887 , n367637 , n367638 , 
 n19890 , n367640 , n367641 , n367642 , n19894 , n367644 , n367645 , n19897 , n367647 , n367648 , 
 n367649 , n19901 , n367651 , n19903 , n19904 , n367654 , n19906 , n367656 , n19908 , n19909 , 
 n367659 , n367660 , n19912 , n367662 , n367663 , n19915 , n367665 , n367666 , n367667 , n19919 , 
 n367669 , n367670 , n19922 , n367672 , n367673 , n367674 , n19926 , n367676 , n19928 , n19929 , 
 n367679 , n19931 , n367681 , n19933 , n19934 , n367684 , n367685 , n19937 , n367687 , n367688 , 
 n19940 , n367690 , n367691 , n367692 , n19944 , n367694 , n367695 , n19947 , n367697 , n367698 , 
 n367699 , n19951 , n367701 , n19953 , n19954 , n367704 , n19956 , n367706 , n19958 , n367708 , 
 n367709 , n19961 , n19962 , n367712 , n19964 , n367714 , n367715 , n19967 , n367717 , n367718 , 
 n367719 , n19971 , n367721 , n367722 , n19974 , n367724 , n367725 , n367726 , n19978 , n367728 , 
 n367729 , n19981 , n367731 , n367732 , n367733 , n367734 , n19988 , n367736 , n19990 , n367738 , 
 n19992 , n19993 , n367741 , n19995 , n367743 , n19997 , n19998 , n367746 , n367747 , n20001 , 
 n367749 , n367750 , n20004 , n367752 , n367753 , n367754 , n20008 , n367756 , n367757 , n20011 , 
 n367759 , n367760 , n20014 , n20016 , n367763 , n367764 , n367765 , n20020 , n367767 , n20022 , 
 n20023 , n367770 , n20025 , n367772 , n20027 , n20028 , n367775 , n367776 , n20031 , n367778 , 
 n367779 , n20034 , n367781 , n367782 , n367783 , n20038 , n367785 , n367786 , n20041 , n367788 , 
 n367789 , n20044 , n20045 , n20046 , n367793 , n367794 , n20049 , n20050 , n20051 , n367798 , 
 n367799 , n20054 , n20055 , n20056 , n367803 , n367804 , n20059 , n20060 , n20061 , n367808 , 
 n367809 , n20064 , n20065 , n20066 , n20067 , n367814 , n20069 , n367816 , n20071 , n20072 , 
 n367819 , n367820 , n20075 , n367822 , n367823 , n20078 , n367825 , n20080 , n20081 , n367828 , 
 n20083 , n20084 , n20085 , n367832 , n367833 , n20088 , n20089 , n20090 , n367837 , n367838 , 
 n20093 , n20094 , n20095 , n367842 , n367843 , n20098 , n20099 , n20100 , n367847 , n367848 , 
 n20103 , n20104 , n20105 , n367852 , n367853 , n20108 , n367855 , n367856 , n20111 , n367858 , 
 n20113 , n20114 , n20115 , n367862 , n367863 , n20118 , n20119 , n367866 , n367867 , n367868 , 
 n20123 , n367870 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n367877 , n367878 , 
 n20133 , n367880 , n367881 , n20136 , n367883 , n367884 , n20139 , n20140 , n367887 , n367888 , 
 n20143 , n367890 , n367891 , n367892 , n20149 , n367894 , n20151 , n20152 , n20153 , n367898 , 
 n20155 , n367900 , n20157 , n20158 , n367903 , n367904 , n20161 , n367906 , n20163 , n367908 , 
 n367909 , n20166 , n367911 , n367912 , n20169 , n367914 , n367915 , n20172 , n367917 , n367918 , 
 n20176 , n20177 , n20178 , n367922 , n20180 , n20183 , n367925 , n367926 , n20189 , n367928 , 
 n20191 , n20192 , n367931 , n20194 , n367933 , n367934 , n367935 , n20198 , n367937 , n20200 , 
 n20201 , n367940 , n20203 , n20206 , n367943 , n367944 , n20212 , n367946 , n367947 , n367948 , 
 n20216 , n367950 , n367951 , n20219 , n367953 , n367954 , n20222 , n367956 , n367957 , n367958 , 
 n367959 , n20227 , n367961 , n20229 , n367963 , n367964 , n20232 , n367966 , n367967 , n367968 , 
 n20236 , n367970 , n20238 , n20239 , n367973 , n367974 , n20242 , n20243 , n367977 , n367978 , 
 n367979 , n20247 , n367981 , n367982 , n20250 , n367984 , n367985 , n20253 , n367987 , n367988 , 
 n20256 , n20257 , n367991 , n367992 , n20260 , n20262 , n367995 , n367996 , n20265 , n20267 , 
 n367999 , n368000 , n20270 , n20271 , n368003 , n368004 , n20274 , n368006 , n20276 , n368008 , 
 n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n368015 , n368016 , n20286 , n368018 , 
 n368019 , n20289 , n368021 , n368022 , n20292 , n20293 , n20294 , n368026 , n368027 , n368028 , 
 n20298 , n368030 , n20300 , n20301 , n368033 , n20303 , n368035 , n20305 , n20306 , n368038 , 
 n368039 , n20309 , n368041 , n368042 , n20312 , n368044 , n368045 , n368046 , n20316 , n368048 , 
 n368049 , n20319 , n368051 , n368052 , n20322 , n20323 , n20324 , n368056 , n368057 , n20327 , 
 n20328 , n20329 , n368061 , n368062 , n368063 , n20333 , n368065 , n20335 , n20336 , n20337 , 
 n20338 , n20339 , n20340 , n368072 , n368073 , n20343 , n368075 , n368076 , n20346 , n368078 , 
 n368079 , n20349 , n368081 , n20351 , n368083 , n20353 , n20354 , n368086 , n368087 , n20357 , 
 n368089 , n368090 , n20360 , n368092 , n20362 , n368094 , n20364 , n368096 , n368097 , n20367 , 
 n20368 , n368100 , n20370 , n368102 , n368103 , n20373 , n368105 , n368106 , n20376 , n20377 , 
 n20378 , n368110 , n368111 , n20381 , n20382 , n20383 , n368115 , n368116 , n20386 , n20387 , 
 n20388 , n368120 , n368121 , n20391 , n20392 , n20393 , n368125 , n368126 , n20396 , n368128 , 
 n368129 , n20399 , n20400 , n368132 , n20402 , n20403 , n368135 , n368136 , n20406 , n20407 , 
 n368139 , n368140 , n368141 , n20411 , n20412 , n368144 , n20414 , n20415 , n368147 , n368148 , 
 n20418 , n368150 , n368151 , n20421 , n368153 , n368154 , n20424 , n368156 , n20426 , n368158 , 
 n20428 , n20429 , n368161 , n20431 , n368163 , n20433 , n20434 , n368166 , n368167 , n20437 , 
 n368169 , n368170 , n20440 , n368172 , n368173 , n368174 , n20444 , n368176 , n368177 , n20447 , 
 n368179 , n368180 , n368181 , n20451 , n368183 , n20453 , n20454 , n368186 , n20456 , n368188 , 
 n20458 , n20459 , n368191 , n368192 , n20462 , n368194 , n368195 , n20465 , n368197 , n368198 , 
 n368199 , n20469 , n368201 , n368202 , n20472 , n368204 , n368205 , n20475 , n20476 , n368208 , 
 n368209 , n20479 , n368211 , n20481 , n368213 , n20483 , n20484 , n368216 , n20486 , n368218 , 
 n20488 , n368220 , n368221 , n20491 , n20492 , n20493 , n368225 , n20495 , n368227 , n368228 , 
 n368229 , n20499 , n368231 , n368232 , n20502 , n368234 , n368235 , n20505 , n20506 , n20507 , 
 n368239 , n368240 , n368241 , n20511 , n368243 , n20513 , n20514 , n20515 , n20516 , n20517 , 
 n20518 , n368250 , n368251 , n20521 , n368253 , n368254 , n20524 , n368256 , n368257 , n20527 , 
 n20528 , n20529 , n368261 , n368262 , n20532 , n20533 , n20534 , n368266 , n368267 , n20537 , 
 n20538 , n20539 , n368271 , n368272 , n20542 , n20543 , n20544 , n368276 , n368277 , n20547 , 
 n20548 , n20549 , n368281 , n368282 , n20552 , n20553 , n20554 , n368286 , n368287 , n20557 , 
 n20558 , n20559 , n368291 , n20561 , n368293 , n20563 , n368295 , n20565 , n20566 , n20567 , 
 n368299 , n368300 , n20570 , n368302 , n368303 , n20573 , n368305 , n20575 , n368307 , n368308 , 
 n20578 , n368310 , n368311 , n20581 , n368313 , n368314 , n368315 , n20585 , n368317 , n368318 , 
 n20588 , n368320 , n368321 , n20591 , n368323 , n368324 , n20594 , n20595 , n20596 , n20597 , 
 n368329 , n368330 , n20600 , n368332 , n368333 , n20603 , n368335 , n368336 , n368337 , n20607 , 
 n368339 , n20609 , n20610 , n368342 , n20612 , n368344 , n20614 , n20615 , n368347 , n368348 , 
 n20618 , n368350 , n368351 , n20621 , n368353 , n368354 , n368355 , n20625 , n368357 , n368358 , 
 n20628 , n368360 , n368361 , n368362 , n20632 , n368364 , n20634 , n20635 , n368367 , n20637 , 
 n368369 , n20639 , n20640 , n368372 , n368373 , n20643 , n368375 , n368376 , n20646 , n368378 , 
 n368379 , n368380 , n20650 , n368382 , n368383 , n20653 , n368385 , n368386 , n20656 , n20657 , 
 n368389 , n368390 , n20660 , n368392 , n20662 , n368394 , n20664 , n20665 , n368397 , n20667 , 
 n368399 , n20669 , n368401 , n368402 , n20672 , n20673 , n368405 , n368406 , n20676 , n368408 , 
 n368409 , n20679 , n368411 , n368412 , n368413 , n20683 , n368415 , n368416 , n20686 , n368418 , 
 n368419 , n20689 , n20690 , n20691 , n368423 , n368424 , n20694 , n20695 , n20696 , n20697 , 
 n20698 , n368430 , n368431 , n20701 , n368433 , n20703 , n368435 , n20705 , n20706 , n20707 , 
 n368439 , n368440 , n20710 , n20711 , n20712 , n368444 , n368445 , n20715 , n20716 , n20717 , 
 n368449 , n368450 , n20720 , n20721 , n20722 , n368454 , n368455 , n20725 , n368457 , n20727 , 
 n20728 , n20729 , n20730 , n20731 , n368463 , n20733 , n20734 , n368466 , n368467 , n20737 , 
 n368469 , n368470 , n20740 , n368472 , n368473 , n20743 , n20744 , n20745 , n368477 , n368478 , 
 n20748 , n20749 , n368481 , n368482 , n20752 , n20753 , n20754 , n368486 , n368487 , n20757 , 
 n20758 , n20759 , n368491 , n368492 , n20762 , n368494 , n368495 , n20765 , n368497 , n20767 , 
 n20768 , n368500 , n368501 , n368502 , n368503 , n368504 , n20776 , n368506 , n20778 , n20779 , 
 n20780 , n20781 , n20782 , n20783 , n368513 , n368514 , n20786 , n368516 , n368517 , n20789 , 
 n368519 , n368520 , n20792 , n368522 , n368523 , n368524 , n20797 , n368526 , n20799 , n20800 , 
 n368529 , n20802 , n20805 , n368532 , n368533 , n20811 , n368535 , n368536 , n368537 , n20815 , 
 n368539 , n368540 , n20818 , n368542 , n368543 , n20821 , n368545 , n368546 , n368547 , n20825 , 
 n368549 , n20827 , n20828 , n368552 , n20830 , n20833 , n368555 , n368556 , n20839 , n368558 , 
 n368559 , n368560 , n20843 , n368562 , n368563 , n20846 , n368565 , n368566 , n20849 , n368568 , 
 n20851 , n368570 , n20853 , n20854 , n368573 , n368574 , n20857 , n20858 , n368577 , n368578 , 
 n368579 , n20862 , n368581 , n368582 , n20865 , n368584 , n368585 , n20868 , n368587 , n368588 , 
 n368589 , n368590 , n20873 , n368592 , n368593 , n368594 , n20877 , n368596 , n368597 , n20880 , 
 n368599 , n368600 , n20883 , n20884 , n368603 , n368604 , n20887 , n20889 , n368607 , n368608 , 
 n20892 , n20894 , n368611 , n368612 , n20897 , n20898 , n368615 , n368616 , n20901 , n368618 , 
 n20903 , n368620 , n20905 , n20906 , n368623 , n20908 , n368625 , n20910 , n20911 , n368628 , 
 n368629 , n20914 , n368631 , n368632 , n20917 , n368634 , n368635 , n368636 , n20921 , n368638 , 
 n368639 , n20924 , n368641 , n368642 , n20927 , n20928 , n20929 , n368646 , n368647 , n20932 , 
 n20933 , n368650 , n368651 , n20936 , n368653 , n20938 , n368655 , n20940 , n20941 , n368658 , 
 n368659 , n20944 , n20945 , n368662 , n20947 , n20948 , n368665 , n368666 , n368667 , n20952 , 
 n368669 , n368670 , n20955 , n368672 , n368673 , n20958 , n20959 , n20960 , n368677 , n368678 , 
 n368679 , n20964 , n368681 , n20966 , n20967 , n20968 , n368685 , n368686 , n20971 , n368688 , 
 n368689 , n20974 , n368691 , n368692 , n20977 , n368694 , n20979 , n20980 , n20981 , n20982 , 
 n20983 , n368700 , n20985 , n20986 , n368703 , n368704 , n20989 , n368706 , n368707 , n20992 , 
 n368709 , n368710 , n20995 , n20996 , n20997 , n368714 , n368715 , n21000 , n21001 , n21002 , 
 n368719 , n368720 , n21005 , n368722 , n21007 , n21008 , n21009 , n368726 , n368727 , n368728 , 
 n21013 , n368730 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n368737 , n368738 , 
 n21023 , n368740 , n368741 , n21026 , n368743 , n368744 , n368745 , n21030 , n368747 , n21032 , 
 n21033 , n368750 , n21035 , n368752 , n21037 , n368754 , n368755 , n21040 , n21041 , n368758 , 
 n368759 , n21044 , n368761 , n368762 , n21047 , n368764 , n368765 , n368766 , n21051 , n368768 , 
 n368769 , n21054 , n368771 , n368772 , n21057 , n21058 , n368775 , n368776 , n21061 , n368778 , 
 n21063 , n368780 , n21065 , n21066 , n368783 , n21068 , n368785 , n21070 , n21071 , n368788 , 
 n368789 , n21074 , n368791 , n368792 , n21077 , n368794 , n368795 , n368796 , n21081 , n368798 , 
 n368799 , n21084 , n368801 , n368802 , n21087 , n21088 , n21089 , n368806 , n368807 , n368808 , 
 n21093 , n368810 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n368817 , n368818 , 
 n21103 , n368820 , n368821 , n21106 , n368823 , n368824 , n21109 , n21110 , n21111 , n368828 , 
 n368829 , n21114 , n21115 , n21116 , n368833 , n368834 , n21119 , n21120 , n21121 , n368838 , 
 n368839 , n21124 , n21125 , n21126 , n368843 , n368844 , n21129 , n21130 , n21131 , n368848 , 
 n368849 , n21134 , n21135 , n21136 , n368853 , n21138 , n21139 , n21140 , n21141 , n368858 , 
 n368859 , n21144 , n21145 , n21146 , n21147 , n368864 , n368865 , n21150 , n368867 , n21152 , 
 n21153 , n21154 , n368871 , n368872 , n21157 , n368874 , n21159 , n368876 , n21161 , n21162 , 
 n21163 , n21164 , n21165 , n21166 , n368883 , n368884 , n21169 , n368886 , n368887 , n21172 , 
 n368889 , n368890 , n368891 , n21176 , n368893 , n21178 , n21179 , n21180 , n21181 , n21182 , 
 n21183 , n368900 , n368901 , n21186 , n368903 , n368904 , n21189 , n368906 , n368907 , n368908 , 
 n21193 , n368910 , n21195 , n21196 , n368913 , n21198 , n368915 , n21200 , n21201 , n368918 , 
 n368919 , n21204 , n368921 , n368922 , n21207 , n368924 , n368925 , n368926 , n21211 , n368928 , 
 n368929 , n21214 , n368931 , n368932 , n21217 , n21218 , n368935 , n368936 , n21221 , n368938 , 
 n368939 , n368940 , n21227 , n368942 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , 
 n368949 , n368950 , n21237 , n368952 , n368953 , n21240 , n368955 , n368956 , n21243 , n368958 , 
 n368959 , n368960 , n21256 , n368962 , n21258 , n21259 , n368965 , n21261 , n21264 , n368968 , 
 n368969 , n21270 , n368971 , n368972 , n368973 , n21274 , n368975 , n368976 , n21277 , n368978 , 
 n368979 , n21280 , n368981 , n368982 , n368983 , n21284 , n368985 , n21286 , n21287 , n368988 , 
 n21289 , n21295 , n368991 , n368992 , n21301 , n368994 , n368995 , n368996 , n21305 , n368998 , 
 n368999 , n21308 , n369001 , n369002 , n21311 , n369004 , n21313 , n369006 , n21315 , n21316 , 
 n369009 , n369010 , n21319 , n21320 , n369013 , n369014 , n369015 , n21324 , n369017 , n369018 , 
 n21327 , n369020 , n369021 , n21330 , n369023 , n369024 , n369025 , n369026 , n21335 , n369028 , 
 n21337 , n369030 , n369031 , n21340 , n369033 , n369034 , n21343 , n369036 , n369037 , n21346 , 
 n369039 , n369040 , n21349 , n21350 , n369043 , n369044 , n21353 , n21355 , n369047 , n369048 , 
 n21358 , n21360 , n369051 , n369052 , n21363 , n21365 , n369055 , n369056 , n369057 , n21369 , 
 n369059 , n21371 , n21372 , n369062 , n21374 , n369064 , n21376 , n21377 , n369067 , n369068 , 
 n21380 , n369070 , n369071 , n21383 , n369073 , n369074 , n369075 , n21387 , n369077 , n369078 , 
 n21390 , n369080 , n369081 , n21393 , n21394 , n21395 , n369085 , n369086 , n21398 , n21399 , 
 n21400 , n369090 , n369091 , n21403 , n21404 , n21405 , n369095 , n369096 , n21408 , n21409 , 
 n21410 , n369100 , n369101 , n21413 , n21414 , n21415 , n369105 , n369106 , n21418 , n21419 , 
 n21420 , n369110 , n369111 , n21423 , n369113 , n369114 , n21426 , n369116 , n369117 , n21429 , 
 n369119 , n21431 , n21432 , n21433 , n21434 , n21435 , n369125 , n21437 , n21438 , n21439 , 
 n21440 , n21441 , n21442 , n369132 , n369133 , n21445 , n369135 , n369136 , n21448 , n369138 , 
 n369139 , n369140 , n21452 , n21453 , n21454 , n21455 , n21456 , n369146 , n21458 , n21459 , 
 n369149 , n21461 , n369151 , n21463 , n21464 , n369154 , n369155 , n21467 , n369157 , n369158 , 
 n21470 , n369160 , n369161 , n369162 , n21474 , n369164 , n369165 , n21477 , n369167 , n369168 , 
 n21480 , n21481 , n369171 , n369172 , n21484 , n369174 , n21486 , n369176 , n21488 , n369178 , 
 n21490 , n21491 , n369181 , n369182 , n21494 , n369184 , n369185 , n21497 , n369187 , n369188 , 
 n21500 , n21501 , n369191 , n21503 , n369193 , n21505 , n21506 , n369196 , n21508 , n369198 , 
 n369199 , n369200 , n21512 , n369202 , n369203 , n21515 , n369205 , n369206 , n369207 , n21519 , 
 n369209 , n369210 , n21522 , n369212 , n369213 , n21525 , n21526 , n21527 , n369217 , n369218 , 
 n369219 , n21531 , n369221 , n21533 , n369223 , n21535 , n21536 , n369226 , n21538 , n369228 , 
 n21540 , n369230 , n369231 , n21543 , n369233 , n369234 , n21546 , n21547 , n21548 , n21549 , 
 n21550 , n21551 , n21552 , n21553 , n21554 , n369244 , n21556 , n369246 , n369247 , n21559 , 
 n369249 , n21561 , n369251 , n21563 , n21564 , n369254 , n369255 , n21567 , n369257 , n369258 , 
 n21570 , n369260 , n369261 , n21573 , n21574 , n369264 , n369265 , n21577 , n369267 , n21579 , 
 n369269 , n21581 , n21582 , n369272 , n369273 , n21585 , n369275 , n369276 , n21588 , n369278 , 
 n369279 , n21591 , n369281 , n369282 , n21594 , n21595 , n21596 , n369286 , n369287 , n21599 , 
 n21600 , n21601 , n21602 , n21603 , n369293 , n369294 , n21606 , n21607 , n369297 , n369298 , 
 n21610 , n369300 , n21612 , n369302 , n21614 , n21615 , n369305 , n369306 , n21618 , n369308 , 
 n369309 , n21621 , n369311 , n369312 , n21624 , n369314 , n369315 , n21627 , n21628 , n21629 , 
 n369319 , n21631 , n21632 , n21633 , n21634 , n21635 , n369325 , n369326 , n369327 , n21639 , 
 n369329 , n21641 , n21642 , n369332 , n369333 , n21645 , n369335 , n369336 , n21648 , n369338 , 
 n369339 , n21651 , n21652 , n21653 , n369343 , n369344 , n21656 , n369346 , n21658 , n21659 , 
 n21660 , n21661 , n369351 , n369352 , n369353 , n21665 , n369355 , n21667 , n21668 , n369358 , 
 n21670 , n369360 , n21672 , n21673 , n369363 , n369364 , n21676 , n369366 , n369367 , n21679 , 
 n369369 , n369370 , n21682 , n369372 , n369373 , n369374 , n21686 , n369376 , n369377 , n21689 , 
 n369379 , n369380 , n369381 , n21693 , n369383 , n21695 , n21696 , n369386 , n21698 , n369388 , 
 n21700 , n21701 , n369391 , n369392 , n21704 , n369394 , n369395 , n21707 , n369397 , n369398 , 
 n369399 , n21711 , n369401 , n369402 , n21714 , n369404 , n369405 , n369406 , n369407 , n21721 , 
 n369409 , n21723 , n369411 , n21725 , n21726 , n369414 , n21728 , n369416 , n21730 , n21731 , 
 n369419 , n369420 , n21734 , n369422 , n369423 , n21737 , n369425 , n369426 , n369427 , n21741 , 
 n369429 , n369430 , n21744 , n369432 , n369433 , n21747 , n21749 , n369436 , n369437 , n21752 , 
 n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n369447 , n21762 , 
 n21763 , n21764 , n369451 , n369452 , n21767 , n21768 , n21769 , n369456 , n369457 , n21772 , 
 n21773 , n21774 , n369461 , n369462 , n21777 , n21778 , n21779 , n369466 , n369467 , n21782 , 
 n369469 , n21784 , n21785 , n21786 , n369473 , n369474 , n21789 , n369476 , n369477 , n369478 , 
 n21795 , n369480 , n21797 , n21798 , n369483 , n21800 , n369485 , n21802 , n21803 , n369488 , 
 n369489 , n21806 , n369491 , n369492 , n21809 , n369494 , n369495 , n369496 , n21813 , n369498 , 
 n369499 , n21816 , n369501 , n369502 , n21819 , n369504 , n369505 , n369506 , n369507 , n369508 , 
 n21832 , n21835 , n369511 , n369512 , n21841 , n369514 , n21843 , n21844 , n21845 , n369518 , 
 n369519 , n21848 , n21852 , n369522 , n369523 , n21855 , n369525 , n21857 , n369527 , n21859 , 
 n369529 , n21861 , n369531 , n369532 , n369533 , n369534 , n21866 , n369536 , n21868 , n369538 , 
 n369539 , n21871 , n369541 , n369542 , n369543 , n369544 , n21876 , n369546 , n369547 , n369548 , 
 n21880 , n369550 , n369551 , n369552 , n21884 , n369554 , n369555 , n21887 , n21888 , n369558 , 
 n369559 , n21891 , n369561 , n369562 , n21894 , n369564 , n369565 , n21897 , n21898 , n369568 , 
 n369569 , n21901 , n369571 , n21903 , n369573 , n21905 , n21906 , n369576 , n369577 , n21909 , 
 n369579 , n369580 , n21912 , n369582 , n369583 , n21915 , n21917 , n369586 , n369587 , n21920 , 
 n21922 , n369590 , n369591 , n21925 , n21926 , n369594 , n369595 , n21929 , n369597 , n21931 , 
 n369599 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n369606 , n369607 , n21941 , 
 n369609 , n369610 , n21944 , n369612 , n369613 , n21947 , n21948 , n21949 , n369617 , n369618 , 
 n21952 , n21953 , n369621 , n369622 , n21956 , n369624 , n21958 , n369626 , n21960 , n21961 , 
 n369629 , n21963 , n369631 , n21965 , n21966 , n369634 , n21968 , n369636 , n21970 , n369638 , 
 n369639 , n21973 , n369641 , n369642 , n369643 , n21977 , n369645 , n369646 , n21980 , n369648 , 
 n369649 , n21983 , n21984 , n21985 , n369653 , n369654 , n21988 , n369656 , n369657 , n21991 , 
 n369659 , n21993 , n369661 , n369662 , n369663 , n21999 , n369665 , n22001 , n369667 , n22003 , 
 n22004 , n369670 , n369671 , n22007 , n369673 , n369674 , n22010 , n369676 , n369677 , n22013 , 
 n22014 , n369680 , n22016 , n369682 , n22018 , n22019 , n369685 , n369686 , n22022 , n369688 , 
 n369689 , n22025 , n369691 , n369692 , n369693 , n22029 , n369695 , n369696 , n22032 , n369698 , 
 n369699 , n22035 , n369701 , n369702 , n369703 , n369704 , n22043 , n22044 , n22045 , n369708 , 
 n22048 , n22051 , n369711 , n369712 , n22057 , n369714 , n22059 , n22060 , n369717 , n22062 , 
 n369719 , n369720 , n369721 , n369722 , n22067 , n369724 , n22069 , n369726 , n369727 , n22072 , 
 n369729 , n369730 , n22075 , n369732 , n369733 , n22078 , n369735 , n369736 , n22081 , n22082 , 
 n369739 , n369740 , n369741 , n22086 , n369743 , n369744 , n22089 , n369746 , n369747 , n22092 , 
 n369749 , n369750 , n22095 , n369752 , n369753 , n22098 , n22099 , n369756 , n369757 , n22102 , 
 n369759 , n22104 , n369761 , n22106 , n22107 , n22108 , n22111 , n22112 , n369767 , n22114 , 
 n369769 , n369770 , n22117 , n22119 , n369773 , n369774 , n22122 , n22124 , n369777 , n369778 , 
 n369779 , n22128 , n369781 , n22130 , n369783 , n22132 , n22133 , n369786 , n369787 , n22136 , 
 n369789 , n369790 , n22139 , n369792 , n369793 , n22142 , n22143 , n369796 , n369797 , n22146 , 
 n369799 , n369800 , n22149 , n369802 , n369803 , n369804 , n369805 , n22156 , n369807 , n22158 , 
 n22159 , n369810 , n22161 , n22162 , n369813 , n22164 , n369815 , n22166 , n22167 , n369818 , 
 n22169 , n369820 , n22171 , n369822 , n369823 , n22174 , n369825 , n369826 , n369827 , n22178 , 
 n369829 , n369830 , n22181 , n369832 , n369833 , n22184 , n369835 , n369836 , n22187 , n369838 , 
 n22189 , n22190 , n22191 , n22192 , n22193 , n369844 , n22195 , n22196 , n369847 , n22198 , 
 n369849 , n22200 , n22201 , n369852 , n22203 , n369854 , n22205 , n369856 , n369857 , n22208 , 
 n369859 , n369860 , n369861 , n22212 , n369863 , n369864 , n22215 , n369866 , n369867 , n22218 , 
 n369869 , n22220 , n369871 , n22222 , n369873 , n22224 , n22225 , n22226 , n22227 , n22228 , 
 n22229 , n369880 , n369881 , n22232 , n369883 , n369884 , n22235 , n369886 , n369887 , n22238 , 
 n22239 , n369890 , n369891 , n22242 , n369893 , n22244 , n369895 , n22246 , n22247 , n22248 , 
 n22249 , n22250 , n22251 , n369902 , n369903 , n22254 , n369905 , n369906 , n22257 , n369908 , 
 n369909 , n22260 , n22261 , n22262 , n369913 , n22264 , n22265 , n369916 , n22267 , n369918 , 
 n369919 , n22271 , n369921 , n22275 , n369923 , n22277 , n22278 , n369926 , n369927 , n22281 , 
 n22282 , n22283 , n22286 , n369932 , n369933 , n22289 , n369935 , n369936 , n22292 , n369938 , 
 n369939 , n369940 , n369941 , n22298 , n369943 , n22300 , n369945 , n22302 , n22303 , n369948 , 
 n22305 , n22306 , n22309 , n22310 , n22311 , n22312 , n369955 , n22314 , n369957 , n369958 , 
 n369959 , n369960 , n22319 , n369962 , n369963 , n369964 , n22323 , n369966 , n369967 , n22326 , 
 n369969 , n369970 , n22329 , n369972 , n22331 , n369974 , n22333 , n22334 , n369977 , n369978 , 
 n22337 , n369980 , n369981 , n22340 , n369983 , n369984 , n22343 , n22344 , n369987 , n369988 , 
 n369989 , n369990 , n22351 , n369992 , n22353 , n369994 , n22355 , n22356 , n369997 , n22358 , 
 n369999 , n22360 , n370001 , n370002 , n22363 , n370004 , n370005 , n22366 , n22367 , n370008 , 
 n370009 , n22370 , n370011 , n22372 , n370013 , n370014 , n22375 , n22376 , n370017 , n22378 , 
 n370019 , n22380 , n370021 , n370022 , n22383 , n370024 , n370025 , n22386 , n370027 , n370028 , 
 n22389 , n370030 , n370031 , n370032 , n370033 , n22396 , n370035 , n22398 , n370037 , n370038 , 
 n22401 , n370040 , n22403 , n370042 , n22405 , n370044 , n22407 , n22408 , n22412 , n370048 , 
 n370049 , n22415 , n370051 , n370052 , n22418 , n370054 , n370055 , n370056 , n370057 , n22434 , 
 n370059 , n370060 , n22437 , n370062 , n22439 , n370064 , n370065 , n22442 , n370067 , n370068 , 
 n22445 , n370070 , n22447 , n370072 , n22449 , n22450 , n370075 , n370076 , n22453 , n370078 , 
 n370079 , n22456 , n370081 , n22458 , n370083 , n22460 , n370085 , n370086 , n22463 , n370088 , 
 n370089 , n22466 , n370091 , n22468 , n370093 , n370094 , n22471 , n22472 , n22473 , n22474 , 
 n22475 , n22476 , n370101 , n22478 , n22479 , n370104 , n22481 , n22493 , n22494 , n22495 , 
 n22497 , n22498 , n370111 , n22500 , n370113 , n22502 , n22503 , n22504 , n370117 , n370118 , 
 n370119 , n22510 , n370121 , n370122 , n22513 , n22514 , n370125 , n22516 , n22517 , n370128 , 
 n370129 , n22520 , n22521 , n370132 , n370133 , n22524 , n370135 , n370136 , n22527 , n370138 , 
 n370139 , n22530 , n22531 , n22532 , n22534 , n370144 , n370145 , n22537 , n370147 , n370148 , 
 n22540 , n22541 , n370151 , n22543 , n22544 , n370154 , n370155 , n22547 , n370157 , n370158 , 
 n22550 , n370160 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n370167 , n22559 , 
 n370169 , n370170 , n370171 , n22563 , n370173 , n22565 , n22566 , n370176 , n370177 , n22569 , 
 n370179 , n370180 , n22572 , n370182 , n370183 , n370184 , n370185 , n22579 , n370187 , n22581 , 
 n370189 , n22583 , n22584 , n370192 , n370193 , n22587 , n370195 , n370196 , n22590 , n370198 , 
 n370199 , n22593 , n370201 , n370202 , n22596 , n370204 , n370205 , n22599 , n22600 , n22602 , 
 n370209 , n370210 , n22605 , n370212 , n370213 , n22608 , n370215 , n370216 , n22611 , n370218 , 
 n370219 , n22614 , n370221 , n370222 , n22617 , n22618 , n22619 , n370226 , n22621 , n22622 , 
 n22623 , n22625 , n370231 , n370232 , n22628 , n370234 , n22630 , n370236 , n22632 , n22633 , 
 n370239 , n370240 , n22636 , n370242 , n370243 , n22639 , n370245 , n370246 , n22642 , n22643 , 
 n370249 , n370250 , n22646 , n370252 , n370253 , n22649 , n370255 , n370256 , n22652 , n22653 , 
 n22654 , n22656 , n370261 , n370262 , n370263 , n22660 , n22661 , n22662 , n22663 , n22664 , 
 n370269 , n22666 , n22667 , n370272 , n370273 , n22670 , n370275 , n370276 , n22673 , n370278 , 
 n370279 , n22676 , n370281 , n22678 , n370283 , n22680 , n22681 , n370286 , n370287 , n22684 , 
 n370289 , n370290 , n22687 , n370292 , n370293 , n22690 , n22691 , n370296 , n370297 , n22694 , 
 n370299 , n22696 , n370301 , n22698 , n22699 , n370304 , n370305 , n22702 , n370307 , n370308 , 
 n22705 , n370310 , n370311 , n22708 , n370313 , n370314 , n22711 , n370316 , n22713 , n22714 , 
 n22715 , n22716 , n370321 , n22718 , n370323 , n22720 , n22721 , n370326 , n370327 , n22724 , 
 n370329 , n370330 , n22727 , n370332 , n22729 , n370334 , n22731 , n370336 , n22733 , n22734 , 
 n370339 , n370340 , n22737 , n370342 , n370343 , n22740 , n370345 , n370346 , n22743 , n22744 , 
 n22745 , n22746 , n370351 , n370352 , n22749 , n22750 , n22751 , n370356 , n370357 , n22754 , 
 n370359 , n370360 , n22757 , n22758 , n22759 , n22760 , n370365 , n370366 , n22763 , n370368 , 
 n22765 , n22766 , n370371 , n370372 , n22769 , n370374 , n22771 , n370376 , n22773 , n22774 , 
 n22775 , n370380 , n22777 , n370382 , n22779 , n22780 , n22781 , n22782 , n370387 , n370388 , 
 n22785 , n370390 , n370391 , n22788 , n370393 , n370394 , n22791 , n22792 , n370397 , n370398 , 
 n22795 , n370400 , n370401 , n22798 , n370403 , n22800 , n22801 , n370406 , n22803 , n370408 , 
 n370409 , n370410 , n22807 , n370412 , n22809 , n22810 , n22811 , n370416 , n22813 , n370418 , 
 n22815 , n370420 , n370421 , n22818 , n370423 , n22820 , n370425 , n22822 , n370427 , n370428 , 
 n370429 , n22826 , n370431 , n370432 , n22829 , n370434 , n22831 , n22832 , n370437 , n370438 , 
 n22835 , n370440 , n22837 , n22838 , n370443 , n22840 , n22841 , n370446 , n370447 , n22844 , 
 n22845 , n22846 , n22847 , n370452 , n370453 , n22850 , n370455 , n370456 , n22853 , n370458 , 
 n370459 , n22856 , n22857 , n370462 , n370463 , n370464 , n22861 , n370466 , n370467 , n22864 , 
 n370469 , n370470 , n22867 , n370472 , n370473 , n22870 , n370475 , n370476 , n22873 , n370478 , 
 n370479 , n22876 , n370481 , n370482 , n22879 , n370484 , n22881 , n370486 , n22883 , n370488 , 
 n22885 , n370490 , n22887 , n370492 , n370493 , n22890 , n370495 , n370496 , n370497 , n370498 , 
 n22895 , n370500 , n370501 , n22898 , n370503 , n22900 , n370505 , n22902 , n370507 , n22904 , 
 n22905 , n22906 , n22907 , n370512 , n22909 , n370514 , n370515 , n370516 , n22913 , n370518 , 
 n370519 , n22916 , n370521 , n370522 , n370523 , n22920 , n370525 , n22922 , n370527 , n370528 , 
 n22925 , n370530 , n370531 , n22928 , n370533 , n370534 , n22931 , n370536 , n370537 , n22934 , 
 n370539 , n22936 , n22937 , n22938 , n370543 , n370544 , n22941 , n370546 , n22943 , n22944 , 
 n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , 
 n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n370565 , n22962 , n22963 , n22964 , 
 n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n370575 , n22972 , n370577 , n370578 , 
 n22975 , n370580 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n370587 , n22984 , 
 n22985 , n370590 , n22987 , n22988 , n22989 , n22990 , n370595 , n370596 , n370597 , n370598 , 
 n22995 , n22996 , n370601 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , 
 n370609 , n370610 , n23007 , n370612 , n370613 , n23010 , n370615 , n370616 , n370617 , n23014 , 
 n370619 , n23016 , n370621 , n370622 , n370623 , n23020 , n370625 , n370626 , n23023 , n370628 , 
 n23025 , n370630 , n23027 , n370632 , n23029 , n370634 , n23031 , n370636 , n370637 , n23034 , 
 n370639 , n370640 , n23037 , n370642 , n23039 , n23040 , n370645 , n370646 , n23043 , n370648 , 
 n370649 , n23046 , n370651 , n370652 , n370653 , n23050 , n370655 , n23052 , n370657 , n23054 , 
 n23055 , n370660 , n370661 , n370662 , n23059 , n370664 , n23061 , n23062 , n23063 , n23064 , 
 n23065 , n23066 , n370671 , n370672 , n23069 , n370674 , n370675 , n23072 , n370677 , n370678 , 
 n23075 , n370680 , n23077 , n370682 , n370683 , n23080 , n370685 , n370686 , n23083 , n23084 , 
 n370689 , n370690 , n23087 , n370692 , n370693 , n23090 , n370695 , n370696 , n23093 , n23094 , 
 n23095 , n370700 , n370701 , n23098 , n370703 , n370704 , n23101 , n23102 , n370707 , n370708 , 
 n370709 , n23106 , n370711 , n23108 , n370713 , n23110 , n23111 , n370716 , n23113 , n23114 , 
 n370719 , n370720 , n23117 , n23118 , n370723 , n370724 , n23121 , n370726 , n370727 , n23124 , 
 n370729 , n370730 , n23127 , n370732 , n23129 , n370734 , n370735 , n23132 , n23133 , n370738 , 
 n23135 , n23136 , n370741 , n370742 , n23139 , n23140 , n370745 , n370746 , n23143 , n370748 , 
 n370749 , n23146 , n370751 , n370752 , n23149 , n23150 , n23151 , n370756 , n370757 , n23154 , 
 n23155 , n370760 , n370761 , n370762 , n23159 , n370764 , n23161 , n23162 , n23163 , n23164 , 
 n370769 , n370770 , n23167 , n370772 , n23169 , n23170 , n23171 , n370776 , n23173 , n370778 , 
 n370779 , n23176 , n23177 , n23178 , n23179 , n23180 , n370785 , n370786 , n23183 , n370788 , 
 n23185 , n23186 , n23187 , n370792 , n370793 , n23190 , n370795 , n23192 , n370797 , n23194 , 
 n370799 , n370800 , n370801 , n23198 , n370803 , n370804 , n23201 , n370806 , n370807 , n23204 , 
 n370809 , n370810 , n370811 , n23208 , n370813 , n23210 , n23211 , n370816 , n23213 , n370818 , 
 n370819 , n23216 , n370821 , n370822 , n370823 , n23220 , n23221 , n370826 , n370827 , n23224 , 
 n370829 , n23226 , n370831 , n370832 , n23229 , n23230 , n23231 , n23232 , n23233 , n370838 , 
 n23235 , n23236 , n370841 , n23238 , n23239 , n370844 , n370845 , n23242 , n370847 , n370848 , 
 n23245 , n370850 , n23247 , n23248 , n370853 , n23250 , n370855 , n370856 , n23253 , n370858 , 
 n370859 , n23256 , n23257 , n23258 , n23259 , n370864 , n370865 , n23262 , n23263 , n23264 , 
 n23265 , n23266 , n23267 , n23268 , n23269 , n370874 , n23271 , n23272 , n23273 , n23274 , 
 n370879 , n370880 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , 
 n23285 , n370890 , n370891 , n23288 , n370893 , n23290 , n23291 , n370896 , n370897 , n23294 , 
 n370899 , n370900 , n23297 , n370902 , n370903 , n23300 , n23301 , n23302 , n23303 , n23304 , 
 n370909 , n370910 , n23307 , n370912 , n370913 , n23310 , n370915 , n370916 , n23313 , n23314 , 
 n23315 , n23316 , n23317 , n370922 , n370923 , n23320 , n23321 , n23322 , n370927 , n370928 , 
 n23325 , n23326 , n23327 , n23328 , n23329 , n370934 , n370935 , n370936 , n23333 , n370938 , 
 n370939 , n23336 , n23337 , n370942 , n23339 , n370944 , n370945 , n23342 , n23343 , n370948 , 
 n370949 , n23346 , n23347 , n370952 , n23349 , n370954 , n23351 , n370956 , n370957 , n23354 , 
 n23355 , n370960 , n23357 , n370962 , n23359 , n370964 , n370965 , n23362 , n370967 , n370968 , 
 n370969 , n23366 , n370971 , n370972 , n23369 , n370974 , n370975 , n23372 , n23373 , n23374 , 
 n23375 , n370980 , n370981 , n23378 , n370983 , n23380 , n23381 , n23382 , n23383 , n23384 , 
 n23385 , n23386 , n23387 , n23388 , n370993 , n23390 , n23391 , n23392 , n23393 , n370998 , 
 n23395 , n371000 , n23397 , n23398 , n23399 , n371004 , n23401 , n371006 , n23403 , n23404 , 
 n23405 , n23406 , n371011 , n371012 , n23409 , n371014 , n23411 , n371016 , n23413 , n371018 , 
 n371019 , n23416 , n371021 , n23418 , n371023 , n23420 , n23421 , n371026 , n371027 , n23424 , 
 n371029 , n371030 , n23427 , n371032 , n371033 , n23430 , n23431 , n23432 , n23433 , n371038 , 
 n371039 , n23436 , n23437 , n23438 , n371043 , n371044 , n23441 , n23442 , n23443 , n371048 , 
 n371049 , n23446 , n371051 , n371052 , n23449 , n371054 , n371055 , n23452 , n23453 , n371058 , 
 n371059 , n23456 , n23457 , n23458 , n23459 , n371064 , n371065 , n23462 , n23463 , n23464 , 
 n371069 , n371070 , n23467 , n23468 , n23469 , n371074 , n371075 , n23472 , n371077 , n371078 , 
 n371079 , n23476 , n371081 , n23478 , n371083 , n23480 , n23481 , n23482 , n371087 , n23484 , 
 n23485 , n23486 , n23487 , n23488 , n371093 , n23490 , n23491 , n371096 , n371097 , n23494 , 
 n371099 , n23496 , n23497 , n371102 , n23499 , n23500 , n23501 , n23502 , n23503 , n371108 , 
 n371109 , n23506 , n371111 , n371112 , n371113 , n23510 , n371115 , n23512 , n371117 , n371118 , 
 n23515 , n371120 , n23517 , n23518 , n371123 , n23520 , n371125 , n371126 , n23523 , n371128 , 
 n371129 , n23526 , n371131 , n23528 , n371133 , n23530 , n23531 , n371136 , n23533 , n23534 , 
 n23535 , n23536 , n371141 , n371142 , n371143 , n23540 , n23541 , n371146 , n23543 , n371148 , 
 n23545 , n371150 , n23547 , n23548 , n23549 , n23550 , n23551 , n371156 , n23553 , n23554 , 
 n371159 , n23556 , n23557 , n23558 , n23559 , n371164 , n371165 , n371166 , n371167 , n23564 , 
 n371169 , n23566 , n371171 , n371172 , n23569 , n371174 , n23571 , n23572 , n371177 , n23574 , 
 n371179 , n371180 , n23577 , n23578 , n371183 , n371184 , n23581 , n23582 , n371187 , n23584 , 
 n23585 , n23586 , n23587 , n371192 , n371193 , n371194 , n23591 , n23592 , n23593 , n371198 , 
 n23595 , n371200 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , 
 n371209 , n23606 , n23607 , n371212 , n23609 , n23610 , n23611 , n23612 , n371217 , n371218 , 
 n371219 , n371220 , n23617 , n371222 , n23619 , n371224 , n23621 , n371226 , n371227 , n371228 , 
 n23625 , n371230 , n371231 , n23628 , n23629 , n371234 , n23631 , n371236 , n23633 , n371238 , 
 n371239 , n23636 , n371241 , n371242 , n23639 , n371244 , n371245 , n23642 , n23643 , n371248 , 
 n23645 , n23646 , n23647 , n23648 , n371253 , n23650 , n371255 , n371256 , n371257 , n23654 , 
 n371259 , n371260 , n23657 , n371262 , n371263 , n23660 , n23661 , n371266 , n23663 , n371268 , 
 n371269 , n371270 , n23667 , n371272 , n371273 , n23670 , n371275 , n371276 , n23673 , n371278 , 
 n371279 , n23676 , n23677 , n371282 , n23679 , n23680 , n23681 , n23682 , n371287 , n371288 , 
 n371289 , n23686 , n371291 , n371292 , n23689 , n371294 , n23691 , n23692 , n371297 , n23694 , 
 n371299 , n23696 , n371301 , n371302 , n23699 , n371304 , n23701 , n371306 , n23703 , n23704 , 
 n371309 , n23706 , n23707 , n23708 , n23709 , n371314 , n371315 , n371316 , n371317 , n371318 , 
 n23715 , n371320 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , 
 n23725 , n371330 , n23727 , n23728 , n371333 , n23730 , n23731 , n23732 , n23733 , n371338 , 
 n371339 , n371340 , n371341 , n23738 , n371343 , n371344 , n371345 , n371346 , n23743 , n371348 , 
 n23745 , n371350 , n23747 , n23748 , n371353 , n23750 , n23751 , n371356 , n371357 , n23754 , 
 n23755 , n371360 , n23757 , n23758 , n23759 , n23760 , n371365 , n371366 , n371367 , n371368 , 
 n371369 , n23766 , n371371 , n371372 , n371373 , n23770 , n371375 , n23772 , n23773 , n23774 , 
 n23775 , n371380 , n23777 , n23778 , n371383 , n23780 , n23781 , n23782 , n23783 , n371388 , 
 n371389 , n371390 , n23787 , n23788 , n23789 , n371394 , n23791 , n371396 , n23793 , n23794 , 
 n371399 , n371400 , n371401 , n23798 , n371403 , n371404 , n23801 , n371406 , n371407 , n23804 , 
 n371409 , n23806 , n23807 , n371412 , n371413 , n23810 , n371415 , n23812 , n23813 , n371418 , 
 n23815 , n371420 , n371421 , n23818 , n23819 , n371424 , n23821 , n23822 , n23823 , n23824 , 
 n371429 , n371430 , n371431 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , 
 n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n371446 , n23843 , n23844 , 
 n371449 , n23846 , n23847 , n23848 , n23849 , n371454 , n371455 , n371456 , n371457 , n23854 , 
 n371459 , n371460 , n371461 , n23858 , n371463 , n371464 , n371465 , n371466 , n23863 , n371468 , 
 n371469 , n23866 , n371471 , n23868 , n371473 , n23870 , n23871 , n371476 , n23873 , n23874 , 
 n23875 , n23876 , n371481 , n371482 , n371483 , n371484 , n371485 , n23882 , n371487 , n23884 , 
 n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n371496 , n23893 , n371498 , 
 n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n371505 , n23902 , n23903 , n371508 , 
 n23905 , n23906 , n23907 , n23908 , n371513 , n371514 , n371515 , n23912 , n371517 , n23914 , 
 n23915 , n371520 , n23917 , n371522 , n371523 , n23920 , n23921 , n371526 , n23923 , n23924 , 
 n23925 , n23926 , n371531 , n371532 , n371533 , n371534 , n23931 , n371536 , n371537 , n23934 , 
 n371539 , n371540 , n23937 , n371542 , n23939 , n23940 , n23941 , n371546 , n23943 , n23944 , 
 n23945 , n23946 , n23947 , n23948 , n23949 , n371554 , n23951 , n23952 , n371557 , n23954 , 
 n371559 , n23956 , n23957 , n23958 , n23959 , n23960 , n371565 , n23962 , n23963 , n371568 , 
 n23965 , n23966 , n23967 , n23968 , n371573 , n371574 , n371575 , n23972 , n371577 , n23974 , 
 n371579 , n23976 , n23977 , n371582 , n23979 , n371584 , n23981 , n23982 , n23983 , n23984 , 
 n23985 , n23986 , n23987 , n23988 , n371593 , n23990 , n23991 , n371596 , n23993 , n23994 , 
 n23995 , n23996 , n371601 , n371602 , n371603 , n371604 , n371605 , n24002 , n371607 , n371608 , 
 n24005 , n24006 , n24007 , n24008 , n371613 , n371614 , n371615 , n24012 , n371617 , n24014 , 
 n24015 , n371620 , n371621 , n24018 , n371623 , n24020 , n24021 , n24022 , n24023 , n24024 , 
 n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n371636 , n371637 , n24034 , 
 n371639 , n371640 , n24037 , n371642 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , 
 n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n371658 , 
 n24055 , n371660 , n24057 , n24058 , n371663 , n24060 , n371665 , n371666 , n24063 , n24064 , 
 n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , 
 n371679 , n24076 , n24077 , n24078 , n371683 , n371684 , n371685 , n24082 , n371687 , n24084 , 
 n24085 , n371690 , n371691 , n24088 , n371693 , n371694 , n24091 , n371696 , n371697 , n24094 , 
 n371699 , n371700 , n24097 , n371702 , n371703 , n24100 , n371705 , n371706 , n24103 , n371708 , 
 n371709 , n24106 , n371711 , n371712 , n371713 , n371714 , n24111 , n371716 , n371717 , n24114 , 
 n371719 , n24116 , n24117 , n24118 , n371723 , n24120 , n24121 , n24122 , n371727 , n371728 , 
 n371729 , n24126 , n371731 , n371732 , n24129 , n371734 , n24131 , n371736 , n371737 , n371738 , 
 n371739 , n24136 , n371741 , n371742 , n24139 , n371744 , n371745 , n24142 , n24143 , n371748 , 
 n24145 , n24146 , n371751 , n371752 , n24149 , n24150 , n24151 , n371756 , n371757 , n24154 , 
 n24155 , n371760 , n371761 , n24158 , n24159 , n24160 , n371765 , n24162 , n24163 , n24164 , 
 n371769 , n24166 , n371771 , n24168 , n371773 , n371774 , n371775 , n371776 , n24173 , n371778 , 
 n371779 , n24176 , n371781 , n371782 , n24179 , n371784 , n371785 , n24182 , n371787 , n24184 , 
 n24185 , n24186 , n24187 , n371792 , n24189 , n24190 , n371795 , n24192 , n371797 , n371798 , 
 n24195 , n371800 , n24197 , n24198 , n24199 , n24200 , n371805 , n24202 , n371807 , n24204 , 
 n371809 , n371810 , n24207 , n371812 , n371813 , n24210 , n371815 , n24212 , n24213 , n24214 , 
 n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , 
 n24225 , n24226 , n24227 , n24228 , n24229 , n371834 , n24231 , n371836 , n371837 , n24234 , 
 n371839 , n371840 , n24237 , n24238 , n24239 , n371844 , n371845 , n24242 , n371847 , n371848 , 
 n24245 , n371850 , n371851 , n371852 , n24249 , n371854 , n24251 , n371856 , n371857 , n371858 , 
 n24255 , n371860 , n24257 , n24258 , n24259 , n371864 , n24261 , n371866 , n371867 , n24264 , 
 n371869 , n24266 , n24267 , n24268 , n24269 , n371874 , n24271 , n371876 , n371877 , n24274 , 
 n371879 , n371880 , n24277 , n24278 , n24279 , n371884 , n371885 , n24282 , n371887 , n371888 , 
 n24285 , n24286 , n24287 , n371892 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , 
 n24295 , n24296 , n24297 , n371902 , n371903 , n24300 , n371905 , n371906 , n371907 , n371908 , 
 n371909 , n24306 , n371911 , n371912 , n24309 , n371914 , n371915 , n371916 , n24313 , n371918 , 
 n371919 , n24316 , n24317 , n371922 , n24319 , n24320 , n371925 , n371926 , n24323 , n24324 , 
 n24325 , n371930 , n371931 , n24328 , n371933 , n24330 , n371935 , n24332 , n24333 , n371938 , 
 n371939 , n24336 , n24337 , n24338 , n371943 , n24340 , n371945 , n371946 , n371947 , n24344 , 
 n371949 , n371950 , n24347 , n371952 , n24349 , n371954 , n371955 , n24352 , n371957 , n371958 , 
 n371959 , n24356 , n24357 , n371962 , n24359 , n371964 , n371965 , n24362 , n371967 , n371968 , 
 n24365 , n371970 , n24367 , n371972 , n24369 , n24370 , n371975 , n24372 , n371977 , n371978 , 
 n24375 , n371980 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , 
 n371989 , n371990 , n371991 , n24388 , n371993 , n371994 , n24391 , n371996 , n371997 , n24394 , 
 n371999 , n372000 , n24397 , n372002 , n372003 , n24400 , n24401 , n24402 , n372007 , n24404 , 
 n24405 , n24406 , n24407 , n24408 , n372013 , n24410 , n372015 , n372016 , n24413 , n372018 , 
 n372019 , n24416 , n372021 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , 
 n372029 , n24426 , n24427 , n372032 , n372033 , n24430 , n372035 , n372036 , n24433 , n372038 , 
 n372039 , n24436 , n24437 , n372042 , n372043 , n24440 , n372045 , n372046 , n24443 , n372048 , 
 n372049 , n24446 , n24447 , n372052 , n372053 , n24450 , n372055 , n372056 , n24453 , n372058 , 
 n372059 , n24456 , n24457 , n372062 , n372063 , n24460 , n372065 , n372066 , n24463 , n372068 , 
 n372069 , n24466 , n24467 , n372072 , n372073 , n24470 , n372075 , n372076 , n24473 , n372078 , 
 n372079 , n24476 , n24477 , n24478 , n372083 , n372084 , n24481 , n24482 , n24483 , n372088 , 
 n372089 , n24486 , n24487 , n24488 , n372093 , n372094 , n24491 , n24492 , n24493 , n372098 , 
 n372099 , n24496 , n24497 , n24498 , n372103 , n372104 , n24501 , n24502 , n24503 , n372108 , 
 n372109 , n24506 , n24507 , n24508 , n372113 , n372114 , n24511 , n24512 , n24513 , n372118 , 
 n372119 , n24516 , n24517 , n24518 , n372123 , n372124 , n24521 , n24522 , n24523 , n372128 , 
 n372129 , n24526 , n24527 , n24528 , n372133 , n372134 , n24531 , n24532 , n24533 , n372138 , 
 n372139 , n372140 , n24537 , n372142 , n372143 , n24540 , n24541 , n24542 , n24543 , n372148 , 
 n24545 , n372150 , n372151 , n24548 , n372153 , n372154 , n24551 , n372156 , n372157 , n24554 , 
 n372159 , n372160 , n24557 , n372162 , n372163 , n372164 , n24561 , n372166 , n24563 , n24564 , 
 n372169 , n24566 , n372171 , n372172 , n24569 , n372174 , n372175 , n372176 , n372177 , n24574 , 
 n372179 , n372180 , n24577 , n24578 , n24579 , n24580 , n372185 , n372186 , n372187 , n24584 , 
 n24585 , n372190 , n24587 , n24588 , n372193 , n372194 , n372195 , n372196 , n372197 , n24594 , 
 n24595 , n24596 , n24597 , n24598 , n372203 , n24600 , n24601 , n372206 , n24603 , n24604 , 
 n372209 , n24606 , n24607 , n372212 , n24609 , n24610 , n372215 , n24612 , n24613 , n372218 , 
 n24615 , n24616 , n372221 , n24618 , n24619 , n372224 , n24621 , n24622 , n372227 , n24624 , 
 n24625 , n372230 , n24627 , n24628 , n372233 , n24630 , n24631 , n372236 , n24633 , n24634 , 
 n372239 , n372240 , n372241 , n372242 , n24639 , n372244 , n372245 , n372246 , n372247 , n24644 , 
 n24645 , n24646 , n24647 , n24648 , n372253 , n372254 , n24651 , n24652 , n24653 , n24654 , 
 n372259 , n372260 , n372261 , n24658 , n24659 , n24660 , n24661 , n24662 , n372267 , n372268 , 
 n372269 , n372270 , n24667 , n372272 , n372273 , n372274 , n372275 , n24672 , n24673 , n24674 , 
 n24675 , n24676 , n372281 , n372282 , n372283 , n372284 , n24681 , n372286 , n372287 , n24684 , 
 n372289 , n372290 , n372291 , n372292 , n24689 , n372294 , n372295 , n24692 , n372297 , n372298 , 
 n372299 , n372300 , n372301 , n24698 , n372303 , n372304 , n24701 , n24702 , n24703 , n24704 , 
 n372309 , n372310 , n372311 , n372312 , n24709 , n372314 , n372315 , n24712 , n372317 , n24714 , 
 n24715 , n372320 , n372321 , n372322 , n24719 , n372324 , n372325 , n372326 , n24723 , n372328 , 
 n24725 , n24726 , n372331 , n372332 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , 
 n24735 , n24736 , n24737 , n372342 , n372343 , n372344 , n24741 , n24742 , n24743 , n24744 , 
 n24745 , n372350 , n24747 , n372352 , n372353 , n372354 , n24751 , n372356 , n372357 , n372358 , 
 n24755 , n372360 , n372361 , n372362 , n24759 , n372364 , n372365 , n372366 , n24763 , n372368 , 
 n372369 , n372370 , n24767 , n24768 , n372373 , n372374 , n24771 , n24772 , n372377 , n24774 , 
 n24775 , n24776 , n24777 , n372382 , n372383 , n372384 , n24781 , n24782 , n24783 , n24784 , 
 n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n372395 , n24792 , n24793 , n372398 , 
 n24795 , n24796 , n24797 , n24798 , n372403 , n372404 , n372405 , n372406 , n24803 , n372408 , 
 n24805 , n372410 , n372411 , n372412 , n24809 , n24810 , n24811 , n372416 , n24813 , n24814 , 
 n372419 , n372420 , n24817 , n24818 , n372423 , n24820 , n24821 , n24822 , n24823 , n372428 , 
 n372429 , n372430 , n24827 , n24828 , n372433 , n24830 , n24831 , n372436 , n24833 , n24834 , 
 n24835 , n24836 , n372441 , n372442 , n372443 , n24840 , n24841 , n372446 , n24843 , n24844 , 
 n372449 , n24846 , n24847 , n24848 , n24849 , n372454 , n372455 , n372456 , n372457 , n372458 , 
 n24855 , n372460 , n372461 , n24858 , n372463 , n24860 , n24861 , n24862 , n24863 , n24864 , 
 n372469 , n24866 , n372471 , n372472 , n24869 , n24870 , n372475 , n24872 , n24873 , n24874 , 
 n24875 , n372480 , n372481 , n372482 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , 
 n24885 , n24886 , n24887 , n372492 , n24889 , n24890 , n372495 , n24892 , n24893 , n24894 , 
 n24895 , n372500 , n372501 , n372502 , n372503 , n24900 , n372505 , n372506 , n24903 , n372508 , 
 n372509 , n24906 , n372511 , n24908 , n372513 , n372514 , n24911 , n24912 , n372517 , n24914 , 
 n372519 , n24916 , n372521 , n372522 , n24919 , n372524 , n372525 , n24922 , n372527 , n372528 , 
 n24925 , n24926 , n372531 , n24928 , n24929 , n24930 , n24931 , n372536 , n372537 , n372538 , 
 n372539 , n24936 , n372541 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n372548 , 
 n24945 , n372550 , n372551 , n24948 , n24949 , n372554 , n24951 , n372556 , n372557 , n24954 , 
 n372559 , n372560 , n372561 , n24958 , n372563 , n372564 , n24961 , n372566 , n372567 , n24964 , 
 n24965 , n372570 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , 
 n24975 , n372580 , n24977 , n372582 , n372583 , n24980 , n24981 , n372586 , n24983 , n372588 , 
 n372589 , n372590 , n24987 , n372592 , n372593 , n24990 , n372595 , n372596 , n372597 , n24994 , 
 n372599 , n372600 , n24997 , n372602 , n372603 , n372604 , n372605 , n25002 , n372607 , n372608 , 
 n372609 , n25006 , n372611 , n25008 , n372613 , n25010 , n25011 , n372616 , n372617 , n25014 , 
 n372619 , n372620 , n25017 , n372622 , n372623 , n25020 , n25021 , n372626 , n25023 , n372628 , 
 n25025 , n25026 , n372631 , n372632 , n25029 , n372634 , n372635 , n25032 , n372637 , n372638 , 
 n372639 , n25036 , n372641 , n372642 , n25039 , n372644 , n372645 , n25042 , n372647 , n25044 , 
 n372649 , n25046 , n372651 , n25048 , n25049 , n372654 , n372655 , n25052 , n372657 , n372658 , 
 n25055 , n372660 , n372661 , n25058 , n25059 , n372664 , n25061 , n372666 , n25063 , n25064 , 
 n25065 , n372670 , n372671 , n25068 , n372673 , n372674 , n25071 , n372676 , n372677 , n372678 , 
 n25075 , n372680 , n372681 , n25078 , n372683 , n372684 , n25081 , n25082 , n25083 , n372688 , 
 n372689 , n372690 , n25087 , n372692 , n25089 , n372694 , n372695 , n372696 , n25093 , n372698 , 
 n25095 , n372700 , n25097 , n25098 , n372703 , n372704 , n25101 , n372706 , n372707 , n25104 , 
 n372709 , n372710 , n25107 , n25108 , n372713 , n372714 , n25111 , n372716 , n372717 , n25114 , 
 n372719 , n372720 , n25117 , n372722 , n25119 , n25120 , n25121 , n25122 , n25123 , n372728 , 
 n25125 , n25126 , n372731 , n372732 , n25129 , n372734 , n372735 , n25132 , n372737 , n372738 , 
 n25135 , n372740 , n372741 , n25138 , n372743 , n25140 , n372745 , n25142 , n372747 , n25144 , 
 n25145 , n25146 , n372751 , n25148 , n372753 , n372754 , n25151 , n25152 , n372757 , n25154 , 
 n372759 , n25156 , n25157 , n372762 , n372763 , n25160 , n372765 , n372766 , n25163 , n372768 , 
 n372769 , n372770 , n25167 , n372772 , n372773 , n25170 , n372775 , n372776 , n25173 , n372778 , 
 n372779 , n25176 , n25177 , n25178 , n372783 , n372784 , n25181 , n25182 , n25183 , n25184 , 
 n25185 , n25186 , n25187 , n25188 , n372793 , n25190 , n25191 , n372796 , n25193 , n25194 , 
 n372799 , n372800 , n25197 , n372802 , n372803 , n25200 , n372805 , n372806 , n372807 , n25204 , 
 n372809 , n25206 , n372811 , n25208 , n25209 , n25210 , n25211 , n25212 , n372817 , n372818 , 
 n25215 , n25216 , n25217 , n372822 , n372823 , n25220 , n372825 , n25222 , n25223 , n372828 , 
 n372829 , n25226 , n372831 , n25228 , n25229 , n25230 , n372835 , n25232 , n372837 , n372838 , 
 n25235 , n372840 , n372841 , n372842 , n25239 , n372844 , n25241 , n372846 , n25243 , n25244 , 
 n372849 , n372850 , n25247 , n372852 , n372853 , n25250 , n372855 , n372856 , n25253 , n25254 , 
 n372859 , n372860 , n25257 , n372862 , n372863 , n25260 , n372865 , n372866 , n25263 , n372868 , 
 n372869 , n25266 , n372871 , n25268 , n372873 , n372874 , n25271 , n372876 , n372877 , n372878 , 
 n25275 , n372880 , n25277 , n25278 , n372883 , n25280 , n372885 , n372886 , n25283 , n372888 , 
 n372889 , n25286 , n25287 , n25288 , n372893 , n372894 , n25291 , n25292 , n25293 , n25294 , 
 n25295 , n372900 , n372901 , n25298 , n25299 , n25300 , n25301 , n372906 , n25303 , n372908 , 
 n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , n372918 , 
 n25315 , n25316 , n25317 , n25318 , n25319 , n372924 , n25321 , n372926 , n25323 , n25324 , 
 n372929 , n372930 , n25327 , n372932 , n372933 , n25330 , n372935 , n372936 , n372937 , n25334 , 
 n372939 , n25336 , n372941 , n25338 , n25339 , n25340 , n25341 , n372946 , n372947 , n25344 , 
 n372949 , n372950 , n25347 , n372952 , n372953 , n372954 , n25351 , n25352 , n25353 , n372958 , 
 n25355 , n25356 , n372961 , n372962 , n25359 , n372964 , n372965 , n25362 , n372967 , n372968 , 
 n25365 , n372970 , n25367 , n372972 , n25369 , n372974 , n25371 , n25372 , n372977 , n372978 , 
 n25375 , n372980 , n372981 , n25378 , n372983 , n372984 , n25381 , n25382 , n372987 , n372988 , 
 n25385 , n372990 , n372991 , n25388 , n25389 , n372994 , n372995 , n25392 , n372997 , n372998 , 
 n25395 , n373000 , n373001 , n25398 , n373003 , n373004 , n25401 , n373006 , n373007 , n25404 , 
 n25405 , n25406 , n373011 , n373012 , n373013 , n25410 , n25411 , n25412 , n25413 , n25414 , 
 n373019 , n25416 , n25417 , n373022 , n25419 , n25420 , n373025 , n25422 , n25423 , n373028 , 
 n373029 , n25426 , n373031 , n373032 , n25429 , n373034 , n373035 , n373036 , n25433 , n373038 , 
 n373039 , n25436 , n373041 , n373042 , n25439 , n373044 , n373045 , n373046 , n25443 , n373048 , 
 n25445 , n25446 , n373051 , n25448 , n373053 , n25450 , n25451 , n373056 , n373057 , n25454 , 
 n373059 , n373060 , n25457 , n373062 , n373063 , n373064 , n25461 , n373066 , n373067 , n25464 , 
 n373069 , n373070 , n25467 , n373072 , n25469 , n373074 , n25471 , n25472 , n373077 , n25474 , 
 n373079 , n25476 , n25477 , n373082 , n373083 , n25480 , n373085 , n373086 , n25483 , n373088 , 
 n373089 , n373090 , n25487 , n373092 , n373093 , n25490 , n373095 , n373096 , n25493 , n25494 , 
 n25495 , n373100 , n373101 , n25498 , n25499 , n373104 , n373105 , n25502 , n373107 , n25504 , 
 n373109 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n373116 , n373117 , n25514 , 
 n373119 , n373120 , n25517 , n373122 , n373123 , n25520 , n25521 , n25522 , n373127 , n373128 , 
 n373129 , n25526 , n373131 , n25528 , n25529 , n373134 , n25531 , n373136 , n25533 , n25534 , 
 n373139 , n373140 , n25537 , n373142 , n373143 , n25540 , n373145 , n373146 , n373147 , n25544 , 
 n373149 , n373150 , n25547 , n373152 , n373153 , n25550 , n25551 , n25552 , n373157 , n373158 , 
 n25555 , n25556 , n25557 , n373162 , n373163 , n25560 , n25561 , n25562 , n25563 , n25564 , 
 n25565 , n25566 , n373171 , n25568 , n373173 , n373174 , n25571 , n373176 , n373177 , n25574 , 
 n373179 , n373180 , n25577 , n25578 , n373183 , n373184 , n373185 , n25582 , n373187 , n373188 , 
 n25585 , n25586 , n373191 , n373192 , n373193 , n25590 , n373195 , n25592 , n25593 , n373198 , 
 n373199 , n25596 , n373201 , n373202 , n25599 , n373204 , n373205 , n373206 , n25603 , n373208 , 
 n373209 , n25606 , n373211 , n373212 , n25609 , n25610 , n25611 , n373216 , n373217 , n373218 , 
 n25615 , n373220 , n25617 , n373222 , n373223 , n373224 , n25621 , n373226 , n25623 , n25624 , 
 n25625 , n25626 , n25627 , n373232 , n25629 , n373234 , n373235 , n373236 , n25633 , n373238 , 
 n373239 , n373240 , n25637 , n373242 , n25639 , n373244 , n25641 , n25642 , n25643 , n373248 , 
 n373249 , n25646 , n373251 , n25648 , n25649 , n373254 , n373255 , n25652 , n373257 , n25654 , 
 n25655 , n25656 , n373261 , n25658 , n25659 , n25660 , n373265 , n25662 , n25663 , n25664 , 
 n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n373277 , n25674 , 
 n25675 , n25676 , n373281 , n25678 , n373283 , n373284 , n25681 , n373286 , n25683 , n373288 , 
 n373289 , n25686 , n373291 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , 
 n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , 
 n25705 , n25706 , n25707 , n25708 , n373313 , n25710 , n373315 , n373316 , n25713 , n373318 , 
 n25715 , n373320 , n25717 , n373322 , n25719 , n25720 , n25721 , n25722 , n373327 , n25724 , 
 n25725 , n373330 , n373331 , n25728 , n373333 , n373334 , n25731 , n373336 , n373337 , n373338 , 
 n25735 , n373340 , n25737 , n25738 , n373343 , n25740 , n25741 , n373346 , n25743 , n25744 , 
 n373349 , n373350 , n25747 , n373352 , n373353 , n25750 , n373355 , n373356 , n373357 , n25754 , 
 n373359 , n373360 , n25757 , n373362 , n373363 , n25760 , n25761 , n25762 , n373367 , n373368 , 
 n25765 , n25766 , n25767 , n373372 , n373373 , n25770 , n25771 , n25772 , n373377 , n373378 , 
 n25775 , n25776 , n25777 , n25778 , n25779 , n373384 , n373385 , n25782 , n25783 , n25784 , 
 n25785 , n25786 , n373391 , n373392 , n25789 , n373394 , n25791 , n25792 , n25793 , n373398 , 
 n25795 , n373400 , n25797 , n25798 , n373403 , n373404 , n25801 , n25802 , n373407 , n25804 , 
 n373409 , n25806 , n373411 , n25808 , n373413 , n25810 , n25811 , n373416 , n25813 , n25814 , 
 n373419 , n373420 , n25817 , n373422 , n373423 , n25820 , n373425 , n373426 , n25823 , n25824 , 
 n373429 , n25826 , n373431 , n25828 , n25829 , n373434 , n373435 , n25832 , n25833 , n373438 , 
 n373439 , n25836 , n373441 , n373442 , n25839 , n373444 , n373445 , n373446 , n25843 , n373448 , 
 n25845 , n373450 , n25847 , n25848 , n373453 , n373454 , n25851 , n373456 , n373457 , n25854 , 
 n373459 , n373460 , n25857 , n25858 , n373463 , n25860 , n373465 , n25862 , n25863 , n25864 , 
 n25865 , n25866 , n25867 , n25868 , n373473 , n25870 , n373475 , n373476 , n25873 , n25874 , 
 n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n373487 , n25884 , 
 n25885 , n373490 , n25887 , n373492 , n25889 , n373494 , n373495 , n25892 , n25893 , n373498 , 
 n373499 , n25896 , n373501 , n373502 , n25899 , n373504 , n25901 , n25902 , n25903 , n25904 , 
 n373509 , n25906 , n373511 , n373512 , n25909 , n25910 , n25911 , n25912 , n25913 , n373518 , 
 n373519 , n373520 , n373521 , n25918 , n373523 , n373524 , n373525 , n25922 , n373527 , n25924 , 
 n373529 , n25926 , n25927 , n373532 , n373533 , n25930 , n373535 , n373536 , n25933 , n373538 , 
 n373539 , n25936 , n25937 , n373542 , n373543 , n25940 , n373545 , n373546 , n25943 , n373548 , 
 n373549 , n25946 , n373551 , n25948 , n25949 , n25950 , n25951 , n25952 , n373557 , n25954 , 
 n25955 , n373560 , n373561 , n25958 , n373563 , n373564 , n25961 , n373566 , n373567 , n25964 , 
 n373569 , n373570 , n25967 , n25968 , n25969 , n25970 , n25971 , n373576 , n373577 , n25974 , 
 n373579 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n373588 , 
 n25985 , n373590 , n373591 , n25988 , n25989 , n25990 , n25991 , n373596 , n373597 , n25994 , 
 n25995 , n25996 , n25997 , n25998 , n373603 , n373604 , n26001 , n373606 , n373607 , n26004 , 
 n373609 , n373610 , n26007 , n373612 , n373613 , n26010 , n373615 , n373616 , n373617 , n26014 , 
 n26015 , n26016 , n26017 , n26018 , n373623 , n26020 , n26021 , n373626 , n26023 , n373628 , 
 n26025 , n26026 , n373631 , n373632 , n26029 , n373634 , n373635 , n26032 , n373637 , n373638 , 
 n373639 , n26036 , n373641 , n373642 , n26039 , n373644 , n373645 , n373646 , n26043 , n373648 , 
 n26045 , n373650 , n373651 , n373652 , n26049 , n373654 , n26051 , n26052 , n373657 , n373658 , 
 n26055 , n373660 , n373661 , n26058 , n373663 , n373664 , n26061 , n26062 , n26063 , n26064 , 
 n26065 , n26066 , n26067 , n373672 , n26069 , n26070 , n26071 , n373676 , n373677 , n26074 , 
 n26075 , n26076 , n373681 , n373682 , n26079 , n26080 , n26081 , n373686 , n373687 , n373688 , 
 n26085 , n373690 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n373697 , n373698 , 
 n26095 , n373700 , n373701 , n26098 , n373703 , n373704 , n26101 , n26102 , n26103 , n373708 , 
 n373709 , n26106 , n26107 , n26108 , n373713 , n373714 , n373715 , n26112 , n373717 , n26114 , 
 n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n373726 , n373727 , n26124 , 
 n373729 , n373730 , n26127 , n373732 , n373733 , n26130 , n26131 , n26132 , n373737 , n373738 , 
 n26135 , n26136 , n26137 , n373742 , n373743 , n26140 , n26141 , n373746 , n373747 , n26144 , 
 n373749 , n26146 , n373751 , n26148 , n373753 , n26150 , n26151 , n373756 , n373757 , n26154 , 
 n373759 , n373760 , n26157 , n373762 , n373763 , n26160 , n26161 , n373766 , n373767 , n26164 , 
 n373769 , n373770 , n26167 , n373772 , n373773 , n373774 , n26171 , n373776 , n26173 , n373778 , 
 n26175 , n26176 , n373781 , n373782 , n26179 , n373784 , n373785 , n26182 , n373787 , n373788 , 
 n26185 , n26186 , n373791 , n373792 , n26189 , n373794 , n373795 , n26192 , n373797 , n373798 , 
 n26195 , n373800 , n26197 , n26198 , n26199 , n373804 , n26201 , n373806 , n26203 , n26204 , 
 n373809 , n26206 , n26207 , n373812 , n373813 , n26210 , n373815 , n373816 , n26213 , n373818 , 
 n373819 , n26216 , n26217 , n26218 , n373823 , n373824 , n26221 , n26222 , n26223 , n373828 , 
 n373829 , n26226 , n26227 , n373832 , n373833 , n26230 , n26231 , n26232 , n373837 , n373838 , 
 n26235 , n26236 , n26237 , n373842 , n373843 , n26240 , n373845 , n373846 , n26243 , n373848 , 
 n26245 , n26246 , n373851 , n26248 , n26249 , n26250 , n373855 , n373856 , n26253 , n26254 , 
 n26255 , n26256 , n373861 , n373862 , n373863 , n26260 , n373865 , n26262 , n26263 , n373868 , 
 n373869 , n26266 , n373871 , n373872 , n26269 , n373874 , n373875 , n26272 , n26273 , n26274 , 
 n373879 , n373880 , n26277 , n26278 , n26279 , n373884 , n373885 , n373886 , n26283 , n373888 , 
 n26285 , n26286 , n373891 , n26288 , n373893 , n26290 , n26291 , n373896 , n373897 , n26294 , 
 n373899 , n373900 , n26297 , n373902 , n373903 , n373904 , n26301 , n373906 , n373907 , n26304 , 
 n373909 , n373910 , n26307 , n26308 , n26309 , n373914 , n373915 , n26312 , n26313 , n26314 , 
 n373919 , n373920 , n26317 , n26318 , n26319 , n373924 , n26321 , n373926 , n26323 , n26324 , 
 n373929 , n373930 , n26327 , n373932 , n373933 , n26330 , n373935 , n26332 , n26333 , n373938 , 
 n26335 , n26336 , n26337 , n373942 , n373943 , n26340 , n26341 , n26342 , n373947 , n373948 , 
 n26345 , n26346 , n373951 , n373952 , n26349 , n373954 , n26351 , n373956 , n26353 , n373958 , 
 n26355 , n26356 , n373961 , n373962 , n26359 , n373964 , n373965 , n26362 , n373967 , n373968 , 
 n26365 , n26366 , n373971 , n373972 , n26369 , n373974 , n373975 , n26372 , n373977 , n373978 , 
 n373979 , n26376 , n373981 , n26378 , n26379 , n373984 , n373985 , n26382 , n26383 , n373988 , 
 n26385 , n26386 , n373991 , n373992 , n373993 , n26390 , n373995 , n373996 , n26393 , n373998 , 
 n373999 , n26396 , n26397 , n26398 , n26399 , n374004 , n374005 , n374006 , n26403 , n374008 , 
 n26405 , n26406 , n374011 , n374012 , n26409 , n374014 , n374015 , n26412 , n374017 , n374018 , 
 n26415 , n26416 , n26417 , n374022 , n374023 , n26420 , n26421 , n26422 , n374027 , n374028 , 
 n26425 , n26426 , n26427 , n374032 , n374033 , n26430 , n26431 , n26432 , n374037 , n374038 , 
 n26435 , n374040 , n26437 , n374042 , n26439 , n26440 , n374045 , n26442 , n374047 , n26444 , 
 n26445 , n26446 , n26447 , n26448 , n374053 , n374054 , n26451 , n374056 , n26453 , n374058 , 
 n26455 , n26456 , n26457 , n374062 , n374063 , n26460 , n26461 , n26462 , n374067 , n374068 , 
 n26465 , n26466 , n26467 , n374072 , n374073 , n26470 , n26471 , n26472 , n374077 , n26474 , 
 n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n374087 , n374088 , 
 n374089 , n26486 , n374091 , n26488 , n374093 , n26490 , n26491 , n374096 , n374097 , n26494 , 
 n374099 , n374100 , n26497 , n374102 , n374103 , n26500 , n26501 , n374106 , n374107 , n26504 , 
 n374109 , n374110 , n26507 , n374112 , n374113 , n26510 , n26511 , n26512 , n26513 , n26514 , 
 n374119 , n374120 , n374121 , n26518 , n374123 , n26520 , n26521 , n374126 , n374127 , n26524 , 
 n374129 , n374130 , n26527 , n374132 , n374133 , n26530 , n26531 , n26532 , n374137 , n374138 , 
 n26535 , n374140 , n374141 , n26538 , n374143 , n374144 , n26541 , n26542 , n26543 , n26544 , 
 n374149 , n374150 , n26547 , n374152 , n26549 , n374154 , n26551 , n374156 , n26553 , n26554 , 
 n374159 , n26556 , n374161 , n26558 , n374163 , n374164 , n26561 , n374166 , n374167 , n26564 , 
 n26565 , n374170 , n374171 , n26568 , n374173 , n374174 , n26571 , n374176 , n374177 , n26574 , 
 n26575 , n26576 , n26577 , n374182 , n374183 , n26580 , n374185 , n26582 , n374187 , n26584 , 
 n374189 , n26586 , n26587 , n374192 , n374193 , n26590 , n374195 , n374196 , n26593 , n374198 , 
 n374199 , n26596 , n26597 , n374202 , n374203 , n26600 , n374205 , n374206 , n26603 , n374208 , 
 n374209 , n26606 , n374211 , n374212 , n26609 , n374214 , n374215 , n26612 , n26613 , n26614 , 
 n26615 , n374220 , n374221 , n26618 , n374223 , n374224 , n26621 , n374226 , n374227 , n26624 , 
 n374229 , n26626 , n26627 , n374232 , n26629 , n374234 , n374235 , n374236 , n26633 , n374238 , 
 n374239 , n26636 , n374241 , n374242 , n374243 , n374244 , n26641 , n374246 , n26643 , n26644 , 
 n374249 , n26646 , n374251 , n374252 , n26649 , n374254 , n374255 , n26652 , n374257 , n374258 , 
 n26655 , n374260 , n26657 , n26658 , n26659 , n26660 , n374265 , n374266 , n26663 , n374268 , 
 n374269 , n26666 , n26667 , n374272 , n374273 , n374274 , n26671 , n374276 , n26673 , n26674 , 
 n374279 , n26676 , n374281 , n26678 , n26679 , n26680 , n26681 , n374286 , n374287 , n26684 , 
 n374289 , n374290 , n26687 , n374292 , n374293 , n26690 , n26691 , n374296 , n374297 , n26694 , 
 n26695 , n26696 , n26697 , n26698 , n374303 , n374304 , n374305 , n26702 , n374307 , n26704 , 
 n26705 , n374310 , n374311 , n26708 , n374313 , n374314 , n26711 , n374316 , n374317 , n26714 , 
 n374319 , n26716 , n374321 , n26718 , n26719 , n374324 , n374325 , n26722 , n374327 , n374328 , 
 n26725 , n374330 , n374331 , n26728 , n26729 , n26730 , n374335 , n374336 , n26733 , n26734 , 
 n26735 , n374340 , n374341 , n26738 , n26739 , n26740 , n374345 , n374346 , n26743 , n26744 , 
 n26745 , n374350 , n374351 , n26748 , n374353 , n374354 , n26751 , n374356 , n374357 , n26754 , 
 n26755 , n374360 , n374361 , n26758 , n26759 , n26760 , n374365 , n374366 , n26763 , n26764 , 
 n374369 , n374370 , n374371 , n26768 , n374373 , n26770 , n26771 , n374376 , n374377 , n26774 , 
 n26775 , n374380 , n26777 , n26778 , n374383 , n374384 , n374385 , n26782 , n374387 , n374388 , 
 n26785 , n374390 , n374391 , n26788 , n26789 , n26790 , n26791 , n26792 , n374397 , n374398 , 
 n26795 , n26796 , n26797 , n374402 , n374403 , n26800 , n26801 , n26802 , n374407 , n374408 , 
 n26805 , n26806 , n26807 , n374412 , n374413 , n26810 , n374415 , n374416 , n26813 , n374418 , 
 n374419 , n26816 , n374421 , n374422 , n26819 , n26820 , n374425 , n26822 , n26823 , n26824 , 
 n26825 , n374430 , n374431 , n26828 , n26829 , n374434 , n374435 , n26832 , n26833 , n26834 , 
 n374439 , n374440 , n26837 , n26838 , n26839 , n374444 , n26841 , n26842 , n26843 , n374448 , 
 n374449 , n26846 , n26847 , n26848 , n26849 , n26850 , n374455 , n374456 , n26853 , n374458 , 
 n374459 , n26856 , n374461 , n26858 , n374463 , n26860 , n374465 , n26862 , n26863 , n374468 , 
 n26865 , n374470 , n374471 , n374472 , n374473 , n26870 , n374475 , n374476 , n374477 , n374478 , 
 n26875 , n374480 , n374481 , n26878 , n374483 , n374484 , n26881 , n374486 , n374487 , n26884 , 
 n374489 , n374490 , n26887 , n374492 , n26889 , n374494 , n374495 , n374496 , n26893 , n374498 , 
 n374499 , n26896 , n374501 , n374502 , n26899 , n374504 , n374505 , n26902 , n26903 , n26904 , 
 n26905 , n374510 , n26907 , n374512 , n374513 , n26910 , n374515 , n26912 , n26913 , n26914 , 
 n26915 , n26916 , n26917 , n374522 , n374523 , n26920 , n374525 , n26922 , n374527 , n374528 , 
 n26925 , n374530 , n374531 , n26928 , n374533 , n26930 , n26931 , n26932 , n26933 , n26934 , 
 n374539 , n374540 , n26937 , n374542 , n374543 , n26940 , n374545 , n26942 , n374547 , n26944 , 
 n26945 , n374550 , n374551 , n26948 , n374553 , n374554 , n26951 , n374556 , n374557 , n26954 , 
 n26955 , n374560 , n374561 , n26958 , n374563 , n374564 , n26961 , n374566 , n374567 , n26964 , 
 n374569 , n26966 , n26967 , n374572 , n26969 , n26970 , n374575 , n374576 , n26973 , n374578 , 
 n374579 , n26976 , n374581 , n374582 , n26979 , n374584 , n374585 , n26982 , n374587 , n26984 , 
 n374589 , n26986 , n26987 , n374592 , n26989 , n374594 , n26991 , n26992 , n374597 , n374598 , 
 n26995 , n374600 , n374601 , n26998 , n374603 , n374604 , n374605 , n27002 , n374607 , n374608 , 
 n27005 , n374610 , n374611 , n27008 , n374613 , n374614 , n27011 , n27012 , n27013 , n27014 , 
 n374619 , n374620 , n27017 , n27018 , n27019 , n27020 , n27021 , n374626 , n374627 , n27024 , 
 n374629 , n374630 , n374631 , n27028 , n374633 , n27030 , n27031 , n374636 , n27033 , n374638 , 
 n27035 , n27036 , n374641 , n374642 , n27039 , n27040 , n374645 , n374646 , n27043 , n374648 , 
 n374649 , n27046 , n27047 , n27048 , n27049 , n374654 , n27051 , n374656 , n27053 , n27054 , 
 n374659 , n27056 , n374661 , n27058 , n374663 , n27060 , n27061 , n27062 , n374667 , n27064 , 
 n374669 , n27066 , n374671 , n374672 , n27069 , n374674 , n374675 , n27072 , n27073 , n374678 , 
 n27075 , n27076 , n374681 , n374682 , n27079 , n27080 , n374685 , n374686 , n27083 , n374688 , 
 n374689 , n27086 , n374691 , n374692 , n27089 , n374694 , n374695 , n374696 , n27093 , n374698 , 
 n27095 , n27096 , n27097 , n27098 , n374703 , n27100 , n374705 , n27102 , n27103 , n374708 , 
 n374709 , n27106 , n374711 , n374712 , n27109 , n374714 , n374715 , n27112 , n27113 , n27114 , 
 n27115 , n374720 , n374721 , n27118 , n374723 , n27120 , n374725 , n27122 , n27123 , n27124 , 
 n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , 
 n27135 , n27136 , n27137 , n27138 , n27139 , n374744 , n374745 , n27142 , n374747 , n374748 , 
 n27145 , n374750 , n374751 , n27148 , n374753 , n374754 , n27151 , n27152 , n27153 , n27154 , 
 n27155 , n374760 , n374761 , n27158 , n374763 , n374764 , n27161 , n27162 , n27163 , n27164 , 
 n27165 , n374770 , n374771 , n27168 , n374773 , n374774 , n27171 , n374776 , n374777 , n27174 , 
 n27175 , n27176 , n27177 , n374782 , n374783 , n27180 , n374785 , n374786 , n27183 , n374788 , 
 n374789 , n374790 , n27187 , n374792 , n27189 , n374794 , n374795 , n27192 , n374797 , n27194 , 
 n27195 , n27196 , n374801 , n27198 , n27199 , n374804 , n27201 , n27202 , n27203 , n27204 , 
 n374809 , n374810 , n374811 , n374812 , n27209 , n27210 , n374815 , n27212 , n27213 , n27214 , 
 n27215 , n374820 , n374821 , n374822 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , 
 n374829 , n27226 , n374831 , n27228 , n27229 , n374834 , n374835 , n27232 , n374837 , n27234 , 
 n374839 , n27236 , n27237 , n374842 , n27239 , n27240 , n27241 , n27242 , n374847 , n374848 , 
 n374849 , n27246 , n374851 , n374852 , n27249 , n374854 , n27251 , n27252 , n374857 , n27254 , 
 n374859 , n27256 , n27257 , n27258 , n374863 , n27260 , n27261 , n374866 , n27263 , n27264 , 
 n27265 , n27266 , n374871 , n374872 , n374873 , n27270 , n374875 , n27272 , n374877 , n27274 , 
 n27275 , n374880 , n27277 , n374882 , n27279 , n27280 , n374885 , n374886 , n27283 , n374888 , 
 n374889 , n374890 , n27287 , n374892 , n27289 , n374894 , n374895 , n27292 , n374897 , n27294 , 
 n27295 , n374900 , n27297 , n374902 , n27299 , n27300 , n27301 , n374906 , n27303 , n27304 , 
 n374909 , n27306 , n27307 , n27308 , n27309 , n374914 , n374915 , n374916 , n27313 , n27314 , 
 n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , n374925 , n27322 , n27323 , n374928 , 
 n27325 , n27326 , n27327 , n27328 , n374933 , n374934 , n374935 , n27332 , n27333 , n27334 , 
 n27335 , n27336 , n27337 , n27338 , n27339 , n374944 , n374945 , n27342 , n374947 , n374948 , 
 n27345 , n374950 , n374951 , n27348 , n27349 , n27350 , n27351 , n374956 , n374957 , n27354 , 
 n27355 , n27356 , n27357 , n374962 , n374963 , n374964 , n27361 , n374966 , n27363 , n27364 , 
 n27365 , n27366 , n27367 , n27368 , n374973 , n374974 , n27371 , n374976 , n374977 , n27374 , 
 n374979 , n374980 , n27377 , n27378 , n27379 , n27380 , n374985 , n27382 , n374987 , n27384 , 
 n27385 , n374990 , n374991 , n27388 , n27389 , n374994 , n27391 , n374996 , n27393 , n374998 , 
 n374999 , n27396 , n27397 , n375002 , n27399 , n375004 , n27401 , n27402 , n375007 , n375008 , 
 n27405 , n375010 , n375011 , n27408 , n375013 , n27410 , n27411 , n27412 , n27413 , n27414 , 
 n27415 , n375020 , n375021 , n375022 , n27419 , n375024 , n375025 , n375026 , n27423 , n375028 , 
 n375029 , n27426 , n375031 , n375032 , n27429 , n27430 , n375035 , n375036 , n27433 , n375038 , 
 n375039 , n27436 , n375041 , n375042 , n27439 , n375044 , n375045 , n27442 , n27443 , n27444 , 
 n27445 , n27446 , n375051 , n375052 , n27449 , n375054 , n27451 , n375056 , n27453 , n375058 , 
 n375059 , n27456 , n375061 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , 
 n375069 , n27466 , n27467 , n375072 , n375073 , n27470 , n375075 , n375076 , n27473 , n375078 , 
 n375079 , n27476 , n375081 , n375082 , n27479 , n375084 , n375085 , n27482 , n27483 , n27484 , 
 n27485 , n375090 , n375091 , n27488 , n27489 , n27490 , n27491 , n27492 , n375097 , n375098 , 
 n375099 , n27496 , n375101 , n27498 , n375103 , n27500 , n375105 , n375106 , n27503 , n27504 , 
 n375109 , n375110 , n27507 , n375112 , n375113 , n27510 , n375115 , n375116 , n27513 , n27514 , 
 n27515 , n27516 , n375121 , n375122 , n27519 , n375124 , n375125 , n27522 , n27523 , n375128 , 
 n375129 , n27526 , n375131 , n375132 , n27529 , n27530 , n27531 , n27532 , n375137 , n375138 , 
 n27535 , n375140 , n27537 , n375142 , n27539 , n27540 , n375145 , n27542 , n27543 , n27544 , 
 n27545 , n27546 , n27547 , n27548 , n375153 , n27550 , n375155 , n27552 , n27553 , n27554 , 
 n375159 , n27556 , n375161 , n375162 , n27559 , n27560 , n375165 , n375166 , n27563 , n375168 , 
 n375169 , n27566 , n375171 , n375172 , n375173 , n27570 , n375175 , n375176 , n27573 , n375178 , 
 n375179 , n27576 , n375181 , n375182 , n27579 , n27580 , n27581 , n27582 , n27583 , n375188 , 
 n375189 , n27586 , n375191 , n375192 , n27589 , n375194 , n375195 , n27592 , n375197 , n375198 , 
 n27595 , n375200 , n375201 , n27598 , n375203 , n375204 , n375205 , n27602 , n375207 , n27604 , 
 n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , n375218 , 
 n27615 , n27616 , n375221 , n27618 , n27619 , n27620 , n27621 , n375226 , n375227 , n375228 , 
 n27625 , n375230 , n27627 , n375232 , n375233 , n375234 , n27631 , n375236 , n375237 , n375238 , 
 n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , 
 n27645 , n27646 , n27647 , n375252 , n375253 , n375254 , n27651 , n375256 , n375257 , n375258 , 
 n27655 , n375260 , n27657 , n375262 , n375263 , n375264 , n375265 , n27662 , n375267 , n375268 , 
 n375269 , n375270 , n27667 , n375272 , n375273 , n27670 , n375275 , n375276 , n27673 , n27674 , 
 n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n375287 , n27684 , 
 n375289 , n375290 , n27687 , n27688 , n27689 , n27690 , n375295 , n375296 , n27693 , n375298 , 
 n27695 , n375300 , n27697 , n27698 , n375303 , n375304 , n27701 , n27702 , n375307 , n375308 , 
 n375309 , n27706 , n375311 , n27708 , n27709 , n375314 , n27711 , n27712 , n27713 , n27714 , 
 n375319 , n375320 , n27717 , n375322 , n375323 , n27720 , n375325 , n375326 , n375327 , n27724 , 
 n375329 , n27726 , n375331 , n27728 , n27729 , n375334 , n375335 , n27732 , n375337 , n375338 , 
 n27735 , n375340 , n375341 , n27738 , n27739 , n375344 , n375345 , n27742 , n375347 , n375348 , 
 n27745 , n375350 , n375351 , n27748 , n375353 , n27750 , n27751 , n27752 , n27753 , n27754 , 
 n375359 , n27756 , n27757 , n27758 , n375363 , n375364 , n27761 , n375366 , n375367 , n27764 , 
 n375369 , n375370 , n27767 , n375372 , n375373 , n27770 , n375375 , n375376 , n27773 , n375378 , 
 n375379 , n27776 , n375381 , n375382 , n27779 , n375384 , n375385 , n27782 , n27783 , n27784 , 
 n27785 , n375390 , n375391 , n27788 , n27789 , n27790 , n27791 , n27792 , n375397 , n375398 , 
 n375399 , n27796 , n27797 , n375402 , n27799 , n27800 , n27801 , n27802 , n375407 , n27804 , 
 n375409 , n27806 , n27807 , n27808 , n27809 , n27810 , n375415 , n27812 , n27813 , n27814 , 
 n27815 , n375420 , n375421 , n27818 , n375423 , n27820 , n375425 , n27822 , n27823 , n27824 , 
 n27825 , n27826 , n27827 , n27828 , n375433 , n27830 , n375435 , n375436 , n27833 , n27834 , 
 n375439 , n27836 , n375441 , n375442 , n375443 , n27840 , n375445 , n375446 , n27843 , n375448 , 
 n375449 , n27846 , n27847 , n375452 , n375453 , n27850 , n375455 , n375456 , n27853 , n375458 , 
 n375459 , n27856 , n375461 , n375462 , n27859 , n27860 , n27861 , n27862 , n27863 , n375468 , 
 n375469 , n27866 , n375471 , n375472 , n27869 , n375474 , n27871 , n27872 , n27873 , n27874 , 
 n375479 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , 
 n27885 , n27886 , n27887 , n27888 , n27889 , n375494 , n375495 , n27892 , n375497 , n375498 , 
 n27895 , n375500 , n27897 , n27898 , n375503 , n27900 , n375505 , n27902 , n27903 , n27904 , 
 n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , 
 n375519 , n375520 , n27917 , n375522 , n375523 , n27920 , n27921 , n375526 , n27923 , n375528 , 
 n375529 , n375530 , n27927 , n375532 , n375533 , n375534 , n375535 , n27932 , n375537 , n375538 , 
 n27935 , n375540 , n375541 , n27938 , n27939 , n27940 , n375545 , n375546 , n27943 , n375548 , 
 n27945 , n375550 , n375551 , n27948 , n375553 , n375554 , n27951 , n375556 , n375557 , n27954 , 
 n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , 
 n375569 , n27966 , n375571 , n375572 , n27969 , n27970 , n27971 , n27972 , n375577 , n375578 , 
 n27975 , n375580 , n27977 , n375582 , n27979 , n27980 , n375585 , n375586 , n27983 , n375588 , 
 n375589 , n27986 , n375591 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , 
 n27995 , n375600 , n27997 , n375602 , n375603 , n375604 , n28001 , n28002 , n28003 , n28004 , 
 n28005 , n375610 , n28007 , n28008 , n375613 , n375614 , n28011 , n375616 , n375617 , n28014 , 
 n375619 , n375620 , n28017 , n375622 , n28019 , n375624 , n28021 , n28022 , n375627 , n375628 , 
 n28025 , n28026 , n375631 , n28028 , n28029 , n375634 , n375635 , n28032 , n375637 , n375638 , 
 n28035 , n375640 , n375641 , n28038 , n375643 , n28040 , n375645 , n28042 , n28043 , n28044 , 
 n375649 , n375650 , n28047 , n375652 , n375653 , n28050 , n375655 , n375656 , n28053 , n375658 , 
 n375659 , n28056 , n375661 , n375662 , n28059 , n28060 , n28061 , n28062 , n375667 , n375668 , 
 n28065 , n28066 , n28067 , n28068 , n375673 , n375674 , n28071 , n28072 , n28073 , n28074 , 
 n375679 , n375680 , n28077 , n375682 , n28079 , n375684 , n28081 , n28082 , n375687 , n375688 , 
 n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n375698 , 
 n28095 , n28096 , n375701 , n375702 , n28099 , n375704 , n375705 , n28102 , n375707 , n375708 , 
 n28105 , n375710 , n375711 , n28108 , n375713 , n375714 , n28111 , n375716 , n375717 , n28114 , 
 n28115 , n28116 , n28117 , n28118 , n375723 , n375724 , n28121 , n375726 , n375727 , n28124 , 
 n28125 , n28126 , n28127 , n28128 , n375733 , n375734 , n28131 , n375736 , n375737 , n28134 , 
 n28135 , n28136 , n28137 , n375742 , n375743 , n28140 , n375745 , n375746 , n28143 , n375748 , 
 n28145 , n375750 , n28147 , n375752 , n375753 , n375754 , n28151 , n375756 , n28153 , n28154 , 
 n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , n375765 , n28162 , n375767 , n375768 , 
 n375769 , n375770 , n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , 
 n375779 , n28176 , n375781 , n375782 , n28179 , n375784 , n28181 , n375786 , n28183 , n28184 , 
 n28185 , n375790 , n375791 , n28188 , n375793 , n28190 , n28191 , n375796 , n375797 , n28194 , 
 n375799 , n375800 , n28197 , n28198 , n375803 , n375804 , n28201 , n375806 , n28203 , n28204 , 
 n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , 
 n28215 , n375820 , n28217 , n375822 , n28219 , n28220 , n28221 , n375826 , n375827 , n28224 , 
 n375829 , n375830 , n28227 , n375832 , n375833 , n28230 , n375835 , n375836 , n28233 , n375838 , 
 n28235 , n375840 , n28237 , n375842 , n375843 , n28240 , n375845 , n28242 , n28243 , n375848 , 
 n375849 , n28246 , n375851 , n28248 , n28249 , n28250 , n375855 , n28252 , n28253 , n28254 , 
 n375859 , n375860 , n28257 , n28258 , n28259 , n28260 , n28261 , n375866 , n28263 , n375868 , 
 n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , n375878 , 
 n28275 , n28276 , n375881 , n375882 , n28279 , n375884 , n28281 , n28282 , n28283 , n28284 , 
 n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , 
 n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , n375905 , n28302 , n375907 , n375908 , 
 n28305 , n375910 , n375911 , n28308 , n28309 , n28310 , n375915 , n28312 , n375917 , n28314 , 
 n375919 , n375920 , n28317 , n375922 , n375923 , n28320 , n375925 , n28322 , n375927 , n28324 , 
 n375929 , n375930 , n28327 , n375932 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , 
 n28335 , n375940 , n28337 , n28338 , n375943 , n28340 , n28341 , n28342 , n28343 , n28344 , 
 n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n375958 , 
 n28355 , n375960 , n375961 , n28358 , n375963 , n28360 , n375965 , n375966 , n28363 , n375968 , 
 n375969 , n28366 , n375971 , n375972 , n375973 , n28370 , n375975 , n28372 , n375977 , n28374 , 
 n375979 , n375980 , n375981 , n28378 , n375983 , n375984 , n28381 , n375986 , n375987 , n28384 , 
 n28385 , n375990 , n28387 , n28388 , n375993 , n28390 , n375995 , n28392 , n28393 , n28394 , 
 n375999 , n376000 , n28397 , n28398 , n28399 , n376004 , n28401 , n376006 , n376007 , n28404 , 
 n376009 , n28406 , n376011 , n28408 , n376013 , n376014 , n28411 , n28412 , n376017 , n28414 , 
 n376019 , n376020 , n28417 , n28418 , n376023 , n28420 , n28421 , n376026 , n28423 , n28424 , 
 n376029 , n376030 , n28427 , n376032 , n376033 , n376034 , n28431 , n376036 , n376037 , n28434 , 
 n376039 , n376040 , n28437 , n376042 , n28439 , n376044 , n28441 , n28442 , n376047 , n376048 , 
 n28445 , n376050 , n376051 , n28448 , n376053 , n376054 , n28451 , n376056 , n376057 , n376058 , 
 n376059 , n28456 , n376061 , n376062 , n28459 , n376064 , n376065 , n28462 , n376067 , n28464 , 
 n28465 , n376070 , n376071 , n28468 , n28469 , n28470 , n376075 , n376076 , n376077 , n28474 , 
 n376079 , n28476 , n28477 , n28478 , n376083 , n376084 , n28481 , n376086 , n28483 , n28484 , 
 n28485 , n376090 , n376091 , n28488 , n376093 , n28490 , n28491 , n28492 , n376097 , n376098 , 
 n28495 , n376100 , n376101 , n376102 , n376103 , n28500 , n376105 , n376106 , n28503 , n376108 , 
 n376109 , n28506 , n376111 , n376112 , n28509 , n376114 , n376115 , n28512 , n376117 , n376118 , 
 n376119 , n376120 , n28517 , n376122 , n376123 , n28520 , n376125 , n376126 , n28523 , n376128 , 
 n376129 , n376130 , n376131 , n28528 , n376133 , n376134 , n28531 , n376136 , n376137 , n28534 , 
 n376139 , n376140 , n28537 , n376142 , n376143 , n28540 , n28541 , n28542 , n376147 , n376148 , 
 n28545 , n376150 , n376151 , n376152 , n28549 , n376154 , n28551 , n376156 , n376157 , n28554 , 
 n376159 , n28556 , n376161 , n28558 , n28559 , n376164 , n376165 , n28562 , n376167 , n376168 , 
 n28565 , n376170 , n28567 , n28568 , n28569 , n28570 , n376175 , n28572 , n28573 , n28574 , 
 n28575 , n28576 , n376181 , n28578 , n376183 , n376184 , n376185 , n376186 , n28583 , n376188 , 
 n376189 , n28586 , n376191 , n376192 , n28589 , n28590 , n376195 , n376196 , n28593 , n376198 , 
 n376199 , n28596 , n376201 , n376202 , n28599 , n376204 , n376205 , n376206 , n28603 , n28604 , 
 n28605 , n28606 , n376211 , n376212 , n28609 , n376214 , n376215 , n28612 , n376217 , n376218 , 
 n28615 , n376220 , n376221 , n28618 , n376223 , n28620 , n28621 , n376226 , n376227 , n28624 , 
 n376229 , n28626 , n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , 
 n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , n28641 , n28642 , n28643 , n28644 , 
 n28645 , n28646 , n28647 , n376252 , n28649 , n376254 , n376255 , n28652 , n376257 , n28654 , 
 n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , n376266 , n28663 , n376268 , 
 n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , n28671 , n376276 , n28673 , n376278 , 
 n28675 , n28676 , n28677 , n376282 , n28679 , n28680 , n376285 , n376286 , n28683 , n376288 , 
 n376289 , n28686 , n376291 , n376292 , n28689 , n376294 , n376295 , n28692 , n28693 , n376298 , 
 n376299 , n28696 , n376301 , n376302 , n28699 , n376304 , n376305 , n28702 , n28703 , n28704 , 
 n376309 , n28706 , n376311 , n28708 , n376313 , n376314 , n28711 , n376316 , n376317 , n28714 , 
 n28715 , n376320 , n376321 , n28718 , n376323 , n376324 , n28721 , n376326 , n376327 , n28724 , 
 n28725 , n28726 , n376331 , n376332 , n28729 , n28730 , n28731 , n376336 , n28733 , n28734 , 
 n28735 , n376340 , n376341 , n28738 , n28739 , n28740 , n376345 , n376346 , n28743 , n28744 , 
 n28745 , n376350 , n376351 , n28748 , n28749 , n28750 , n376355 , n376356 , n28753 , n28754 , 
 n28755 , n376360 , n376361 , n376362 , n376363 , n28760 , n376365 , n376366 , n376367 , n28764 , 
 n376369 , n376370 , n28767 , n376372 , n376373 , n28770 , n376375 , n28772 , n28773 , n28774 , 
 n376379 , n28776 , n376381 , n28778 , n28779 , n376384 , n28781 , n376386 , n376387 , n28784 , 
 n376389 , n28786 , n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , 
 n28795 , n28796 , n376401 , n376402 , n28799 , n376404 , n28801 , n376406 , n28803 , n28804 , 
 n376409 , n376410 , n28807 , n376412 , n376413 , n28810 , n376415 , n376416 , n28813 , n28814 , 
 n28815 , n376420 , n376421 , n28818 , n376423 , n28820 , n376425 , n28822 , n376427 , n376428 , 
 n28825 , n376430 , n28827 , n376432 , n28829 , n28830 , n376435 , n28832 , n376437 , n28834 , 
 n28835 , n376440 , n376441 , n28838 , n376443 , n376444 , n28841 , n376446 , n376447 , n376448 , 
 n28845 , n376450 , n376451 , n28848 , n376453 , n376454 , n28851 , n376456 , n376457 , n28854 , 
 n28855 , n28856 , n28857 , n376462 , n376463 , n28860 , n376465 , n28862 , n376467 , n376468 , 
 n28865 , n28866 , n376471 , n28868 , n28869 , n376474 , n376475 , n28872 , n28873 , n376478 , 
 n376479 , n28876 , n376481 , n376482 , n28879 , n28880 , n376485 , n376486 , n28883 , n376488 , 
 n376489 , n28886 , n28887 , n28888 , n28889 , n376494 , n376495 , n28892 , n376497 , n28894 , 
 n376499 , n28896 , n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , 
 n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , n376518 , 
 n28915 , n376520 , n376521 , n28918 , n28919 , n376524 , n28921 , n376526 , n376527 , n28924 , 
 n28925 , n376530 , n376531 , n28928 , n28929 , n376534 , n376535 , n28932 , n376537 , n376538 , 
 n28935 , n376540 , n376541 , n28938 , n376543 , n376544 , n28941 , n376546 , n376547 , n28944 , 
 n28945 , n28946 , n28947 , n376552 , n376553 , n28950 , n28951 , n28952 , n28953 , n28954 , 
 n376559 , n376560 , n376561 , n28958 , n28959 , n28960 , n376565 , n28962 , n376567 , n28964 , 
 n28965 , n376570 , n28967 , n28968 , n376573 , n376574 , n28971 , n376576 , n376577 , n28974 , 
 n376579 , n376580 , n376581 , n376582 , n28979 , n376584 , n376585 , n376586 , n28983 , n376588 , 
 n28985 , n376590 , n28987 , n28988 , n376593 , n376594 , n28991 , n376596 , n376597 , n28994 , 
 n376599 , n376600 , n28997 , n28998 , n376603 , n376604 , n29001 , n376606 , n376607 , n29004 , 
 n376609 , n376610 , n29007 , n376612 , n29009 , n29010 , n29011 , n29012 , n376617 , n376618 , 
 n29015 , n376620 , n29017 , n376622 , n29019 , n29020 , n29021 , n376626 , n29023 , n376628 , 
 n376629 , n29026 , n376631 , n376632 , n29029 , n29030 , n29031 , n29032 , n29033 , n376638 , 
 n376639 , n29036 , n376641 , n376642 , n29039 , n29040 , n29041 , n29042 , n29043 , n376648 , 
 n376649 , n29046 , n376651 , n376652 , n29049 , n376654 , n376655 , n29052 , n29053 , n29054 , 
 n29055 , n29056 , n376661 , n376662 , n29059 , n376664 , n376665 , n29062 , n376667 , n376668 , 
 n29065 , n376670 , n376671 , n376672 , n29069 , n376674 , n29071 , n29072 , n29073 , n29074 , 
 n29075 , n29076 , n29077 , n29078 , n376683 , n29080 , n376685 , n376686 , n29083 , n376688 , 
 n376689 , n29086 , n29087 , n29088 , n29089 , n376694 , n376695 , n29092 , n376697 , n376698 , 
 n29095 , n376700 , n376701 , n29098 , n376703 , n376704 , n29101 , n376706 , n376707 , n29104 , 
 n376709 , n376710 , n376711 , n376712 , n29109 , n376714 , n29111 , n376716 , n376717 , n29114 , 
 n376719 , n376720 , n29117 , n29118 , n29119 , n29120 , n376725 , n376726 , n376727 , n29124 , 
 n376729 , n376730 , n29127 , n29128 , n29129 , n29130 , n376735 , n376736 , n376737 , n29134 , 
 n29135 , n376740 , n29137 , n29138 , n376743 , n376744 , n376745 , n376746 , n376747 , n29144 , 
 n29145 , n29146 , n29147 , n29148 , n376753 , n29150 , n29151 , n376756 , n29153 , n29154 , 
 n376759 , n29156 , n29157 , n376762 , n29159 , n29160 , n376765 , n376766 , n376767 , n376768 , 
 n29165 , n29166 , n376771 , n29168 , n29169 , n376774 , n376775 , n376776 , n376777 , n29174 , 
 n29175 , n29176 , n29177 , n29178 , n376783 , n376784 , n376785 , n376786 , n376787 , n29184 , 
 n376789 , n376790 , n29187 , n29188 , n29189 , n29190 , n376795 , n376796 , n376797 , n29194 , 
 n29195 , n376800 , n29197 , n29198 , n376803 , n376804 , n376805 , n376806 , n376807 , n29204 , 
 n29205 , n29206 , n29207 , n29208 , n376813 , n376814 , n376815 , n376816 , n29213 , n376818 , 
 n376819 , n376820 , n376821 , n29218 , n29219 , n29220 , n29221 , n29222 , n376827 , n376828 , 
 n376829 , n29226 , n376831 , n376832 , n376833 , n376834 , n376835 , n29232 , n29233 , n29234 , 
 n29235 , n29236 , n376841 , n376842 , n376843 , n376844 , n376845 , n29242 , n376847 , n376848 , 
 n29245 , n29246 , n29247 , n29248 , n376853 , n29250 , n29251 , n376856 , n376857 , n376858 , 
 n29255 , n376860 , n376861 , n376862 , n29259 , n376864 , n376865 , n376866 , n29263 , n376868 , 
 n376869 , n376870 , n29267 , n376872 , n376873 , n376874 , n29271 , n376876 , n376877 , n376878 , 
 n29275 , n376880 , n376881 , n376882 , n376883 , n376884 , n29281 , n376886 , n376887 , n29284 , 
 n29285 , n29286 , n29287 , n376892 , n29289 , n29290 , n376895 , n29292 , n29293 , n376898 , 
 n29295 , n29296 , n376901 , n29298 , n29299 , n376904 , n376905 , n376906 , n376907 , n29304 , 
 n29305 , n29306 , n29307 , n376912 , n376913 , n376914 , n376915 , n29312 , n29313 , n29314 , 
 n29315 , n376920 , n376921 , n376922 , n376923 , n29320 , n29321 , n29322 , n29323 , n376928 , 
 n376929 , n376930 , n376931 , n29328 , n29329 , n29330 , n29331 , n376936 , n376937 , n376938 , 
 n376939 , n29336 , n29337 , n29338 , n29339 , n376944 , n376945 , n376946 , n376947 , n29344 , 
 n29345 , n29346 , n29347 , n376952 , n29349 , n29350 , n29351 , n29352 , n376957 , n376958 , 
 n29355 , n376960 , n376961 , n376962 , n29359 , n376964 , n29361 , n29362 , n29363 , n29364 , 
 n376969 , n376970 , n29367 , n376972 , n376973 , n376974 , n29371 , n376976 , n376977 , n376978 , 
 n29375 , n376980 , n376981 , n376982 , n29379 , n376984 , n376985 , n29382 , n376987 , n29384 , 
 n376989 , n29386 , n376991 , n376992 , n29389 , n376994 , n376995 , n29392 , n29393 , n376998 , 
 n376999 , n29396 , n377001 , n377002 , n29399 , n377004 , n377005 , n29402 , n29403 , n377008 , 
 n29405 , n377010 , n29407 , n29408 , n377013 , n377014 , n29411 , n377016 , n377017 , n29414 , 
 n377019 , n377020 , n377021 , n29418 , n377023 , n377024 , n29421 , n377026 , n377027 , n29424 , 
 n377029 , n377030 , n377031 , n377032 , n29429 , n377034 , n29431 , n377036 , n377037 , n29434 , 
 n29435 , n377040 , n29437 , n377042 , n377043 , n377044 , n29441 , n377046 , n377047 , n29444 , 
 n377049 , n377050 , n29447 , n377052 , n29449 , n377054 , n29451 , n377056 , n377057 , n29454 , 
 n377059 , n29456 , n29457 , n377062 , n377063 , n29460 , n377065 , n29462 , n29463 , n29464 , 
 n377069 , n29466 , n377071 , n29468 , n377073 , n377074 , n29471 , n377076 , n377077 , n29474 , 
 n377079 , n29476 , n377081 , n377082 , n29479 , n377084 , n377085 , n377086 , n29483 , n377088 , 
 n29485 , n29486 , n29487 , n29488 , n377093 , n29490 , n29491 , n377096 , n377097 , n29494 , 
 n377099 , n377100 , n29497 , n377102 , n377103 , n29500 , n29501 , n377106 , n29503 , n377108 , 
 n29505 , n29506 , n377111 , n377112 , n29509 , n377114 , n377115 , n29512 , n377117 , n377118 , 
 n377119 , n29516 , n377121 , n377122 , n29519 , n377124 , n377125 , n377126 , n29523 , n377128 , 
 n29525 , n29526 , n377131 , n29528 , n377133 , n29530 , n377135 , n377136 , n377137 , n377138 , 
 n377139 , n29536 , n377141 , n377142 , n377143 , n377144 , n377145 , n377146 , n377147 , n29544 , 
 n377149 , n377150 , n377151 , n377152 , n377153 , n29550 , n377155 , n377156 , n377157 , n377158 , 
 n377159 , n29556 , n377161 , n29558 , n377163 , n29560 , n377165 , n29562 , n377167 , n377168 , 
 n377169 , n377170 , n377171 , n377172 , n377173 , n29570 , n377175 , n29572 , n377177 , n29574 , 
 n377179 , n377180 , n377181 , n29578 , n377183 , n377184 , n377185 , n377186 , n377187 , n377188 , 
 n377189 , n377190 , n377191 , n29588 , n377193 , n377194 , n377195 , n29592 , n377197 , n29594 , 
 n377199 , n377200 , n377201 , n377202 , n377203 , n29600 , n377205 , n377206 , n377207 , n377208 , 
 n377209 , n29606 , n377211 , n377212 , n377213 , n29610 , n377215 , n377216 , n377217 , n377218 , 
 n377219 , n29616 , n377221 , n29618 , n377223 , n29620 , n377225 , n377226 , n377227 , n29624 , 
 n377229 , n377230 , n377231 , n29628 , n377233 , n377234 , n377235 , n29632 , n377237 , n377238 , 
 n377239 , n377240 , n377241 , n377242 , n377243 , n377244 , n377245 , n29642 , n377247 , n377248 , 
 n377249 , n377250 , n377251 , n29648 , n377253 , n377254 , n377255 , n29652 , n377257 , n377258 , 
 n377259 , n377260 , n377261 , n29658 , n377263 , n377264 , n377265 , n29662 , n377267 , n29664 , 
 n377269 , n377270 , n377271 , n377272 , n377273 , n29670 , n377275 , n377276 , n377277 , n377278 , 
 n377279 , n29676 , n377281 , n377282 , n377283 , n29680 , n377285 , n377286 , n377287 , n377288 , 
 n377289 , n29686 , n377291 , n29688 , n377293 , n29690 , n377295 , n29692 , n377297 , n377298 , 
 n377299 , n29696 , n377301 , n377302 , n377303 , n377304 , n377305 , n29702 , n377307 , n377308 , 
 n377309 , n29706 , n377311 , n377312 , n377313 , n377314 , n377315 , n29712 , n377317 , n29714 , 
 n377319 , n377320 , n377321 , n377322 , n377323 , n377324 , n377325 , n29722 , n377327 , n29724 , 
 n377329 , n29726 , n377331 , n377332 , n377333 , n29730 , n377335 , n377336 , n377337 , n377338 , 
 n377339 , n377340 , n377341 , n377342 , n377343 , n29740 , n377345 , n377346 , n377347 , n29744 , 
 n377349 , n377350 , n377351 , n377352 , n377353 , n377354 , n377355 , n29752 , n377357 , n377358 , 
 n377359 , n377360 , n377361 , n29758 , n377363 , n29760 , n377365 , n29762 , n377367 , n377368 , 
 n377369 , n377370 , n377371 , n29768 , n377373 , n377374 , n377375 , n377376 , n377377 , n29774 , 
 n377379 , n377380 , n377381 , n29778 , n377383 , n377384 , n377385 , n377386 , n377387 , n377388 , 
 n377389 , n29783 , n377391 , n377392 , n29786 , n29787 , n29788 , n377396 , n377397 , n29791 , 
 n29792 , n29793 , n377401 , n377402 , n29796 , n377404 , n29798 , n377406 , n29800 , n377408 , 
 n377409 , n29803 , n377411 , n377412 , n377413 , n29807 , n377415 , n377416 , n377417 , n29811 , 
 n377419 , n29813 , n377421 , n29815 , n377423 , n29817 , n377425 , n377426 , n29820 , n29821 , 
 n377429 , n377430 , n377431 , n377432 , n377433 , n29827 , n377435 , n377436 , n377437 , n29831 , 
 n377439 , n29833 , n377441 , n29835 , n29836 , n377444 , n29838 , n377446 , n29840 , n377448 , 
 n377449 , n29843 , n377451 , n377452 , n29846 , n29847 , n377455 , n377456 , n29850 , n377458 , 
 n377459 , n29853 , n377461 , n377462 , n29856 , n29857 , n29858 , n377466 , n377467 , n377468 , 
 n29862 , n377470 , n377471 , n29865 , n29866 , n29867 , n377475 , n377476 , n29870 , n29871 , 
 n377479 , n377480 , n377481 , n29875 , n377483 , n377484 , n29878 , n377486 , n29880 , n377488 , 
 n29882 , n377490 , n377491 , n29885 , n377493 , n29887 , n377495 , n377496 , n377497 , n377498 , 
 n29892 , n377500 , n377501 , n29895 , n29896 , n377504 , n377505 , n377506 , n377507 , n377508 , 
 n29902 , n377510 , n377511 , n377512 , n377513 , n29907 , n377515 , n377516 , n377517 , n29911 , 
 n29912 , n377520 , n377521 , n29915 , n377523 , n377524 , n29918 , n377526 , n377527 , n29921 , 
 n29922 , n377530 , n377531 , n29925 , n377533 , n377534 , n29928 , n377536 , n377537 , n29931 , 
 n377539 , n29933 , n377541 , n29935 , n29936 , n377544 , n29938 , n377546 , n29940 , n29941 , 
 n377549 , n377550 , n377551 , n377552 , n377553 , n29947 , n377555 , n377556 , n377557 , n377558 , 
 n29952 , n377560 , n377561 , n29955 , n377563 , n377564 , n29958 , n377566 , n29960 , n377568 , 
 n377569 , n29963 , n377571 , n29965 , n377573 , n377574 , n29968 , n377576 , n29970 , n377578 , 
 n377579 , n29973 , n377581 , n29975 , n377583 , n377584 , n29978 , n377586 , n29980 , n377588 , 
 n29982 , n29983 , n377591 , n29985 , n377593 , n377594 , n29988 , n377596 , n377597 , n377598 , 
 n29992 , n29993 , n377601 , n29995 , n29996 , n29997 , n377605 , n377606 , n377607 , n30001 , 
 n30002 , n377610 , n377611 , n30005 , n377613 , n377614 , n30008 , n377616 , n30010 , n30011 , 
 n377619 , n30013 , n377621 , n377622 , n377623 , n30017 , n377625 , n377626 , n30020 , n377628 , 
 n377629 , n30023 , n377631 , n30025 , n377633 , n377634 , n377635 , n377636 , n377637 , n30031 , 
 n30032 , n30033 , n377641 , n30035 , n377643 , n377644 , n30038 , n377646 , n30040 , n377648 , 
 n377649 , n30043 , n377651 , n377652 , n30046 , n377654 , n377655 , n377656 , n30050 , n30051 , 
 n30052 , n30053 , n377661 , n30055 , n30056 , n30057 , n30058 , n377666 , n377667 , n30061 , 
 n377669 , n30063 , n377671 , n30065 , n30066 , n30067 , n377675 , n377676 , n30070 , n30071 , 
 n377679 , n377680 , n377681 , n30075 , n30076 , n377684 , n377685 , n377686 , n30080 , n30081 , 
 n377689 , n377690 , n377691 , n30085 , n30086 , n377694 , n30088 , n377696 , n377697 , n30091 , 
 n30092 , n377700 , n377701 , n30095 , n30096 , n30097 , n377705 , n377706 , n30100 , n377708 , 
 n377709 , n30103 , n377711 , n30105 , n30106 , n377714 , n377715 , n377716 , n30110 , n377718 , 
 n30112 , n30113 , n377721 , n30115 , n377723 , n30117 , n30118 , n377726 , n377727 , n377728 , 
 n30122 , n377730 , n377731 , n30125 , n377733 , n377734 , n377735 , n377736 , n377737 , n377738 , 
 n30132 , n377740 , n377741 , n377742 , n30136 , n377744 , n377745 , n377746 , n30140 , n377748 , 
 n377749 , n30143 , n377751 , n377752 , n377753 , n30147 , n377755 , n377756 , n377757 , n377758 , 
 n30152 , n30153 , n377761 , n30155 , n377763 , n377764 , n30158 , n377766 , n30160 , n377768 , 
 n377769 , n30163 , n377771 , n377772 , n30166 , n30167 , n377775 , n377776 , n30170 , n377778 , 
 n377779 , n30173 , n377781 , n377782 , n30176 , n377784 , n377785 , n377786 , n377787 , n377788 , 
 n30182 , n30183 , n377791 , n30185 , n30186 , n377794 , n377795 , n377796 , n377797 , n377798 , 
 n30192 , n377800 , n377801 , n30195 , n377803 , n377804 , n30198 , n377806 , n377807 , n30201 , 
 n377809 , n30203 , n377811 , n30205 , n377813 , n30207 , n30208 , n377816 , n30210 , n377818 , 
 n30212 , n30213 , n377821 , n377822 , n30216 , n377824 , n377825 , n377826 , n377827 , n377828 , 
 n377829 , n30223 , n377831 , n377832 , n30226 , n377834 , n377835 , n377836 , n30230 , n377838 , 
 n30232 , n30233 , n377841 , n377842 , n30236 , n377844 , n30238 , n377846 , n30240 , n30241 , 
 n30242 , n377850 , n377851 , n377852 , n377853 , n377854 , n30248 , n377856 , n30250 , n377858 , 
 n30252 , n30253 , n377861 , n30255 , n377863 , n30257 , n377865 , n377866 , n30260 , n377868 , 
 n377869 , n30263 , n377871 , n377872 , n377873 , n30267 , n377875 , n377876 , n30270 , n377878 , 
 n377879 , n30273 , n377881 , n30275 , n377883 , n30277 , n377885 , n377886 , n30280 , n377888 , 
 n30282 , n377890 , n377891 , n377892 , n377893 , n30287 , n377895 , n377896 , n30290 , n30291 , 
 n377899 , n377900 , n377901 , n377902 , n377903 , n30297 , n377905 , n377906 , n30300 , n30301 , 
 n30302 , n377910 , n377911 , n30305 , n30306 , n30307 , n377915 , n377916 , n30310 , n377918 , 
 n377919 , n377920 , n377921 , n377922 , n30316 , n30317 , n377925 , n377926 , n30320 , n377928 , 
 n377929 , n30323 , n377931 , n30325 , n30326 , n377934 , n377935 , n377936 , n30330 , n30331 , 
 n30332 , n377940 , n377941 , n30335 , n377943 , n30337 , n377945 , n377946 , n30340 , n377948 , 
 n377949 , n30343 , n377951 , n377952 , n30346 , n377954 , n377955 , n377956 , n30350 , n30351 , 
 n377959 , n377960 , n377961 , n30355 , n30356 , n377964 , n377965 , n377966 , n30360 , n377968 , 
 n377969 , n30363 , n377971 , n30365 , n377973 , n30367 , n30368 , n377976 , n30370 , n377978 , 
 n30372 , n377980 , n377981 , n377982 , n30376 , n30377 , n377985 , n377986 , n30380 , n377988 , 
 n377989 , n377990 , n377991 , n377992 , n30386 , n377994 , n377995 , n377996 , n377997 , n30391 , 
 n30392 , n30393 , n378001 , n378002 , n30396 , n378004 , n378005 , n378006 , n378007 , n378008 , 
 n30402 , n378010 , n378011 , n30405 , n30406 , n30407 , n378015 , n378016 , n30410 , n30411 , 
 n30412 , n378020 , n378021 , n30415 , n30416 , n378024 , n378025 , n30419 , n378027 , n30421 , 
 n378029 , n30423 , n378031 , n30425 , n30426 , n378034 , n378035 , n30429 , n378037 , n378038 , 
 n30432 , n378040 , n378041 , n30435 , n30436 , n378044 , n30438 , n378046 , n30440 , n30441 , 
 n378049 , n30443 , n378051 , n378052 , n378053 , n30447 , n378055 , n378056 , n30450 , n378058 , 
 n378059 , n378060 , n30454 , n378062 , n30456 , n30457 , n378065 , n30459 , n378067 , n30461 , 
 n30462 , n378070 , n378071 , n30465 , n378073 , n378074 , n30468 , n378076 , n378077 , n378078 , 
 n30472 , n378080 , n378081 , n30475 , n378083 , n378084 , n30478 , n378086 , n30480 , n378088 , 
 n30482 , n378090 , n30484 , n30485 , n378093 , n378094 , n30488 , n378096 , n378097 , n30491 , 
 n378099 , n378100 , n30494 , n30495 , n378103 , n378104 , n30498 , n378106 , n378107 , n30501 , 
 n378109 , n378110 , n30504 , n30505 , n30506 , n378114 , n378115 , n30509 , n30510 , n30511 , 
 n378119 , n378120 , n30514 , n378122 , n378123 , n30517 , n30518 , n30519 , n378127 , n378128 , 
 n378129 , n30523 , n378131 , n30525 , n378133 , n30527 , n30528 , n378136 , n378137 , n30531 , 
 n378139 , n378140 , n30534 , n378142 , n378143 , n30537 , n30538 , n378146 , n378147 , n30541 , 
 n378149 , n378150 , n30544 , n378152 , n378153 , n378154 , n30548 , n378156 , n30550 , n30551 , 
 n378159 , n30553 , n378161 , n30555 , n30556 , n378164 , n378165 , n30559 , n378167 , n378168 , 
 n30562 , n378170 , n378171 , n378172 , n30566 , n378174 , n378175 , n30569 , n378177 , n378178 , 
 n30572 , n378180 , n30574 , n378182 , n30576 , n30577 , n378185 , n30579 , n378187 , n30581 , 
 n30582 , n378190 , n378191 , n30585 , n378193 , n378194 , n30588 , n378196 , n378197 , n378198 , 
 n30592 , n378200 , n378201 , n30595 , n378203 , n378204 , n378205 , n30599 , n30600 , n30601 , 
 n30602 , n30603 , n378211 , n30605 , n30606 , n378214 , n378215 , n30609 , n378217 , n378218 , 
 n30612 , n378220 , n378221 , n30615 , n378223 , n30617 , n378225 , n30619 , n30620 , n378228 , 
 n30622 , n30623 , n378231 , n30625 , n30626 , n378234 , n378235 , n30629 , n378237 , n378238 , 
 n30632 , n378240 , n378241 , n378242 , n30636 , n378244 , n378245 , n30639 , n378247 , n378248 , 
 n30642 , n30643 , n30644 , n378252 , n378253 , n30647 , n30648 , n30649 , n378257 , n378258 , 
 n30652 , n30653 , n30654 , n378262 , n378263 , n30657 , n30658 , n30659 , n30660 , n30661 , 
 n378269 , n378270 , n30664 , n378272 , n30666 , n378274 , n30668 , n30669 , n378277 , n378278 , 
 n30672 , n378280 , n378281 , n30675 , n378283 , n30677 , n30678 , n30679 , n30680 , n378288 , 
 n30682 , n378290 , n30684 , n30685 , n30686 , n378294 , n378295 , n30689 , n30690 , n378298 , 
 n378299 , n30693 , n378301 , n30695 , n378303 , n30697 , n30698 , n30699 , n30700 , n30701 , 
 n30702 , n378310 , n378311 , n30705 , n378313 , n378314 , n30708 , n378316 , n378317 , n30711 , 
 n30712 , n30713 , n378321 , n378322 , n30716 , n30717 , n30718 , n378326 , n378327 , n30721 , 
 n30722 , n30723 , n378331 , n378332 , n30726 , n30727 , n30728 , n378336 , n378337 , n30731 , 
 n378339 , n30733 , n30734 , n30735 , n378343 , n378344 , n30738 , n30739 , n378347 , n378348 , 
 n30742 , n30743 , n30744 , n378352 , n378353 , n378354 , n30748 , n378356 , n30750 , n30751 , 
 n378359 , n30753 , n378361 , n30755 , n30756 , n378364 , n30758 , n378366 , n30760 , n378368 , 
 n378369 , n30763 , n378371 , n378372 , n30766 , n378374 , n378375 , n378376 , n30770 , n378378 , 
 n30772 , n378380 , n30774 , n30775 , n378383 , n378384 , n30778 , n378386 , n378387 , n30781 , 
 n378389 , n378390 , n30784 , n30785 , n378393 , n378394 , n30788 , n378396 , n378397 , n30791 , 
 n378399 , n378400 , n30794 , n378402 , n30796 , n378404 , n30798 , n30799 , n30800 , n30801 , 
 n30802 , n30803 , n378411 , n378412 , n30806 , n378414 , n378415 , n30809 , n378417 , n378418 , 
 n378419 , n30813 , n378421 , n30815 , n30816 , n378424 , n30818 , n378426 , n30820 , n30821 , 
 n378429 , n378430 , n30824 , n378432 , n378433 , n30827 , n378435 , n378436 , n378437 , n30831 , 
 n378439 , n378440 , n30834 , n378442 , n378443 , n30837 , n378445 , n378446 , n30840 , n378448 , 
 n378449 , n30843 , n378451 , n30845 , n378453 , n30847 , n378455 , n30849 , n30850 , n378458 , 
 n30852 , n378460 , n30854 , n30855 , n378463 , n378464 , n30858 , n378466 , n378467 , n30861 , 
 n378469 , n378470 , n378471 , n30865 , n378473 , n378474 , n30868 , n378476 , n378477 , n30871 , 
 n30872 , n30873 , n378481 , n378482 , n30876 , n30877 , n30878 , n378486 , n378487 , n30881 , 
 n30882 , n30883 , n378491 , n378492 , n30886 , n30887 , n378495 , n30889 , n378497 , n30891 , 
 n30892 , n378500 , n378501 , n30895 , n378503 , n378504 , n30898 , n378506 , n30900 , n30901 , 
 n30902 , n30903 , n30904 , n30905 , n30906 , n30907 , n378515 , n30909 , n30910 , n378518 , 
 n378519 , n30913 , n378521 , n30915 , n378523 , n30917 , n30918 , n378526 , n30920 , n378528 , 
 n30922 , n378530 , n378531 , n30925 , n378533 , n30927 , n378535 , n30929 , n378537 , n378538 , 
 n30932 , n30933 , n378541 , n30935 , n378543 , n378544 , n30938 , n378546 , n378547 , n30941 , 
 n30942 , n30943 , n378551 , n378552 , n30946 , n30947 , n378555 , n378556 , n30950 , n30951 , 
 n30952 , n378560 , n378561 , n30955 , n30956 , n30957 , n378565 , n378566 , n30960 , n30961 , 
 n30962 , n378570 , n378571 , n30965 , n30966 , n30967 , n378575 , n30969 , n30970 , n30971 , 
 n30972 , n378580 , n30974 , n30975 , n378583 , n378584 , n30978 , n30979 , n378587 , n378588 , 
 n30982 , n30983 , n30984 , n378592 , n378593 , n378594 , n30988 , n30989 , n30990 , n30991 , 
 n30992 , n378600 , n30994 , n30995 , n378603 , n378604 , n30998 , n378606 , n378607 , n31001 , 
 n378609 , n378610 , n378611 , n31005 , n378613 , n31007 , n31008 , n378616 , n31010 , n378618 , 
 n31012 , n31013 , n378621 , n31015 , n378623 , n378624 , n378625 , n31019 , n31020 , n378628 , 
 n378629 , n31023 , n378631 , n31025 , n378633 , n378634 , n31028 , n378636 , n378637 , n31031 , 
 n378639 , n31033 , n378641 , n31035 , n31036 , n378644 , n31038 , n378646 , n31040 , n31041 , 
 n378649 , n378650 , n31044 , n378652 , n378653 , n31047 , n378655 , n378656 , n378657 , n31051 , 
 n378659 , n378660 , n31054 , n378662 , n378663 , n378664 , n31058 , n378666 , n31060 , n31061 , 
 n31062 , n378670 , n31064 , n378672 , n378673 , n31067 , n378675 , n378676 , n31070 , n378678 , 
 n31072 , n378680 , n31074 , n31075 , n31076 , n31077 , n31078 , n31079 , n378687 , n31081 , 
 n378689 , n378690 , n31084 , n31085 , n31086 , n378694 , n378695 , n31089 , n378697 , n31091 , 
 n31092 , n378700 , n378701 , n31095 , n378703 , n31097 , n378705 , n31099 , n31100 , n378708 , 
 n378709 , n31103 , n378711 , n378712 , n31106 , n378714 , n378715 , n31109 , n31110 , n31111 , 
 n378719 , n378720 , n31114 , n31115 , n31116 , n378724 , n378725 , n31119 , n378727 , n31121 , 
 n378729 , n31123 , n378731 , n378732 , n378733 , n31127 , n378735 , n31129 , n378737 , n378738 , 
 n378739 , n378740 , n31134 , n378742 , n378743 , n378744 , n378745 , n31139 , n378747 , n378748 , 
 n31142 , n378750 , n378751 , n31145 , n31146 , n378754 , n378755 , n31149 , n378757 , n31151 , 
 n378759 , n378760 , n31154 , n31155 , n378763 , n31157 , n31158 , n378766 , n378767 , n31161 , 
 n31162 , n378770 , n378771 , n31165 , n31166 , n378774 , n378775 , n31169 , n31170 , n31171 , 
 n378779 , n378780 , n31174 , n31175 , n378783 , n378784 , n31178 , n31179 , n31180 , n378788 , 
 n378789 , n31183 , n31184 , n31185 , n378793 , n378794 , n31188 , n31189 , n31190 , n378798 , 
 n378799 , n31193 , n31194 , n31195 , n378803 , n31197 , n31198 , n31199 , n31200 , n31201 , 
 n31202 , n378810 , n378811 , n31205 , n31206 , n378814 , n378815 , n31209 , n31210 , n31211 , 
 n31212 , n31213 , n378821 , n378822 , n31216 , n378824 , n31218 , n31219 , n31220 , n31221 , 
 n31222 , n378830 , n31224 , n31225 , n31226 , n31227 , n378835 , n31229 , n31230 , n31231 , 
 n31232 , n31233 , n378841 , n31235 , n31236 , n31237 , n31238 , n378846 , n31240 , n378848 , 
 n31242 , n31243 , n31244 , n378852 , n378853 , n378854 , n31248 , n378856 , n31250 , n31251 , 
 n378859 , n378860 , n31254 , n378862 , n378863 , n31257 , n378865 , n378866 , n378867 , n31261 , 
 n31262 , n378870 , n31264 , n31265 , n378873 , n378874 , n31268 , n378876 , n378877 , n31271 , 
 n378879 , n378880 , n31274 , n378882 , n31276 , n378884 , n31278 , n31279 , n31280 , n378888 , 
 n378889 , n31283 , n378891 , n378892 , n31286 , n378894 , n378895 , n31289 , n31290 , n31291 , 
 n378899 , n378900 , n378901 , n31295 , n378903 , n31297 , n31298 , n378906 , n31300 , n378908 , 
 n378909 , n378910 , n31304 , n378912 , n31306 , n31307 , n378915 , n378916 , n31310 , n378918 , 
 n378919 , n31313 , n378921 , n378922 , n31316 , n31317 , n31318 , n31319 , n378927 , n378928 , 
 n31322 , n31323 , n31324 , n378932 , n378933 , n31327 , n31328 , n31329 , n378937 , n378938 , 
 n31332 , n378940 , n31334 , n378942 , n31336 , n31337 , n378945 , n378946 , n31340 , n378948 , 
 n378949 , n31343 , n378951 , n378952 , n31346 , n378954 , n378955 , n31349 , n31350 , n31351 , 
 n378959 , n378960 , n31354 , n31355 , n31356 , n31357 , n378965 , n378966 , n31360 , n378968 , 
 n31362 , n378970 , n378971 , n31365 , n31366 , n378974 , n31368 , n31369 , n378977 , n378978 , 
 n31372 , n31373 , n378981 , n31375 , n378983 , n31377 , n31378 , n378986 , n378987 , n31381 , 
 n378989 , n378990 , n31384 , n378992 , n378993 , n378994 , n31388 , n378996 , n378997 , n31391 , 
 n378999 , n379000 , n31394 , n31395 , n31396 , n31397 , n31398 , n31399 , n31400 , n31401 , 
 n31402 , n379010 , n31404 , n31405 , n31406 , n31407 , n379015 , n379016 , n379017 , n31411 , 
 n379019 , n379020 , n31414 , n31415 , n31416 , n379024 , n379025 , n31419 , n31420 , n31421 , 
 n379029 , n379030 , n31424 , n31425 , n31426 , n31427 , n31428 , n379036 , n379037 , n31431 , 
 n31432 , n379040 , n379041 , n31435 , n31436 , n31437 , n379045 , n379046 , n31440 , n31441 , 
 n31442 , n31443 , n379051 , n379052 , n31446 , n31447 , n31448 , n379056 , n379057 , n31451 , 
 n31452 , n31453 , n379061 , n379062 , n31456 , n379064 , n379065 , n31459 , n379067 , n379068 , 
 n31462 , n31463 , n379071 , n379072 , n31466 , n31467 , n379075 , n379076 , n31470 , n31471 , 
 n31472 , n31473 , n31474 , n379082 , n379083 , n31477 , n31478 , n379086 , n379087 , n31481 , 
 n31482 , n31483 , n31484 , n31485 , n379093 , n379094 , n31488 , n31489 , n31490 , n379098 , 
 n379099 , n31493 , n31494 , n31495 , n379103 , n379104 , n31498 , n379106 , n31500 , n31501 , 
 n379109 , n379110 , n31504 , n31505 , n379113 , n379114 , n31508 , n31509 , n379117 , n379118 , 
 n31512 , n31513 , n31514 , n31515 , n31516 , n379124 , n379125 , n31519 , n31520 , n31521 , 
 n379129 , n379130 , n31524 , n379132 , n31526 , n379134 , n379135 , n31529 , n379137 , n31531 , 
 n31532 , n31533 , n379141 , n379142 , n31536 , n31537 , n379145 , n379146 , n31540 , n31541 , 
 n31542 , n31543 , n31544 , n379152 , n379153 , n31547 , n379155 , n31549 , n31550 , n31551 , 
 n31552 , n31553 , n379161 , n379162 , n31556 , n379164 , n31558 , n31559 , n31560 , n379168 , 
 n31562 , n31563 , n31564 , n31565 , n31566 , n379174 , n31568 , n31569 , n31570 , n31571 , 
 n31572 , n31573 , n31574 , n31575 , n379183 , n31577 , n379185 , n31579 , n31580 , n31581 , 
 n31582 , n31583 , n31584 , n379192 , n31586 , n379194 , n31588 , n31589 , n31590 , n31591 , 
 n31592 , n31593 , n31594 , n31595 , n31596 , n31597 , n31598 , n31599 , n31600 , n31601 , 
 n379209 , n379210 , n31604 , n31605 , n31606 , n31607 , n379215 , n379216 , n31610 , n379218 , 
 n31612 , n31613 , n31614 , n31615 , n379223 , n31617 , n379225 , n31619 , n31620 , n379228 , 
 n379229 , n31623 , n379231 , n379232 , n31626 , n379234 , n31628 , n31629 , n31630 , n379238 , 
 n31632 , n379240 , n379241 , n31635 , n379243 , n31637 , n379245 , n379246 , n379247 , n31641 , 
 n379249 , n379250 , n31644 , n379252 , n379253 , n31647 , n379255 , n31649 , n31650 , n379258 , 
 n379259 , n31653 , n379261 , n31655 , n31656 , n31657 , n379265 , n31659 , n379267 , n379268 , 
 n31662 , n379270 , n31664 , n379272 , n31666 , n379274 , n379275 , n31669 , n379277 , n31671 , 
 n31672 , n379280 , n31674 , n379282 , n379283 , n31677 , n379285 , n31679 , n379287 , n379288 , 
 n31682 , n379290 , n379291 , n379292 , n31686 , n379294 , n31688 , n31689 , n31690 , n379298 , 
 n31692 , n379300 , n379301 , n31695 , n379303 , n31697 , n31698 , n379306 , n379307 , n31701 , 
 n379309 , n379310 , n31704 , n379312 , n379313 , n31707 , n379315 , n379316 , n379317 , n31711 , 
 n379319 , n31713 , n379321 , n379322 , n31716 , n379324 , n31718 , n379326 , n31720 , n31721 , 
 n379329 , n31723 , n379331 , n31725 , n379333 , n379334 , n31728 , n379336 , n379337 , n31731 , 
 n379339 , n31733 , n31734 , n31735 , n31736 , n31737 , n379345 , n379346 , n31740 , n31741 , 
 n31742 , n31743 , n379351 , n379352 , n379353 , n31747 , n379355 , n31749 , n379357 , n31751 , 
 n31752 , n379360 , n379361 , n31755 , n379363 , n379364 , n31758 , n379366 , n379367 , n31761 , 
 n31762 , n379370 , n379371 , n31765 , n379373 , n379374 , n31768 , n379376 , n379377 , n379378 , 
 n31772 , n379380 , n31774 , n31775 , n379383 , n31777 , n379385 , n31779 , n31780 , n379388 , 
 n379389 , n31783 , n379391 , n379392 , n31786 , n379394 , n379395 , n379396 , n31790 , n379398 , 
 n379399 , n31793 , n379401 , n379402 , n31796 , n379404 , n379405 , n31799 , n379407 , n379408 , 
 n31802 , n379410 , n379411 , n31805 , n31806 , n31807 , n31808 , n31809 , n379417 , n379418 , 
 n31812 , n379420 , n379421 , n31815 , n379423 , n379424 , n31818 , n379426 , n31820 , n379428 , 
 n379429 , n31823 , n379431 , n31825 , n31826 , n31827 , n31828 , n31829 , n31830 , n31831 , 
 n31832 , n31833 , n31834 , n31835 , n31836 , n31837 , n31838 , n31839 , n31840 , n31841 , 
 n31842 , n31843 , n31844 , n31845 , n31846 , n31847 , n31848 , n31849 , n31850 , n379458 , 
 n31852 , n379460 , n379461 , n31855 , n379463 , n379464 , n31858 , n379466 , n379467 , n31861 , 
 n379469 , n31863 , n379471 , n379472 , n379473 , n31867 , n379475 , n379476 , n31870 , n379478 , 
 n31872 , n31873 , n379481 , n31875 , n379483 , n379484 , n31878 , n379486 , n379487 , n31881 , 
 n379489 , n31883 , n379491 , n379492 , n31886 , n379494 , n379495 , n31889 , n31890 , n379498 , 
 n379499 , n31893 , n379501 , n379502 , n31896 , n379504 , n379505 , n31899 , n379507 , n379508 , 
 n31902 , n31903 , n31904 , n31905 , n31906 , n379514 , n379515 , n31909 , n379517 , n31911 , 
 n31912 , n31913 , n31914 , n379522 , n31916 , n379524 , n379525 , n31919 , n379527 , n31921 , 
 n379529 , n31923 , n379531 , n31925 , n379533 , n379534 , n31928 , n379536 , n379537 , n31931 , 
 n379539 , n379540 , n31934 , n379542 , n379543 , n31937 , n379545 , n379546 , n379547 , n379548 , 
 n31942 , n379550 , n31944 , n379552 , n379553 , n31947 , n379555 , n379556 , n31950 , n379558 , 
 n379559 , n31953 , n379561 , n31955 , n31956 , n379564 , n379565 , n31959 , n379567 , n31961 , 
 n31962 , n31963 , n31964 , n379572 , n31966 , n379574 , n379575 , n31969 , n379577 , n379578 , 
 n31972 , n379580 , n31974 , n379582 , n31976 , n379584 , n31978 , n379586 , n379587 , n31981 , 
 n31982 , n379590 , n379591 , n31985 , n379593 , n379594 , n31988 , n379596 , n379597 , n31991 , 
 n31992 , n379600 , n31994 , n379602 , n31996 , n379604 , n379605 , n31999 , n379607 , n379608 , 
 n32002 , n32003 , n379611 , n379612 , n32006 , n379614 , n379615 , n32009 , n379617 , n379618 , 
 n379619 , n32013 , n379621 , n379622 , n32016 , n379624 , n379625 , n379626 , n32020 , n379628 , 
 n32022 , n379630 , n32024 , n32025 , n379633 , n379634 , n32028 , n379636 , n379637 , n32031 , 
 n379639 , n379640 , n32034 , n32035 , n379643 , n32037 , n379645 , n32039 , n379647 , n379648 , 
 n32042 , n32043 , n379651 , n379652 , n32046 , n379654 , n379655 , n32049 , n379657 , n379658 , 
 n379659 , n32053 , n379661 , n379662 , n32056 , n379664 , n379665 , n379666 , n379667 , n32061 , 
 n379669 , n379670 , n32064 , n379672 , n379673 , n32067 , n379675 , n32069 , n379677 , n32071 , 
 n379679 , n379680 , n32074 , n32075 , n379683 , n379684 , n32078 , n379686 , n379687 , n32081 , 
 n379689 , n379690 , n379691 , n32085 , n379693 , n32087 , n379695 , n379696 , n32090 , n379698 , 
 n379699 , n32093 , n32094 , n32095 , n379703 , n379704 , n32098 , n32099 , n379707 , n32101 , 
 n379709 , n32103 , n32104 , n379712 , n32106 , n379714 , n379715 , n379716 , n32110 , n379718 , 
 n379719 , n32113 , n379721 , n32115 , n32116 , n379724 , n32118 , n379726 , n32120 , n32121 , 
 n379729 , n32123 , n379731 , n379732 , n379733 , n32127 , n379735 , n379736 , n32130 , n379738 , 
 n32132 , n32133 , n379741 , n379742 , n32136 , n379744 , n32138 , n379746 , n32140 , n379748 , 
 n379749 , n32143 , n32144 , n379752 , n379753 , n32147 , n379755 , n379756 , n32150 , n379758 , 
 n379759 , n32153 , n32154 , n32155 , n32156 , n32157 , n379765 , n379766 , n32160 , n379768 , 
 n32162 , n32163 , n379771 , n32165 , n379773 , n379774 , n32168 , n379776 , n379777 , n32171 , 
 n379779 , n379780 , n32174 , n379782 , n379783 , n32177 , n379785 , n379786 , n379787 , n32181 , 
 n379789 , n32183 , n379791 , n32185 , n379793 , n379794 , n32188 , n32189 , n379797 , n32191 , 
 n379799 , n379800 , n379801 , n32195 , n379803 , n379804 , n32198 , n379806 , n379807 , n32201 , 
 n32202 , n379810 , n32204 , n32205 , n379813 , n32207 , n32208 , n379816 , n379817 , n32211 , 
 n379819 , n379820 , n32214 , n379822 , n379823 , n379824 , n32218 , n379826 , n379827 , n32221 , 
 n379829 , n379830 , n32224 , n32225 , n32226 , n32227 , n32228 , n32229 , n379837 , n379838 , 
 n32232 , n379840 , n32234 , n379842 , n32236 , n379844 , n379845 , n32239 , n379847 , n379848 , 
 n379849 , n32243 , n379851 , n32245 , n32246 , n379854 , n32248 , n379856 , n32250 , n32251 , 
 n379859 , n379860 , n32254 , n379862 , n379863 , n32257 , n379865 , n379866 , n379867 , n32261 , 
 n379869 , n379870 , n32264 , n379872 , n379873 , n32267 , n379875 , n32269 , n379877 , n32271 , 
 n32272 , n379880 , n32274 , n379882 , n32276 , n379884 , n379885 , n32279 , n32280 , n379888 , 
 n379889 , n32283 , n379891 , n379892 , n32286 , n379894 , n379895 , n379896 , n32290 , n379898 , 
 n379899 , n32293 , n379901 , n379902 , n32296 , n32297 , n32298 , n379906 , n379907 , n32301 , 
 n379909 , n379910 , n379911 , n32305 , n379913 , n32307 , n32308 , n379916 , n32310 , n379918 , 
 n32312 , n32313 , n379921 , n379922 , n32316 , n379924 , n379925 , n32319 , n379927 , n379928 , 
 n379929 , n32323 , n379931 , n379932 , n32326 , n379934 , n379935 , n379936 , n32330 , n379938 , 
 n32332 , n32333 , n379941 , n32335 , n379943 , n379944 , n379945 , n32339 , n379947 , n32341 , 
 n379949 , n379950 , n379951 , n32345 , n32346 , n379954 , n379955 , n32349 , n379957 , n379958 , 
 n32352 , n32353 , n32354 , n32355 , n379963 , n32357 , n379965 , n32359 , n32360 , n379968 , 
 n379969 , n32363 , n379971 , n379972 , n32366 , n379974 , n379975 , n379976 , n32370 , n379978 , 
 n32372 , n379980 , n379981 , n32375 , n379983 , n32377 , n379985 , n32379 , n32380 , n379988 , 
 n379989 , n32383 , n379991 , n379992 , n32386 , n379994 , n379995 , n32389 , n32390 , n379998 , 
 n379999 , n32393 , n380001 , n380002 , n32396 , n380004 , n380005 , n32399 , n380007 , n32401 , 
 n380009 , n32403 , n380011 , n32405 , n32406 , n380014 , n380015 , n32409 , n380017 , n380018 , 
 n32412 , n380020 , n380021 , n32415 , n32416 , n380024 , n380025 , n32419 , n380027 , n380028 , 
 n32422 , n380030 , n380031 , n32425 , n32426 , n32427 , n380035 , n380036 , n32430 , n32431 , 
 n32432 , n380040 , n380041 , n32435 , n32436 , n32437 , n380045 , n380046 , n32440 , n32441 , 
 n380049 , n380050 , n32444 , n380052 , n380053 , n32447 , n380055 , n32449 , n32450 , n380058 , 
 n32452 , n380060 , n32454 , n380062 , n380063 , n32457 , n380065 , n380066 , n380067 , n32461 , 
 n380069 , n380070 , n380071 , n380072 , n32466 , n380074 , n380075 , n380076 , n380077 , n32471 , 
 n380079 , n380080 , n32474 , n380082 , n380083 , n32477 , n380085 , n32479 , n380087 , n32481 , 
 n32482 , n380090 , n32484 , n380092 , n32486 , n32487 , n380095 , n380096 , n32490 , n380098 , 
 n380099 , n32493 , n380101 , n380102 , n380103 , n32497 , n380105 , n380106 , n32500 , n380108 , 
 n380109 , n32503 , n32504 , n32505 , n380113 , n380114 , n32508 , n32509 , n32510 , n380118 , 
 n380119 , n32513 , n380121 , n380122 , n32516 , n32517 , n32518 , n380126 , n380127 , n32521 , 
 n32522 , n32523 , n32524 , n32525 , n32526 , n32527 , n32528 , n380136 , n380137 , n32531 , 
 n380139 , n32533 , n32534 , n32535 , n32536 , n32537 , n380145 , n380146 , n32540 , n380148 , 
 n32542 , n380150 , n380151 , n32545 , n380153 , n380154 , n32548 , n380156 , n380157 , n380158 , 
 n380159 , n32553 , n380161 , n380162 , n32556 , n380164 , n32558 , n380166 , n32560 , n32561 , 
 n380169 , n32563 , n380171 , n32565 , n32566 , n380174 , n380175 , n32569 , n380177 , n380178 , 
 n32572 , n380180 , n380181 , n380182 , n32576 , n380184 , n380185 , n32579 , n380187 , n380188 , 
 n32582 , n32583 , n32584 , n380192 , n380193 , n32587 , n380195 , n32589 , n380197 , n32591 , 
 n32592 , n380200 , n32594 , n380202 , n32596 , n32597 , n380205 , n380206 , n32600 , n380208 , 
 n380209 , n32603 , n380211 , n380212 , n380213 , n32607 , n380215 , n380216 , n32610 , n380218 , 
 n380219 , n32613 , n32614 , n32615 , n32616 , n380224 , n380225 , n32619 , n380227 , n32621 , 
 n32622 , n32623 , n380231 , n380232 , n32626 , n380234 , n32628 , n380236 , n32630 , n32631 , 
 n32632 , n32633 , n380241 , n380242 , n32636 , n380244 , n32638 , n32639 , n32640 , n32641 , 
 n380249 , n32643 , n32644 , n32645 , n380253 , n380254 , n32648 , n32649 , n32650 , n380258 , 
 n380259 , n32653 , n32654 , n32655 , n380263 , n380264 , n32658 , n32659 , n380267 , n380268 , 
 n32662 , n380270 , n32664 , n32665 , n32666 , n32667 , n32668 , n380276 , n32670 , n32671 , 
 n32672 , n32673 , n32674 , n32675 , n380283 , n32677 , n380285 , n380286 , n32680 , n380288 , 
 n380289 , n32683 , n380291 , n32685 , n380293 , n380294 , n32688 , n380296 , n380297 , n32691 , 
 n32692 , n32693 , n380301 , n380302 , n32696 , n32697 , n32698 , n380306 , n380307 , n32701 , 
 n32702 , n32703 , n380311 , n380312 , n32706 , n32707 , n32708 , n380316 , n380317 , n32711 , 
 n380319 , n32713 , n32714 , n32715 , n380323 , n380324 , n32718 , n32719 , n380327 , n380328 , 
 n32722 , n32723 , n32724 , n380332 , n380333 , n380334 , n32728 , n380336 , n32730 , n32731 , 
 n380339 , n380340 , n32734 , n380342 , n380343 , n32737 , n380345 , n380346 , n380347 , n32741 , 
 n380349 , n380350 , n380351 , n32745 , n380353 , n380354 , n380355 , n32749 , n380357 , n380358 , 
 n380359 , n32753 , n380361 , n380362 , n32756 , n380364 , n380365 , n380366 , n32760 , n380368 , 
 n380369 , n32763 , n380371 , n380372 , n380373 , n32767 , n32768 , n380376 , n380377 , n32771 , 
 n32772 , n380380 , n380381 , n32775 , n380383 , n380384 , n32778 , n380386 , n380387 , n380388 , 
 n380389 , n32783 , n380391 , n380392 , n32786 , n380394 , n32788 , n32789 , n32790 , n32791 , 
 n32792 , n380400 , n32794 , n32795 , n380403 , n380404 , n32798 , n380406 , n380407 , n32801 , 
 n380409 , n380410 , n32804 , n32805 , n32806 , n380414 , n380415 , n32809 , n32810 , n32811 , 
 n380419 , n32813 , n380421 , n380422 , n380423 , n32817 , n380425 , n380426 , n32820 , n380428 , 
 n32822 , n380430 , n32824 , n32825 , n380433 , n32827 , n380435 , n32829 , n32830 , n380438 , 
 n380439 , n32833 , n380441 , n380442 , n32836 , n380444 , n380445 , n380446 , n32840 , n380448 , 
 n380449 , n32843 , n380451 , n380452 , n32846 , n32847 , n32848 , n380456 , n380457 , n32851 , 
 n32852 , n32853 , n380461 , n380462 , n32856 , n32857 , n32858 , n380466 , n380467 , n32861 , 
 n32862 , n380470 , n380471 , n32865 , n380473 , n32867 , n380475 , n32869 , n32870 , n380478 , 
 n32872 , n380480 , n32874 , n32875 , n380483 , n380484 , n32878 , n380486 , n380487 , n32881 , 
 n380489 , n380490 , n380491 , n32885 , n380493 , n380494 , n32888 , n380496 , n380497 , n380498 , 
 n32892 , n380500 , n32894 , n32895 , n380503 , n32897 , n380505 , n32899 , n32900 , n380508 , 
 n380509 , n32903 , n380511 , n380512 , n32906 , n380514 , n380515 , n380516 , n32910 , n380518 , 
 n380519 , n32913 , n380521 , n380522 , n32916 , n32917 , n32918 , n380526 , n380527 , n32921 , 
 n32922 , n32923 , n380531 , n380532 , n32926 , n32927 , n32928 , n380536 , n380537 , n32931 , 
 n32932 , n32933 , n380541 , n380542 , n32936 , n32937 , n32938 , n380546 , n32940 , n32941 , 
 n32942 , n32943 , n380551 , n380552 , n32946 , n32947 , n380555 , n380556 , n32950 , n32951 , 
 n32952 , n380560 , n380561 , n380562 , n32956 , n380564 , n380565 , n32959 , n32960 , n380568 , 
 n32962 , n32963 , n380571 , n380572 , n32966 , n32967 , n380575 , n380576 , n32970 , n380578 , 
 n380579 , n32973 , n380581 , n380582 , n380583 , n32977 , n380585 , n32979 , n380587 , n32981 , 
 n32982 , n380590 , n380591 , n32985 , n380593 , n380594 , n32988 , n380596 , n380597 , n32991 , 
 n32992 , n32993 , n380601 , n32995 , n380603 , n380604 , n380605 , n32999 , n380607 , n33001 , 
 n33002 , n33003 , n380611 , n380612 , n380613 , n33007 , n380615 , n380616 , n33010 , n380618 , 
 n380619 , n33013 , n380621 , n33015 , n380623 , n33017 , n33018 , n380626 , n33020 , n380628 , 
 n33022 , n33023 , n380631 , n380632 , n33026 , n380634 , n380635 , n33029 , n380637 , n380638 , 
 n380639 , n33033 , n380641 , n380642 , n33036 , n380644 , n380645 , n33039 , n33040 , n33041 , 
 n380649 , n380650 , n33044 , n380652 , n380653 , n33047 , n380655 , n33049 , n33050 , n380658 , 
 n33052 , n380660 , n33054 , n33055 , n380663 , n380664 , n33058 , n380666 , n380667 , n33061 , 
 n380669 , n380670 , n380671 , n33065 , n380673 , n380674 , n33068 , n380676 , n380677 , n33071 , 
 n380679 , n33073 , n33074 , n33075 , n33076 , n33077 , n380685 , n33079 , n33080 , n380688 , 
 n380689 , n33083 , n380691 , n380692 , n33086 , n380694 , n380695 , n33089 , n33090 , n33091 , 
 n380699 , n380700 , n33094 , n33095 , n33096 , n380704 , n380705 , n33099 , n33100 , n33101 , 
 n380709 , n380710 , n380711 , n33105 , n33106 , n380714 , n33108 , n33109 , n380717 , n33111 , 
 n380719 , n33113 , n33114 , n380722 , n33116 , n380724 , n380725 , n380726 , n33120 , n380728 , 
 n380729 , n33123 , n380731 , n380732 , n380733 , n380734 , n33128 , n380736 , n380737 , n380738 , 
 n33132 , n380740 , n33134 , n380742 , n33136 , n33137 , n380745 , n380746 , n33140 , n380748 , 
 n380749 , n33143 , n380751 , n380752 , n33146 , n33147 , n380755 , n380756 , n33150 , n380758 , 
 n380759 , n33153 , n380761 , n380762 , n33156 , n380764 , n33158 , n380766 , n33160 , n33161 , 
 n380769 , n33163 , n380771 , n33165 , n33166 , n380774 , n380775 , n33169 , n380777 , n380778 , 
 n33172 , n380780 , n380781 , n380782 , n33176 , n380784 , n380785 , n33179 , n380787 , n380788 , 
 n33182 , n33183 , n33184 , n380792 , n380793 , n33187 , n380795 , n33189 , n380797 , n33191 , 
 n33192 , n380800 , n380801 , n33195 , n380803 , n380804 , n33198 , n380806 , n380807 , n380808 , 
 n33202 , n380810 , n33204 , n380812 , n380813 , n33207 , n380815 , n380816 , n33210 , n33211 , 
 n33212 , n380820 , n380821 , n33215 , n33216 , n33217 , n380825 , n380826 , n33220 , n33221 , 
 n33222 , n380830 , n380831 , n33225 , n33226 , n33227 , n380835 , n380836 , n33230 , n33231 , 
 n33232 , n380840 , n380841 , n33235 , n33236 , n380844 , n380845 , n33239 , n380847 , n33241 , 
 n33242 , n33243 , n33244 , n33245 , n380853 , n380854 , n33248 , n33249 , n33250 , n33251 , 
 n380859 , n380860 , n380861 , n33255 , n380863 , n33257 , n380865 , n33259 , n33260 , n380868 , 
 n380869 , n33263 , n380871 , n380872 , n33266 , n380874 , n380875 , n33269 , n33270 , n33271 , 
 n380879 , n33273 , n380881 , n380882 , n380883 , n33277 , n380885 , n33279 , n380887 , n380888 , 
 n33282 , n33283 , n380891 , n33285 , n380893 , n380894 , n33288 , n380896 , n33290 , n380898 , 
 n33292 , n33293 , n380901 , n33295 , n380903 , n33297 , n33298 , n33299 , n380907 , n380908 , 
 n33302 , n380910 , n380911 , n33305 , n380913 , n380914 , n380915 , n33309 , n380917 , n380918 , 
 n33312 , n380920 , n380921 , n33315 , n380923 , n380924 , n33318 , n380926 , n33320 , n380928 , 
 n33322 , n380930 , n33324 , n33325 , n380933 , n380934 , n33328 , n380936 , n380937 , n33331 , 
 n380939 , n380940 , n33334 , n33335 , n380943 , n380944 , n33338 , n380946 , n380947 , n33341 , 
 n380949 , n380950 , n33344 , n33345 , n33346 , n33347 , n380955 , n380956 , n33350 , n380958 , 
 n33352 , n380960 , n380961 , n33355 , n380963 , n380964 , n33358 , n380966 , n380967 , n33361 , 
 n33362 , n380970 , n380971 , n33365 , n380973 , n380974 , n33368 , n380976 , n380977 , n380978 , 
 n380979 , n33373 , n380981 , n380982 , n33376 , n380984 , n33378 , n380986 , n380987 , n33381 , 
 n380989 , n380990 , n33384 , n380992 , n380993 , n33387 , n380995 , n380996 , n33390 , n33391 , 
 n33392 , n33393 , n33394 , n381002 , n381003 , n33397 , n381005 , n33399 , n33400 , n33401 , 
 n33402 , n33403 , n381011 , n33405 , n33406 , n33407 , n381015 , n33409 , n381017 , n33411 , 
 n381019 , n33413 , n33414 , n381022 , n33416 , n381024 , n381025 , n381026 , n33420 , n381028 , 
 n381029 , n33423 , n381031 , n381032 , n33426 , n33427 , n381035 , n381036 , n33430 , n381038 , 
 n381039 , n33433 , n381041 , n381042 , n381043 , n33437 , n381045 , n33439 , n33440 , n381048 , 
 n33442 , n381050 , n33444 , n33445 , n381053 , n381054 , n33448 , n381056 , n381057 , n33451 , 
 n381059 , n381060 , n381061 , n33455 , n381063 , n381064 , n33458 , n381066 , n381067 , n33461 , 
 n33462 , n33463 , n33464 , n33465 , n381073 , n381074 , n33468 , n381076 , n381077 , n33471 , 
 n33472 , n33473 , n33474 , n381082 , n381083 , n381084 , n33478 , n381086 , n33480 , n381088 , 
 n33482 , n33483 , n381091 , n381092 , n33486 , n381094 , n381095 , n33489 , n381097 , n381098 , 
 n33492 , n33493 , n381101 , n381102 , n33496 , n381104 , n381105 , n33499 , n381107 , n381108 , 
 n33502 , n381110 , n33504 , n381112 , n33506 , n33507 , n33508 , n33509 , n33510 , n33511 , 
 n33512 , n33513 , n381121 , n33515 , n381123 , n381124 , n33518 , n381126 , n381127 , n33521 , 
 n381129 , n381130 , n33524 , n381132 , n381133 , n33527 , n33528 , n33529 , n33530 , n33531 , 
 n381139 , n381140 , n33534 , n381142 , n381143 , n33537 , n33538 , n33539 , n33540 , n33541 , 
 n381149 , n381150 , n33544 , n381152 , n33546 , n33547 , n33548 , n33549 , n381157 , n33551 , 
 n33552 , n33553 , n33554 , n381162 , n381163 , n33557 , n381165 , n381166 , n381167 , n33561 , 
 n381169 , n33563 , n381171 , n381172 , n33566 , n33567 , n381175 , n33569 , n381177 , n33571 , 
 n33572 , n381180 , n381181 , n33575 , n381183 , n381184 , n33578 , n381186 , n381187 , n33581 , 
 n381189 , n381190 , n33584 , n381192 , n33586 , n381194 , n381195 , n33589 , n381197 , n381198 , 
 n33592 , n33593 , n381201 , n33595 , n381203 , n33597 , n33598 , n381206 , n381207 , n33601 , 
 n381209 , n381210 , n33604 , n381212 , n381213 , n381214 , n33608 , n381216 , n381217 , n33611 , 
 n381219 , n381220 , n33614 , n33615 , n33616 , n381224 , n381225 , n381226 , n33620 , n33621 , 
 n33622 , n33623 , n33624 , n381232 , n33626 , n33627 , n381235 , n381236 , n33630 , n381238 , 
 n381239 , n33633 , n381241 , n381242 , n381243 , n33637 , n381245 , n33639 , n381247 , n33641 , 
 n33642 , n381250 , n33644 , n381252 , n381253 , n381254 , n33648 , n381256 , n381257 , n33651 , 
 n381259 , n381260 , n33654 , n33655 , n381263 , n33657 , n381265 , n33659 , n33660 , n381268 , 
 n381269 , n33663 , n381271 , n381272 , n33666 , n381274 , n381275 , n381276 , n33670 , n381278 , 
 n381279 , n33673 , n381281 , n381282 , n33676 , n381284 , n381285 , n33679 , n381287 , n381288 , 
 n33682 , n381290 , n381291 , n33685 , n381293 , n33687 , n381295 , n33689 , n33690 , n33691 , 
 n33692 , n33693 , n381301 , n381302 , n33696 , n381304 , n33698 , n33699 , n381307 , n33701 , 
 n381309 , n381310 , n381311 , n381312 , n33706 , n381314 , n381315 , n33709 , n381317 , n381318 , 
 n33712 , n33713 , n33714 , n381322 , n381323 , n33717 , n33718 , n33719 , n381327 , n381328 , 
 n33722 , n381330 , n33724 , n381332 , n33726 , n381334 , n33728 , n33729 , n33730 , n381338 , 
 n381339 , n381340 , n33734 , n381342 , n381343 , n33737 , n381345 , n381346 , n381347 , n33741 , 
 n381349 , n33743 , n33744 , n381352 , n381353 , n33747 , n381355 , n381356 , n33750 , n381358 , 
 n33752 , n33753 , n33754 , n33755 , n33756 , n33757 , n381365 , n33759 , n381367 , n33761 , 
 n381369 , n33763 , n381371 , n33765 , n33766 , n381374 , n381375 , n33769 , n381377 , n381378 , 
 n33772 , n381380 , n381381 , n33775 , n33776 , n381384 , n381385 , n33779 , n381387 , n381388 , 
 n33782 , n381390 , n381391 , n33785 , n33786 , n33787 , n381395 , n381396 , n33790 , n33791 , 
 n381399 , n381400 , n33794 , n381402 , n33796 , n381404 , n381405 , n381406 , n33800 , n381408 , 
 n33802 , n33803 , n381411 , n381412 , n33806 , n381414 , n381415 , n33809 , n381417 , n381418 , 
 n33812 , n381420 , n381421 , n33815 , n381423 , n33817 , n381425 , n381426 , n33820 , n381428 , 
 n381429 , n33823 , n33824 , n33825 , n381433 , n381434 , n33828 , n33829 , n33830 , n381438 , 
 n381439 , n33833 , n33834 , n33835 , n381443 , n381444 , n33838 , n33839 , n33840 , n381448 , 
 n33842 , n33843 , n33844 , n33845 , n33846 , n33847 , n381455 , n33849 , n33850 , n33851 , 
 n33852 , n381460 , n381461 , n33855 , n33856 , n381464 , n381465 , n33859 , n33860 , n33861 , 
 n33862 , n381470 , n381471 , n33865 , n381473 , n33867 , n33868 , n33869 , n381477 , n381478 , 
 n33872 , n381480 , n33874 , n381482 , n33876 , n381484 , n33878 , n381486 , n33880 , n33881 , 
 n381489 , n381490 , n33884 , n381492 , n381493 , n33887 , n381495 , n381496 , n33890 , n381498 , 
 n381499 , n33893 , n381501 , n381502 , n33896 , n33897 , n33898 , n33899 , n33900 , n381508 , 
 n381509 , n33903 , n381511 , n33905 , n381513 , n33907 , n33908 , n33909 , n33910 , n381518 , 
 n381519 , n33913 , n33914 , n33915 , n33916 , n381524 , n381525 , n33919 , n33920 , n381528 , 
 n381529 , n33923 , n33924 , n33925 , n33926 , n33927 , n381535 , n381536 , n33930 , n381538 , 
 n381539 , n33933 , n381541 , n381542 , n33936 , n381544 , n381545 , n33939 , n33940 , n33941 , 
 n33942 , n381550 , n33944 , n33945 , n381553 , n33947 , n381555 , n33949 , n381557 , n33951 , 
 n381559 , n33953 , n381561 , n33955 , n33956 , n33957 , n381565 , n381566 , n33960 , n33961 , 
 n381569 , n381570 , n33964 , n33965 , n381573 , n381574 , n33968 , n33969 , n33970 , n381578 , 
 n381579 , n33973 , n33974 , n381582 , n381583 , n381584 , n33978 , n381586 , n33980 , n33981 , 
 n381589 , n33983 , n381591 , n33985 , n33986 , n381594 , n381595 , n33989 , n381597 , n381598 , 
 n33992 , n381600 , n381601 , n381602 , n33996 , n381604 , n381605 , n33999 , n381607 , n381608 , 
 n34002 , n381610 , n34004 , n381612 , n34006 , n381614 , n34008 , n34009 , n381617 , n381618 , 
 n34012 , n381620 , n381621 , n34015 , n381623 , n381624 , n34018 , n34019 , n381627 , n381628 , 
 n34022 , n381630 , n381631 , n34025 , n381633 , n381634 , n381635 , n34029 , n34030 , n34031 , 
 n34032 , n34033 , n381641 , n34035 , n34036 , n381644 , n381645 , n34039 , n381647 , n381648 , 
 n34042 , n381650 , n381651 , n34045 , n381653 , n34047 , n381655 , n34049 , n381657 , n34051 , 
 n34052 , n381660 , n381661 , n34055 , n381663 , n381664 , n34058 , n381666 , n381667 , n34061 , 
 n34062 , n381670 , n381671 , n34065 , n381673 , n381674 , n34068 , n381676 , n381677 , n34071 , 
 n34072 , n34073 , n381681 , n381682 , n34076 , n34077 , n34078 , n381686 , n381687 , n34081 , 
 n34082 , n34083 , n381691 , n381692 , n381693 , n381694 , n34088 , n381696 , n381697 , n381698 , 
 n34092 , n381700 , n34094 , n34095 , n34096 , n34097 , n34098 , n34099 , n34100 , n381708 , 
 n34102 , n381710 , n381711 , n34105 , n34106 , n34107 , n34108 , n34109 , n34110 , n381718 , 
 n34112 , n34113 , n34114 , n381722 , n381723 , n381724 , n34118 , n381726 , n34120 , n34121 , 
 n34122 , n34123 , n34124 , n34125 , n381733 , n381734 , n34128 , n381736 , n381737 , n34131 , 
 n381739 , n381740 , n34134 , n381742 , n34136 , n381744 , n34138 , n34139 , n381747 , n34141 , 
 n381749 , n34143 , n34144 , n381752 , n381753 , n34147 , n34148 , n381756 , n381757 , n34151 , 
 n381759 , n381760 , n34154 , n34155 , n34156 , n381764 , n381765 , n34159 , n34160 , n34161 , 
 n381769 , n381770 , n34164 , n34165 , n34166 , n381774 , n381775 , n34169 , n34170 , n34171 , 
 n381779 , n381780 , n34174 , n34175 , n34176 , n381784 , n381785 , n34179 , n381787 , n381788 , 
 n34182 , n34183 , n381791 , n381792 , n34186 , n34187 , n381795 , n381796 , n34190 , n34191 , 
 n381799 , n381800 , n34194 , n34195 , n34196 , n381804 , n381805 , n381806 , n34200 , n381808 , 
 n381809 , n34203 , n34204 , n381812 , n34206 , n34207 , n381815 , n381816 , n34210 , n34211 , 
 n381819 , n381820 , n34214 , n381822 , n381823 , n34217 , n381825 , n381826 , n34220 , n381828 , 
 n34222 , n381830 , n34224 , n34225 , n381833 , n381834 , n34228 , n381836 , n381837 , n34231 , 
 n381839 , n381840 , n381841 , n34235 , n381843 , n34237 , n34238 , n34239 , n381847 , n34241 , 
 n381849 , n381850 , n34244 , n381852 , n34246 , n381854 , n34248 , n34249 , n381857 , n381858 , 
 n34252 , n381860 , n381861 , n34255 , n381863 , n381864 , n34258 , n34259 , n34260 , n381868 , 
 n381869 , n34263 , n34264 , n34265 , n381873 , n381874 , n34268 , n34269 , n381877 , n381878 , 
 n34272 , n34273 , n34274 , n381882 , n381883 , n381884 , n34278 , n381886 , n381887 , n34281 , 
 n34282 , n381890 , n34284 , n34285 , n381893 , n381894 , n34288 , n34289 , n381897 , n381898 , 
 n34292 , n381900 , n381901 , n34295 , n34296 , n381904 , n381905 , n34299 , n381907 , n381908 , 
 n34302 , n34303 , n381911 , n381912 , n34306 , n381914 , n34308 , n381916 , n34310 , n34311 , 
 n381919 , n381920 , n34314 , n381922 , n381923 , n34317 , n381925 , n381926 , n34320 , n34321 , 
 n34322 , n381930 , n381931 , n34325 , n34326 , n34327 , n381935 , n381936 , n34330 , n34331 , 
 n381939 , n381940 , n381941 , n34335 , n34336 , n34337 , n381945 , n381946 , n34340 , n34341 , 
 n34342 , n381950 , n381951 , n34345 , n381953 , n381954 , n34348 , n381956 , n34350 , n34351 , 
 n34352 , n381960 , n381961 , n34355 , n34356 , n381964 , n381965 , n34359 , n34360 , n381968 , 
 n381969 , n34363 , n34364 , n34365 , n34366 , n34367 , n381975 , n381976 , n34370 , n34371 , 
 n34372 , n34373 , n381981 , n381982 , n34376 , n381984 , n34378 , n381986 , n34380 , n34381 , 
 n381989 , n34383 , n381991 , n34385 , n381993 , n381994 , n34388 , n381996 , n381997 , n34391 , 
 n34392 , n34393 , n382001 , n382002 , n34396 , n34397 , n382005 , n382006 , n34400 , n34401 , 
 n34402 , n382010 , n382011 , n34405 , n34406 , n34407 , n34408 , n382016 , n382017 , n34411 , 
 n34412 , n34413 , n382021 , n382022 , n34416 , n34417 , n34418 , n382026 , n382027 , n34421 , 
 n34422 , n34423 , n382031 , n382032 , n34426 , n34427 , n34428 , n382036 , n382037 , n34431 , 
 n382039 , n382040 , n34434 , n34435 , n382043 , n382044 , n34438 , n34439 , n382047 , n382048 , 
 n34442 , n34443 , n34444 , n34445 , n382053 , n382054 , n34448 , n34449 , n382057 , n382058 , 
 n34452 , n34453 , n34454 , n34455 , n34456 , n382064 , n382065 , n34459 , n34460 , n34461 , 
 n382069 , n382070 , n34464 , n34465 , n34466 , n382074 , n382075 , n34469 , n34470 , n34471 , 
 n382079 , n382080 , n34474 , n382082 , n382083 , n34477 , n382085 , n382086 , n34480 , n382088 , 
 n382089 , n34483 , n382091 , n34485 , n34486 , n382094 , n382095 , n34489 , n382097 , n382098 , 
 n34492 , n34493 , n382101 , n34495 , n34496 , n382104 , n382105 , n34499 , n382107 , n382108 , 
 n34502 , n382110 , n34504 , n34505 , n34506 , n382114 , n382115 , n34509 , n382117 , n34511 , 
 n34512 , n34513 , n34514 , n382122 , n382123 , n34517 , n34518 , n382126 , n382127 , n34521 , 
 n34522 , n34523 , n34524 , n34525 , n382133 , n382134 , n34528 , n382136 , n382137 , n34531 , 
 n382139 , n382140 , n34534 , n34535 , n34536 , n34537 , n382145 , n382146 , n34540 , n382148 , 
 n382149 , n34543 , n382151 , n34545 , n34546 , n382154 , n382155 , n34549 , n34550 , n34551 , 
 n34552 , n34553 , n382161 , n382162 , n34556 , n382164 , n382165 , n34559 , n382167 , n34561 , 
 n34562 , n34563 , n34564 , n34565 , n382173 , n382174 , n34568 , n382176 , n34570 , n34571 , 
 n382179 , n382180 , n34574 , n382182 , n382183 , n382184 , n34578 , n382186 , n34580 , n34581 , 
 n382189 , n382190 , n34584 , n382192 , n382193 , n382194 , n382195 , n34589 , n382197 , n382198 , 
 n34592 , n382200 , n34594 , n34595 , n34596 , n34597 , n34598 , n34599 , n382207 , n34601 , 
 n382209 , n34603 , n34604 , n34605 , n34606 , n34607 , n34608 , n382216 , n382217 , n34611 , 
 n382219 , n34613 , n382221 , n382222 , n34616 , n382224 , n34618 , n34619 , n34620 , n382228 , 
 n34622 , n382230 , n34624 , n34625 , n34626 , n34627 , n34628 , n34629 , n34630 , n34631 , 
 n34632 , n34633 , n34634 , n34635 , n34636 , n34637 , n34638 , n34639 , n34640 , n382248 , 
 n34642 , n382250 , n34644 , n34645 , n34646 , n34647 , n34648 , n34649 , n34650 , n34651 , 
 n34652 , n34653 , n34654 , n34655 , n34656 , n34657 , n382265 , n34659 , n382267 , n34661 , 
 n382269 , n382270 , n34664 , n382272 , n382273 , n34667 , n34668 , n382276 , n34670 , n382278 , 
 n34672 , n34673 , n382281 , n382282 , n34676 , n382284 , n382285 , n34679 , n382287 , n382288 , 
 n382289 , n34683 , n382291 , n382292 , n34686 , n382294 , n382295 , n382296 , n382297 , n34691 , 
 n382299 , n382300 , n34694 , n382302 , n34696 , n382304 , n34698 , n34699 , n382307 , n34701 , 
 n382309 , n382310 , n34704 , n382312 , n382313 , n34707 , n382315 , n34709 , n382317 , n34711 , 
 n34712 , n382320 , n382321 , n34715 , n382323 , n382324 , n34718 , n382326 , n382327 , n34721 , 
 n34722 , n34723 , n382331 , n382332 , n34726 , n34727 , n34728 , n382336 , n382337 , n34731 , 
 n382339 , n34733 , n382341 , n382342 , n34736 , n34737 , n382345 , n34739 , n382347 , n382348 , 
 n34742 , n382350 , n382351 , n34745 , n382353 , n34747 , n382355 , n382356 , n34750 , n382358 , 
 n34752 , n34753 , n382361 , n34755 , n34756 , n34757 , n34758 , n382366 , n382367 , n382368 , 
 n34763 , n382370 , n382371 , n382372 , n34769 , n382374 , n382375 , n34772 , n382377 , n34774 , 
 n382379 , n382380 , n34777 , n34778 , n382383 , n382384 , n34781 , n34782 , n34783 , n34784 , 
 n34785 , n382390 , n382391 , n34788 , n382393 , n34790 , n34791 , n34792 , n34793 , n382398 , 
 n34795 , n382400 , n34797 , n34798 , n34799 , n34800 , n382405 , n382406 , n34803 , n34804 , 
 n382409 , n382410 , n34807 , n382412 , n382413 , n34810 , n382415 , n382416 , n34813 , n382418 , 
 n382419 , n34816 , n382421 , n382422 , n34819 , n34820 , n34821 , n382426 , n382427 , n34824 , 
 n382429 , n382430 , n382431 , n382432 , n34829 , n382434 , n382435 , n34832 , n382437 , n382438 , 
 n34835 , n382440 , n382441 , n34838 , n382443 , n34840 , n34841 , n382446 , n34843 , n34844 , 
 n382449 , n382450 , n34847 , n382452 , n382453 , n34850 , n34851 , n382456 , n34853 , n382458 , 
 n382459 , n34856 , n382461 , n34858 , n34859 , n34860 , n34861 , n34862 , n34863 , n382468 , 
 n34865 , n34866 , n382471 , n34868 , n382473 , n382474 , n382475 , n34872 , n382477 , n382478 , 
 n34875 , n382480 , n382481 , n34878 , n34879 , n382484 , n34881 , n34882 , n34883 , n34884 , 
 n382489 , n34886 , n382491 , n34888 , n34889 , n34890 , n34891 , n34892 , n34893 , n382498 , 
 n382499 , n34896 , n382501 , n34898 , n34899 , n34900 , n34901 , n34902 , n34903 , n34904 , 
 n34905 , n34906 , n34907 , n34908 , n34909 , n34910 , n34911 , n34912 , n34913 , n34914 , 
 n382519 , n382520 , n34917 , n382522 , n34919 , n382524 , n34921 , n382526 , n382527 , n34924 , 
 n382529 , n382530 , n34927 , n382532 , n382533 , n34930 , n382535 , n382536 , n34933 , n382538 , 
 n382539 , n34936 , n34937 , n382542 , n382543 , n34940 , n382545 , n382546 , n34943 , n382548 , 
 n382549 , n34946 , n382551 , n382552 , n34949 , n382554 , n382555 , n34952 , n382557 , n382558 , 
 n382559 , n382560 , n34957 , n382562 , n34959 , n34960 , n382565 , n34962 , n382567 , n382568 , 
 n34965 , n382570 , n382571 , n34968 , n382573 , n34970 , n34971 , n34972 , n34973 , n34974 , 
 n34975 , n382580 , n382581 , n34978 , n382583 , n382584 , n34981 , n382586 , n382587 , n34984 , 
 n382589 , n382590 , n34987 , n382592 , n382593 , n34990 , n382595 , n382596 , n34993 , n382598 , 
 n382599 , n34996 , n382601 , n382602 , n34999 , n382604 , n382605 , n35002 , n382607 , n382608 , 
 n35005 , n382610 , n382611 , n35008 , n382613 , n382614 , n35011 , n382616 , n35013 , n382618 , 
 n35015 , n35016 , n35017 , n35018 , n382623 , n382624 , n382625 , n35022 , n382627 , n35024 , 
 n35025 , n382630 , n35027 , n382632 , n35029 , n35030 , n382635 , n382636 , n35033 , n382638 , 
 n382639 , n35036 , n382641 , n382642 , n382643 , n35040 , n382645 , n382646 , n35043 , n382648 , 
 n382649 , n382650 , n382651 , n382652 , n382653 , n382654 , n35051 , n35052 , n35053 , n35054 , 
 n35055 , n382660 , n382661 , n35058 , n382663 , n382664 , n35061 , n382666 , n35063 , n382668 , 
 n35065 , n35066 , n35067 , n35068 , n382673 , n382674 , n382675 , n35072 , n382677 , n35074 , 
 n382679 , n382680 , n35077 , n35078 , n382683 , n35080 , n382685 , n382686 , n35083 , n382688 , 
 n382689 , n35086 , n382691 , n35088 , n382693 , n382694 , n35091 , n382696 , n382697 , n35094 , 
 n382699 , n382700 , n35097 , n382702 , n382703 , n35100 , n382705 , n382706 , n35103 , n382708 , 
 n35105 , n35106 , n35107 , n382712 , n35109 , n382714 , n35111 , n35112 , n382717 , n35114 , 
 n382719 , n35116 , n35117 , n35118 , n35119 , n35120 , n35121 , n35122 , n35123 , n35124 , 
 n35125 , n35126 , n35127 , n35128 , n382733 , n35130 , n382735 , n382736 , n35133 , n382738 , 
 n382739 , n35136 , n382741 , n35138 , n382743 , n382744 , n382745 , n35142 , n382747 , n382748 , 
 n35145 , n382750 , n382751 , n35148 , n382753 , n382754 , n35151 , n382756 , n382757 , n35154 , 
 n382759 , n382760 , n35157 , n35158 , n382763 , n382764 , n35161 , n382766 , n382767 , n35164 , 
 n382769 , n35166 , n35167 , n35168 , n35169 , n382774 , n382775 , n382776 , n35173 , n382778 , 
 n35175 , n382780 , n382781 , n35178 , n382783 , n35180 , n382785 , n382786 , n35183 , n382788 , 
 n35185 , n35186 , n35187 , n35188 , n35189 , n35190 , n35191 , n35192 , n382797 , n35194 , 
 n382799 , n35196 , n382801 , n382802 , n35199 , n382804 , n35201 , n35202 , n382807 , n35204 , 
 n382809 , n382810 , n35207 , n382812 , n382813 , n382814 , n35211 , n382816 , n382817 , n35214 , 
 n382819 , n35216 , n35217 , n35218 , n35219 , n382824 , n35221 , n382826 , n35223 , n35224 , 
 n35225 , n35226 , n35227 , n35231 , n35232 , n35233 , n35234 , n382836 , n35236 , n382838 , 
 n35238 , n35239 , n382841 , n35241 , n382843 , n382844 , n382845 , n35245 , n382847 , n35247 , 
 n382849 , n35249 , n35262 , n382852 , n35264 , n382854 , n382855 , n35267 , n382857 , n382858 , 
 n35270 , n35271 , n35272 , n382862 , n35274 , n382864 , n382865 , n35277 , n382867 , n35279 , 
 n35280 , n35281 , n35282 , n35283 , n35284 , n35285 , n35286 , n382876 , n35288 , n382878 , 
 n35290 , n35291 , n35292 , n35293 , n35294 , n35295 , n35296 , n35297 , n35298 , n35299 , 
 n35300 , n35301 , n382891 , n35303 , n382893 , n382894 , n35306 , n382896 , n382897 , n35309 , 
 n35310 , n382900 , n382901 , n35313 , n382903 , n382904 , n35316 , n382906 , n382907 , n35319 , 
 n382909 , n382910 , n35325 , n35326 , n35327 , n35328 , n35329 , n35330 , n35331 , n35332 , 
 n382919 , n35334 , n382921 , n382922 , n35337 , n382924 , n382925 , n35340 , n35341 , n382928 , 
 n382929 , n35344 , n382931 , n382932 , n35347 , n382934 , n382935 , n382936 , n35351 , n382938 , 
 n382939 , n35354 , n382941 , n382942 , n35357 , n382944 , n382945 , n35360 , n382947 , n382948 , 
 n35363 , n382950 , n382951 , n35366 , n382953 , n382954 , n35369 , n382956 , n382957 , n35372 , 
 n382959 , n382960 , n35375 , n35376 , n35377 , n35378 , n35379 , n35380 , n35381 , n382968 , 
 n382969 , n35384 , n382971 , n382972 , n35387 , n382974 , n35389 , n35390 , n35391 , n35392 , 
 n382979 , n35394 , n382981 , n382982 , n35397 , n382984 , n35399 , n35400 , n382987 , n35402 , 
 n382989 , n35404 , n35405 , n382992 , n35407 , n382994 , n382995 , n382996 , n382997 , n35412 , 
 n35413 , n383000 , n35415 , n35416 , n383003 , n383004 , n35419 , n35420 , n383007 , n35422 , 
 n35423 , n383010 , n35425 , n383012 , n35427 , n383014 , n383015 , n35430 , n383017 , n35432 , 
 n383019 , n35434 , n35435 , n383022 , n35437 , n383024 , n383025 , n35440 , n383027 , n383028 , 
 n35443 , n35444 , n35445 , n383032 , n35447 , n383034 , n35449 , n383036 , n35451 , n35452 , 
 n35453 , n35454 , n35455 , n35456 , n35457 , n35458 , n35459 , n35460 , n35461 , n35462 , 
 n35463 , n35464 , n383051 , n35466 , n383053 , n383054 , n35469 , n383056 , n383057 , n35472 , 
 n383059 , n383060 , n35475 , n383062 , n383063 , n35478 , n35479 , n383066 , n35481 , n383068 , 
 n383069 , n383070 , n35485 , n383072 , n383073 , n35488 , n383075 , n383076 , n35491 , n383078 , 
 n383079 , n35494 , n35495 , n383082 , n35497 , n35498 , n35499 , n35500 , n35501 , n383088 , 
 n35503 , n383090 , n35505 , n383092 , n383093 , n35508 , n383095 , n35510 , n383097 , n35512 , 
 n35513 , n35514 , n35515 , n35516 , n35517 , n35518 , n35519 , n383106 , n35521 , n383108 , 
 n383109 , n35524 , n383111 , n383112 , n35527 , n383114 , n383115 , n35530 , n383117 , n383118 , 
 n35533 , n35534 , n383121 , n35536 , n383123 , n383124 , n383125 , n35540 , n383127 , n383128 , 
 n35543 , n383130 , n383131 , n383132 , n35547 , n383134 , n383135 , n35550 , n383137 , n383138 , 
 n35553 , n383140 , n383141 , n35556 , n383143 , n383144 , n35559 , n383146 , n383147 , n383148 , 
 n383149 , n35564 , n383151 , n383152 , n35567 , n383154 , n383155 , n35570 , n383157 , n383158 , 
 n35573 , n383160 , n383161 , n383162 , n35577 , n383164 , n35579 , n383166 , n35581 , n383168 , 
 n35583 , n35584 , n383171 , n383172 , n35587 , n383174 , n383175 , n35590 , n383177 , n383178 , 
 n35593 , n383180 , n35595 , n383182 , n383183 , n35598 , n383185 , n383186 , n383187 , n35602 , 
 n383189 , n35604 , n35605 , n383192 , n383193 , n35608 , n35609 , n383196 , n383197 , n383198 , 
 n35613 , n383200 , n383201 , n35616 , n383203 , n383204 , n35619 , n383206 , n383207 , n383208 , 
 n383209 , n35626 , n383211 , n383212 , n383213 , n35636 , n35637 , n383216 , n35639 , n35640 , 
 n383219 , n383220 , n383221 , n35644 , n383223 , n383224 , n35647 , n383226 , n383227 , n35650 , 
 n383229 , n35652 , n383231 , n35654 , n35655 , n383234 , n383235 , n35658 , n383237 , n383238 , 
 n35661 , n383240 , n383241 , n35664 , n383243 , n35666 , n383245 , n383246 , n35669 , n383248 , 
 n35671 , n35672 , n383251 , n35674 , n383253 , n383254 , n35677 , n383256 , n383257 , n35680 , 
 n383259 , n383260 , n35683 , n383262 , n35685 , n383264 , n35687 , n383266 , n383267 , n35690 , 
 n35691 , n35695 , n383271 , n383272 , n35698 , n383274 , n383275 , n35701 , n35702 , n383278 , 
 n383279 , n35705 , n383281 , n383282 , n35708 , n383284 , n383285 , n35711 , n383287 , n35713 , 
 n383289 , n35715 , n383291 , n35717 , n35718 , n383294 , n35720 , n383296 , n35722 , n383298 , 
 n35724 , n35725 , n383301 , n383302 , n35728 , n35729 , n383305 , n383306 , n35732 , n35733 , 
 n383309 , n383310 , n35736 , n35737 , n383313 , n383314 , n35740 , n383316 , n383317 , n35743 , 
 n383319 , n35745 , n35746 , n383322 , n35748 , n35749 , n383325 , n383326 , n35752 , n383328 , 
 n383329 , n35755 , n383331 , n383332 , n383333 , n35759 , n383335 , n383336 , n383337 , n35763 , 
 n383339 , n35765 , n35766 , n383342 , n35768 , n383344 , n35770 , n35771 , n383347 , n383348 , 
 n35774 , n35775 , n383351 , n383352 , n35778 , n383354 , n35780 , n383356 , n383357 , n35783 , 
 n383359 , n383360 , n35786 , n35787 , n383363 , n35789 , n383365 , n35791 , n35792 , n35793 , 
 n35794 , n35795 , n35796 , n35797 , n35798 , n35799 , n35800 , n383376 , n35802 , n383378 , 
 n35804 , n383380 , n35806 , n35807 , n383383 , n35809 , n383385 , n35811 , n35812 , n383388 , 
 n35814 , n383390 , n35816 , n35817 , n35818 , n35819 , n35820 , n35821 , n35822 , n35823 , 
 n35824 , n35825 , n383401 , n35827 , n383403 , n383404 , n35830 , n383406 , n383407 , n35833 , 
 n383409 , n383410 , n35836 , n383412 , n35838 , n383414 , n383415 , n35841 , n383417 , n383418 , 
 n35844 , n383420 , n383421 , n35847 , n383423 , n383424 , n35850 , n383426 , n383427 , n35853 , 
 n383429 , n35855 , n35856 , n35857 , n35858 , n383434 , n35860 , n35861 , n383437 , n35863 , 
 n383439 , n35865 , n35866 , n383442 , n383443 , n35869 , n383445 , n383446 , n35872 , n383448 , 
 n383449 , n35875 , n383451 , n383452 , n383453 , n383454 , n383455 , n35881 , n35882 , n383458 , 
 n35884 , n383460 , n383461 , n35887 , n35888 , n383464 , n383465 , n35891 , n383467 , n383468 , 
 n35894 , n383470 , n383471 , n35897 , n383473 , n383474 , n35900 , n383476 , n383477 , n35903 , 
 n383479 , n383480 , n35906 , n383482 , n383483 , n35909 , n383485 , n383486 , n35912 , n383488 , 
 n383489 , n35915 , n35916 , n383492 , n383493 , n35919 , n383495 , n383496 , n383497 , n35923 , 
 n383499 , n383500 , n35926 , n383502 , n383503 , n35929 , n383505 , n383506 , n35932 , n383508 , 
 n383509 , n35935 , n383511 , n383512 , n35938 , n383514 , n383515 , n383516 , n35942 , n383518 , 
 n35944 , n35945 , n383521 , n383522 , n35948 , n35949 , n383525 , n35951 , n35952 , n35953 , 
 n35954 , n383530 , n35956 , n383532 , n35958 , n383534 , n35960 , n383536 , n35962 , n35963 , 
 n383539 , n383540 , n35966 , n383542 , n383543 , n35969 , n383545 , n383546 , n35972 , n35973 , 
 n383549 , n383550 , n35976 , n383552 , n383553 , n35979 , n383555 , n383556 , n35982 , n35983 , 
 n383559 , n35985 , n35986 , n35987 , n35988 , n35989 , n35990 , n35991 , n35992 , n35993 , 
 n35994 , n35995 , n35996 , n35997 , n383573 , n35999 , n383575 , n383576 , n36002 , n383578 , 
 n383579 , n36005 , n36006 , n383582 , n36008 , n383584 , n383585 , n383586 , n36012 , n383588 , 
 n383589 , n36015 , n383591 , n36018 , n383593 , n36020 , n383595 , n383596 , n36023 , n36024 , 
 n36025 , n36026 , n383601 , n36028 , n383603 , n36030 , n36031 , n383606 , n383607 , n36034 , 
 n383609 , n383610 , n36037 , n383612 , n36039 , n36040 , n383615 , n36042 , n383617 , n383618 , 
 n36045 , n383620 , n36047 , n383622 , n36049 , n36050 , n383625 , n36052 , n36053 , n36054 , 
 n36055 , n36056 , n36057 , n36058 , n36059 , n36060 , n36061 , n36062 , n36063 , n36064 , 
 n36065 , n36066 , n36067 , n36068 , n36069 , n383644 , n36071 , n36072 , n36073 , n383648 , 
 n383649 , n36076 , n383651 , n383652 , n36079 , n383654 , n383655 , n383656 , n36086 , n383658 , 
 n383659 , n36089 , n36090 , n383662 , n36092 , n383664 , n383665 , n383666 , n36096 , n383668 , 
 n383669 , n383670 , n36100 , n383672 , n36102 , n383674 , n36104 , n36105 , n383677 , n383678 , 
 n36108 , n383680 , n383681 , n36111 , n383683 , n383684 , n36114 , n36115 , n383687 , n383688 , 
 n36118 , n383690 , n383691 , n36121 , n383693 , n383694 , n36124 , n383696 , n383697 , n36127 , 
 n383699 , n383700 , n36130 , n36131 , n383703 , n36133 , n383705 , n36135 , n383707 , n383708 , 
 n36138 , n383710 , n383711 , n36141 , n36142 , n36143 , n383715 , n36145 , n383717 , n36147 , 
 n383719 , n36149 , n36150 , n383722 , n383723 , n36153 , n383725 , n383726 , n36156 , n383728 , 
 n383729 , n383730 , n36160 , n36161 , n383733 , n36163 , n36164 , n383736 , n36166 , n36167 , 
 n383739 , n383740 , n36170 , n383742 , n36172 , n36173 , n36174 , n383746 , n383747 , n36177 , 
 n383749 , n36179 , n36180 , n36181 , n36182 , n36183 , n36184 , n36185 , n36186 , n36187 , 
 n36188 , n383760 , n36190 , n383762 , n383763 , n36193 , n383765 , n383766 , n36196 , n36197 , 
 n383769 , n36199 , n36200 , n383772 , n36202 , n36203 , n383775 , n36205 , n383777 , n383778 , 
 n383779 , n36209 , n383781 , n36211 , n36212 , n36213 , n36214 , n36215 , n36216 , n36217 , 
 n36218 , n36219 , n36220 , n36221 , n36222 , n36223 , n36224 , n36225 , n36226 , n36227 , 
 n36228 , n383800 , n383801 , n36231 , n383803 , n36233 , n383805 , n383806 , n36236 , n383808 , 
 n36238 , n36239 , n36240 , n36241 , n36242 , n36243 , n36244 , n36245 , n36246 , n36247 , 
 n36248 , n36249 , n36250 , n36251 , n36252 , n36253 , n36254 , n36255 , n36256 , n36257 , 
 n36258 , n36259 , n383831 , n36261 , n383833 , n36263 , n383835 , n383836 , n383837 , n36267 , 
 n383839 , n383840 , n36270 , n383842 , n36272 , n36273 , n36274 , n383846 , n383847 , n36277 , 
 n383849 , n36279 , n383851 , n36281 , n383853 , n383854 , n36284 , n383856 , n383857 , n36287 , 
 n383859 , n36289 , n383861 , n36291 , n383863 , n383864 , n36294 , n383866 , n36296 , n36297 , 
 n36298 , n36299 , n36300 , n36301 , n36302 , n36303 , n36304 , n36305 , n36306 , n36307 , 
 n36308 , n36309 , n36310 , n383882 , n36312 , n383884 , n36314 , n383886 , n36316 , n36317 , 
 n383889 , n36319 , n383891 , n383892 , n36322 , n383894 , n383895 , n36325 , n383897 , n383898 , 
 n36328 , n383900 , n36330 , n383902 , n36332 , n383904 , n383905 , n36335 , n383907 , n383908 , 
 n36338 , n383910 , n36340 , n36341 , n383913 , n36343 , n383915 , n36345 , n36346 , n36347 , 
 n36348 , n36349 , n36350 , n36351 , n36352 , n36353 , n36354 , n36355 , n36356 , n36357 , 
 n36358 , n36359 , n36360 , n36361 , n36362 , n36363 , n383935 , n36365 , n383937 , n383938 , 
 n36368 , n383940 , n383941 , n36371 , n383943 , n383944 , n36374 , n383946 , n36376 , n36377 , 
 n383949 , n36379 , n383951 , n36381 , n383953 , n36383 , n383955 , n36385 , n383957 , n36387 , 
 n36388 , n383960 , n383961 , n36391 , n383963 , n36393 , n36394 , n36395 , n36396 , n36397 , 
 n36398 , n36399 , n36400 , n36401 , n383973 , n36403 , n383975 , n36405 , n36406 , n36407 , 
 n36408 , n383980 , n36410 , n383982 , n36412 , n36413 , n383985 , n383986 , n36416 , n383988 , 
 n383989 , n36419 , n383991 , n383992 , n36422 , n36423 , n36424 , n36425 , n36426 , n36427 , 
 n36428 , n36429 , n384001 , n36431 , n384003 , n36433 , n36434 , n384006 , n36436 , n384008 , 
 n384009 , n36439 , n384011 , n384012 , n36442 , n384014 , n36444 , n36445 , n36446 , n36447 , 
 n36448 , n36449 , n36450 , n36451 , n36452 , n36453 , n36454 , n36455 , n36456 , n384028 , 
 n36458 , n384030 , n36460 , n384032 , n384033 , n36463 , n384035 , n36465 , n384037 , n384038 , 
 n36468 , n384040 , n36470 , n384042 , n384043 , n36473 , n384045 , n384046 , n36476 , n36477 , 
 n384049 , n384050 , n36480 , n384052 , n384053 , n36483 , n384055 , n384056 , n36486 , n384058 , 
 n36488 , n384060 , n384061 , n36491 , n384063 , n384064 , n36494 , n384066 , n36496 , n384068 , 
 n384069 , n36499 , n384071 , n384072 , n36502 , n384074 , n36504 , n36505 , n36506 , n36507 , 
 n36508 , n36509 , n384081 , n36511 , n384083 , n384084 , n36514 , n36515 , n384087 , n36517 , 
 n384089 , n384090 , n36520 , n384092 , n384093 , n384094 , n36524 , n384096 , n384097 , n36527 , 
 n384099 , n384100 , n36530 , n384102 , n36532 , n36533 , n384105 , n36535 , n384107 , n36537 , 
 n384109 , n36539 , n384111 , n36541 , n384113 , n36543 , n384115 , n36545 , n36546 , n36547 , 
 n36548 , n384120 , n384121 , n36551 , n384123 , n36553 , n36554 , n36555 , n36556 , n36557 , 
 n36558 , n36559 , n36560 , n36561 , n36562 , n36563 , n36564 , n36565 , n384137 , n36567 , 
 n36568 , n384140 , n384141 , n36571 , n384143 , n384144 , n36574 , n384146 , n384147 , n36577 , 
 n384149 , n384150 , n36583 , n384152 , n384153 , n36586 , n36587 , n36588 , n36589 , n36590 , 
 n36591 , n36592 , n36593 , n36594 , n36595 , n36596 , n36597 , n36598 , n36599 , n36600 , 
 n36601 , n36602 , n384171 , n36604 , n36605 , n36606 , n384175 , n36608 , n384177 , n384178 , 
 n36611 , n384180 , n384181 , n36614 , n384183 , n384184 , n36617 , n384186 , n384187 , n36620 , 
 n384189 , n384190 , n36623 , n384192 , n36625 , n36626 , n384195 , n36628 , n384197 , n36630 , 
 n384199 , n384200 , n36633 , n384202 , n384203 , n36636 , n384205 , n384206 , n36639 , n384208 , 
 n384209 , n36642 , n384211 , n384212 , n384213 , n36646 , n384215 , n36648 , n384217 , n36650 , 
 n36651 , n384220 , n384221 , n36654 , n36655 , n36656 , n36657 , n36658 , n36659 , n36660 , 
 n36661 , n36662 , n36663 , n36664 , n36665 , n36666 , n36667 , n36668 , n384237 , n36670 , 
 n384239 , n36672 , n384241 , n36674 , n36675 , n36676 , n384245 , n384246 , n36679 , n384248 , 
 n384249 , n36682 , n384251 , n384252 , n36685 , n384254 , n384255 , n36688 , n384257 , n384258 , 
 n36691 , n36692 , n384261 , n36694 , n36695 , n36696 , n36697 , n36698 , n36699 , n36700 , 
 n36701 , n36702 , n36703 , n36704 , n36705 , n36706 , n36707 , n36708 , n36709 , n384278 , 
 n36711 , n384280 , n384281 , n36714 , n36715 , n384284 , n36717 , n384286 , n384287 , n384288 , 
 n36721 , n384290 , n384291 , n36724 , n384293 , n36726 , n36727 , n384296 , n36732 , n384298 , 
 n36734 , n36735 , n36736 , n384302 , n36738 , n384304 , n36740 , n36741 , n36742 , n36743 , 
 n36744 , n384310 , n384311 , n36747 , n384313 , n384314 , n384315 , n36751 , n384317 , n36753 , 
 n36754 , n36755 , n36756 , n36757 , n36758 , n36759 , n36760 , n384326 , n36762 , n384328 , 
 n384329 , n36765 , n384331 , n36767 , n384333 , n36769 , n36770 , n36771 , n36772 , n36773 , 
 n36774 , n36775 , n384341 , n36777 , n384343 , n36779 , n36780 , n36781 , n36782 , n384348 , 
 n384349 , n36785 , n384351 , n36787 , n36788 , n36789 , n36790 , n36791 , n36792 , n36793 , 
 n36794 , n36795 , n36796 , n36797 , n36798 , n36799 , n36800 , n36801 , n384367 , n36803 , 
 n384369 , n384370 , n36806 , n36807 , n36808 , n36809 , n36810 , n36811 , n384377 , n36813 , 
 n384379 , n36815 , n384381 , n384382 , n36818 , n36819 , n384385 , n36821 , n36822 , n384388 , 
 n36824 , n384390 , n384391 , n36827 , n384393 , n384394 , n36830 , n36831 , n384397 , n36833 , 
 n384399 , n36835 , n36836 , n384402 , n384403 , n36839 , n384405 , n384406 , n36842 , n384408 , 
 n384409 , n36845 , n384411 , n36847 , n384413 , n384414 , n36850 , n384416 , n384417 , n36853 , 
 n384419 , n384420 , n36856 , n384422 , n384423 , n36859 , n36860 , n36861 , n384427 , n36863 , 
 n384429 , n36865 , n384431 , n36867 , n384433 , n36869 , n36870 , n384436 , n384437 , n36873 , 
 n384439 , n384440 , n36876 , n384442 , n384443 , n36879 , n36880 , n384446 , n36882 , n384448 , 
 n384449 , n36885 , n384451 , n384452 , n36888 , n384454 , n36890 , n36891 , n36892 , n384458 , 
 n384459 , n36895 , n384461 , n36897 , n36898 , n36899 , n36900 , n384466 , n36902 , n36903 , 
 n384469 , n36905 , n384471 , n384472 , n384473 , n36909 , n384475 , n384476 , n36912 , n384478 , 
 n384479 , n384480 , n36916 , n384482 , n384483 , n36919 , n384485 , n384486 , n384487 , n36923 , 
 n384489 , n36925 , n36926 , n384492 , n36928 , n384494 , n36930 , n36931 , n384497 , n384498 , 
 n36934 , n384500 , n384501 , n36937 , n384503 , n384504 , n384505 , n36941 , n384507 , n384508 , 
 n36944 , n384510 , n384511 , n36947 , n384513 , n36949 , n36950 , n36951 , n36952 , n36953 , 
 n36954 , n384520 , n384521 , n384522 , n36958 , n384524 , n384525 , n36961 , n384527 , n36963 , 
 n36964 , n36965 , n36966 , n36967 , n384533 , n36969 , n384535 , n36971 , n36972 , n36973 , 
 n36974 , n36975 , n36976 , n36977 , n384543 , n36979 , n384545 , n384546 , n36982 , n384548 , 
 n384549 , n36985 , n384551 , n384552 , n36988 , n384554 , n384555 , n36991 , n384557 , n384558 , 
 n36994 , n384560 , n36996 , n384562 , n384563 , n36999 , n384565 , n384566 , n37002 , n384568 , 
 n384569 , n37005 , n384571 , n37007 , n37008 , n384574 , n384575 , n37011 , n384577 , n384578 , 
 n37014 , n384580 , n384581 , n37017 , n384583 , n384584 , n37020 , n37021 , n384587 , n37023 , 
 n384589 , n37025 , n37026 , n37027 , n384593 , n37029 , n384595 , n37031 , n384597 , n384598 , 
 n37034 , n384600 , n384601 , n37037 , n384603 , n384604 , n37040 , n384606 , n384607 , n37043 , 
 n384609 , n384610 , n384611 , n384612 , n37048 , n384614 , n37050 , n384616 , n37052 , n384618 , 
 n384619 , n37055 , n384621 , n384622 , n37058 , n384624 , n384625 , n37061 , n384627 , n384628 , 
 n37064 , n384630 , n384631 , n37067 , n384633 , n384634 , n37070 , n384636 , n384637 , n37073 , 
 n384639 , n37075 , n384641 , n384642 , n37078 , n384644 , n384645 , n37081 , n384647 , n37083 , 
 n384649 , n37085 , n37086 , n384652 , n384653 , n37089 , n384655 , n384656 , n37092 , n384658 , 
 n384659 , n37095 , n37096 , n384662 , n37098 , n384664 , n37100 , n384666 , n37102 , n37103 , 
 n384669 , n384670 , n37106 , n384672 , n384673 , n37109 , n384675 , n384676 , n37112 , n384678 , 
 n384679 , n37115 , n384681 , n384682 , n384683 , n37119 , n384685 , n37121 , n384687 , n37123 , 
 n384689 , n37125 , n37126 , n37127 , n384693 , n37129 , n384695 , n37131 , n37132 , n37133 , 
 n384699 , n384700 , n37136 , n384702 , n37138 , n37139 , n37140 , n37141 , n37142 , n37143 , 
 n37144 , n37145 , n37146 , n37147 , n384713 , n37149 , n384715 , n384716 , n37152 , n37153 , 
 n384719 , n37155 , n384721 , n384722 , n384723 , n37159 , n384725 , n384726 , n37162 , n384728 , 
 n384729 , n37165 , n37166 , n37167 , n37168 , n37169 , n37170 , n37171 , n37172 , n37173 , 
 n384739 , n37175 , n384741 , n384742 , n37178 , n384744 , n37180 , n37181 , n37182 , n384748 , 
 n384749 , n37185 , n384751 , n384752 , n37188 , n384754 , n384755 , n37191 , n384757 , n37193 , 
 n384759 , n37195 , n384761 , n37197 , n37198 , n384764 , n384765 , n37201 , n384767 , n384768 , 
 n37204 , n384770 , n384771 , n37207 , n37208 , n384774 , n37210 , n37211 , n384777 , n37213 , 
 n37214 , n37215 , n37216 , n384782 , n384783 , n37219 , n384785 , n384786 , n37222 , n384788 , 
 n384789 , n384790 , n37226 , n384792 , n384793 , n37229 , n384795 , n384796 , n37232 , n37233 , 
 n37234 , n384800 , n384801 , n37242 , n384803 , n384804 , n37245 , n384806 , n384807 , n37248 , 
 n384809 , n384810 , n384811 , n37252 , n384813 , n37254 , n37255 , n384816 , n384817 , n37258 , 
 n384819 , n384820 , n37261 , n384822 , n384823 , n37264 , n384825 , n37266 , n384827 , n37268 , 
 n37269 , n384830 , n384831 , n37272 , n384833 , n384834 , n37275 , n384836 , n384837 , n37278 , 
 n384839 , n384840 , n37281 , n37282 , n37283 , n37284 , n384845 , n384846 , n37287 , n384848 , 
 n384849 , n37290 , n384851 , n37292 , n37293 , n37294 , n37295 , n37296 , n37297 , n37298 , 
 n37299 , n37300 , n37301 , n37302 , n37303 , n37304 , n37305 , n384866 , n37307 , n384868 , 
 n37309 , n37310 , n37311 , n37312 , n37313 , n37314 , n37315 , n37316 , n37317 , n384878 , 
 n37319 , n384880 , n37321 , n384882 , n37323 , n37324 , n384885 , n37326 , n384887 , n384888 , 
 n384889 , n37330 , n384891 , n37332 , n37333 , n37334 , n37335 , n37336 , n37337 , n37338 , 
 n384899 , n37340 , n384901 , n384902 , n37343 , n37344 , n37345 , n37346 , n37347 , n384908 , 
 n37349 , n384910 , n37351 , n37352 , n384913 , n37354 , n384915 , n37356 , n384917 , n384918 , 
 n37359 , n384920 , n384921 , n37362 , n384923 , n384924 , n384925 , n37366 , n37367 , n37368 , 
 n37369 , n37370 , n37371 , n37372 , n384933 , n37374 , n37375 , n384936 , n37377 , n384938 , 
 n37379 , n37380 , n37381 , n384942 , n384943 , n37384 , n384945 , n384946 , n37387 , n384948 , 
 n384949 , n384950 , n37391 , n384952 , n384953 , n37394 , n384955 , n384956 , n37397 , n37398 , 
 n384959 , n384960 , n37401 , n37402 , n384963 , n37404 , n384965 , n384966 , n37407 , n384968 , 
 n37409 , n37410 , n37411 , n384972 , n37413 , n384974 , n384975 , n384976 , n37417 , n384978 , 
 n384979 , n37420 , n384981 , n384982 , n37423 , n37424 , n384985 , n384986 , n37427 , n384988 , 
 n384989 , n37430 , n384991 , n384992 , n37433 , n384994 , n37435 , n384996 , n37437 , n37438 , 
 n384999 , n385000 , n37441 , n37442 , n385003 , n37444 , n37445 , n385006 , n385007 , n385008 , 
 n37449 , n385010 , n385011 , n37452 , n385013 , n385014 , n37455 , n37456 , n37457 , n385018 , 
 n385019 , n37460 , n37461 , n37462 , n385023 , n385024 , n37465 , n37466 , n37467 , n385028 , 
 n385029 , n37470 , n37471 , n37472 , n37473 , n37474 , n37475 , n385036 , n385037 , n37478 , 
 n385039 , n37480 , n37481 , n385042 , n37483 , n385044 , n37485 , n37486 , n385047 , n385048 , 
 n37489 , n385050 , n385051 , n37492 , n385053 , n385054 , n385055 , n37496 , n385057 , n385058 , 
 n37499 , n385060 , n385061 , n37502 , n385063 , n37504 , n385065 , n37506 , n37507 , n385068 , 
 n385069 , n37510 , n385071 , n385072 , n37513 , n385074 , n385075 , n37516 , n37517 , n37518 , 
 n385079 , n37520 , n37521 , n37522 , n37523 , n385084 , n37525 , n385086 , n37527 , n385088 , 
 n37529 , n385090 , n37531 , n37532 , n385093 , n385094 , n37535 , n385096 , n385097 , n37538 , 
 n385099 , n385100 , n37541 , n37542 , n385103 , n385104 , n37545 , n385106 , n385107 , n37548 , 
 n385109 , n385110 , n385111 , n37552 , n385113 , n385114 , n37555 , n385116 , n37557 , n385118 , 
 n37559 , n37560 , n37561 , n37562 , n37563 , n385124 , n37568 , n385126 , n37570 , n385128 , 
 n37572 , n37573 , n385131 , n37575 , n37576 , n385134 , n37578 , n37579 , n385137 , n385138 , 
 n37582 , n37583 , n37584 , n385142 , n385143 , n37587 , n37588 , n385146 , n385147 , n37591 , 
 n385149 , n37593 , n385151 , n37595 , n37596 , n37597 , n37598 , n37599 , n37600 , n37601 , 
 n37602 , n37603 , n385161 , n37605 , n385163 , n385164 , n385165 , n37609 , n385167 , n37611 , 
 n385169 , n37613 , n37614 , n385172 , n385173 , n37617 , n385175 , n385176 , n37620 , n385178 , 
 n385179 , n37623 , n37624 , n385182 , n385183 , n37627 , n385185 , n385186 , n37630 , n385188 , 
 n385189 , n37633 , n37634 , n37635 , n385193 , n385194 , n37638 , n37639 , n37640 , n385198 , 
 n385199 , n37643 , n37644 , n37645 , n385203 , n385204 , n37648 , n37649 , n385207 , n385208 , 
 n37652 , n37653 , n385211 , n385212 , n37656 , n37657 , n385215 , n385216 , n37660 , n37661 , 
 n385219 , n37663 , n37664 , n385222 , n37666 , n37667 , n385225 , n37669 , n385227 , n37671 , 
 n37672 , n37673 , n385231 , n385232 , n37676 , n37677 , n37678 , n37679 , n37680 , n37681 , 
 n37682 , n385240 , n37684 , n37685 , n385243 , n385244 , n37688 , n385246 , n385247 , n37691 , 
 n385249 , n385250 , n37694 , n37695 , n385253 , n37697 , n385255 , n37699 , n37700 , n385258 , 
 n385259 , n37703 , n37704 , n385262 , n37706 , n37707 , n385265 , n385266 , n385267 , n37711 , 
 n385269 , n385270 , n37714 , n385272 , n385273 , n37717 , n385275 , n385276 , n37720 , n37721 , 
 n37722 , n385280 , n385281 , n37725 , n37726 , n385284 , n385285 , n37729 , n37730 , n37731 , 
 n37732 , n385290 , n37739 , n385292 , n385293 , n37742 , n37743 , n37744 , n37745 , n37746 , 
 n385299 , n385300 , n385301 , n37750 , n385303 , n385304 , n37753 , n385306 , n37755 , n37756 , 
 n37757 , n37758 , n37759 , n37760 , n37761 , n37762 , n37763 , n385316 , n37765 , n385318 , 
 n385319 , n37768 , n37769 , n385322 , n37771 , n385324 , n385325 , n385326 , n37775 , n385328 , 
 n385329 , n37778 , n385331 , n385332 , n37781 , n385334 , n385335 , n37784 , n385337 , n385338 , 
 n37789 , n385340 , n37791 , n385342 , n385343 , n37794 , n385345 , n385346 , n37797 , n385348 , 
 n385349 , n37800 , n385351 , n37802 , n37803 , n385354 , n37805 , n385356 , n385357 , n37808 , 
 n385359 , n385360 , n385361 , n37812 , n37813 , n385364 , n385365 , n385366 , n37823 , n385368 , 
 n37825 , n37826 , n37827 , n37828 , n37829 , n385374 , n385375 , n37832 , n385377 , n37834 , 
 n37835 , n385380 , n385381 , n37838 , n385383 , n385384 , n37841 , n385386 , n385387 , n37844 , 
 n385389 , n37846 , n37847 , n37848 , n37849 , n37850 , n37851 , n385396 , n385397 , n37854 , 
 n385399 , n37856 , n37857 , n385402 , n385403 , n37860 , n385405 , n385406 , n37863 , n385408 , 
 n385409 , n385410 , n37867 , n385412 , n37869 , n37870 , n37871 , n385416 , n37873 , n385418 , 
 n37875 , n37876 , n385421 , n385422 , n37879 , n385424 , n385425 , n37882 , n385427 , n37884 , 
 n37885 , n385430 , n385431 , n37888 , n385433 , n37890 , n37891 , n37892 , n37893 , n385438 , 
 n37895 , n37896 , n37897 , n385442 , n385443 , n37900 , n37901 , n385446 , n385447 , n37904 , 
 n37905 , n37906 , n385451 , n385452 , n37909 , n37910 , n385455 , n385456 , n37913 , n37914 , 
 n37915 , n37916 , n37917 , n37918 , n37919 , n37920 , n37921 , n37922 , n37923 , n37924 , 
 n385469 , n37926 , n385471 , n37928 , n385473 , n37930 , n37931 , n37932 , n385477 , n37934 , 
 n385479 , n385480 , n37937 , n385482 , n385483 , n37940 , n37941 , n385486 , n37943 , n385488 , 
 n385489 , n37946 , n385491 , n385492 , n37949 , n385494 , n385495 , n37952 , n385497 , n37954 , 
 n385499 , n385500 , n37957 , n385502 , n385503 , n37960 , n37961 , n385506 , n385507 , n37964 , 
 n385509 , n385510 , n37967 , n385512 , n385513 , n37970 , n385515 , n37972 , n37973 , n37974 , 
 n385519 , n37976 , n385521 , n37978 , n37979 , n385524 , n385525 , n37982 , n385527 , n385528 , 
 n37985 , n385530 , n385531 , n385532 , n37989 , n385534 , n37991 , n37992 , n385537 , n37994 , 
 n385539 , n37996 , n37997 , n385542 , n385543 , n38000 , n38001 , n385546 , n38003 , n38004 , 
 n385549 , n385550 , n385551 , n38008 , n385553 , n385554 , n38011 , n385556 , n38013 , n38014 , 
 n38015 , n385560 , n38017 , n38018 , n38019 , n38020 , n385565 , n385566 , n38023 , n385568 , 
 n38025 , n38026 , n38027 , n38028 , n385573 , n385574 , n38031 , n385576 , n38033 , n385578 , 
 n38035 , n38036 , n38037 , n385582 , n385583 , n38040 , n38041 , n38042 , n385587 , n385588 , 
 n38045 , n38046 , n38047 , n385592 , n385593 , n38050 , n38051 , n38052 , n385597 , n385598 , 
 n38055 , n385600 , n385601 , n38058 , n385603 , n385604 , n38061 , n38062 , n385607 , n38064 , 
 n38065 , n385610 , n38067 , n38068 , n38069 , n38070 , n385615 , n385616 , n385617 , n38074 , 
 n385619 , n38076 , n38077 , n385622 , n38079 , n385624 , n38081 , n38082 , n385627 , n385628 , 
 n38085 , n385630 , n385631 , n38088 , n385633 , n385634 , n38091 , n385636 , n385637 , n38094 , 
 n385639 , n385640 , n385641 , n38098 , n385643 , n385644 , n38101 , n385646 , n385647 , n385648 , 
 n38105 , n385650 , n38107 , n38108 , n385653 , n385654 , n38111 , n38112 , n385657 , n38114 , 
 n38115 , n385660 , n385661 , n385662 , n38119 , n385664 , n385665 , n38122 , n385667 , n385668 , 
 n38125 , n38126 , n38127 , n385672 , n38129 , n38130 , n38131 , n385676 , n385677 , n38134 , 
 n38135 , n385680 , n385681 , n38138 , n38139 , n38140 , n385685 , n38142 , n38143 , n38144 , 
 n385689 , n385690 , n38147 , n385692 , n38149 , n385694 , n385695 , n385696 , n38153 , n38154 , 
 n38155 , n385700 , n38157 , n38158 , n38159 , n385704 , n38161 , n38162 , n385707 , n385708 , 
 n38165 , n385710 , n38167 , n38168 , n385713 , n385714 , n38171 , n385716 , n385717 , n38174 , 
 n385719 , n385720 , n38177 , n385722 , n38179 , n385724 , n38181 , n38182 , n385727 , n38184 , 
 n385729 , n385730 , n38187 , n385732 , n38189 , n385734 , n385735 , n38192 , n38193 , n385738 , 
 n38195 , n385740 , n385741 , n385742 , n38199 , n385744 , n385745 , n38202 , n385747 , n385748 , 
 n385749 , n38206 , n385751 , n385752 , n38209 , n385754 , n385755 , n38212 , n385757 , n385758 , 
 n38215 , n38216 , n38217 , n385762 , n385763 , n385764 , n38221 , n385766 , n38223 , n38224 , 
 n385769 , n38226 , n38227 , n385772 , n38229 , n385774 , n385775 , n38232 , n38233 , n385778 , 
 n385779 , n38236 , n385781 , n385782 , n38239 , n385784 , n385785 , n385786 , n38243 , n385788 , 
 n385789 , n38246 , n385791 , n385792 , n38249 , n385794 , n38251 , n385796 , n38253 , n385798 , 
 n38255 , n38256 , n385801 , n385802 , n38259 , n385804 , n385805 , n38262 , n385807 , n385808 , 
 n38265 , n38266 , n385811 , n385812 , n38269 , n385814 , n385815 , n38272 , n385817 , n385818 , 
 n38275 , n38276 , n38277 , n385822 , n385823 , n38280 , n38281 , n38282 , n385827 , n38284 , 
 n385829 , n38286 , n38287 , n385832 , n38289 , n385834 , n385835 , n385836 , n38293 , n385838 , 
 n385839 , n38296 , n385841 , n385842 , n385843 , n38300 , n385845 , n38302 , n385847 , n385848 , 
 n38305 , n385850 , n38307 , n385852 , n38309 , n38310 , n38311 , n38312 , n385857 , n38314 , 
 n38315 , n385860 , n385861 , n38318 , n385863 , n385864 , n38321 , n385866 , n385867 , n38324 , 
 n385869 , n38326 , n385871 , n38328 , n38329 , n385874 , n38331 , n385876 , n38333 , n38334 , 
 n385879 , n385880 , n38337 , n385882 , n385883 , n38340 , n385885 , n385886 , n385887 , n38344 , 
 n385889 , n385890 , n38347 , n385892 , n385893 , n38350 , n385895 , n385896 , n38353 , n385898 , 
 n38355 , n38356 , n38357 , n38358 , n38359 , n38360 , n38361 , n385906 , n38363 , n38364 , 
 n385909 , n385910 , n38367 , n385912 , n385913 , n38370 , n385915 , n385916 , n38373 , n38374 , 
 n38375 , n385920 , n385921 , n38378 , n38379 , n38380 , n385925 , n38382 , n38383 , n38384 , 
 n385929 , n385930 , n38387 , n38388 , n38389 , n385934 , n385935 , n38392 , n38393 , n38394 , 
 n385939 , n385940 , n38397 , n38398 , n38399 , n385944 , n385945 , n38402 , n385947 , n38404 , 
 n38405 , n385950 , n385951 , n38408 , n385953 , n38410 , n385955 , n38412 , n385957 , n385958 , 
 n38415 , n38416 , n38417 , n385962 , n385963 , n385964 , n38421 , n385966 , n38423 , n38424 , 
 n38425 , n385970 , n38427 , n385972 , n385973 , n38430 , n385975 , n385976 , n38433 , n385978 , 
 n38435 , n38436 , n385981 , n38438 , n385983 , n385984 , n385985 , n38442 , n385987 , n385988 , 
 n38445 , n385990 , n385991 , n38448 , n385993 , n385994 , n385995 , n38452 , n385997 , n385998 , 
 n38455 , n386000 , n386001 , n386002 , n38459 , n386004 , n38461 , n38462 , n386007 , n386008 , 
 n38465 , n386010 , n38467 , n386012 , n386013 , n38470 , n38471 , n38472 , n386017 , n386018 , 
 n38475 , n386020 , n386021 , n38478 , n386023 , n386024 , n38481 , n386026 , n386027 , n38484 , 
 n386029 , n386030 , n38487 , n386032 , n38489 , n386034 , n38491 , n38492 , n386037 , n38494 , 
 n386039 , n38496 , n38497 , n38498 , n386043 , n38500 , n386045 , n386046 , n386047 , n38504 , 
 n386049 , n386050 , n38507 , n386052 , n386053 , n38510 , n38511 , n38512 , n386057 , n386058 , 
 n38515 , n38516 , n38517 , n386062 , n386063 , n38520 , n38521 , n386066 , n386067 , n38524 , 
 n386069 , n38526 , n386071 , n38528 , n38529 , n386074 , n38531 , n38532 , n386077 , n38534 , 
 n38535 , n386080 , n386081 , n386082 , n386083 , n386084 , n38541 , n386086 , n386087 , n386088 , 
 n38545 , n386090 , n386091 , n38548 , n386093 , n386094 , n38551 , n386096 , n38553 , n386098 , 
 n38555 , n38556 , n386101 , n386102 , n38559 , n386104 , n386105 , n38562 , n386107 , n386108 , 
 n386109 , n38566 , n386111 , n38568 , n386113 , n38570 , n38571 , n386116 , n386117 , n38574 , 
 n386119 , n386120 , n38577 , n386122 , n386123 , n38580 , n386125 , n38582 , n386127 , n386128 , 
 n38585 , n386130 , n386131 , n38588 , n386133 , n386134 , n38591 , n386136 , n386137 , n38594 , 
 n38595 , n386140 , n386141 , n38598 , n386143 , n38606 , n386145 , n38608 , n386147 , n386148 , 
 n38611 , n386150 , n386151 , n38614 , n38615 , n386154 , n386155 , n38618 , n38619 , n386158 , 
 n386159 , n38625 , n386161 , n386162 , n386163 , n38629 , n38630 , n38631 , n386167 , n38633 , 
 n38634 , n386170 , n38636 , n386172 , n386173 , n386174 , n38640 , n386176 , n386177 , n38643 , 
 n386179 , n386180 , n38646 , n386182 , n386183 , n38649 , n38650 , n386186 , n386187 , n38653 , 
 n386189 , n386190 , n38656 , n386192 , n386193 , n38659 , n38660 , n38661 , n38662 , n386198 , 
 n386199 , n38665 , n386201 , n38667 , n38668 , n38669 , n38670 , n386206 , n386207 , n38673 , 
 n386209 , n386210 , n38676 , n386212 , n386213 , n38679 , n386215 , n38681 , n386217 , n38683 , 
 n386219 , n38685 , n386221 , n38687 , n386223 , n386224 , n386225 , n38691 , n38692 , n386228 , 
 n38694 , n38695 , n386231 , n386232 , n38698 , n386234 , n38700 , n386236 , n386237 , n386238 , 
 n38704 , n386240 , n386241 , n38707 , n38708 , n386244 , n386245 , n386246 , n38712 , n38713 , 
 n386249 , n386250 , n38716 , n38717 , n38718 , n386254 , n386255 , n38721 , n386257 , n386258 , 
 n38724 , n386260 , n386261 , n38727 , n386263 , n386264 , n38730 , n386266 , n386267 , n38733 , 
 n38734 , n38735 , n386271 , n386272 , n38738 , n386274 , n386275 , n38741 , n38742 , n38743 , 
 n386279 , n386280 , n386281 , n386282 , n38751 , n38752 , n386285 , n386286 , n386287 , n38756 , 
 n386289 , n386290 , n38759 , n386292 , n38761 , n386294 , n386295 , n38764 , n38765 , n386298 , 
 n38767 , n386300 , n386301 , n38770 , n38771 , n386304 , n386305 , n38774 , n386307 , n386308 , 
 n38777 , n386310 , n386311 , n38780 , n386313 , n386314 , n38783 , n386316 , n386317 , n38786 , 
 n38787 , n38788 , n386321 , n386322 , n386323 , n38792 , n386325 , n38794 , n38795 , n386328 , 
 n386329 , n38798 , n386331 , n386332 , n38801 , n386334 , n386335 , n38804 , n38805 , n38806 , 
 n386339 , n386340 , n38809 , n38810 , n38811 , n386344 , n386345 , n38814 , n386347 , n38816 , 
 n386349 , n38818 , n38819 , n386352 , n38821 , n38822 , n38823 , n386356 , n38825 , n38826 , 
 n386359 , n386360 , n38829 , n386362 , n386363 , n38832 , n386365 , n386366 , n386367 , n38836 , 
 n386369 , n386370 , n38839 , n386372 , n386373 , n38842 , n386375 , n386376 , n38845 , n386378 , 
 n386379 , n38848 , n386381 , n38850 , n386383 , n38852 , n386385 , n386386 , n38855 , n38856 , 
 n386389 , n38858 , n386391 , n386392 , n38861 , n386394 , n38863 , n386396 , n386397 , n38866 , 
 n386399 , n386400 , n38869 , n386402 , n38871 , n386404 , n386405 , n38874 , n386407 , n386408 , 
 n38877 , n38878 , n386411 , n38880 , n386413 , n38882 , n38883 , n386416 , n38885 , n386418 , 
 n386419 , n38888 , n386421 , n386422 , n38891 , n386424 , n386425 , n38894 , n386427 , n38896 , 
 n386429 , n386430 , n38899 , n386432 , n386433 , n386434 , n38903 , n386436 , n38905 , n386438 , 
 n38907 , n386440 , n386441 , n38910 , n386443 , n386444 , n38913 , n386446 , n386447 , n38916 , 
 n386449 , n386450 , n386451 , n38920 , n386453 , n386454 , n386455 , n38924 , n386457 , n386458 , 
 n38927 , n386460 , n386461 , n38930 , n386463 , n386464 , n38933 , n38934 , n38935 , n38936 , 
 n38937 , n38938 , n38939 , n386472 , n38941 , n386474 , n386475 , n38944 , n386477 , n386478 , 
 n38947 , n386480 , n386481 , n38950 , n386483 , n386484 , n38953 , n38954 , n38955 , n38956 , 
 n38957 , n38958 , n38959 , n38960 , n38961 , n386494 , n38963 , n386496 , n386497 , n38966 , 
 n386499 , n386500 , n38969 , n38970 , n38971 , n38972 , n386505 , n38974 , n386507 , n38976 , 
 n38977 , n386510 , n386511 , n38980 , n386513 , n386514 , n38983 , n386516 , n386517 , n38986 , 
 n386519 , n386520 , n38989 , n38990 , n386523 , n386524 , n38993 , n386526 , n38995 , n386528 , 
 n38997 , n38998 , n386531 , n386532 , n39001 , n39002 , n386535 , n39004 , n39005 , n386538 , 
 n386539 , n386540 , n39009 , n386542 , n386543 , n39012 , n386545 , n386546 , n39015 , n39016 , 
 n39017 , n386550 , n386551 , n39020 , n39021 , n386554 , n386555 , n39024 , n386557 , n39026 , 
 n386559 , n39028 , n386561 , n39030 , n39031 , n39032 , n39033 , n386566 , n39035 , n39036 , 
 n386569 , n386570 , n39039 , n386572 , n386573 , n39042 , n386575 , n386576 , n39045 , n386578 , 
 n386579 , n39048 , n39049 , n39050 , n39051 , n39052 , n39053 , n39054 , n39055 , n39056 , 
 n39057 , n39058 , n39059 , n39060 , n386593 , n39062 , n39063 , n39064 , n39065 , n386598 , 
 n386599 , n39068 , n386601 , n386602 , n39071 , n386604 , n386605 , n39074 , n386607 , n386608 , 
 n39077 , n386610 , n386611 , n39080 , n39081 , n39082 , n386615 , n386616 , n39085 , n386618 , 
 n386619 , n39088 , n386621 , n386622 , n39091 , n39092 , n386625 , n386626 , n39095 , n386628 , 
 n386629 , n39098 , n386631 , n39100 , n39101 , n39102 , n386635 , n386636 , n39105 , n39106 , 
 n39107 , n39108 , n386641 , n386642 , n39111 , n39112 , n39113 , n386646 , n386647 , n39116 , 
 n386649 , n39118 , n39119 , n39120 , n39121 , n39122 , n386655 , n39124 , n39125 , n39126 , 
 n39127 , n386660 , n386661 , n39130 , n386663 , n39132 , n39133 , n39134 , n39135 , n386668 , 
 n39137 , n39138 , n39139 , n39140 , n386673 , n39142 , n39143 , n39144 , n386677 , n39146 , 
 n39147 , n39148 , n39149 , n39150 , n39151 , n39152 , n39153 , n386686 , n386687 , n386688 , 
 n39157 , n39158 , n386691 , n39160 , n39161 , n386694 , n39163 , n39164 , n39165 , n386698 , 
 n39167 , n386700 , n386701 , n386702 , n39171 , n386704 , n39173 , n386706 , n386707 , n39176 , 
 n386709 , n39178 , n39179 , n386712 , n386713 , n39182 , n386715 , n386716 , n39185 , n386718 , 
 n386719 , n39188 , n39189 , n39190 , n39191 , n39192 , n39193 , n39194 , n386727 , n39211 , 
 n39212 , n386730 , n39214 , n386732 , n39216 , n386734 , n386735 , n39219 , n386737 , n386738 , 
 n39222 , n386740 , n386741 , n39225 , n386743 , n386744 , n39228 , n39229 , n386747 , n386748 , 
 n39232 , n386750 , n386751 , n39235 , n386753 , n39237 , n39238 , n39239 , n39240 , n39241 , 
 n386759 , n386760 , n39244 , n39245 , n39246 , n39247 , n39248 , n386766 , n39250 , n386768 , 
 n39252 , n386770 , n386771 , n39255 , n386773 , n386774 , n39258 , n386776 , n386777 , n39261 , 
 n386779 , n39263 , n39264 , n39265 , n39266 , n386784 , n39268 , n386786 , n39270 , n386788 , 
 n39272 , n39273 , n386791 , n386792 , n39276 , n386794 , n386795 , n39279 , n386797 , n386798 , 
 n39282 , n39283 , n386801 , n386802 , n39286 , n386804 , n386805 , n39289 , n386807 , n386808 , 
 n39292 , n386810 , n39294 , n386812 , n39296 , n386814 , n386815 , n39299 , n39300 , n386818 , 
 n39302 , n386820 , n39304 , n39305 , n386823 , n386824 , n39308 , n386826 , n386827 , n39311 , 
 n386829 , n386830 , n386831 , n39315 , n386833 , n386834 , n39318 , n386836 , n386837 , n39321 , 
 n386839 , n386840 , n39324 , n39325 , n386843 , n39327 , n386845 , n386846 , n386847 , n39331 , 
 n386849 , n386850 , n39334 , n386852 , n386853 , n386854 , n39338 , n386856 , n39340 , n39341 , 
 n39342 , n39343 , n39344 , n386862 , n386863 , n39347 , n386865 , n39349 , n386867 , n386868 , 
 n39352 , n386870 , n386871 , n39355 , n386873 , n386874 , n39358 , n386876 , n39360 , n386878 , 
 n386879 , n39363 , n386881 , n39365 , n386883 , n386884 , n386885 , n386886 , n39370 , n386888 , 
 n386889 , n39373 , n386891 , n39375 , n386893 , n39377 , n386895 , n386896 , n39380 , n39381 , 
 n386899 , n39383 , n39384 , n386902 , n386903 , n386904 , n39388 , n386906 , n39390 , n39391 , 
 n386909 , n39393 , n386911 , n386912 , n39396 , n386914 , n39398 , n386916 , n39400 , n39401 , 
 n39402 , n39403 , n39404 , n386922 , n386923 , n39407 , n386925 , n39409 , n386927 , n39411 , 
 n39412 , n386930 , n386931 , n39415 , n386933 , n386934 , n39418 , n386936 , n386937 , n39421 , 
 n39422 , n386940 , n386941 , n39425 , n386943 , n386944 , n39428 , n386946 , n386947 , n39431 , 
 n39432 , n39433 , n39434 , n39435 , n386953 , n386954 , n39438 , n386956 , n39440 , n39441 , 
 n39442 , n39443 , n39444 , n386962 , n39446 , n386964 , n39448 , n39449 , n39450 , n39451 , 
 n39452 , n39453 , n386971 , n39455 , n39456 , n386974 , n39458 , n386976 , n386977 , n39461 , 
 n39462 , n386980 , n386981 , n39465 , n39466 , n39467 , n39468 , n386986 , n386987 , n39471 , 
 n386989 , n386990 , n39474 , n386992 , n386993 , n386994 , n39478 , n386996 , n39480 , n386998 , 
 n39482 , n39483 , n387001 , n387002 , n39486 , n387004 , n387005 , n39489 , n387007 , n387008 , 
 n39492 , n39493 , n387011 , n39495 , n387013 , n39497 , n39498 , n387016 , n387017 , n39501 , 
 n387019 , n387020 , n39504 , n387022 , n387023 , n387024 , n39508 , n387026 , n387027 , n39511 , 
 n387029 , n387030 , n387031 , n39515 , n387033 , n39517 , n387035 , n387036 , n39520 , n39521 , 
 n387039 , n39523 , n387041 , n39525 , n39526 , n387044 , n387045 , n39529 , n387047 , n387048 , 
 n39532 , n387050 , n387051 , n39535 , n387053 , n387054 , n387055 , n39539 , n387057 , n39541 , 
 n387059 , n39543 , n39544 , n387062 , n387063 , n39547 , n387065 , n387066 , n39550 , n387068 , 
 n387069 , n39553 , n39554 , n39555 , n39556 , n39557 , n39558 , n387076 , n387077 , n39564 , 
 n387079 , n387080 , n39567 , n387082 , n39569 , n387084 , n39571 , n387086 , n39573 , n39574 , 
 n387089 , n387090 , n39577 , n387092 , n387093 , n39580 , n387095 , n387096 , n39583 , n39584 , 
 n387099 , n39586 , n387101 , n39588 , n39589 , n387104 , n387105 , n39592 , n387107 , n387108 , 
 n39595 , n387110 , n387111 , n387112 , n39599 , n387114 , n387115 , n39602 , n387117 , n387118 , 
 n39605 , n387120 , n387121 , n39608 , n387123 , n39610 , n387125 , n39612 , n387127 , n39614 , 
 n39615 , n387130 , n387131 , n39618 , n387133 , n387134 , n39621 , n387136 , n387137 , n39624 , 
 n39625 , n387140 , n387141 , n39628 , n387143 , n387144 , n39631 , n387146 , n39635 , n39636 , 
 n39637 , n39638 , n387151 , n387152 , n39644 , n387154 , n387155 , n39647 , n387157 , n39649 , 
 n387159 , n39651 , n387161 , n39653 , n39654 , n387164 , n387165 , n39657 , n387167 , n387168 , 
 n39660 , n387170 , n387171 , n387172 , n39664 , n387174 , n39666 , n39667 , n39668 , n39669 , 
 n39670 , n387180 , n39672 , n387182 , n387183 , n39675 , n39676 , n39677 , n39678 , n387188 , 
 n39680 , n387190 , n39682 , n387192 , n39684 , n39685 , n387195 , n387196 , n39688 , n387198 , 
 n387199 , n39691 , n387201 , n387202 , n39694 , n39695 , n387205 , n387206 , n39698 , n387208 , 
 n39700 , n387210 , n39702 , n387212 , n387213 , n39705 , n387215 , n387216 , n39708 , n387218 , 
 n39710 , n387220 , n39712 , n387222 , n387223 , n39715 , n387225 , n387226 , n39718 , n387228 , 
 n387229 , n39721 , n387231 , n39723 , n39724 , n39725 , n39726 , n39727 , n387237 , n387238 , 
 n387239 , n39731 , n387241 , n387242 , n39734 , n39735 , n387245 , n39737 , n39738 , n387248 , 
 n387249 , n39741 , n387251 , n387252 , n39744 , n39745 , n387255 , n387256 , n39748 , n387258 , 
 n387259 , n39751 , n387261 , n387262 , n39754 , n387264 , n39756 , n387266 , n39758 , n39759 , 
 n387269 , n387270 , n39765 , n387272 , n387273 , n39768 , n39769 , n39770 , n387277 , n387278 , 
 n39773 , n39774 , n387281 , n39776 , n387283 , n387284 , n39779 , n387286 , n387287 , n39782 , 
 n39783 , n387290 , n39785 , n39786 , n387293 , n39788 , n39789 , n39790 , n387297 , n387298 , 
 n39793 , n387300 , n39795 , n39796 , n39797 , n39798 , n39799 , n387306 , n387307 , n39802 , 
 n387309 , n387310 , n39805 , n39806 , n387313 , n39808 , n39809 , n39810 , n39811 , n39812 , 
 n39813 , n387320 , n39815 , n39816 , n39817 , n39818 , n39819 , n387326 , n39821 , n39822 , 
 n39823 , n39824 , n39825 , n39826 , n387333 , n387334 , n39829 , n387336 , n387337 , n39832 , 
 n387339 , n39834 , n39835 , n39836 , n39837 , n39838 , n387345 , n39840 , n387347 , n39842 , 
 n387349 , n39844 , n39845 , n387352 , n387353 , n39848 , n387355 , n387356 , n39851 , n387358 , 
 n387359 , n39854 , n39855 , n387362 , n39857 , n387364 , n39859 , n387366 , n387367 , n39862 , 
 n387369 , n39864 , n387371 , n39866 , n387373 , n39868 , n39869 , n39870 , n39871 , n39872 , 
 n39873 , n387380 , n387381 , n39876 , n387383 , n387384 , n39879 , n387386 , n39881 , n39882 , 
 n39883 , n39884 , n39885 , n387392 , n39887 , n39888 , n387395 , n387396 , n39891 , n387398 , 
 n387399 , n387400 , n39895 , n387402 , n39897 , n387404 , n39899 , n39900 , n387407 , n39902 , 
 n387409 , n387410 , n387411 , n39906 , n387413 , n39908 , n387415 , n387416 , n39911 , n387418 , 
 n39913 , n39914 , n39915 , n39916 , n39917 , n387424 , n387425 , n39920 , n387427 , n39922 , 
 n39923 , n387430 , n39925 , n39926 , n387433 , n39928 , n387435 , n387436 , n39931 , n387438 , 
 n39933 , n39934 , n387441 , n387442 , n39937 , n39938 , n387445 , n387446 , n39941 , n387448 , 
 n39943 , n387450 , n39945 , n39946 , n387453 , n387454 , n39949 , n387456 , n387457 , n39952 , 
 n387459 , n387460 , n39955 , n387462 , n387463 , n39958 , n39959 , n387466 , n387467 , n39962 , 
 n387469 , n39964 , n39965 , n39966 , n39967 , n39968 , n387475 , n39970 , n387477 , n387478 , 
 n39973 , n387480 , n39975 , n387482 , n39977 , n39978 , n39979 , n39980 , n39981 , n39982 , 
 n39983 , n387490 , n39985 , n387492 , n39987 , n39988 , n39989 , n39990 , n39991 , n39992 , 
 n39993 , n39994 , n39995 , n39996 , n39997 , n39998 , n39999 , n40000 , n40001 , n40002 , 
 n40003 , n40004 , n387511 , n387512 , n40007 , n387514 , n40009 , n387516 , n387517 , n387518 , 
 n387519 , n40014 , n387521 , n387522 , n40017 , n387524 , n40019 , n40020 , n40021 , n40022 , 
 n387529 , n40024 , n40025 , n40026 , n40027 , n387534 , n40029 , n387536 , n40031 , n40032 , 
 n40033 , n387540 , n40035 , n387542 , n40037 , n40038 , n40039 , n40040 , n387547 , n40042 , 
 n40043 , n387550 , n40045 , n387552 , n40047 , n387554 , n387555 , n40050 , n40051 , n40052 , 
 n40053 , n387560 , n40055 , n387562 , n387563 , n387564 , n40059 , n387566 , n40061 , n40062 , 
 n387569 , n387570 , n40065 , n387572 , n40067 , n387574 , n387575 , n40070 , n387577 , n387578 , 
 n40073 , n387580 , n40075 , n387582 , n40077 , n387584 , n387585 , n40080 , n40081 , n387588 , 
 n40083 , n387590 , n387591 , n387592 , n40087 , n387594 , n40089 , n387596 , n387597 , n40092 , 
 n387599 , n387600 , n387601 , n40096 , n387603 , n40098 , n40099 , n387606 , n40101 , n387608 , 
 n40103 , n40104 , n387611 , n387612 , n40107 , n387614 , n387615 , n40110 , n387617 , n387618 , 
 n387619 , n40114 , n387621 , n387622 , n40117 , n387624 , n387625 , n40125 , n40126 , n40127 , 
 n40128 , n387630 , n387631 , n40131 , n387633 , n387634 , n40134 , n387636 , n387637 , n40137 , 
 n387639 , n387640 , n40140 , n387642 , n40142 , n387644 , n40144 , n40145 , n387647 , n40147 , 
 n387649 , n40149 , n40150 , n387652 , n387653 , n40153 , n387655 , n387656 , n40156 , n387658 , 
 n387659 , n387660 , n40160 , n387662 , n387663 , n40163 , n387665 , n387666 , n40166 , n387668 , 
 n387669 , n40169 , n387671 , n40171 , n387673 , n40173 , n387675 , n40175 , n40176 , n387678 , 
 n387679 , n40179 , n387681 , n387682 , n40182 , n387684 , n387685 , n40185 , n40186 , n387688 , 
 n387689 , n40189 , n387691 , n387692 , n40192 , n387694 , n387695 , n40195 , n40196 , n40197 , 
 n40198 , n387700 , n387701 , n40201 , n387703 , n40203 , n387705 , n40205 , n40206 , n40207 , 
 n40208 , n40209 , n40210 , n387712 , n387713 , n40213 , n387715 , n387716 , n40216 , n387718 , 
 n387719 , n40219 , n387721 , n387722 , n40222 , n387724 , n387725 , n40225 , n387727 , n387728 , 
 n40228 , n40229 , n387731 , n387732 , n40232 , n387734 , n387735 , n40235 , n387737 , n387738 , 
 n40238 , n387740 , n387741 , n40241 , n40242 , n387744 , n387745 , n40245 , n40246 , n40247 , 
 n40248 , n387750 , n387751 , n40251 , n387753 , n387754 , n40254 , n387756 , n387757 , n40257 , 
 n40258 , n387760 , n40260 , n40261 , n387763 , n40263 , n40264 , n40265 , n40266 , n40267 , 
 n40268 , n387770 , n40270 , n387772 , n387773 , n40273 , n387775 , n387776 , n40276 , n387778 , 
 n40278 , n40279 , n387781 , n387782 , n40282 , n387784 , n387785 , n40285 , n387787 , n387788 , 
 n40288 , n40289 , n40290 , n387792 , n387793 , n40293 , n387795 , n40295 , n40296 , n40297 , 
 n40298 , n387800 , n40300 , n387802 , n40302 , n40303 , n387805 , n40305 , n387807 , n40307 , 
 n40308 , n40309 , n387811 , n40311 , n40312 , n387814 , n40314 , n387816 , n387817 , n40317 , 
 n387819 , n387820 , n40320 , n387822 , n40322 , n40323 , n387825 , n40325 , n387827 , n387828 , 
 n387829 , n387830 , n40330 , n387832 , n387833 , n40333 , n387835 , n387836 , n387837 , n40337 , 
 n387839 , n40339 , n40340 , n387842 , n387843 , n40346 , n387845 , n387846 , n387847 , n40350 , 
 n387849 , n40352 , n40353 , n387852 , n387853 , n40356 , n387855 , n387856 , n40359 , n387858 , 
 n387859 , n40362 , n387861 , n40364 , n387863 , n40366 , n40367 , n387866 , n387867 , n40370 , 
 n387869 , n387870 , n40373 , n387872 , n387873 , n40376 , n387875 , n387876 , n40379 , n40380 , 
 n40381 , n40382 , n387881 , n387882 , n387883 , n40386 , n387885 , n40388 , n40389 , n387888 , 
 n40391 , n387890 , n387891 , n387892 , n40395 , n387894 , n40397 , n40398 , n387897 , n387898 , 
 n40401 , n387900 , n387901 , n40404 , n387903 , n387904 , n40407 , n387906 , n40409 , n387908 , 
 n387909 , n40412 , n40413 , n40414 , n40415 , n40416 , n387915 , n387916 , n40419 , n387918 , 
 n387919 , n40422 , n40423 , n40424 , n40425 , n40426 , n387925 , n387926 , n40429 , n387928 , 
 n387929 , n40432 , n387931 , n387932 , n40435 , n40436 , n40437 , n40438 , n387937 , n387938 , 
 n40441 , n40442 , n40443 , n40444 , n387943 , n387944 , n40447 , n40448 , n40449 , n40450 , 
 n40451 , n387950 , n40453 , n387952 , n40455 , n387954 , n40457 , n40458 , n387957 , n387958 , 
 n40461 , n387960 , n387961 , n40464 , n387963 , n387964 , n387965 , n40468 , n387967 , n40470 , 
 n387969 , n40472 , n387971 , n387972 , n40475 , n40476 , n40477 , n40478 , n387977 , n387978 , 
 n40481 , n387980 , n387981 , n40484 , n387983 , n387984 , n40487 , n387986 , n40489 , n40490 , 
 n40491 , n40492 , n387991 , n387992 , n40495 , n387994 , n40497 , n387996 , n40499 , n40500 , 
 n387999 , n388000 , n40503 , n40504 , n388003 , n40506 , n388005 , n388006 , n40509 , n388008 , 
 n40511 , n40512 , n388011 , n388012 , n40515 , n40516 , n388015 , n40518 , n388017 , n40520 , 
 n388019 , n388020 , n40523 , n388022 , n388023 , n388024 , n40527 , n388026 , n388027 , n40530 , 
 n388029 , n388030 , n40533 , n388032 , n388033 , n40536 , n388035 , n388036 , n40539 , n388038 , 
 n388039 , n40542 , n40543 , n388042 , n388043 , n40546 , n40547 , n40548 , n40549 , n40550 , 
 n388049 , n388050 , n40553 , n388052 , n388053 , n40556 , n388055 , n40558 , n40559 , n388058 , 
 n40561 , n388060 , n40563 , n388062 , n40565 , n388064 , n40567 , n388066 , n40569 , n388068 , 
 n388069 , n40572 , n388071 , n388072 , n40575 , n388074 , n40577 , n388076 , n388077 , n388078 , 
 n40581 , n388080 , n388081 , n40584 , n40585 , n388084 , n40587 , n40588 , n388087 , n40590 , 
 n40591 , n40592 , n388091 , n40594 , n388093 , n388094 , n40597 , n40598 , n40599 , n40600 , 
 n40601 , n388100 , n40603 , n388102 , n388103 , n40606 , n388105 , n388106 , n40609 , n388108 , 
 n40611 , n40612 , n388111 , n40614 , n388113 , n388114 , n388115 , n40618 , n388117 , n388118 , 
 n40621 , n388120 , n388121 , n40624 , n388123 , n388124 , n40627 , n388126 , n40629 , n388128 , 
 n40631 , n40632 , n40633 , n40634 , n40635 , n40636 , n40637 , n40638 , n40639 , n40640 , 
 n388139 , n40642 , n388141 , n388142 , n40645 , n40646 , n40647 , n40648 , n40649 , n40650 , 
 n40651 , n40652 , n40653 , n388152 , n40655 , n388154 , n388155 , n40658 , n388157 , n388158 , 
 n40661 , n388160 , n388161 , n40664 , n388163 , n40666 , n40667 , n388166 , n388167 , n40670 , 
 n388169 , n388170 , n40673 , n388172 , n388173 , n40676 , n40677 , n388176 , n40679 , n388178 , 
 n40681 , n40682 , n388181 , n388182 , n40685 , n388184 , n388185 , n40688 , n388187 , n388188 , 
 n40691 , n388190 , n40693 , n388192 , n40695 , n40696 , n40697 , n40698 , n40699 , n40700 , 
 n40701 , n388200 , n40703 , n388202 , n388203 , n40706 , n388205 , n388206 , n40709 , n40710 , 
 n40711 , n40712 , n40713 , n40714 , n388213 , n40716 , n388215 , n40718 , n40719 , n40720 , 
 n388219 , n40722 , n388221 , n40724 , n40725 , n388224 , n388225 , n40728 , n388227 , n388228 , 
 n40731 , n388230 , n388231 , n40734 , n388233 , n40736 , n388235 , n388236 , n40739 , n40740 , 
 n388239 , n388240 , n40743 , n388242 , n388243 , n40746 , n388245 , n388246 , n40749 , n388248 , 
 n388249 , n40752 , n388251 , n388252 , n40755 , n388254 , n388255 , n40758 , n40759 , n40760 , 
 n388259 , n40762 , n388261 , n40764 , n388263 , n388264 , n40767 , n388266 , n388267 , n40770 , 
 n40771 , n388270 , n40773 , n388272 , n40775 , n388274 , n40777 , n40778 , n40779 , n388278 , 
 n40781 , n388280 , n388281 , n40784 , n388283 , n388284 , n40787 , n388286 , n40789 , n40790 , 
 n40791 , n40792 , n388291 , n40794 , n388293 , n40796 , n40797 , n388296 , n388297 , n40800 , 
 n388299 , n388300 , n40803 , n388302 , n40805 , n40806 , n388305 , n40808 , n388307 , n388308 , 
 n388309 , n40812 , n40813 , n40814 , n40815 , n40816 , n40817 , n40818 , n40819 , n388318 , 
 n388319 , n40822 , n40823 , n40824 , n388323 , n40826 , n40827 , n388326 , n388327 , n40830 , 
 n40831 , n40832 , n40833 , n388332 , n40835 , n388334 , n40837 , n40838 , n40839 , n40840 , 
 n388339 , n40842 , n40843 , n388342 , n388343 , n388344 , n40847 , n388346 , n388347 , n40850 , 
 n388349 , n388350 , n40853 , n40854 , n388353 , n388354 , n40857 , n40858 , n388357 , n40860 , 
 n388359 , n388360 , n40863 , n40864 , n40865 , n40866 , n388365 , n40868 , n388367 , n388368 , 
 n40871 , n388370 , n388371 , n40874 , n388373 , n388374 , n40877 , n388376 , n388377 , n40880 , 
 n40881 , n40882 , n40883 , n40884 , n40885 , n40886 , n388385 , n40888 , n40889 , n40890 , 
 n40891 , n40892 , n388391 , n40894 , n388393 , n388394 , n40897 , n388396 , n388397 , n40900 , 
 n40901 , n388400 , n40903 , n388402 , n388403 , n388404 , n40907 , n388406 , n388407 , n40910 , 
 n388409 , n388410 , n40913 , n388412 , n388413 , n388414 , n40917 , n40918 , n388417 , n40920 , 
 n388419 , n388420 , n40923 , n40924 , n388423 , n388424 , n40927 , n40928 , n388427 , n388428 , 
 n40931 , n40932 , n40933 , n388432 , n388433 , n40936 , n40937 , n388436 , n40939 , n388438 , 
 n40941 , n40942 , n40943 , n388442 , n388443 , n40946 , n388445 , n388446 , n40949 , n388448 , 
 n388449 , n40952 , n388451 , n40954 , n40955 , n40956 , n40957 , n40958 , n388457 , n388458 , 
 n40961 , n388460 , n388461 , n40964 , n388463 , n388464 , n388465 , n40968 , n40969 , n388468 , 
 n40971 , n40972 , n40973 , n40974 , n40975 , n40976 , n40977 , n40978 , n40979 , n40980 , 
 n388479 , n40982 , n40983 , n388482 , n388483 , n40986 , n388485 , n388486 , n40990 , n388488 , 
 n388489 , n40993 , n40994 , n388492 , n40996 , n40997 , n388495 , n388496 , n41002 , n388498 , 
 n388499 , n388500 , n41006 , n388502 , n388503 , n41009 , n388505 , n41011 , n41012 , n388508 , 
 n388509 , n41015 , n388511 , n388512 , n41018 , n388514 , n388515 , n41021 , n388517 , n388518 , 
 n41024 , n388520 , n388521 , n41027 , n41028 , n388524 , n388525 , n41031 , n388527 , n388528 , 
 n41034 , n41035 , n41036 , n388532 , n388533 , n41039 , n388535 , n388536 , n388537 , n41043 , 
 n388539 , n388540 , n388541 , n41047 , n388543 , n388544 , n41050 , n388546 , n388547 , n41053 , 
 n388549 , n388550 , n388551 , n41057 , n41058 , n388554 , n41060 , n388556 , n388557 , n41063 , 
 n41064 , n388560 , n388561 , n41067 , n388563 , n388564 , n41070 , n388566 , n388567 , n41073 , 
 n388569 , n388570 , n388571 , n41077 , n41078 , n388574 , n41080 , n388576 , n388577 , n41083 , 
 n41084 , n388580 , n388581 , n41087 , n41088 , n388584 , n41090 , n388586 , n41092 , n388588 , 
 n388589 , n41095 , n388591 , n41097 , n41098 , n388594 , n388595 , n41101 , n41102 , n388598 , 
 n41104 , n41105 , n41106 , n41107 , n41108 , n41109 , n41110 , n388606 , n41112 , n388608 , 
 n388609 , n388610 , n41116 , n41117 , n41118 , n388614 , n41120 , n41121 , n388617 , n388618 , 
 n41124 , n388620 , n41126 , n41127 , n388623 , n388624 , n41130 , n388626 , n388627 , n41133 , 
 n388629 , n388630 , n41136 , n388632 , n388633 , n41139 , n388635 , n388636 , n41142 , n41143 , 
 n41144 , n41145 , n388641 , n41147 , n388643 , n388644 , n41150 , n388646 , n388647 , n41153 , 
 n388649 , n41155 , n41156 , n388652 , n41158 , n388654 , n388655 , n388656 , n41162 , n388658 , 
 n388659 , n41165 , n388661 , n388662 , n41168 , n388664 , n41170 , n41171 , n388667 , n41173 , 
 n388669 , n388670 , n388671 , n41177 , n388673 , n388674 , n41180 , n388676 , n388677 , n41183 , 
 n388679 , n388680 , n41186 , n388682 , n388683 , n41189 , n388685 , n41191 , n41192 , n388688 , 
 n41194 , n41195 , n388691 , n41197 , n388693 , n388694 , n41200 , n388696 , n388697 , n41203 , 
 n388699 , n388700 , n41206 , n388702 , n41208 , n388704 , n388705 , n388706 , n41212 , n41213 , 
 n388709 , n388710 , n41216 , n41217 , n41218 , n388714 , n41220 , n41221 , n388717 , n41223 , 
 n388719 , n388720 , n41226 , n388722 , n41228 , n388724 , n388725 , n388726 , n41232 , n388728 , 
 n388729 , n388730 , n41236 , n388732 , n41238 , n388734 , n388735 , n41241 , n388737 , n388738 , 
 n41244 , n388740 , n388741 , n41247 , n388743 , n388744 , n41250 , n388746 , n388747 , n41253 , 
 n388749 , n41255 , n388751 , n388752 , n41258 , n388754 , n388755 , n41261 , n388757 , n388758 , 
 n41264 , n388760 , n388761 , n41267 , n388763 , n41269 , n388765 , n388766 , n41272 , n41273 , 
 n388769 , n41275 , n388771 , n388772 , n41278 , n388774 , n388775 , n388776 , n41282 , n388778 , 
 n388779 , n41285 , n388781 , n388782 , n41288 , n41289 , n388785 , n41291 , n388787 , n41293 , 
 n41294 , n388790 , n388791 , n41297 , n388793 , n388794 , n41300 , n388796 , n388797 , n388798 , 
 n41304 , n388800 , n388801 , n41307 , n388803 , n388804 , n41310 , n388806 , n388807 , n41313 , 
 n388809 , n388810 , n41316 , n388812 , n388813 , n41319 , n388815 , n388816 , n41322 , n41323 , 
 n41324 , n41325 , n41326 , n41327 , n41328 , n41329 , n41330 , n41331 , n41332 , n388828 , 
 n41334 , n388830 , n388831 , n41337 , n388833 , n388834 , n41340 , n41341 , n41342 , n388838 , 
 n41344 , n388840 , n41346 , n41347 , n388843 , n41349 , n388845 , n41351 , n388847 , n388848 , 
 n41354 , n388850 , n388851 , n41357 , n41358 , n41359 , n41360 , n41361 , n41362 , n41363 , 
 n388859 , n41365 , n41366 , n388862 , n388863 , n41369 , n388865 , n41371 , n41372 , n41373 , 
 n41374 , n388870 , n41376 , n388872 , n388873 , n41379 , n388875 , n388876 , n41382 , n388878 , 
 n388879 , n41385 , n41386 , n41387 , n388883 , n388884 , n41390 , n41391 , n41392 , n388888 , 
 n388889 , n388890 , n41396 , n388892 , n388893 , n41399 , n388895 , n41401 , n388897 , n388898 , 
 n41404 , n41405 , n388901 , n41407 , n388903 , n41409 , n388905 , n388906 , n41412 , n388908 , 
 n388909 , n41415 , n41416 , n388912 , n41418 , n41419 , n41420 , n388916 , n388917 , n41423 , 
 n388919 , n388920 , n41426 , n388922 , n388923 , n41429 , n41430 , n388926 , n41432 , n388928 , 
 n388929 , n41435 , n388931 , n388932 , n41438 , n41439 , n388935 , n388936 , n388937 , n41443 , 
 n388939 , n41445 , n388941 , n41447 , n388943 , n41449 , n388945 , n41451 , n388947 , n41453 , 
 n388949 , n388950 , n41456 , n388952 , n388953 , n41459 , n388955 , n388956 , n41462 , n41463 , 
 n388959 , n388960 , n41466 , n388962 , n388963 , n41469 , n388965 , n388966 , n41472 , n388968 , 
 n388969 , n41475 , n388971 , n388972 , n41478 , n41479 , n388975 , n41481 , n388977 , n41483 , 
 n388979 , n388980 , n41486 , n41487 , n41488 , n388984 , n41490 , n388986 , n388987 , n388988 , 
 n41494 , n388990 , n388991 , n41497 , n388993 , n388994 , n41500 , n388996 , n41502 , n388998 , 
 n388999 , n41505 , n389001 , n41507 , n41508 , n389004 , n389005 , n41511 , n389007 , n389008 , 
 n41514 , n389010 , n389011 , n41517 , n389013 , n41519 , n389015 , n389016 , n41522 , n41523 , 
 n389019 , n41525 , n389021 , n389022 , n41528 , n389024 , n389025 , n389026 , n41532 , n389028 , 
 n41534 , n41535 , n389031 , n389032 , n41538 , n389034 , n389035 , n41541 , n389037 , n389038 , 
 n41544 , n389040 , n389041 , n41547 , n389043 , n389044 , n41550 , n41551 , n41552 , n389048 , 
 n389049 , n41555 , n41556 , n41557 , n41558 , n41559 , n41560 , n41561 , n41562 , n41563 , 
 n41564 , n41565 , n389061 , n41567 , n389063 , n41569 , n389065 , n41571 , n389067 , n389068 , 
 n41574 , n41575 , n389071 , n41577 , n389073 , n41579 , n389075 , n389076 , n41582 , n389078 , 
 n389079 , n41585 , n389081 , n389082 , n41588 , n41589 , n389085 , n41591 , n41592 , n41593 , 
 n41594 , n41595 , n41596 , n389092 , n41598 , n41599 , n389095 , n389096 , n41602 , n389098 , 
 n389099 , n41605 , n389101 , n389102 , n389103 , n41609 , n389105 , n41611 , n389107 , n389108 , 
 n41614 , n389110 , n389111 , n389112 , n41618 , n389114 , n41620 , n389116 , n389117 , n41623 , 
 n389119 , n389120 , n41626 , n389122 , n389123 , n41629 , n389125 , n389126 , n41632 , n389128 , 
 n389129 , n41635 , n389131 , n389132 , n41638 , n41639 , n41640 , n389136 , n389137 , n41643 , 
 n41644 , n41645 , n389141 , n389142 , n41648 , n41649 , n389145 , n389146 , n41652 , n41653 , 
 n389149 , n41655 , n41656 , n389152 , n41658 , n41659 , n41660 , n41661 , n41662 , n41663 , 
 n41664 , n389160 , n41666 , n389162 , n389163 , n41669 , n41670 , n41671 , n389167 , n41673 , 
 n389169 , n41675 , n41676 , n389172 , n41678 , n389174 , n41680 , n389176 , n389177 , n41683 , 
 n389179 , n389180 , n41686 , n41687 , n389183 , n41689 , n389185 , n41691 , n41692 , n389188 , 
 n389189 , n41695 , n389191 , n389192 , n41698 , n389194 , n389195 , n389196 , n389197 , n41703 , 
 n389199 , n41705 , n41706 , n41707 , n41708 , n41709 , n41710 , n41711 , n389207 , n41713 , 
 n389209 , n389210 , n41716 , n389212 , n389213 , n41719 , n41720 , n41721 , n389217 , n389218 , 
 n41724 , n389220 , n389221 , n41727 , n389223 , n41729 , n41730 , n389226 , n41732 , n389228 , 
 n41734 , n389230 , n389231 , n41737 , n389233 , n389234 , n389235 , n41741 , n389237 , n41743 , 
 n389239 , n41745 , n389241 , n389242 , n41748 , n389244 , n389245 , n41751 , n389247 , n389248 , 
 n41754 , n389250 , n41756 , n389252 , n41758 , n41759 , n389255 , n41761 , n389257 , n41763 , 
 n41764 , n389260 , n389261 , n41767 , n389263 , n389264 , n41770 , n389266 , n389267 , n389268 , 
 n41774 , n389270 , n389271 , n41777 , n389273 , n389274 , n41780 , n41781 , n389277 , n389278 , 
 n41784 , n389280 , n41786 , n389282 , n41788 , n41789 , n389285 , n41791 , n389287 , n41793 , 
 n389289 , n389290 , n41796 , n41797 , n389293 , n389294 , n41800 , n389296 , n389297 , n41803 , 
 n389299 , n389300 , n389301 , n41807 , n389303 , n389304 , n41810 , n389306 , n389307 , n389308 , 
 n41814 , n389310 , n41816 , n41817 , n389313 , n389314 , n41820 , n389316 , n389317 , n41823 , 
 n389319 , n389320 , n41826 , n389322 , n41828 , n41829 , n389325 , n389326 , n41832 , n389328 , 
 n389329 , n41835 , n389331 , n389332 , n41838 , n389334 , n389335 , n389336 , n41842 , n389338 , 
 n389339 , n41845 , n389341 , n41847 , n41848 , n41849 , n41850 , n389346 , n41858 , n389348 , 
 n389349 , n41861 , n389351 , n41863 , n389353 , n389354 , n41866 , n389356 , n389357 , n41869 , 
 n389359 , n389360 , n41872 , n389362 , n41874 , n41875 , n389365 , n389366 , n389367 , n389368 , 
 n389369 , n41881 , n389371 , n41883 , n389373 , n41885 , n41886 , n389376 , n389377 , n41889 , 
 n389379 , n41891 , n389381 , n389382 , n41894 , n389384 , n41896 , n41897 , n41898 , n389388 , 
 n41900 , n41901 , n389391 , n41903 , n41904 , n389394 , n41906 , n41907 , n41908 , n41909 , 
 n389399 , n41911 , n389401 , n389402 , n389403 , n41915 , n389405 , n389406 , n41918 , n389408 , 
 n389409 , n41921 , n41922 , n41923 , n389413 , n389414 , n41926 , n389416 , n41928 , n389418 , 
 n41930 , n389420 , n389421 , n41933 , n389423 , n41935 , n389425 , n41937 , n41938 , n389428 , 
 n41940 , n389430 , n41942 , n41943 , n389433 , n41945 , n389435 , n389436 , n389437 , n41949 , 
 n389439 , n389440 , n41952 , n389442 , n389443 , n389444 , n41956 , n389446 , n389447 , n41959 , 
 n389449 , n389450 , n41962 , n41963 , n41964 , n389454 , n389455 , n41967 , n389457 , n389458 , 
 n41970 , n389460 , n389461 , n41973 , n389463 , n41975 , n389465 , n41977 , n389467 , n389468 , 
 n41980 , n41981 , n389471 , n389472 , n41984 , n389474 , n389475 , n41987 , n389477 , n389478 , 
 n41990 , n41991 , n389481 , n41993 , n389483 , n41995 , n389485 , n389486 , n41998 , n41999 , 
 n389489 , n389490 , n42002 , n389492 , n389493 , n42005 , n389495 , n389496 , n389497 , n42009 , 
 n389499 , n389500 , n42012 , n389502 , n389503 , n389504 , n42016 , n389506 , n42018 , n389508 , 
 n42020 , n42021 , n389511 , n389512 , n42024 , n389514 , n389515 , n42027 , n389517 , n389518 , 
 n42030 , n42031 , n389521 , n42033 , n389523 , n42035 , n389525 , n389526 , n42038 , n42039 , 
 n389529 , n389530 , n42042 , n389532 , n389533 , n42045 , n389535 , n389536 , n389537 , n42049 , 
 n389539 , n389540 , n42052 , n389542 , n389543 , n42055 , n389545 , n42062 , n389547 , n389548 , 
 n42065 , n42066 , n389551 , n42068 , n389553 , n42070 , n42071 , n389556 , n42073 , n42074 , 
 n389559 , n42076 , n389561 , n389562 , n42079 , n389564 , n389565 , n42082 , n389567 , n389568 , 
 n42085 , n389570 , n389571 , n389572 , n42089 , n389574 , n42091 , n42092 , n42093 , n42094 , 
 n42095 , n42096 , n389581 , n42098 , n389583 , n389584 , n42101 , n389586 , n389587 , n42104 , 
 n389589 , n389590 , n389591 , n42108 , n389593 , n389594 , n42111 , n389596 , n42113 , n389598 , 
 n389599 , n389600 , n42117 , n389602 , n389603 , n42120 , n42121 , n389606 , n389607 , n42124 , 
 n389609 , n389610 , n42127 , n42128 , n389613 , n389614 , n42131 , n42132 , n42133 , n389618 , 
 n389619 , n42136 , n389621 , n42138 , n42139 , n42140 , n389625 , n42142 , n42143 , n42144 , 
 n42145 , n42146 , n389631 , n389632 , n389633 , n42150 , n42151 , n42152 , n42153 , n42154 , 
 n42155 , n389640 , n389641 , n42158 , n389643 , n42160 , n389645 , n42162 , n42163 , n389648 , 
 n389649 , n42166 , n389651 , n389652 , n42169 , n389654 , n389655 , n42172 , n42173 , n42174 , 
 n389659 , n389660 , n42177 , n389662 , n389663 , n389664 , n389665 , n42182 , n389667 , n389668 , 
 n42185 , n389670 , n42187 , n42188 , n42189 , n42190 , n42191 , n42192 , n42193 , n389678 , 
 n389679 , n389680 , n42197 , n389682 , n42199 , n42200 , n389685 , n42202 , n389687 , n42204 , 
 n42205 , n389690 , n42207 , n389692 , n389693 , n389694 , n42211 , n389696 , n389697 , n42214 , 
 n389699 , n389700 , n389701 , n42218 , n389703 , n389704 , n42221 , n389706 , n389707 , n389708 , 
 n42225 , n389710 , n42227 , n42228 , n389713 , n42230 , n389715 , n42232 , n42233 , n42234 , 
 n389719 , n42236 , n389721 , n42238 , n389723 , n389724 , n42241 , n389726 , n389727 , n389728 , 
 n42245 , n389730 , n389731 , n42248 , n389733 , n389734 , n42251 , n389736 , n42253 , n389738 , 
 n389739 , n389740 , n42257 , n389742 , n42259 , n389744 , n389745 , n42262 , n42263 , n389748 , 
 n389749 , n42266 , n389751 , n42268 , n389753 , n389754 , n42271 , n42272 , n389757 , n42274 , 
 n389759 , n389760 , n389761 , n42278 , n389763 , n389764 , n42281 , n389766 , n389767 , n42284 , 
 n389769 , n389770 , n42287 , n389772 , n389773 , n42290 , n389775 , n42301 , n389777 , n389778 , 
 n389779 , n42305 , n42306 , n389782 , n389783 , n42309 , n42310 , n42311 , n389787 , n389788 , 
 n42314 , n389790 , n389791 , n42317 , n389793 , n42319 , n389795 , n42321 , n389797 , n42323 , 
 n42324 , n389800 , n42326 , n389802 , n389803 , n42329 , n389805 , n389806 , n42332 , n389808 , 
 n389809 , n389810 , n42336 , n389812 , n389813 , n42339 , n389815 , n389816 , n42342 , n42343 , 
 n389819 , n42345 , n389821 , n42347 , n389823 , n389824 , n42350 , n389826 , n389827 , n389828 , 
 n42354 , n389830 , n42356 , n389832 , n42358 , n42359 , n389835 , n389836 , n42362 , n389838 , 
 n389839 , n42365 , n389841 , n389842 , n42368 , n42369 , n389845 , n389846 , n42372 , n389848 , 
 n389849 , n42375 , n389851 , n389852 , n42378 , n389854 , n42380 , n389856 , n389857 , n42383 , 
 n389859 , n389860 , n42386 , n389862 , n389863 , n42389 , n42390 , n389866 , n42392 , n42393 , 
 n389869 , n389870 , n42396 , n389872 , n389873 , n42399 , n389875 , n389876 , n42402 , n389878 , 
 n42404 , n389880 , n389881 , n42407 , n389883 , n389884 , n42410 , n42411 , n389887 , n42413 , 
 n389889 , n42415 , n42416 , n389892 , n42418 , n389894 , n389895 , n42421 , n389897 , n389898 , 
 n389899 , n42425 , n389901 , n389902 , n42428 , n389904 , n389905 , n389906 , n42432 , n389908 , 
 n389909 , n42435 , n389911 , n389912 , n42438 , n389914 , n389915 , n42441 , n42442 , n42443 , 
 n389919 , n389920 , n389921 , n42447 , n389923 , n42449 , n42450 , n389926 , n42452 , n389928 , 
 n389929 , n42455 , n389931 , n42457 , n42458 , n389934 , n42460 , n389936 , n389937 , n389938 , 
 n42464 , n389940 , n389941 , n42467 , n389943 , n389944 , n42470 , n389946 , n389947 , n389948 , 
 n42474 , n389950 , n389951 , n42477 , n389953 , n389954 , n42480 , n389956 , n389957 , n389958 , 
 n389959 , n42485 , n42486 , n389962 , n42488 , n389964 , n389965 , n42491 , n42492 , n389968 , 
 n389969 , n42495 , n389971 , n42497 , n42498 , n389974 , n389975 , n42501 , n42502 , n389978 , 
 n389979 , n42505 , n389981 , n389982 , n42508 , n389984 , n42510 , n389986 , n42512 , n42513 , 
 n389989 , n389990 , n42516 , n389992 , n42518 , n42519 , n389995 , n42521 , n389997 , n389998 , 
 n389999 , n42525 , n390001 , n390002 , n390003 , n390004 , n390005 , n42531 , n390007 , n390008 , 
 n42534 , n390010 , n390011 , n42537 , n390013 , n390014 , n42540 , n390016 , n42542 , n390018 , 
 n42544 , n42545 , n390021 , n390022 , n42548 , n390024 , n390025 , n42551 , n390027 , n390028 , 
 n42554 , n390030 , n390031 , n42557 , n390033 , n42559 , n42560 , n42561 , n42562 , n390038 , 
 n42564 , n390040 , n42566 , n42567 , n42568 , n42569 , n390045 , n42571 , n390047 , n390048 , 
 n42574 , n42575 , n42576 , n42577 , n390053 , n390054 , n390055 , n42581 , n390057 , n42583 , 
 n42584 , n390060 , n42586 , n390062 , n42588 , n42589 , n390065 , n390066 , n42592 , n390068 , 
 n390069 , n42595 , n390071 , n390072 , n390073 , n42599 , n390075 , n390076 , n42602 , n390078 , 
 n390079 , n42605 , n42606 , n42607 , n42608 , n42609 , n390085 , n390086 , n42612 , n390088 , 
 n390089 , n42615 , n42616 , n42617 , n390093 , n390094 , n42620 , n390096 , n42622 , n390098 , 
 n42624 , n390100 , n390101 , n42627 , n390103 , n42629 , n42630 , n42631 , n390107 , n42633 , 
 n42634 , n390110 , n42636 , n390112 , n42638 , n390114 , n42640 , n42641 , n390117 , n42643 , 
 n390119 , n390120 , n390121 , n42647 , n390123 , n390124 , n42650 , n390126 , n390127 , n390128 , 
 n42654 , n390130 , n42656 , n390132 , n42658 , n390134 , n390135 , n42661 , n390137 , n390138 , 
 n390139 , n42665 , n390141 , n42667 , n42668 , n390144 , n42670 , n390146 , n390147 , n390148 , 
 n42674 , n390150 , n42676 , n390152 , n390153 , n42679 , n390155 , n390156 , n42682 , n390158 , 
 n390159 , n42685 , n42686 , n390162 , n390163 , n42689 , n42690 , n390166 , n42692 , n390168 , 
 n42694 , n390170 , n42696 , n390172 , n390173 , n42699 , n42700 , n390176 , n42702 , n390178 , 
 n390179 , n390180 , n42706 , n390182 , n390183 , n42709 , n390185 , n390186 , n390187 , n42713 , 
 n390189 , n42715 , n390191 , n42717 , n42718 , n390194 , n390195 , n42721 , n390197 , n390198 , 
 n42724 , n390200 , n390201 , n42727 , n390203 , n42729 , n390205 , n390206 , n42732 , n390208 , 
 n390209 , n42735 , n390211 , n42737 , n390213 , n390214 , n42740 , n390216 , n42742 , n390218 , 
 n390219 , n42745 , n42746 , n390222 , n390223 , n390224 , n42750 , n42751 , n390227 , n42753 , 
 n42754 , n390230 , n390231 , n42757 , n390233 , n390234 , n42760 , n390236 , n390237 , n42763 , 
 n390239 , n390240 , n42766 , n42767 , n390243 , n42769 , n390245 , n390246 , n390247 , n42773 , 
 n390249 , n390250 , n42776 , n390252 , n390253 , n390254 , n42780 , n390256 , n42782 , n390258 , 
 n42784 , n390260 , n390261 , n42787 , n42788 , n390264 , n42790 , n390266 , n42792 , n42793 , 
 n390269 , n42795 , n390271 , n390272 , n42798 , n42799 , n390275 , n42801 , n390277 , n390278 , 
 n42804 , n390280 , n390281 , n390282 , n42808 , n390284 , n390285 , n42811 , n390287 , n390288 , 
 n42814 , n390290 , n42816 , n390292 , n390293 , n390294 , n42820 , n390296 , n390297 , n42823 , 
 n390299 , n42825 , n390301 , n390302 , n42828 , n42829 , n390305 , n42831 , n390307 , n390308 , 
 n42834 , n42835 , n390311 , n390312 , n42838 , n42839 , n390315 , n390316 , n42842 , n390318 , 
 n390319 , n42845 , n390321 , n42847 , n390323 , n42849 , n390325 , n42851 , n42852 , n390328 , 
 n390329 , n42855 , n42856 , n390332 , n42858 , n42859 , n390335 , n390336 , n42862 , n390338 , 
 n42864 , n42865 , n390341 , n42867 , n390343 , n42869 , n390345 , n390346 , n42872 , n42873 , 
 n390349 , n42875 , n390351 , n390352 , n390353 , n42879 , n390355 , n390356 , n42882 , n390358 , 
 n390359 , n390360 , n42886 , n390362 , n390363 , n42889 , n42890 , n390366 , n390367 , n42893 , 
 n390369 , n42895 , n390371 , n42897 , n390373 , n390374 , n42900 , n42901 , n390377 , n42903 , 
 n390379 , n390380 , n390381 , n42907 , n390383 , n390384 , n42910 , n390386 , n390387 , n42913 , 
 n390389 , n42915 , n42916 , n390392 , n390393 , n42919 , n390395 , n42921 , n42922 , n42923 , 
 n42924 , n42925 , n390401 , n42927 , n390403 , n42929 , n390405 , n42931 , n390407 , n42933 , 
 n42934 , n390410 , n390411 , n42937 , n390413 , n390414 , n42940 , n390416 , n42942 , n42943 , 
 n42944 , n390420 , n42946 , n390422 , n42948 , n42949 , n42950 , n42951 , n390427 , n42953 , 
 n390429 , n390430 , n42956 , n390432 , n390433 , n42959 , n390435 , n42961 , n42962 , n390438 , 
 n42964 , n390440 , n390441 , n42967 , n42968 , n390444 , n390445 , n42971 , n42972 , n390448 , 
 n390449 , n42975 , n390451 , n42977 , n390453 , n390454 , n42980 , n42981 , n390457 , n390458 , 
 n42984 , n390460 , n390461 , n42987 , n390463 , n390464 , n42990 , n390466 , n390467 , n42993 , 
 n390469 , n42995 , n42996 , n390472 , n42998 , n390474 , n43000 , n390476 , n390477 , n43003 , 
 n390479 , n390480 , n43006 , n390482 , n390483 , n43009 , n390485 , n390486 , n43012 , n390488 , 
 n43014 , n390490 , n390491 , n43017 , n390493 , n43019 , n43020 , n390496 , n43022 , n390498 , 
 n390499 , n390500 , n43026 , n390502 , n390503 , n43029 , n390505 , n390506 , n43032 , n43033 , 
 n390509 , n390510 , n43036 , n390512 , n390513 , n43039 , n390515 , n43041 , n390517 , n43043 , 
 n43044 , n390520 , n43046 , n43047 , n390523 , n43049 , n390525 , n43051 , n390527 , n390528 , 
 n43054 , n390530 , n390531 , n43057 , n43058 , n390534 , n43060 , n390536 , n390537 , n43063 , 
 n43064 , n390540 , n43066 , n390542 , n43068 , n43069 , n390545 , n390546 , n43072 , n390548 , 
 n390549 , n43075 , n390551 , n390552 , n43078 , n390554 , n390555 , n390556 , n43082 , n390558 , 
 n390559 , n43085 , n390561 , n390562 , n390563 , n43089 , n390565 , n43091 , n390567 , n390568 , 
 n43094 , n43095 , n390571 , n43097 , n390573 , n43099 , n390575 , n390576 , n43102 , n390578 , 
 n390579 , n43105 , n390581 , n43107 , n390583 , n43109 , n43110 , n390586 , n390587 , n43113 , 
 n390589 , n390590 , n43116 , n390592 , n390593 , n43119 , n390595 , n43121 , n43122 , n390598 , 
 n390599 , n43125 , n390601 , n390602 , n43128 , n390604 , n390605 , n43131 , n43132 , n43133 , 
 n390609 , n43135 , n43136 , n43137 , n43138 , n43139 , n43140 , n43141 , n43142 , n390618 , 
 n43144 , n390620 , n43146 , n390622 , n43148 , n390624 , n43150 , n390626 , n390627 , n43153 , 
 n390629 , n390630 , n43156 , n43157 , n390633 , n43159 , n390635 , n390636 , n390637 , n43163 , 
 n390639 , n390640 , n43166 , n390642 , n390643 , n43169 , n43170 , n43171 , n390647 , n43173 , 
 n390649 , n43175 , n390651 , n390652 , n43178 , n43179 , n390655 , n43181 , n390657 , n390658 , 
 n390659 , n43185 , n390661 , n390662 , n43188 , n390664 , n43190 , n43191 , n390667 , n43193 , 
 n43194 , n43195 , n390671 , n43197 , n390673 , n43199 , n43200 , n43201 , n43202 , n43203 , 
 n43204 , n390680 , n390681 , n43207 , n390683 , n43209 , n43210 , n390686 , n43212 , n390688 , 
 n43214 , n43215 , n390691 , n390692 , n43218 , n390694 , n390695 , n43221 , n390697 , n43223 , 
 n43224 , n390700 , n43226 , n390702 , n43228 , n390704 , n390705 , n43231 , n43232 , n390708 , 
 n390709 , n43235 , n390711 , n390712 , n43238 , n390714 , n43240 , n43241 , n43242 , n43243 , 
 n390719 , n43245 , n390721 , n43247 , n43248 , n390724 , n390725 , n43251 , n390727 , n390728 , 
 n43254 , n390730 , n43256 , n43257 , n43258 , n390734 , n43260 , n390736 , n43262 , n43263 , 
 n390739 , n390740 , n43266 , n390742 , n390743 , n43269 , n390745 , n390746 , n43272 , n390748 , 
 n43274 , n390750 , n43276 , n43277 , n43278 , n43279 , n390755 , n43281 , n43282 , n43283 , 
 n390759 , n43285 , n43286 , n390762 , n43288 , n390764 , n43290 , n390766 , n43292 , n43293 , 
 n390769 , n390770 , n43296 , n390772 , n390773 , n43299 , n390775 , n390776 , n43302 , n43303 , 
 n390779 , n43305 , n390781 , n43307 , n390783 , n390784 , n43310 , n390786 , n43312 , n43313 , 
 n43314 , n390790 , n43316 , n390792 , n43318 , n390794 , n390795 , n43321 , n43322 , n390798 , 
 n390799 , n43325 , n390801 , n390802 , n43328 , n390804 , n43330 , n390806 , n43332 , n390808 , 
 n43334 , n390810 , n390811 , n43337 , n43338 , n390814 , n390815 , n43341 , n390817 , n390818 , 
 n43344 , n390820 , n43346 , n43347 , n43348 , n390824 , n43350 , n390826 , n43352 , n390828 , 
 n43354 , n390830 , n43356 , n390832 , n390833 , n43359 , n43360 , n390836 , n390837 , n43363 , 
 n390839 , n390840 , n43366 , n390842 , n390843 , n43369 , n43370 , n43371 , n43372 , n43373 , 
 n390849 , n390850 , n43376 , n390852 , n43378 , n43379 , n390855 , n43381 , n43382 , n390858 , 
 n43384 , n390860 , n43386 , n43387 , n390863 , n43389 , n390865 , n390866 , n43392 , n43393 , 
 n390869 , n390870 , n390871 , n43397 , n390873 , n43399 , n390875 , n390876 , n43402 , n43403 , 
 n390879 , n390880 , n43406 , n390882 , n390883 , n43409 , n390885 , n390886 , n43412 , n390888 , 
 n43414 , n43415 , n390891 , n390892 , n43418 , n390894 , n390895 , n43421 , n390897 , n390898 , 
 n43424 , n390900 , n390901 , n43427 , n43428 , n390904 , n43430 , n43431 , n390907 , n390908 , 
 n43434 , n390910 , n43436 , n43437 , n390913 , n43439 , n390915 , n43441 , n43442 , n390918 , 
 n43444 , n390920 , n390921 , n390922 , n43448 , n390924 , n43450 , n43451 , n390927 , n43453 , 
 n390929 , n390930 , n390931 , n43457 , n390933 , n390934 , n43460 , n390936 , n390937 , n43463 , 
 n390939 , n43465 , n43466 , n390942 , n390943 , n43469 , n390945 , n390946 , n43472 , n390948 , 
 n390949 , n43475 , n43476 , n43477 , n43478 , n43479 , n390955 , n43481 , n390957 , n43483 , 
 n43484 , n390960 , n390961 , n43487 , n390963 , n390964 , n43490 , n390966 , n390967 , n43493 , 
 n43494 , n43495 , n390971 , n390972 , n43498 , n390974 , n43500 , n43501 , n43502 , n43503 , 
 n43504 , n43505 , n43506 , n43507 , n390983 , n43509 , n390985 , n390986 , n43512 , n390988 , 
 n43514 , n43515 , n43516 , n390992 , n43518 , n43519 , n390995 , n43521 , n390997 , n43523 , 
 n43524 , n43525 , n43526 , n43527 , n43528 , n43529 , n43530 , n43531 , n43532 , n43533 , 
 n43534 , n43535 , n43536 , n43537 , n391013 , n43539 , n43540 , n391016 , n43542 , n391018 , 
 n391019 , n43545 , n391021 , n391022 , n43548 , n391024 , n391025 , n43551 , n391027 , n391028 , 
 n43554 , n391030 , n43556 , n391032 , n391033 , n43559 , n43560 , n391036 , n391037 , n43563 , 
 n391039 , n391040 , n43566 , n391042 , n391043 , n43569 , n391045 , n391046 , n43572 , n43573 , 
 n391049 , n391050 , n43576 , n43577 , n43578 , n391054 , n391055 , n43581 , n391057 , n43583 , 
 n43584 , n391060 , n43586 , n391062 , n43588 , n391064 , n43590 , n43591 , n43592 , n43593 , 
 n43594 , n43595 , n43596 , n43597 , n43598 , n43599 , n43600 , n391076 , n43602 , n391078 , 
 n43604 , n391080 , n391081 , n43607 , n391083 , n43609 , n43610 , n391086 , n43612 , n391088 , 
 n43614 , n43615 , n391091 , n391092 , n43618 , n391094 , n391095 , n43621 , n391097 , n391098 , 
 n391099 , n43625 , n391101 , n391102 , n43628 , n391104 , n391105 , n391106 , n43632 , n391108 , 
 n43634 , n43635 , n391111 , n391112 , n43638 , n391114 , n391115 , n43641 , n391117 , n391118 , 
 n43644 , n391120 , n43646 , n391122 , n43648 , n43649 , n391125 , n43651 , n391127 , n43653 , 
 n391129 , n391130 , n43656 , n43657 , n391133 , n391134 , n43660 , n391136 , n391137 , n43663 , 
 n391139 , n391140 , n391141 , n43667 , n391143 , n391144 , n43670 , n391146 , n391147 , n391148 , 
 n43674 , n391150 , n43676 , n43677 , n391153 , n391154 , n43680 , n391156 , n391157 , n43683 , 
 n391159 , n391160 , n43686 , n391162 , n43688 , n391164 , n391165 , n391166 , n43692 , n391168 , 
 n43694 , n391170 , n391171 , n43697 , n391173 , n391174 , n43700 , n391176 , n391177 , n391178 , 
 n391179 , n43705 , n391181 , n43707 , n391183 , n391184 , n391185 , n43711 , n43712 , n391188 , 
 n391189 , n43715 , n43716 , n391192 , n391193 , n43719 , n391195 , n391196 , n43722 , n391198 , 
 n43724 , n391200 , n43726 , n43727 , n391203 , n43729 , n391205 , n43731 , n391207 , n43733 , 
 n43734 , n391210 , n43736 , n391212 , n391213 , n391214 , n43740 , n391216 , n391217 , n43743 , 
 n391219 , n391220 , n43746 , n43747 , n391223 , n391224 , n43750 , n391226 , n391227 , n43753 , 
 n391229 , n391230 , n43756 , n391232 , n43758 , n43759 , n391235 , n391236 , n43762 , n391238 , 
 n391239 , n43765 , n391241 , n391242 , n43768 , n391244 , n43770 , n43771 , n391247 , n391248 , 
 n43774 , n391250 , n391251 , n43777 , n391253 , n391254 , n391255 , n391256 , n43782 , n43783 , 
 n391259 , n43785 , n43786 , n391262 , n391263 , n43789 , n391265 , n391266 , n43792 , n391268 , 
 n43794 , n391270 , n391271 , n43797 , n43798 , n391274 , n43800 , n391276 , n43802 , n391278 , 
 n391279 , n43805 , n391281 , n391282 , n43808 , n43809 , n391285 , n391286 , n391287 , n43813 , 
 n43814 , n43815 , n391291 , n43817 , n391293 , n43819 , n391295 , n43821 , n391297 , n43823 , 
 n43824 , n391300 , n391301 , n43827 , n391303 , n391304 , n43830 , n391306 , n391307 , n43833 , 
 n43834 , n391310 , n391311 , n43837 , n391313 , n391314 , n43840 , n391316 , n43842 , n43843 , 
 n43844 , n391320 , n43846 , n43847 , n391323 , n43849 , n391325 , n391326 , n43852 , n43853 , 
 n43854 , n43855 , n43856 , n43857 , n43858 , n391334 , n43860 , n391336 , n43862 , n43863 , 
 n391339 , n391340 , n43866 , n391342 , n391343 , n43869 , n391345 , n391346 , n43872 , n391348 , 
 n391349 , n391350 , n43876 , n391352 , n43878 , n391354 , n43880 , n391356 , n391357 , n43883 , 
 n43884 , n391360 , n391361 , n43887 , n391363 , n391364 , n43890 , n391366 , n391367 , n43893 , 
 n391369 , n391370 , n43896 , n391372 , n391373 , n43899 , n43900 , n391376 , n391377 , n43903 , 
 n43904 , n391380 , n43906 , n391382 , n43908 , n43909 , n43910 , n43911 , n391387 , n43913 , 
 n43914 , n391390 , n391391 , n43917 , n43918 , n391394 , n391395 , n43921 , n391397 , n43923 , 
 n391399 , n43925 , n43926 , n43927 , n43928 , n391404 , n391405 , n43931 , n43932 , n391408 , 
 n43934 , n391410 , n391411 , n43937 , n43938 , n391414 , n391415 , n391416 , n43942 , n391418 , 
 n43944 , n43945 , n391421 , n391422 , n43948 , n43949 , n391425 , n43951 , n43952 , n391428 , 
 n391429 , n391430 , n43956 , n391432 , n391433 , n43959 , n391435 , n391436 , n43962 , n391438 , 
 n43964 , n391440 , n391441 , n43967 , n391443 , n391444 , n43970 , n391446 , n391447 , n43973 , 
 n391449 , n43975 , n43976 , n391452 , n391453 , n43979 , n391455 , n391456 , n43982 , n391458 , 
 n391459 , n43985 , n391461 , n391462 , n391463 , n43994 , n391465 , n391466 , n43997 , n391468 , 
 n391469 , n391470 , n44001 , n391472 , n44003 , n44004 , n391475 , n44006 , n44007 , n391478 , 
 n44009 , n44010 , n391481 , n44012 , n391483 , n391484 , n44015 , n391486 , n391487 , n391488 , 
 n44019 , n391490 , n391491 , n44022 , n391493 , n391494 , n391495 , n44026 , n391497 , n391498 , 
 n44029 , n391500 , n391501 , n44032 , n391503 , n44034 , n391505 , n44036 , n391507 , n44038 , 
 n44039 , n391510 , n391511 , n44042 , n391513 , n391514 , n44045 , n391516 , n391517 , n44048 , 
 n44049 , n391520 , n391521 , n44052 , n391523 , n391524 , n44055 , n391526 , n391527 , n44058 , 
 n391529 , n391530 , n391531 , n391532 , n44063 , n391534 , n391535 , n44066 , n391537 , n391538 , 
 n44069 , n44070 , n391541 , n391542 , n44073 , n44074 , n44075 , n44076 , n44077 , n391548 , 
 n44079 , n391550 , n391551 , n44082 , n391553 , n44084 , n44085 , n44086 , n44087 , n44088 , 
 n44089 , n391560 , n391561 , n44092 , n391563 , n44094 , n44095 , n44096 , n391567 , n44098 , 
 n391569 , n44100 , n44101 , n44102 , n44103 , n44104 , n391575 , n391576 , n44107 , n391578 , 
 n44109 , n391580 , n44111 , n391582 , n44113 , n391584 , n44115 , n44116 , n391587 , n391588 , 
 n44119 , n391590 , n391591 , n44122 , n391593 , n391594 , n44125 , n391596 , n44127 , n44128 , 
 n391599 , n391600 , n44131 , n391602 , n391603 , n44134 , n391605 , n391606 , n44137 , n391608 , 
 n391609 , n44140 , n44141 , n44142 , n391613 , n391614 , n391615 , n44146 , n391617 , n44148 , 
 n44149 , n391620 , n391621 , n44152 , n391623 , n391624 , n44155 , n391626 , n391627 , n44158 , 
 n391629 , n44160 , n44161 , n391632 , n391633 , n44164 , n391635 , n391636 , n44167 , n391638 , 
 n391639 , n44170 , n391641 , n391642 , n44173 , n391644 , n391645 , n44176 , n391647 , n44178 , 
 n391649 , n391650 , n44181 , n391652 , n391653 , n44184 , n391655 , n391656 , n391657 , n391658 , 
 n44189 , n44190 , n391661 , n44192 , n44193 , n391664 , n391665 , n44196 , n391667 , n391668 , 
 n44199 , n44200 , n391671 , n391672 , n44203 , n44204 , n44205 , n391676 , n391677 , n44208 , 
 n44209 , n44210 , n391681 , n391682 , n44213 , n44214 , n44215 , n391686 , n391687 , n44218 , 
 n44219 , n44220 , n391691 , n391692 , n44223 , n44224 , n44225 , n391696 , n391697 , n44228 , 
 n391699 , n391700 , n44231 , n44232 , n44233 , n44234 , n44235 , n44236 , n44237 , n44238 , 
 n44239 , n391710 , n391711 , n391712 , n44243 , n391714 , n44245 , n391716 , n44247 , n44248 , 
 n391719 , n44250 , n391721 , n391722 , n391723 , n44254 , n391725 , n391726 , n44257 , n391728 , 
 n391729 , n44260 , n44261 , n391732 , n391733 , n44264 , n391735 , n391736 , n44267 , n391738 , 
 n391739 , n391740 , n391741 , n44277 , n391743 , n44279 , n44280 , n391746 , n391747 , n44283 , 
 n391749 , n391750 , n44286 , n391752 , n391753 , n44289 , n391755 , n391756 , n44292 , n391758 , 
 n391759 , n391760 , n44296 , n391762 , n44298 , n391764 , n44300 , n391766 , n44302 , n44303 , 
 n391769 , n391770 , n44306 , n391772 , n391773 , n44309 , n391775 , n391776 , n44312 , n391778 , 
 n44314 , n391780 , n44316 , n391782 , n391783 , n44319 , n44320 , n391786 , n391787 , n44323 , 
 n391789 , n44325 , n44326 , n391792 , n391793 , n44329 , n391795 , n391796 , n44332 , n391798 , 
 n391799 , n44335 , n391801 , n391802 , n44338 , n391804 , n391805 , n44341 , n391807 , n391808 , 
 n44344 , n44345 , n44346 , n44347 , n44348 , n391814 , n391815 , n44351 , n391817 , n391818 , 
 n44354 , n391820 , n44356 , n391822 , n44358 , n391824 , n44360 , n44361 , n391827 , n391828 , 
 n44364 , n391830 , n391831 , n44367 , n391833 , n391834 , n44370 , n44371 , n391837 , n391838 , 
 n44374 , n391840 , n391841 , n44377 , n391843 , n391844 , n44380 , n44381 , n44382 , n44383 , 
 n44384 , n44385 , n44386 , n391852 , n391853 , n44389 , n391855 , n44391 , n391857 , n44393 , 
 n391859 , n44395 , n391861 , n44397 , n44398 , n44399 , n44400 , n44401 , n44402 , n391868 , 
 n44404 , n391870 , n391871 , n391872 , n44408 , n391874 , n44410 , n391876 , n391877 , n44413 , 
 n391879 , n391880 , n44416 , n391882 , n391883 , n391884 , n44420 , n391886 , n44422 , n44423 , 
 n391889 , n44425 , n44426 , n391892 , n391893 , n44429 , n391895 , n391896 , n44432 , n391898 , 
 n391899 , n44435 , n391901 , n391902 , n44438 , n44439 , n391905 , n44441 , n391907 , n44443 , 
 n391909 , n391910 , n44446 , n391912 , n391913 , n44449 , n391915 , n44451 , n391917 , n391918 , 
 n44454 , n391920 , n391921 , n391922 , n44458 , n391924 , n391925 , n391926 , n44462 , n391928 , 
 n391929 , n44465 , n44466 , n391932 , n391933 , n44469 , n44470 , n391936 , n391937 , n44473 , 
 n391939 , n391940 , n44476 , n391942 , n391943 , n44479 , n391945 , n44481 , n44482 , n44483 , 
 n44484 , n44485 , n391951 , n44487 , n391953 , n44489 , n391955 , n44491 , n44492 , n391958 , 
 n44494 , n391960 , n391961 , n44497 , n44498 , n391964 , n391965 , n44501 , n44502 , n44503 , 
 n391969 , n391970 , n44506 , n44507 , n44508 , n391974 , n44510 , n391976 , n44512 , n44513 , 
 n44514 , n44515 , n44516 , n391982 , n44518 , n391984 , n44520 , n44521 , n391987 , n44523 , 
 n391989 , n391990 , n44526 , n391992 , n44528 , n391994 , n391995 , n44531 , n44532 , n391998 , 
 n391999 , n44535 , n392001 , n44537 , n392003 , n392004 , n44540 , n44541 , n392007 , n392008 , 
 n44544 , n392010 , n44546 , n392012 , n44548 , n44549 , n44550 , n44551 , n44552 , n44553 , 
 n392019 , n392020 , n44556 , n392022 , n392023 , n44559 , n392025 , n392026 , n392027 , n44563 , 
 n392029 , n44565 , n44566 , n392032 , n392033 , n44569 , n392035 , n392036 , n44572 , n392038 , 
 n392039 , n44575 , n392041 , n44577 , n44578 , n392044 , n392045 , n44581 , n392047 , n392048 , 
 n44584 , n392050 , n392051 , n44587 , n44588 , n44589 , n392055 , n392056 , n44592 , n392058 , 
 n44594 , n44595 , n44596 , n44597 , n44598 , n44599 , n392065 , n392066 , n44602 , n392068 , 
 n44604 , n44605 , n392071 , n392072 , n44608 , n392074 , n392075 , n44611 , n392077 , n392078 , 
 n44614 , n392080 , n44616 , n44617 , n392083 , n392084 , n44620 , n392086 , n392087 , n44623 , 
 n392089 , n392090 , n44626 , n392092 , n44628 , n392094 , n44630 , n44631 , n392097 , n392098 , 
 n44634 , n392100 , n392101 , n44637 , n392103 , n392104 , n44640 , n392106 , n44642 , n44643 , 
 n392109 , n44645 , n392111 , n392112 , n392113 , n44649 , n392115 , n392116 , n44652 , n392118 , 
 n392119 , n44655 , n44656 , n44657 , n392123 , n392124 , n44660 , n44661 , n44662 , n392128 , 
 n44664 , n44665 , n44666 , n392132 , n392133 , n44669 , n392135 , n44671 , n392137 , n44673 , 
 n44674 , n392140 , n44676 , n392142 , n44678 , n392144 , n392145 , n44681 , n44682 , n392148 , 
 n392149 , n44685 , n392151 , n392152 , n44688 , n392154 , n392155 , n392156 , n44692 , n392158 , 
 n392159 , n44695 , n392161 , n392162 , n44698 , n44699 , n44700 , n392166 , n392167 , n44703 , 
 n44704 , n44705 , n392171 , n392172 , n44708 , n392174 , n392175 , n392176 , n44712 , n392178 , 
 n392179 , n392180 , n44716 , n392182 , n392183 , n44719 , n392185 , n392186 , n44722 , n392188 , 
 n44724 , n44725 , n392191 , n44727 , n44728 , n44729 , n44730 , n44731 , n44732 , n44733 , 
 n44734 , n44735 , n44736 , n44737 , n44738 , n44739 , n44740 , n44741 , n44742 , n392208 , 
 n44744 , n392210 , n44746 , n392212 , n44748 , n392214 , n392215 , n44751 , n392217 , n392218 , 
 n392219 , n44755 , n392221 , n392222 , n44758 , n392224 , n392225 , n44761 , n44762 , n44763 , 
 n392229 , n44765 , n392231 , n44767 , n44768 , n44769 , n44770 , n44771 , n392237 , n44773 , 
 n44774 , n44775 , n44776 , n392242 , n44778 , n392244 , n392245 , n44781 , n392247 , n392248 , 
 n44784 , n392250 , n44786 , n44787 , n392253 , n392254 , n44790 , n392256 , n392257 , n44793 , 
 n392259 , n392260 , n44796 , n392262 , n392263 , n44799 , n392265 , n392266 , n44802 , n392268 , 
 n392269 , n44805 , n44806 , n44807 , n392273 , n392274 , n44810 , n44811 , n44812 , n392278 , 
 n44814 , n392280 , n44816 , n392282 , n392283 , n44819 , n392285 , n44821 , n392287 , n44823 , 
 n44824 , n44825 , n44826 , n44827 , n44828 , n392294 , n44830 , n392296 , n392297 , n44833 , 
 n392299 , n44835 , n392301 , n44837 , n44838 , n392304 , n392305 , n44841 , n392307 , n392308 , 
 n44844 , n392310 , n392311 , n392312 , n44848 , n44849 , n44850 , n392316 , n44852 , n392318 , 
 n392319 , n44855 , n392321 , n392322 , n44858 , n392324 , n44860 , n392326 , n44862 , n44863 , 
 n392329 , n44865 , n392331 , n44867 , n392333 , n392334 , n44870 , n44871 , n392337 , n392338 , 
 n44874 , n392340 , n392341 , n44877 , n392343 , n392344 , n392345 , n44881 , n392347 , n392348 , 
 n44884 , n392350 , n392351 , n44887 , n44888 , n392354 , n392355 , n44891 , n44892 , n44893 , 
 n392359 , n44895 , n392361 , n392362 , n44898 , n392364 , n392365 , n44901 , n44902 , n44903 , 
 n392369 , n44905 , n44906 , n392372 , n392373 , n44909 , n44910 , n44911 , n392377 , n392378 , 
 n44914 , n44915 , n392381 , n44917 , n392383 , n44919 , n392385 , n392386 , n44922 , n44923 , 
 n392389 , n44925 , n44926 , n392392 , n392393 , n44929 , n44930 , n392396 , n392397 , n44933 , 
 n392399 , n392400 , n44936 , n392402 , n392403 , n44939 , n392405 , n44941 , n392407 , n44943 , 
 n44944 , n44945 , n392411 , n392412 , n44948 , n392414 , n392415 , n44951 , n392417 , n392418 , 
 n44954 , n44955 , n392421 , n392422 , n44958 , n392424 , n392425 , n44961 , n392427 , n44963 , 
 n44964 , n44965 , n44966 , n44967 , n392433 , n44969 , n392435 , n44971 , n392437 , n44973 , 
 n44974 , n392440 , n44976 , n392442 , n44978 , n44979 , n392445 , n392446 , n44982 , n392448 , 
 n392449 , n44985 , n392451 , n392452 , n392453 , n44989 , n392455 , n392456 , n44992 , n392458 , 
 n392459 , n44995 , n44996 , n44997 , n392463 , n392464 , n45000 , n392466 , n392467 , n45003 , 
 n392469 , n392470 , n45006 , n45007 , n392473 , n45009 , n392475 , n392476 , n45012 , n392478 , 
 n45014 , n45015 , n45016 , n45017 , n392483 , n45019 , n392485 , n392486 , n45022 , n392488 , 
 n392489 , n45025 , n45026 , n45027 , n392493 , n392494 , n45030 , n392496 , n392497 , n45033 , 
 n392499 , n45035 , n45036 , n45037 , n392503 , n392504 , n45040 , n392506 , n392507 , n45043 , 
 n392509 , n45045 , n392511 , n392512 , n45048 , n392514 , n392515 , n45051 , n45052 , n392518 , 
 n45054 , n392520 , n392521 , n45057 , n392523 , n45059 , n45060 , n45061 , n45062 , n392528 , 
 n392529 , n45065 , n45066 , n45067 , n392533 , n45069 , n45070 , n392536 , n392537 , n45073 , 
 n392539 , n45075 , n45076 , n45077 , n45078 , n45079 , n392545 , n392546 , n45082 , n392548 , 
 n45084 , n392550 , n392551 , n45087 , n392553 , n45089 , n45090 , n45091 , n392557 , n45093 , 
 n392559 , n45095 , n45096 , n392562 , n45098 , n392564 , n45100 , n45101 , n45102 , n45103 , 
 n45104 , n45105 , n45106 , n392572 , n392573 , n45109 , n392575 , n392576 , n45112 , n392578 , 
 n392579 , n392580 , n45116 , n392582 , n45118 , n45119 , n392585 , n392586 , n45122 , n392588 , 
 n392589 , n45125 , n392591 , n392592 , n45128 , n392594 , n45130 , n45131 , n392597 , n392598 , 
 n45134 , n392600 , n392601 , n45137 , n392603 , n392604 , n45140 , n392606 , n45143 , n392608 , 
 n392609 , n45146 , n392611 , n392612 , n45149 , n392614 , n45151 , n45152 , n392617 , n392618 , 
 n45155 , n392620 , n392621 , n45158 , n392623 , n392624 , n45161 , n392626 , n392627 , n392628 , 
 n45170 , n392630 , n392631 , n45173 , n45174 , n392634 , n392635 , n45177 , n45178 , n45179 , 
 n392639 , n45181 , n45182 , n392642 , n392643 , n45185 , n392645 , n45187 , n45188 , n392648 , 
 n392649 , n45191 , n392651 , n392652 , n45194 , n392654 , n392655 , n45197 , n392657 , n45199 , 
 n392659 , n392660 , n45202 , n45203 , n392663 , n392664 , n45206 , n392666 , n392667 , n45209 , 
 n392669 , n392670 , n45212 , n392672 , n392673 , n45215 , n392675 , n392676 , n45218 , n45219 , 
 n45220 , n45221 , n45222 , n45223 , n45224 , n45225 , n392685 , n45227 , n45228 , n392688 , 
 n392689 , n392690 , n45232 , n45233 , n392693 , n45235 , n45236 , n392696 , n392697 , n45239 , 
 n392699 , n392700 , n45242 , n45243 , n392703 , n392704 , n45246 , n392706 , n392707 , n392708 , 
 n45250 , n392710 , n392711 , n392712 , n45254 , n392714 , n392715 , n45257 , n392717 , n392718 , 
 n45260 , n392720 , n45262 , n392722 , n45264 , n392724 , n45266 , n45267 , n392727 , n392728 , 
 n45270 , n392730 , n392731 , n45273 , n392733 , n392734 , n45276 , n45277 , n392737 , n392738 , 
 n45280 , n392740 , n392741 , n45283 , n392743 , n392744 , n45286 , n392746 , n392747 , n45289 , 
 n45290 , n45291 , n392751 , n392752 , n45294 , n45295 , n45296 , n392756 , n392757 , n45299 , 
 n45300 , n45301 , n392761 , n392762 , n45304 , n45305 , n45306 , n392766 , n392767 , n45309 , 
 n392769 , n45311 , n45312 , n45313 , n45314 , n45315 , n392775 , n45317 , n45318 , n392778 , 
 n392779 , n45321 , n392781 , n392782 , n45324 , n392784 , n392785 , n392786 , n45328 , n392788 , 
 n392789 , n45331 , n392791 , n45333 , n45334 , n392794 , n45336 , n392796 , n45338 , n45339 , 
 n392799 , n392800 , n45342 , n392802 , n392803 , n45345 , n392805 , n392806 , n392807 , n45349 , 
 n392809 , n392810 , n45352 , n392812 , n392813 , n45355 , n392815 , n45357 , n392817 , n45359 , 
 n392819 , n45361 , n45362 , n392822 , n392823 , n45365 , n392825 , n392826 , n45368 , n392828 , 
 n392829 , n45371 , n392831 , n392832 , n45374 , n392834 , n392835 , n45377 , n45378 , n392838 , 
 n45380 , n392840 , n45382 , n392842 , n392843 , n45385 , n392845 , n392846 , n45388 , n392848 , 
 n45390 , n45391 , n392851 , n392852 , n45394 , n45395 , n392855 , n45397 , n45398 , n392858 , 
 n392859 , n45401 , n45402 , n392862 , n392863 , n45405 , n392865 , n392866 , n45408 , n392868 , 
 n392869 , n45411 , n392871 , n392872 , n45414 , n392874 , n392875 , n392876 , n45418 , n392878 , 
 n392879 , n45421 , n392881 , n392882 , n45424 , n392884 , n392885 , n45427 , n392887 , n392888 , 
 n392889 , n45431 , n45432 , n392892 , n45434 , n45435 , n392895 , n392896 , n392897 , n45446 , 
 n392899 , n392900 , n45449 , n392902 , n392903 , n45452 , n392905 , n392906 , n45455 , n392908 , 
 n392909 , n45458 , n392911 , n45460 , n45461 , n392914 , n45463 , n392916 , n45465 , n392918 , 
 n45467 , n45468 , n392921 , n392922 , n45471 , n392924 , n392925 , n45474 , n392927 , n45476 , 
 n45477 , n45478 , n45479 , n45480 , n392933 , n45482 , n392935 , n392936 , n45485 , n45486 , 
 n392939 , n392940 , n45489 , n392942 , n45491 , n45492 , n392945 , n392946 , n45495 , n45496 , 
 n392949 , n392950 , n45499 , n392952 , n45501 , n392954 , n392955 , n392956 , n45505 , n45506 , 
 n392959 , n392960 , n45509 , n392962 , n392963 , n392964 , n45513 , n392966 , n45515 , n392968 , 
 n392969 , n45518 , n392971 , n45520 , n45521 , n45522 , n392975 , n392976 , n45525 , n392978 , 
 n45527 , n392980 , n392981 , n45530 , n392983 , n45532 , n392985 , n45534 , n392987 , n45536 , 
 n45537 , n45538 , n392991 , n392992 , n45541 , n45542 , n45543 , n392996 , n392997 , n392998 , 
 n45547 , n393000 , n45549 , n393002 , n45551 , n393004 , n45553 , n45554 , n45555 , n393008 , 
 n393009 , n45558 , n45559 , n45560 , n393013 , n393014 , n45563 , n45564 , n45565 , n393018 , 
 n393019 , n45568 , n393021 , n393022 , n45571 , n393024 , n45573 , n45574 , n393027 , n393028 , 
 n45577 , n393030 , n45579 , n45580 , n393033 , n393034 , n393035 , n45584 , n393037 , n45586 , 
 n45587 , n45588 , n45589 , n45590 , n45591 , n393044 , n393045 , n393046 , n45595 , n45596 , 
 n393049 , n45598 , n45599 , n393052 , n393053 , n45602 , n393055 , n45604 , n45605 , n45606 , 
 n45607 , n45608 , n45609 , n393062 , n393063 , n393064 , n393065 , n45614 , n393067 , n45616 , 
 n393069 , n393070 , n45619 , n393072 , n45621 , n45622 , n45623 , n45624 , n45625 , n45626 , 
 n393079 , n45628 , n45629 , n393082 , n393083 , n45632 , n393085 , n393086 , n45635 , n393088 , 
 n393089 , n393090 , n393091 , n45640 , n45641 , n393094 , n45643 , n45644 , n393097 , n393098 , 
 n45647 , n393100 , n45649 , n45650 , n45651 , n45652 , n45653 , n393106 , n393107 , n45656 , 
 n393109 , n393110 , n45659 , n393112 , n45661 , n45662 , n393115 , n45664 , n393117 , n45666 , 
 n45667 , n45668 , n45669 , n45670 , n45671 , n45672 , n393125 , n45674 , n393127 , n45676 , 
 n45677 , n45678 , n393131 , n45680 , n393133 , n45682 , n393135 , n393136 , n45685 , n45686 , 
 n393139 , n393140 , n45689 , n393142 , n393143 , n45692 , n393145 , n45694 , n45695 , n45696 , 
 n45697 , n45698 , n45699 , n393152 , n45701 , n393154 , n393155 , n45704 , n393157 , n45706 , 
 n45707 , n45708 , n45709 , n393162 , n45711 , n393164 , n45713 , n45714 , n45715 , n393168 , 
 n45717 , n393170 , n45719 , n393172 , n45721 , n45722 , n45723 , n45724 , n393177 , n45726 , 
 n393179 , n45728 , n45729 , n393182 , n393183 , n45732 , n393185 , n393186 , n45735 , n393188 , 
 n393189 , n45738 , n393191 , n45740 , n45741 , n45742 , n45743 , n45744 , n45745 , n45746 , 
 n393199 , n45748 , n393201 , n393202 , n45751 , n45752 , n393205 , n45754 , n45755 , n45756 , 
 n45757 , n393210 , n393211 , n45760 , n393213 , n45762 , n393215 , n45764 , n393217 , n45766 , 
 n393219 , n45768 , n393221 , n45770 , n45771 , n393224 , n393225 , n45774 , n393227 , n393228 , 
 n45777 , n393230 , n393231 , n45780 , n45781 , n393234 , n393235 , n45784 , n393237 , n393238 , 
 n45787 , n393240 , n393241 , n45790 , n45791 , n45792 , n393245 , n393246 , n45795 , n45796 , 
 n393249 , n393250 , n45799 , n45800 , n45801 , n393254 , n45803 , n393256 , n45805 , n393258 , 
 n45807 , n45808 , n393261 , n45810 , n393263 , n45812 , n45813 , n393266 , n393267 , n45816 , 
 n393269 , n393270 , n45819 , n393272 , n393273 , n393274 , n45823 , n393276 , n393277 , n45826 , 
 n393279 , n45828 , n45829 , n45830 , n45831 , n45832 , n393285 , n45834 , n45835 , n45836 , 
 n45837 , n45838 , n45839 , n45840 , n45841 , n393294 , n45843 , n393296 , n45845 , n45846 , 
 n393299 , n393300 , n45849 , n393302 , n393303 , n45852 , n393305 , n45854 , n45855 , n393308 , 
 n393309 , n45858 , n393311 , n45860 , n45861 , n45862 , n45863 , n393316 , n45865 , n45866 , 
 n45867 , n393320 , n393321 , n45870 , n45871 , n45872 , n393325 , n393326 , n45875 , n393328 , 
 n45877 , n45878 , n45879 , n45880 , n393333 , n45882 , n45883 , n45884 , n393337 , n393338 , 
 n45887 , n393340 , n45889 , n45890 , n393343 , n45892 , n45893 , n393346 , n45895 , n45896 , 
 n45897 , n393350 , n393351 , n45900 , n393353 , n393354 , n45903 , n393356 , n393357 , n393358 , 
 n45907 , n393360 , n393361 , n45910 , n393363 , n45912 , n393365 , n45914 , n393367 , n45916 , 
 n393369 , n393370 , n45919 , n393372 , n45921 , n393374 , n393375 , n45924 , n45925 , n393378 , 
 n393379 , n45928 , n393381 , n393382 , n45931 , n393384 , n393385 , n45934 , n393387 , n393388 , 
 n45937 , n393390 , n393391 , n45940 , n45941 , n45942 , n393395 , n45944 , n393397 , n45946 , 
 n45947 , n45948 , n45949 , n393402 , n45951 , n393404 , n393405 , n45954 , n393407 , n45956 , 
 n393409 , n393410 , n45959 , n393412 , n393413 , n45962 , n393415 , n393416 , n45965 , n393418 , 
 n393419 , n45968 , n45969 , n393422 , n45971 , n393424 , n45973 , n45974 , n393427 , n45976 , 
 n393429 , n45978 , n45979 , n393432 , n393433 , n45982 , n393435 , n393436 , n45985 , n393438 , 
 n393439 , n393440 , n45989 , n393442 , n393443 , n45992 , n393445 , n393446 , n45995 , n393448 , 
 n393449 , n393450 , n393451 , n46000 , n393453 , n393454 , n46003 , n393456 , n393457 , n46006 , 
 n393459 , n393460 , n46009 , n393462 , n46011 , n393464 , n393465 , n46014 , n393467 , n393468 , 
 n46017 , n46018 , n393471 , n46020 , n393473 , n46022 , n46023 , n46024 , n46025 , n46026 , 
 n46027 , n46028 , n46029 , n46030 , n46031 , n393484 , n393485 , n46034 , n393487 , n46036 , 
 n393489 , n46038 , n46039 , n46040 , n46041 , n46042 , n46043 , n393496 , n46045 , n46046 , 
 n393499 , n393500 , n46049 , n393502 , n393503 , n46052 , n393505 , n393506 , n46055 , n46056 , 
 n393509 , n46058 , n46059 , n46060 , n46061 , n46062 , n393515 , n46064 , n393517 , n46066 , 
 n393519 , n46068 , n46069 , n393522 , n393523 , n46072 , n393525 , n393526 , n46075 , n393528 , 
 n393529 , n46078 , n393531 , n393532 , n46081 , n393534 , n393535 , n46084 , n393537 , n393538 , 
 n46087 , n46088 , n46089 , n393542 , n46091 , n393544 , n393545 , n393546 , n46095 , n393548 , 
 n46097 , n393550 , n46099 , n46100 , n46101 , n46102 , n393555 , n46104 , n393557 , n393558 , 
 n46107 , n393560 , n46109 , n393562 , n393563 , n46112 , n393565 , n46114 , n46115 , n46116 , 
 n46117 , n46118 , n393571 , n46120 , n46121 , n46122 , n393575 , n393576 , n46125 , n393578 , 
 n46127 , n46128 , n393581 , n393582 , n46131 , n393584 , n393585 , n46134 , n393587 , n393588 , 
 n46137 , n393590 , n46139 , n393592 , n393593 , n46142 , n393595 , n393596 , n46145 , n46146 , 
 n393599 , n393600 , n46149 , n393602 , n393603 , n46152 , n393605 , n393606 , n46155 , n393608 , 
 n46157 , n46158 , n393611 , n46160 , n46161 , n393614 , n46163 , n46164 , n393617 , n393618 , 
 n46167 , n393620 , n393621 , n46170 , n393623 , n46172 , n46173 , n46174 , n46175 , n46176 , 
 n46177 , n46178 , n46179 , n393632 , n393633 , n46182 , n393635 , n46184 , n46185 , n393638 , 
 n393639 , n46188 , n393641 , n393642 , n46191 , n393644 , n393645 , n46194 , n393647 , n46196 , 
 n46197 , n46198 , n46199 , n46200 , n393653 , n46202 , n393655 , n393656 , n46205 , n46206 , 
 n46207 , n393660 , n393661 , n46210 , n46211 , n46212 , n393665 , n393666 , n46215 , n393668 , 
 n393669 , n46218 , n46219 , n393672 , n46221 , n393674 , n46223 , n46224 , n46225 , n46226 , 
 n393679 , n46228 , n393681 , n46230 , n46231 , n393684 , n393685 , n46234 , n393687 , n393688 , 
 n46237 , n393690 , n46239 , n46240 , n46241 , n46242 , n46243 , n46244 , n393697 , n46246 , 
 n393699 , n393700 , n46249 , n393702 , n393703 , n46252 , n46253 , n393706 , n46255 , n46256 , 
 n393709 , n46258 , n393711 , n46260 , n46261 , n46262 , n393715 , n393716 , n46265 , n393718 , 
 n393719 , n46268 , n46269 , n393722 , n393723 , n393724 , n393725 , n46274 , n393727 , n46276 , 
 n393729 , n46278 , n46279 , n393732 , n393733 , n46282 , n46283 , n46284 , n393737 , n393738 , 
 n46287 , n46288 , n393741 , n393742 , n46291 , n46292 , n46293 , n393746 , n46295 , n46296 , 
 n46297 , n393750 , n46299 , n46300 , n46301 , n393754 , n46303 , n46304 , n46305 , n46306 , 
 n393759 , n393760 , n393761 , n46310 , n46311 , n393764 , n46313 , n46314 , n393767 , n393768 , 
 n46317 , n393770 , n393771 , n393772 , n393773 , n46322 , n393775 , n46324 , n393777 , n393778 , 
 n46327 , n393780 , n46329 , n393782 , n46331 , n46332 , n393785 , n46334 , n393787 , n46336 , 
 n46337 , n393790 , n393791 , n46340 , n393793 , n393794 , n46343 , n393796 , n393797 , n393798 , 
 n46347 , n393800 , n393801 , n46350 , n393803 , n393804 , n46353 , n46354 , n46355 , n393808 , 
 n46357 , n46358 , n46359 , n46360 , n46361 , n46362 , n46363 , n46364 , n46365 , n46366 , 
 n46367 , n46368 , n46369 , n46370 , n393823 , n46372 , n393825 , n393826 , n46375 , n393828 , 
 n46377 , n393830 , n46379 , n46380 , n393833 , n393834 , n46383 , n393836 , n393837 , n46386 , 
 n393839 , n393840 , n46389 , n46390 , n393843 , n393844 , n46393 , n393846 , n393847 , n46396 , 
 n393849 , n46398 , n46399 , n46400 , n46401 , n46402 , n46403 , n46404 , n46405 , n46406 , 
 n46407 , n46408 , n46409 , n393862 , n46411 , n393864 , n393865 , n46414 , n393867 , n393868 , 
 n46417 , n393870 , n46419 , n46420 , n46421 , n393874 , n393875 , n46424 , n393877 , n393878 , 
 n46427 , n46428 , n393881 , n393882 , n393883 , n393884 , n46433 , n46434 , n393887 , n46436 , 
 n46437 , n393890 , n393891 , n46440 , n393893 , n393894 , n46443 , n393896 , n46445 , n46446 , 
 n393899 , n46448 , n393901 , n46450 , n393903 , n393904 , n46453 , n393906 , n393907 , n46456 , 
 n393909 , n393910 , n46459 , n46460 , n46461 , n46462 , n46463 , n46464 , n393917 , n46466 , 
 n393919 , n393920 , n393921 , n46470 , n393923 , n46472 , n46473 , n46474 , n46475 , n46476 , 
 n46477 , n46478 , n46479 , n46480 , n46481 , n46482 , n46483 , n393936 , n46485 , n393938 , 
 n46487 , n46488 , n393941 , n393942 , n46491 , n393944 , n393945 , n46494 , n393947 , n393948 , 
 n46497 , n393950 , n46499 , n393952 , n46501 , n393954 , n46503 , n46504 , n393957 , n46506 , 
 n393959 , n46508 , n46509 , n393962 , n46511 , n393964 , n46513 , n46514 , n393967 , n393968 , 
 n46517 , n393970 , n46519 , n393972 , n393973 , n46522 , n393975 , n393976 , n46525 , n393978 , 
 n46527 , n46528 , n46529 , n46530 , n46531 , n46532 , n393985 , n46534 , n393987 , n393988 , 
 n46537 , n46538 , n393991 , n46540 , n46541 , n393994 , n393995 , n46544 , n46545 , n393998 , 
 n393999 , n46548 , n394001 , n394002 , n46551 , n394004 , n46553 , n394006 , n394007 , n46556 , 
 n394009 , n46558 , n394011 , n46560 , n394013 , n394014 , n46563 , n394016 , n394017 , n46566 , 
 n394019 , n394020 , n46569 , n394022 , n46571 , n394024 , n46573 , n46574 , n394027 , n46576 , 
 n394029 , n46578 , n46579 , n394032 , n394033 , n46582 , n394035 , n394036 , n46585 , n394038 , 
 n394039 , n394040 , n46589 , n394042 , n394043 , n46592 , n394045 , n394046 , n46595 , n394048 , 
 n394049 , n46598 , n46599 , n46600 , n46601 , n46602 , n46603 , n46604 , n46605 , n46606 , 
 n46607 , n46608 , n46609 , n394062 , n46611 , n394064 , n394065 , n394066 , n46615 , n394068 , 
 n46617 , n394070 , n394071 , n46620 , n394073 , n394074 , n46623 , n46624 , n46625 , n394078 , 
 n394079 , n46628 , n46629 , n46630 , n394083 , n46632 , n46633 , n46634 , n394087 , n46636 , 
 n46637 , n46638 , n394091 , n394092 , n394093 , n46642 , n394095 , n46644 , n46645 , n394098 , 
 n46647 , n394100 , n46649 , n394102 , n394103 , n46652 , n394105 , n46654 , n46655 , n46656 , 
 n394109 , n394110 , n46659 , n394112 , n46661 , n394114 , n394115 , n46664 , n394117 , n394118 , 
 n46667 , n394120 , n394121 , n46670 , n46671 , n394124 , n46673 , n46674 , n394127 , n394128 , 
 n46677 , n46678 , n394131 , n394132 , n46681 , n394134 , n394135 , n46684 , n394137 , n394138 , 
 n46687 , n394140 , n394141 , n46690 , n394143 , n46692 , n394145 , n46694 , n46695 , n46696 , 
 n46697 , n46698 , n46699 , n46700 , n46701 , n46702 , n46703 , n46704 , n46705 , n46706 , 
 n46707 , n46708 , n46709 , n46710 , n46711 , n394164 , n46713 , n394166 , n46715 , n394168 , 
 n394169 , n46718 , n394171 , n394172 , n46721 , n394174 , n46723 , n394176 , n46725 , n46726 , 
 n394179 , n394180 , n46729 , n394182 , n394183 , n46732 , n394185 , n394186 , n46735 , n394188 , 
 n46737 , n46738 , n394191 , n394192 , n46741 , n394194 , n394195 , n46744 , n394197 , n394198 , 
 n46747 , n394200 , n394201 , n46750 , n394203 , n46752 , n394205 , n46754 , n394207 , n394208 , 
 n46757 , n394210 , n394211 , n46760 , n394213 , n46762 , n46763 , n394216 , n394217 , n46766 , 
 n394219 , n394220 , n46769 , n394222 , n394223 , n46772 , n394225 , n46781 , n46782 , n46783 , 
 n46784 , n394230 , n394231 , n46787 , n394233 , n46789 , n394235 , n46791 , n46792 , n46793 , 
 n394239 , n394240 , n46796 , n46797 , n46798 , n46799 , n46800 , n46801 , n46802 , n46803 , 
 n46804 , n46805 , n394251 , n46807 , n46808 , n46809 , n46810 , n46811 , n46812 , n46813 , 
 n46814 , n46815 , n46816 , n46817 , n394263 , n46819 , n46820 , n46821 , n394267 , n394268 , 
 n46824 , n394270 , n46826 , n394272 , n46828 , n394274 , n46830 , n46831 , n394277 , n394278 , 
 n46834 , n394280 , n394281 , n46837 , n394283 , n394284 , n46840 , n46841 , n394287 , n394288 , 
 n46844 , n394290 , n394291 , n46847 , n394293 , n394294 , n394295 , n46851 , n394297 , n46853 , 
 n46854 , n394300 , n46856 , n394302 , n46858 , n46859 , n394305 , n46861 , n394307 , n394308 , 
 n46864 , n394310 , n46866 , n394312 , n394313 , n46869 , n394315 , n394316 , n394317 , n46873 , 
 n394319 , n394320 , n46876 , n394322 , n394323 , n46879 , n46880 , n46881 , n46882 , n394328 , 
 n46884 , n394330 , n394331 , n394332 , n46888 , n46889 , n394335 , n46891 , n46892 , n394338 , 
 n46894 , n46895 , n46896 , n46897 , n46898 , n46899 , n394345 , n46901 , n394347 , n46903 , 
 n46904 , n394350 , n46906 , n394352 , n46908 , n394354 , n394355 , n46911 , n394357 , n46913 , 
 n46914 , n46915 , n46916 , n46917 , n46918 , n46919 , n46920 , n46921 , n46922 , n46923 , 
 n46924 , n46925 , n394371 , n46927 , n394373 , n46929 , n46930 , n394376 , n394377 , n46933 , 
 n394379 , n394380 , n46936 , n394382 , n46938 , n46939 , n46940 , n46941 , n394387 , n394388 , 
 n46944 , n394390 , n46946 , n394392 , n394393 , n46949 , n46950 , n394396 , n394397 , n46953 , 
 n394399 , n394400 , n46956 , n394402 , n394403 , n46959 , n394405 , n46961 , n46962 , n394408 , 
 n394409 , n46965 , n394411 , n394412 , n46968 , n394414 , n394415 , n46971 , n394417 , n46973 , 
 n394419 , n46975 , n46976 , n394422 , n46978 , n394424 , n46980 , n394426 , n394427 , n46983 , 
 n46984 , n394430 , n394431 , n46987 , n394433 , n394434 , n46990 , n394436 , n394437 , n394438 , 
 n46994 , n394440 , n394441 , n46997 , n394443 , n394444 , n47000 , n47001 , n47002 , n394448 , 
 n394449 , n47005 , n394451 , n394452 , n47008 , n394454 , n47010 , n394456 , n47012 , n394458 , 
 n47014 , n47015 , n394461 , n47017 , n394463 , n394464 , n394465 , n47021 , n394467 , n394468 , 
 n47024 , n394470 , n394471 , n47027 , n47028 , n394474 , n394475 , n47031 , n394477 , n394478 , 
 n47034 , n394480 , n394481 , n47037 , n47038 , n394484 , n394485 , n47041 , n394487 , n47043 , 
 n394489 , n47045 , n47046 , n394492 , n394493 , n47049 , n394495 , n394496 , n47052 , n394498 , 
 n394499 , n47055 , n394501 , n47057 , n47058 , n394504 , n394505 , n47061 , n394507 , n394508 , 
 n47064 , n394510 , n394511 , n47067 , n47068 , n394514 , n394515 , n47071 , n394517 , n47073 , 
 n394519 , n47075 , n47076 , n394522 , n394523 , n47079 , n394525 , n394526 , n47082 , n394528 , 
 n394529 , n47085 , n394531 , n47087 , n47088 , n394534 , n47090 , n394536 , n47092 , n394538 , 
 n394539 , n47095 , n394541 , n394542 , n47098 , n47099 , n47100 , n394546 , n394547 , n47103 , 
 n394549 , n394550 , n47106 , n394552 , n394553 , n47109 , n47110 , n47111 , n394557 , n394558 , 
 n47114 , n47115 , n47116 , n394562 , n394563 , n47119 , n394565 , n47121 , n47122 , n47123 , 
 n394569 , n394570 , n47126 , n394572 , n47128 , n394574 , n47130 , n394576 , n394577 , n47133 , 
 n394579 , n47135 , n47136 , n394582 , n394583 , n47139 , n394585 , n47141 , n47142 , n47143 , 
 n47144 , n47145 , n47146 , n47147 , n47148 , n394594 , n47150 , n394596 , n394597 , n47153 , 
 n47154 , n394600 , n394601 , n47157 , n47158 , n394604 , n47160 , n47161 , n394607 , n394608 , 
 n394609 , n47165 , n394611 , n394612 , n47168 , n47169 , n394615 , n47171 , n47172 , n394618 , 
 n394619 , n47175 , n47176 , n47177 , n47178 , n47179 , n47180 , n47181 , n47182 , n47183 , 
 n394629 , n47185 , n394631 , n394632 , n47188 , n394634 , n47190 , n394636 , n394637 , n47193 , 
 n47194 , n394640 , n394641 , n47197 , n394643 , n394644 , n47200 , n394646 , n47202 , n47203 , 
 n47204 , n394650 , n394651 , n47207 , n394653 , n47209 , n47210 , n47211 , n394657 , n47213 , 
 n394659 , n47215 , n394661 , n47217 , n394663 , n394664 , n47220 , n394666 , n394667 , n394668 , 
 n47224 , n47225 , n394671 , n47227 , n47228 , n394674 , n47230 , n47231 , n47232 , n394678 , 
 n47234 , n394680 , n47236 , n47237 , n394683 , n394684 , n47240 , n47241 , n394687 , n47243 , 
 n47244 , n47245 , n394691 , n47247 , n394693 , n47249 , n47250 , n394696 , n394697 , n394698 , 
 n47254 , n47255 , n47256 , n394702 , n47258 , n47259 , n394705 , n394706 , n47262 , n394708 , 
 n394709 , n47265 , n47266 , n394712 , n394713 , n47269 , n394715 , n394716 , n394717 , n47273 , 
 n394719 , n47275 , n394721 , n394722 , n47278 , n394724 , n394725 , n47281 , n394727 , n394728 , 
 n394729 , n47285 , n394731 , n47287 , n47288 , n394734 , n47290 , n394736 , n47292 , n394738 , 
 n394739 , n47295 , n394741 , n394742 , n47298 , n394744 , n47300 , n47301 , n394747 , n47303 , 
 n394749 , n47305 , n394751 , n394752 , n47308 , n394754 , n394755 , n47311 , n394757 , n47313 , 
 n394759 , n47315 , n394761 , n47317 , n47318 , n394764 , n394765 , n47321 , n47322 , n394768 , 
 n394769 , n47325 , n47326 , n394772 , n394773 , n47329 , n47330 , n394776 , n394777 , n47333 , 
 n47334 , n47335 , n394781 , n394782 , n47338 , n394784 , n394785 , n47341 , n394787 , n47343 , 
 n394789 , n47345 , n394791 , n47347 , n47348 , n394794 , n394795 , n47351 , n394797 , n394798 , 
 n47354 , n394800 , n394801 , n47357 , n47358 , n394804 , n394805 , n47361 , n394807 , n394808 , 
 n47364 , n394810 , n47366 , n394812 , n47368 , n394814 , n394815 , n47371 , n394817 , n394818 , 
 n47374 , n394820 , n47376 , n47377 , n394823 , n394824 , n47380 , n394826 , n394827 , n47383 , 
 n394829 , n394830 , n394831 , n47393 , n394833 , n394834 , n47396 , n394836 , n47398 , n47399 , 
 n394839 , n394840 , n47402 , n394842 , n394843 , n47405 , n394845 , n47407 , n394847 , n47409 , 
 n47410 , n47411 , n47412 , n394852 , n47414 , n394854 , n47416 , n394856 , n394857 , n47419 , 
 n394859 , n394860 , n47422 , n47423 , n394863 , n394864 , n47426 , n394866 , n394867 , n47429 , 
 n394869 , n394870 , n47432 , n394872 , n47434 , n47435 , n394875 , n47437 , n394877 , n47439 , 
 n394879 , n47441 , n47442 , n394882 , n47444 , n394884 , n394885 , n47447 , n394887 , n47449 , 
 n47450 , n394890 , n394891 , n47453 , n394893 , n394894 , n47456 , n394896 , n394897 , n394898 , 
 n47460 , n394900 , n394901 , n47463 , n394903 , n394904 , n47466 , n394906 , n394907 , n47469 , 
 n47470 , n394910 , n47472 , n47473 , n394913 , n394914 , n47476 , n394916 , n47478 , n47479 , 
 n394919 , n394920 , n47482 , n47483 , n394923 , n394924 , n47486 , n394926 , n394927 , n47489 , 
 n47490 , n394930 , n47492 , n394932 , n47494 , n394934 , n394935 , n47497 , n394937 , n394938 , 
 n47500 , n394940 , n394941 , n47503 , n394943 , n394944 , n47506 , n47507 , n47508 , n394948 , 
 n47510 , n394950 , n394951 , n394952 , n394953 , n394954 , n394955 , n47517 , n394957 , n394958 , 
 n47520 , n394960 , n394961 , n47523 , n394963 , n394964 , n47526 , n394966 , n394967 , n47529 , 
 n47530 , n394970 , n47532 , n47533 , n394973 , n394974 , n394975 , n47537 , n394977 , n394978 , 
 n47540 , n47541 , n394981 , n47543 , n394983 , n47545 , n394985 , n47547 , n47548 , n394988 , 
 n394989 , n47551 , n394991 , n394992 , n47554 , n394994 , n394995 , n47557 , n47558 , n394998 , 
 n394999 , n47561 , n395001 , n395002 , n47564 , n395004 , n395005 , n47567 , n395007 , n47569 , 
 n395009 , n47571 , n47572 , n395012 , n395013 , n47575 , n47576 , n395016 , n395017 , n47579 , 
 n395019 , n47581 , n47582 , n395022 , n395023 , n47585 , n47586 , n395026 , n395027 , n47589 , 
 n395029 , n395030 , n47592 , n47593 , n395033 , n395034 , n47596 , n47597 , n47598 , n395038 , 
 n395039 , n47601 , n395041 , n395042 , n47604 , n395044 , n395045 , n47607 , n395047 , n395048 , 
 n395049 , n47611 , n395051 , n47613 , n395053 , n395054 , n47616 , n395056 , n47618 , n47619 , 
 n47620 , n395060 , n47622 , n47623 , n47624 , n47625 , n47626 , n47627 , n47628 , n395068 , 
 n395069 , n47631 , n395071 , n395072 , n47634 , n395074 , n395075 , n47637 , n47638 , n395078 , 
 n47640 , n47641 , n395081 , n395082 , n47644 , n47645 , n395085 , n395086 , n47648 , n395088 , 
 n47650 , n395090 , n47652 , n395092 , n47654 , n47655 , n395095 , n395096 , n47658 , n395098 , 
 n395099 , n47661 , n395101 , n395102 , n47664 , n47665 , n395105 , n395106 , n47668 , n395108 , 
 n395109 , n47671 , n395111 , n395112 , n47674 , n47675 , n395115 , n395116 , n47678 , n47679 , 
 n47680 , n395120 , n395121 , n47683 , n395123 , n47685 , n47686 , n395126 , n395127 , n47689 , 
 n395129 , n395130 , n47692 , n395132 , n395133 , n47695 , n395135 , n47697 , n47698 , n395138 , 
 n395139 , n47701 , n395141 , n395142 , n47704 , n395144 , n395145 , n47707 , n395147 , n47709 , 
 n395149 , n47711 , n395151 , n47713 , n47714 , n395154 , n395155 , n47717 , n395157 , n395158 , 
 n47720 , n395160 , n395161 , n47723 , n47724 , n395164 , n47726 , n395166 , n47728 , n395168 , 
 n395169 , n47731 , n395171 , n395172 , n47734 , n47735 , n395175 , n395176 , n47738 , n47739 , 
 n395179 , n47741 , n395181 , n47743 , n47744 , n395184 , n395185 , n47747 , n395187 , n395188 , 
 n47750 , n395190 , n47752 , n47753 , n47754 , n47755 , n47756 , n47757 , n395197 , n47759 , 
 n395199 , n47761 , n47762 , n395202 , n395203 , n47765 , n395205 , n47767 , n47768 , n395208 , 
 n47770 , n395210 , n47772 , n47773 , n395213 , n395214 , n47776 , n47777 , n395217 , n395218 , 
 n47780 , n395220 , n47782 , n395222 , n395223 , n47785 , n395225 , n395226 , n47788 , n47789 , 
 n47790 , n47791 , n47792 , n47793 , n395233 , n47795 , n395235 , n47797 , n47798 , n395238 , 
 n47800 , n395240 , n47802 , n395242 , n395243 , n47805 , n395245 , n395246 , n47808 , n47809 , 
 n47810 , n395250 , n395251 , n47813 , n395253 , n395254 , n47816 , n395256 , n395257 , n47819 , 
 n395259 , n47821 , n395261 , n47823 , n47824 , n395264 , n47826 , n395266 , n47828 , n47829 , 
 n395269 , n395270 , n47832 , n395272 , n395273 , n47835 , n395275 , n395276 , n395277 , n47839 , 
 n395279 , n395280 , n47842 , n395282 , n395283 , n47845 , n47846 , n47847 , n395287 , n395288 , 
 n47850 , n395290 , n395291 , n47853 , n395293 , n395294 , n47856 , n47857 , n47858 , n395298 , 
 n47860 , n395300 , n47862 , n47863 , n395303 , n47865 , n395305 , n47867 , n47868 , n395308 , 
 n47870 , n395310 , n47872 , n395312 , n395313 , n47875 , n395315 , n395316 , n47878 , n395318 , 
 n395319 , n47881 , n395321 , n395322 , n395323 , n47885 , n395325 , n395326 , n47888 , n395328 , 
 n47890 , n47891 , n395331 , n47893 , n395333 , n395334 , n395335 , n47897 , n395337 , n395338 , 
 n395339 , n47901 , n395341 , n47903 , n47904 , n395344 , n47906 , n395346 , n395347 , n47909 , 
 n395349 , n395350 , n47912 , n395352 , n395353 , n395354 , n47916 , n395356 , n395357 , n47919 , 
 n395359 , n395360 , n47922 , n395362 , n395363 , n47925 , n395365 , n395366 , n47928 , n395368 , 
 n395369 , n47931 , n395371 , n395372 , n395373 , n47935 , n395375 , n47937 , n47938 , n395378 , 
 n47940 , n395380 , n47942 , n47943 , n395383 , n395384 , n47946 , n395386 , n395387 , n47949 , 
 n395389 , n395390 , n395391 , n47953 , n395393 , n395394 , n47956 , n395396 , n395397 , n47959 , 
 n47960 , n47961 , n47962 , n395402 , n47964 , n395404 , n47966 , n47967 , n395407 , n395408 , 
 n47970 , n395410 , n395411 , n47973 , n395413 , n395414 , n395415 , n47977 , n395417 , n47979 , 
 n395419 , n47981 , n47982 , n47983 , n395423 , n47985 , n47986 , n395426 , n47988 , n395428 , 
 n47990 , n47991 , n47992 , n395432 , n47994 , n395434 , n47996 , n47997 , n395437 , n395438 , 
 n48000 , n395440 , n48002 , n48003 , n395443 , n395444 , n48006 , n395446 , n395447 , n48009 , 
 n395449 , n395450 , n48012 , n395452 , n395453 , n48015 , n395455 , n395456 , n48018 , n395458 , 
 n395459 , n48021 , n48022 , n48023 , n48024 , n48025 , n48026 , n48027 , n395467 , n48029 , 
 n395469 , n48031 , n48032 , n395472 , n48034 , n48035 , n395475 , n395476 , n48038 , n395478 , 
 n395479 , n48041 , n395481 , n48043 , n48044 , n395484 , n395485 , n48047 , n48048 , n395488 , 
 n395489 , n48051 , n395491 , n395492 , n48054 , n48055 , n395495 , n395496 , n48058 , n395498 , 
 n395499 , n395500 , n48062 , n395502 , n48064 , n395504 , n395505 , n48067 , n395507 , n395508 , 
 n48070 , n395510 , n48072 , n48073 , n395513 , n395514 , n48076 , n395516 , n395517 , n48079 , 
 n395519 , n48081 , n48082 , n48083 , n395523 , n395524 , n48086 , n395526 , n48088 , n48089 , 
 n48090 , n48091 , n48092 , n48093 , n48094 , n48095 , n48096 , n48097 , n48098 , n48099 , 
 n48100 , n48101 , n48102 , n48103 , n48104 , n48105 , n48106 , n48107 , n395547 , n48109 , 
 n48110 , n48111 , n48112 , n48113 , n395553 , n48115 , n48116 , n48117 , n48118 , n48119 , 
 n48120 , n395560 , n48122 , n48123 , n48124 , n395564 , n48126 , n395566 , n395567 , n48129 , 
 n48130 , n395570 , n48132 , n48133 , n395573 , n48135 , n48136 , n48137 , n48138 , n48139 , 
 n48140 , n395580 , n48142 , n48143 , n395583 , n48145 , n48146 , n48147 , n48148 , n395588 , 
 n48150 , n48151 , n48152 , n48153 , n48154 , n48155 , n48156 , n48157 , n48158 , n48159 , 
 n48160 , n48161 , n48162 , n48163 , n395603 , n48165 , n395605 , n48167 , n395607 , n48169 , 
 n395609 , n395610 , n48172 , n395612 , n395613 , n48175 , n48176 , n48177 , n395617 , n395618 , 
 n48180 , n48181 , n48182 , n395622 , n48184 , n395624 , n48186 , n48187 , n48188 , n48189 , 
 n48190 , n48191 , n395631 , n48193 , n48194 , n48195 , n48196 , n48197 , n395637 , n48199 , 
 n48200 , n48201 , n48202 , n48203 , n48204 , n48205 , n48206 , n48207 , n395647 , n48209 , 
 n48210 , n48211 , n48212 , n48213 , n48214 , n48215 , n48216 , n48217 , n395657 , n395658 , 
 n48220 , n48221 , n48222 , n48223 , n395663 , n395664 , n395665 , n48227 , n395667 , n48229 , 
 n395669 , n48231 , n48232 , n48233 , n48234 , n395674 , n395675 , n48237 , n395677 , n395678 , 
 n48240 , n395680 , n395681 , n48243 , n48244 , n395684 , n395685 , n48247 , n395687 , n395688 , 
 n48250 , n395690 , n395691 , n48253 , n48254 , n48255 , n48256 , n395696 , n395697 , n48259 , 
 n48260 , n395700 , n48262 , n395702 , n48264 , n48265 , n395705 , n395706 , n48268 , n48269 , 
 n395709 , n48271 , n48272 , n48275 , n395713 , n48277 , n395715 , n48279 , n48280 , n395718 , 
 n395719 , n395720 , n48284 , n395722 , n395723 , n48287 , n48288 , n395726 , n48290 , n48291 , 
 n395729 , n395730 , n48294 , n395732 , n395733 , n48297 , n395735 , n395736 , n48300 , n395738 , 
 n395739 , n395740 , n48304 , n395742 , n48306 , n48307 , n395745 , n395746 , n48310 , n395748 , 
 n48312 , n48313 , n395751 , n395752 , n48316 , n395754 , n395755 , n48319 , n395757 , n395758 , 
 n48322 , n395760 , n395761 , n48325 , n395763 , n395764 , n48328 , n395766 , n48330 , n48331 , 
 n395769 , n48333 , n395771 , n395772 , n48336 , n395774 , n48338 , n395776 , n48340 , n395778 , 
 n48342 , n48343 , n395781 , n395782 , n48346 , n395784 , n395785 , n48349 , n395787 , n395788 , 
 n48352 , n48353 , n395791 , n395792 , n48356 , n395794 , n395795 , n48359 , n395797 , n395798 , 
 n395799 , n48363 , n395801 , n48365 , n48366 , n48367 , n48368 , n48369 , n48370 , n395808 , 
 n48372 , n395810 , n48374 , n395812 , n395813 , n48377 , n395815 , n395816 , n48380 , n395818 , 
 n395819 , n48383 , n395821 , n48385 , n395823 , n48387 , n48388 , n395826 , n48390 , n395828 , 
 n48392 , n395830 , n395831 , n48395 , n48396 , n395834 , n395835 , n48399 , n395837 , n395838 , 
 n48402 , n395840 , n395841 , n395842 , n48406 , n395844 , n395845 , n48409 , n395847 , n395848 , 
 n48412 , n395850 , n395851 , n395852 , n48416 , n395854 , n48418 , n48419 , n48420 , n48421 , 
 n48422 , n48423 , n395861 , n395862 , n48426 , n395864 , n395865 , n48429 , n395867 , n395868 , 
 n48432 , n395870 , n395871 , n48435 , n395873 , n395874 , n48438 , n395876 , n395877 , n48441 , 
 n395879 , n395880 , n48444 , n48445 , n395883 , n48447 , n395885 , n395886 , n48450 , n48451 , 
 n395889 , n395890 , n395891 , n48455 , n48456 , n395894 , n395895 , n395896 , n48460 , n395898 , 
 n48462 , n48463 , n48464 , n48465 , n48466 , n48467 , n48468 , n48469 , n48470 , n48471 , 
 n395909 , n48473 , n395911 , n395912 , n48476 , n395914 , n395915 , n48479 , n395917 , n48481 , 
 n395919 , n395920 , n48484 , n48485 , n395923 , n395924 , n48488 , n395926 , n395927 , n48491 , 
 n395929 , n395930 , n48494 , n395932 , n395933 , n48497 , n48498 , n395936 , n395937 , n48501 , 
 n395939 , n395940 , n48504 , n395942 , n395943 , n48507 , n395945 , n395946 , n48510 , n48511 , 
 n48512 , n48513 , n48514 , n395952 , n395953 , n48517 , n395955 , n48519 , n395957 , n48521 , 
 n395959 , n48523 , n48524 , n48525 , n48526 , n395964 , n395965 , n48529 , n395967 , n48531 , 
 n48532 , n48533 , n48534 , n395972 , n48536 , n395974 , n48538 , n48539 , n395977 , n395978 , 
 n48542 , n395980 , n395981 , n48545 , n395983 , n395984 , n395985 , n48549 , n395987 , n48551 , 
 n48552 , n48553 , n48554 , n48555 , n48556 , n395994 , n48558 , n395996 , n48560 , n48561 , 
 n395999 , n396000 , n48564 , n396002 , n396003 , n48567 , n396005 , n48569 , n48570 , n48571 , 
 n396009 , n48573 , n48574 , n48575 , n48576 , n48577 , n396015 , n396016 , n48580 , n396018 , 
 n396019 , n48583 , n396021 , n48585 , n48586 , n48587 , n48588 , n48589 , n48590 , n396028 , 
 n396029 , n48593 , n48594 , n48595 , n48596 , n396034 , n396035 , n48599 , n396037 , n48601 , 
 n396039 , n48603 , n48604 , n396042 , n48606 , n396044 , n48608 , n48609 , n396047 , n48611 , 
 n396049 , n396050 , n48614 , n396052 , n396053 , n48617 , n48618 , n48619 , n48620 , n48621 , 
 n48622 , n48623 , n48624 , n48625 , n48626 , n396064 , n48628 , n396066 , n48630 , n396068 , 
 n48632 , n396070 , n48634 , n48635 , n48636 , n396074 , n48638 , n396076 , n396077 , n48641 , 
 n48642 , n396080 , n396081 , n48645 , n396083 , n396084 , n48648 , n396086 , n396087 , n48651 , 
 n396089 , n396090 , n396091 , n48655 , n396093 , n48657 , n48658 , n396096 , n48660 , n396098 , 
 n396099 , n396100 , n396101 , n48665 , n396103 , n396104 , n48668 , n396106 , n396107 , n48671 , 
 n48672 , n48673 , n48674 , n48675 , n396113 , n396114 , n396115 , n48679 , n396117 , n48681 , 
 n48682 , n396120 , n48684 , n396122 , n48686 , n48687 , n396125 , n396126 , n48690 , n396128 , 
 n396129 , n48693 , n396131 , n396132 , n396133 , n48697 , n396135 , n396136 , n48700 , n396138 , 
 n396139 , n48703 , n48704 , n48705 , n48706 , n48707 , n396145 , n396146 , n48710 , n396148 , 
 n396149 , n48713 , n48714 , n48715 , n48716 , n48717 , n396155 , n48719 , n48720 , n396158 , 
 n396159 , n48723 , n396161 , n396162 , n48726 , n396164 , n48728 , n48729 , n48730 , n48731 , 
 n48732 , n396170 , n48734 , n396172 , n48736 , n396174 , n396175 , n48739 , n396177 , n48741 , 
 n396179 , n48743 , n396181 , n396182 , n48746 , n396184 , n396185 , n48749 , n396187 , n48751 , 
 n48752 , n48753 , n396191 , n48755 , n396193 , n48757 , n48758 , n396196 , n396197 , n48761 , 
 n396199 , n396200 , n48764 , n396202 , n396203 , n48767 , n396205 , n48769 , n48770 , n48771 , 
 n48772 , n48773 , n48774 , n48775 , n48776 , n48777 , n48778 , n48779 , n48780 , n396218 , 
 n48782 , n396220 , n48784 , n396222 , n48786 , n396224 , n48788 , n48789 , n396227 , n396228 , 
 n48792 , n396230 , n396231 , n48795 , n396233 , n396234 , n48798 , n396236 , n48800 , n48801 , 
 n396239 , n48803 , n396241 , n48805 , n396243 , n396244 , n48808 , n396246 , n396247 , n48811 , 
 n396249 , n48813 , n396251 , n48815 , n48816 , n396254 , n396255 , n48819 , n396257 , n396258 , 
 n48822 , n396260 , n396261 , n48825 , n396263 , n48827 , n48828 , n48829 , n48830 , n396268 , 
 n48832 , n396270 , n396271 , n48835 , n48836 , n396274 , n396275 , n48839 , n48840 , n48841 , 
 n396279 , n48843 , n396281 , n396282 , n48846 , n396284 , n396285 , n48849 , n48850 , n396288 , 
 n396289 , n48853 , n396291 , n48855 , n396293 , n48857 , n48858 , n396296 , n48860 , n396298 , 
 n396299 , n396300 , n48864 , n396302 , n396303 , n48867 , n396305 , n48869 , n48870 , n48871 , 
 n48872 , n48873 , n396311 , n48875 , n48876 , n48877 , n396315 , n48879 , n48880 , n396318 , 
 n48882 , n396320 , n48884 , n396322 , n396323 , n48887 , n48888 , n396326 , n396327 , n48891 , 
 n396329 , n48893 , n396331 , n396332 , n48896 , n396334 , n396335 , n48899 , n396337 , n48901 , 
 n396339 , n48903 , n396341 , n48905 , n48906 , n396344 , n396345 , n48909 , n396347 , n396348 , 
 n48912 , n396350 , n396351 , n48915 , n48916 , n396354 , n48918 , n396356 , n48920 , n396358 , 
 n396359 , n48923 , n396361 , n396362 , n396363 , n396364 , n48928 , n396366 , n396367 , n396368 , 
 n48932 , n48933 , n396371 , n48935 , n396373 , n396374 , n48938 , n48939 , n396377 , n48941 , 
 n48942 , n48943 , n396381 , n396382 , n48946 , n396384 , n48948 , n48949 , n396387 , n396388 , 
 n48952 , n396390 , n396391 , n48955 , n396393 , n48957 , n48958 , n48959 , n396397 , n48961 , 
 n396399 , n48963 , n396401 , n48965 , n396403 , n48967 , n396405 , n48969 , n396407 , n48971 , 
 n396409 , n48973 , n48974 , n396412 , n396413 , n48977 , n396415 , n396416 , n48980 , n396418 , 
 n396419 , n48983 , n48984 , n396422 , n396423 , n48987 , n396425 , n396426 , n48990 , n396428 , 
 n396429 , n48993 , n396431 , n396432 , n48996 , n48997 , n48998 , n48999 , n49000 , n49001 , 
 n49002 , n49003 , n396441 , n49005 , n396443 , n396444 , n49008 , n396446 , n49010 , n396448 , 
 n49012 , n49013 , n396451 , n49015 , n396453 , n49017 , n49018 , n396456 , n396457 , n49021 , 
 n396459 , n396460 , n49024 , n396462 , n396463 , n396464 , n49028 , n396466 , n396467 , n49031 , 
 n396469 , n396470 , n49034 , n49035 , n49036 , n396474 , n396475 , n49039 , n49040 , n396478 , 
 n49042 , n396480 , n49044 , n396482 , n396483 , n49047 , n49048 , n49049 , n49050 , n396488 , 
 n49052 , n396490 , n49054 , n396492 , n49056 , n396494 , n49058 , n49059 , n396497 , n49061 , 
 n396499 , n49063 , n396501 , n396502 , n49066 , n396504 , n396505 , n49069 , n49070 , n396508 , 
 n396509 , n49073 , n396511 , n396512 , n49076 , n396514 , n396515 , n49079 , n49080 , n396518 , 
 n396519 , n49083 , n396521 , n49085 , n396523 , n49087 , n49088 , n396526 , n396527 , n49091 , 
 n396529 , n49093 , n49094 , n396532 , n49096 , n396534 , n396535 , n49099 , n396537 , n396538 , 
 n49102 , n396540 , n49104 , n396542 , n396543 , n49107 , n396545 , n396546 , n49110 , n396548 , 
 n396549 , n49113 , n396551 , n396552 , n49116 , n49117 , n396555 , n49119 , n396557 , n49121 , 
 n49122 , n396560 , n49124 , n396562 , n49126 , n396564 , n396565 , n49129 , n396567 , n396568 , 
 n396569 , n49138 , n396571 , n396572 , n49141 , n396574 , n396575 , n49144 , n396577 , n49146 , 
 n396579 , n49148 , n49149 , n396582 , n396583 , n49152 , n396585 , n396586 , n49155 , n396588 , 
 n396589 , n49158 , n396591 , n396592 , n49161 , n396594 , n49163 , n49164 , n396597 , n49166 , 
 n396599 , n49168 , n396601 , n396602 , n49171 , n396604 , n396605 , n49174 , n396607 , n49176 , 
 n396609 , n49178 , n49179 , n396612 , n396613 , n49182 , n396615 , n396616 , n49185 , n396618 , 
 n396619 , n396620 , n49189 , n396622 , n396623 , n49192 , n396625 , n396626 , n49195 , n396628 , 
 n396629 , n49198 , n396631 , n396632 , n49201 , n396634 , n396635 , n49204 , n49205 , n396638 , 
 n49207 , n396640 , n396641 , n49210 , n396643 , n49212 , n49213 , n49214 , n396647 , n49216 , 
 n396649 , n49218 , n49219 , n396652 , n396653 , n49222 , n49223 , n396656 , n49225 , n49226 , 
 n49227 , n396660 , n49229 , n396662 , n49231 , n396664 , n49233 , n396666 , n49235 , n396668 , 
 n396669 , n49238 , n396671 , n396672 , n49241 , n49242 , n49243 , n396676 , n396677 , n49246 , 
 n396679 , n396680 , n49249 , n396682 , n396683 , n49252 , n396685 , n396686 , n49255 , n396688 , 
 n396689 , n49258 , n396691 , n49260 , n49261 , n49262 , n49263 , n49264 , n49265 , n49266 , 
 n49267 , n49268 , n49269 , n49270 , n49271 , n49272 , n49273 , n49274 , n49275 , n396708 , 
 n49277 , n49278 , n49279 , n49280 , n49281 , n396714 , n49283 , n396716 , n49285 , n396718 , 
 n49287 , n49288 , n49289 , n49290 , n49291 , n49292 , n49293 , n396726 , n49295 , n396728 , 
 n49297 , n49298 , n396731 , n396732 , n49301 , n49302 , n49303 , n396736 , n49305 , n396738 , 
 n49307 , n396740 , n49309 , n396742 , n49311 , n49312 , n396745 , n396746 , n49315 , n396748 , 
 n396749 , n49318 , n396751 , n396752 , n49321 , n49322 , n396755 , n49324 , n396757 , n49326 , 
 n396759 , n396760 , n49329 , n396762 , n396763 , n49332 , n396765 , n49334 , n49335 , n396768 , 
 n49337 , n396770 , n49339 , n49340 , n396773 , n49342 , n396775 , n49344 , n396777 , n396778 , 
 n49347 , n396780 , n396781 , n396782 , n49351 , n396784 , n396785 , n49354 , n396787 , n49356 , 
 n49357 , n49358 , n396791 , n396792 , n49361 , n396794 , n49363 , n396796 , n49365 , n396798 , 
 n49367 , n49368 , n49369 , n49370 , n49371 , n49372 , n49373 , n49374 , n49375 , n49376 , 
 n49377 , n49378 , n49379 , n49380 , n49381 , n49382 , n49383 , n49384 , n49385 , n49386 , 
 n396819 , n396820 , n49389 , n396822 , n49391 , n396824 , n396825 , n396826 , n49395 , n396828 , 
 n49397 , n396830 , n49399 , n49400 , n396833 , n396834 , n49403 , n396836 , n396837 , n49406 , 
 n396839 , n396840 , n49409 , n49410 , n396843 , n396844 , n49413 , n396846 , n396847 , n49416 , 
 n396849 , n396850 , n49419 , n49420 , n49421 , n396854 , n396855 , n49424 , n49425 , n49426 , 
 n396859 , n396860 , n49429 , n396862 , n49431 , n396864 , n49433 , n396866 , n49435 , n396868 , 
 n396869 , n49438 , n49439 , n396872 , n396873 , n49442 , n396875 , n396876 , n49445 , n396878 , 
 n396879 , n49448 , n396881 , n49450 , n396883 , n49452 , n49453 , n396886 , n49455 , n396888 , 
 n49457 , n49458 , n396891 , n396892 , n49461 , n396894 , n396895 , n49464 , n396897 , n396898 , 
 n396899 , n49468 , n396901 , n396902 , n49471 , n396904 , n396905 , n49474 , n49475 , n49476 , 
 n396909 , n396910 , n49479 , n49480 , n396913 , n396914 , n49483 , n49484 , n49485 , n396918 , 
 n49487 , n396920 , n396921 , n49490 , n396923 , n49492 , n396925 , n49494 , n396927 , n49496 , 
 n49497 , n396930 , n49499 , n396932 , n49501 , n49502 , n396935 , n396936 , n49505 , n396938 , 
 n396939 , n49508 , n396941 , n396942 , n396943 , n49512 , n396945 , n396946 , n49515 , n396948 , 
 n49517 , n396950 , n49519 , n396952 , n49521 , n396954 , n49523 , n49524 , n49525 , n396958 , 
 n396959 , n49528 , n396961 , n396962 , n49531 , n396964 , n396965 , n49534 , n49535 , n396968 , 
 n396969 , n49538 , n396971 , n396972 , n49541 , n396974 , n396975 , n49544 , n396977 , n49546 , 
 n49547 , n396980 , n396981 , n49550 , n49551 , n396984 , n49553 , n49554 , n396987 , n396988 , 
 n49557 , n396990 , n49559 , n49560 , n396993 , n396994 , n49563 , n396996 , n396997 , n49566 , 
 n396999 , n49568 , n49569 , n397002 , n49571 , n397004 , n49573 , n397006 , n49575 , n49576 , 
 n397009 , n397010 , n49579 , n397012 , n397013 , n49582 , n397015 , n397016 , n49585 , n397018 , 
 n49587 , n49588 , n397021 , n397022 , n49591 , n397024 , n397025 , n49594 , n397027 , n397028 , 
 n49597 , n49598 , n397031 , n49600 , n397033 , n397034 , n49603 , n397036 , n49605 , n49606 , 
 n397039 , n49608 , n397041 , n49610 , n49611 , n397044 , n397045 , n49614 , n397047 , n397048 , 
 n49617 , n397050 , n397051 , n49620 , n397053 , n49622 , n49623 , n397056 , n49625 , n397058 , 
 n49627 , n397060 , n397061 , n49630 , n397063 , n49632 , n49633 , n49634 , n397067 , n49636 , 
 n397069 , n397070 , n49639 , n397072 , n49641 , n49642 , n397075 , n49644 , n397077 , n397078 , 
 n397079 , n49648 , n397081 , n49650 , n49651 , n49652 , n49653 , n397086 , n49655 , n397088 , 
 n49657 , n49658 , n397091 , n49660 , n49661 , n397094 , n49663 , n397096 , n397097 , n49666 , 
 n397099 , n397100 , n49669 , n397102 , n49671 , n49672 , n397105 , n397106 , n49675 , n397108 , 
 n49677 , n49678 , n49679 , n397112 , n49681 , n397114 , n397115 , n49684 , n397117 , n49686 , 
 n397119 , n49688 , n397121 , n49690 , n49691 , n397124 , n397125 , n49694 , n397127 , n397128 , 
 n49697 , n397130 , n397131 , n49700 , n397133 , n397134 , n49703 , n397136 , n49705 , n397138 , 
 n397139 , n397140 , n49709 , n49710 , n397143 , n397144 , n49713 , n49714 , n49715 , n397148 , 
 n397149 , n49718 , n397151 , n49720 , n49721 , n397154 , n397155 , n49724 , n397157 , n397158 , 
 n49727 , n397160 , n397161 , n49730 , n397163 , n49732 , n397165 , n397166 , n49735 , n49736 , 
 n397169 , n397170 , n49739 , n397172 , n397173 , n49742 , n397175 , n49744 , n49745 , n49746 , 
 n49747 , n49748 , n397181 , n49750 , n397183 , n397184 , n49753 , n397186 , n49755 , n49756 , 
 n397189 , n397190 , n49759 , n397192 , n49761 , n49762 , n397195 , n397196 , n49765 , n49766 , 
 n49767 , n49768 , n397201 , n397202 , n49771 , n397204 , n49773 , n49774 , n397207 , n49776 , 
 n397209 , n397210 , n49779 , n397212 , n49781 , n397214 , n397215 , n49784 , n49785 , n397218 , 
 n49787 , n49788 , n397221 , n397222 , n397223 , n49792 , n397225 , n397226 , n49795 , n49796 , 
 n397229 , n49798 , n49799 , n397232 , n397233 , n49802 , n397235 , n49804 , n49805 , n49806 , 
 n49807 , n49808 , n397241 , n49810 , n397243 , n397244 , n397245 , n49814 , n397247 , n49816 , 
 n49817 , n397250 , n397251 , n49820 , n397253 , n397254 , n49823 , n397256 , n397257 , n49826 , 
 n397259 , n49828 , n49829 , n49830 , n397263 , n49832 , n397265 , n397266 , n49835 , n397268 , 
 n49837 , n397270 , n49839 , n397272 , n49841 , n49842 , n397275 , n49844 , n397277 , n397278 , 
 n397279 , n49848 , n397281 , n397282 , n49851 , n397284 , n397285 , n49854 , n49855 , n397288 , 
 n397289 , n49858 , n397291 , n397292 , n49861 , n397294 , n397295 , n49864 , n49865 , n49866 , 
 n397299 , n49868 , n49869 , n397302 , n49871 , n49872 , n397305 , n49874 , n49875 , n49876 , 
 n397309 , n49878 , n49879 , n49880 , n397313 , n397314 , n49883 , n397316 , n49885 , n49886 , 
 n49887 , n49888 , n49889 , n49890 , n397323 , n49892 , n49893 , n49894 , n49895 , n49896 , 
 n49897 , n49898 , n49899 , n49900 , n397333 , n49902 , n49903 , n49904 , n397337 , n49906 , 
 n49907 , n49908 , n49909 , n49910 , n49911 , n49912 , n49913 , n397346 , n397347 , n49916 , 
 n397349 , n49918 , n397351 , n397352 , n49921 , n49922 , n49923 , n49924 , n397357 , n49926 , 
 n49927 , n397360 , n49929 , n397362 , n49931 , n49932 , n49933 , n49934 , n49935 , n397368 , 
 n49937 , n49938 , n397371 , n49940 , n397373 , n49942 , n397375 , n49944 , n49945 , n397378 , 
 n397379 , n49948 , n397381 , n397382 , n49951 , n397384 , n397385 , n49954 , n397387 , n397388 , 
 n49957 , n397390 , n49959 , n49960 , n49961 , n49962 , n49963 , n397396 , n49965 , n49966 , 
 n397399 , n397400 , n49969 , n397402 , n397403 , n49972 , n397405 , n49974 , n397407 , n49976 , 
 n49977 , n397410 , n49979 , n397412 , n49981 , n49982 , n397415 , n49984 , n397417 , n49986 , 
 n397419 , n397420 , n49989 , n49990 , n397423 , n397424 , n49993 , n397426 , n397427 , n49996 , 
 n397429 , n397430 , n397431 , n50000 , n397433 , n397434 , n50003 , n397436 , n50005 , n397438 , 
 n397439 , n50008 , n397441 , n50010 , n397443 , n397444 , n50013 , n397446 , n50015 , n50016 , 
 n397449 , n50018 , n397451 , n50020 , n50021 , n50022 , n397455 , n50024 , n397457 , n50026 , 
 n50027 , n397460 , n50029 , n397462 , n50031 , n50032 , n397465 , n397466 , n50035 , n397468 , 
 n397469 , n50038 , n397471 , n397472 , n50041 , n397474 , n50043 , n397476 , n397477 , n50046 , 
 n397479 , n397480 , n50049 , n397482 , n397483 , n397484 , n50053 , n397486 , n397487 , n50056 , 
 n397489 , n397490 , n50059 , n397492 , n397493 , n50062 , n397495 , n397496 , n50065 , n397498 , 
 n397499 , n50068 , n397501 , n50070 , n50071 , n397504 , n397505 , n50074 , n397507 , n397508 , 
 n50077 , n397510 , n397511 , n397512 , n50086 , n397514 , n397515 , n50089 , n397517 , n397518 , 
 n50092 , n50093 , n50094 , n397522 , n50096 , n397524 , n50098 , n50099 , n397527 , n50101 , 
 n397529 , n50103 , n50104 , n397532 , n397533 , n50107 , n397535 , n397536 , n50110 , n397538 , 
 n397539 , n50113 , n50114 , n50115 , n397543 , n50117 , n50118 , n397546 , n50120 , n397548 , 
 n397549 , n50123 , n397551 , n397552 , n397553 , n397554 , n50128 , n397556 , n397557 , n50131 , 
 n397559 , n397560 , n50134 , n50135 , n50136 , n50137 , n397565 , n50139 , n397567 , n50141 , 
 n397569 , n397570 , n50144 , n397572 , n50146 , n397574 , n50148 , n50149 , n50150 , n397578 , 
 n50152 , n397580 , n397581 , n50155 , n397583 , n50157 , n50158 , n50159 , n50160 , n397588 , 
 n50162 , n397590 , n397591 , n50165 , n397593 , n50167 , n50168 , n397596 , n50170 , n50171 , 
 n50172 , n397600 , n50174 , n397602 , n397603 , n50177 , n397605 , n50179 , n397607 , n50181 , 
 n50182 , n50183 , n50184 , n397612 , n397613 , n50187 , n50188 , n50189 , n397617 , n397618 , 
 n50192 , n397620 , n397621 , n50195 , n397623 , n397624 , n50198 , n50199 , n50200 , n50201 , 
 n50202 , n397630 , n397631 , n50205 , n397633 , n397634 , n50208 , n397636 , n397637 , n50211 , 
 n50212 , n397640 , n397641 , n397642 , n50216 , n50217 , n397645 , n50219 , n50220 , n397648 , 
 n397649 , n50223 , n397651 , n50225 , n397653 , n397654 , n397655 , n50229 , n397657 , n397658 , 
 n50232 , n50233 , n397661 , n397662 , n397663 , n397664 , n50238 , n397666 , n50240 , n397668 , 
 n397669 , n50243 , n397671 , n50245 , n50246 , n50247 , n50248 , n397676 , n50250 , n397678 , 
 n397679 , n50253 , n397681 , n397682 , n50256 , n50257 , n397685 , n397686 , n50260 , n50261 , 
 n50262 , n397690 , n397691 , n50265 , n397693 , n397694 , n397695 , n50269 , n397697 , n397698 , 
 n397699 , n50273 , n397701 , n397702 , n50276 , n397704 , n397705 , n50279 , n50280 , n397708 , 
 n50282 , n397710 , n397711 , n50285 , n50286 , n397714 , n50288 , n50289 , n397717 , n50291 , 
 n397719 , n50293 , n50294 , n397722 , n397723 , n50297 , n50298 , n397726 , n397727 , n397728 , 
 n50302 , n397730 , n397731 , n50305 , n50306 , n397734 , n50308 , n50309 , n397737 , n50311 , 
 n50312 , n50313 , n50314 , n397742 , n50316 , n50317 , n397745 , n50319 , n50320 , n397748 , 
 n397749 , n50323 , n397751 , n397752 , n50326 , n397754 , n397755 , n397756 , n50330 , n397758 , 
 n50332 , n50333 , n50334 , n50335 , n397763 , n50337 , n397765 , n50339 , n50340 , n397768 , 
 n397769 , n50343 , n397771 , n397772 , n50346 , n397774 , n50348 , n50349 , n50350 , n50351 , 
 n397779 , n50353 , n397781 , n50355 , n50356 , n50357 , n397785 , n50359 , n397787 , n50361 , 
 n50362 , n397790 , n50364 , n397792 , n50366 , n397794 , n397795 , n50369 , n397797 , n50371 , 
 n50372 , n397800 , n397801 , n50375 , n397803 , n50377 , n50378 , n397806 , n397807 , n50381 , 
 n397809 , n50383 , n397811 , n397812 , n50386 , n50387 , n50388 , n50389 , n397817 , n397818 , 
 n50392 , n397820 , n50394 , n50395 , n50396 , n397824 , n50398 , n397826 , n50400 , n397828 , 
 n50402 , n397830 , n50404 , n50405 , n397833 , n397834 , n50408 , n397836 , n397837 , n50411 , 
 n397839 , n397840 , n50414 , n397842 , n397843 , n50417 , n397845 , n50419 , n50420 , n50421 , 
 n50422 , n397850 , n50424 , n397852 , n50426 , n50427 , n50428 , n50429 , n50430 , n397858 , 
 n397859 , n50433 , n397861 , n50435 , n50436 , n50437 , n397865 , n397866 , n50440 , n397868 , 
 n50442 , n50443 , n50444 , n50445 , n397873 , n50447 , n397875 , n397876 , n50450 , n397878 , 
 n397879 , n50453 , n397881 , n50455 , n50456 , n397884 , n50458 , n397886 , n50460 , n397888 , 
 n50462 , n397890 , n50464 , n397892 , n397893 , n50467 , n397895 , n50469 , n397897 , n397898 , 
 n50472 , n50473 , n50474 , n50475 , n50476 , n50477 , n397905 , n50479 , n50480 , n397908 , 
 n50482 , n397910 , n50484 , n50485 , n397913 , n397914 , n50488 , n50489 , n397917 , n50491 , 
 n50492 , n397920 , n397921 , n397922 , n50496 , n397924 , n397925 , n50499 , n397927 , n50501 , 
 n397929 , n397930 , n50504 , n397932 , n50506 , n397934 , n50508 , n50509 , n397937 , n397938 , 
 n50512 , n397940 , n397941 , n50515 , n397943 , n397944 , n50518 , n397946 , n50520 , n397948 , 
 n397949 , n50523 , n397951 , n50525 , n50526 , n397954 , n50530 , n397956 , n50532 , n50533 , 
 n50547 , n50553 , n50554 , n50555 , n50557 , n50561 , n50562 , n50563 , n50564 , n397968 , 
 n50566 , n50567 , n50568 , n50569 , n50570 , n50571 , n50572 , n50573 , n50574 , n50575 , 
 n50576 , n50577 , n50578 , n50579 , n50580 , n397984 , n50582 , n50583 , n50584 , n397988 , 
 n50586 , n397990 , n397991 , n50589 , n397993 , n50591 , n50592 , n397996 , n397997 , n50595 , 
 n397999 , n398000 , n50598 , n398002 , n398003 , n50601 , n398005 , n50603 , n50604 , n398008 , 
 n50606 , n398010 , n50608 , n398012 , n50610 , n398014 , n50612 , n398016 , n398017 , n50615 , 
 n398019 , n50617 , n398021 , n398022 , n50620 , n398024 , n398025 , n50623 , n50624 , n398028 , 
 n50626 , n398030 , n398031 , n50629 , n398033 , n50631 , n50632 , n50633 , n50634 , n398038 , 
 n398039 , n50637 , n398041 , n398042 , n50640 , n398044 , n398045 , n50643 , n398047 , n50645 , 
 n398049 , n50647 , n398051 , n50649 , n50650 , n398054 , n50652 , n398056 , n398057 , n50655 , 
 n398059 , n398060 , n50658 , n50659 , n398063 , n398064 , n50662 , n398066 , n398067 , n50665 , 
 n398069 , n398070 , n50668 , n398072 , n398073 , n50671 , n50672 , n50673 , n398077 , n50675 , 
 n398079 , n398080 , n50678 , n398082 , n50680 , n398084 , n50682 , n50683 , n50684 , n398088 , 
 n50686 , n50687 , n50688 , n50689 , n50690 , n50691 , n50692 , n398096 , n398097 , n50695 , 
 n398099 , n50697 , n398101 , n50699 , n50700 , n50701 , n398105 , n398106 , n50704 , n398108 , 
 n398109 , n50707 , n398111 , n50709 , n50710 , n398114 , n50712 , n398116 , n398117 , n50715 , 
 n398119 , n50717 , n50718 , n398122 , n398123 , n50721 , n398125 , n398126 , n50724 , n398128 , 
 n398129 , n398130 , n50728 , n50729 , n398133 , n398134 , n50732 , n398136 , n50734 , n398138 , 
 n50736 , n50737 , n398141 , n398142 , n50740 , n398144 , n398145 , n50743 , n398147 , n398148 , 
 n50746 , n398150 , n50748 , n50749 , n50750 , n50751 , n50752 , n398156 , n50754 , n50755 , 
 n398159 , n50757 , n398161 , n50759 , n50760 , n398164 , n50762 , n398166 , n50764 , n50765 , 
 n398169 , n398170 , n50768 , n398172 , n398173 , n50771 , n398175 , n398176 , n398177 , n50775 , 
 n398179 , n398180 , n50778 , n398182 , n398183 , n50781 , n398185 , n398186 , n50784 , n398188 , 
 n50786 , n398190 , n50788 , n398192 , n50790 , n398194 , n398195 , n50793 , n398197 , n398198 , 
 n50796 , n50797 , n398201 , n398202 , n50800 , n50801 , n398205 , n398206 , n398207 , n50805 , 
 n398209 , n50807 , n50808 , n398212 , n50810 , n398214 , n50812 , n50813 , n398217 , n398218 , 
 n50816 , n398220 , n398221 , n50819 , n398223 , n398224 , n398225 , n50823 , n398227 , n398228 , 
 n50826 , n398230 , n398231 , n50829 , n398233 , n398234 , n50832 , n398236 , n50834 , n50835 , 
 n398239 , n398240 , n50838 , n398242 , n398243 , n50841 , n398245 , n398246 , n50844 , n398248 , 
 n50846 , n50847 , n50848 , n398252 , n50850 , n398254 , n50852 , n398256 , n398257 , n398258 , 
 n50856 , n398260 , n50858 , n50859 , n398263 , n398264 , n50862 , n398266 , n398267 , n50865 , 
 n398269 , n398270 , n50868 , n398272 , n50870 , n50871 , n398275 , n398276 , n50874 , n398278 , 
 n398279 , n50877 , n398281 , n398282 , n50880 , n398284 , n50882 , n398286 , n50884 , n50885 , 
 n50886 , n398290 , n50888 , n398292 , n50890 , n50891 , n398295 , n398296 , n50894 , n398298 , 
 n398299 , n50897 , n398301 , n50899 , n398303 , n398304 , n50902 , n398306 , n398307 , n50905 , 
 n398309 , n398310 , n50908 , n50909 , n50910 , n398314 , n398315 , n50913 , n50914 , n50915 , 
 n398319 , n398320 , n50918 , n398322 , n50920 , n398324 , n398325 , n50923 , n398327 , n398328 , 
 n50926 , n50927 , n398331 , n50929 , n50930 , n398334 , n398335 , n50933 , n50934 , n398338 , 
 n398339 , n50937 , n398341 , n398342 , n50940 , n398344 , n398345 , n50943 , n50944 , n50945 , 
 n398349 , n398350 , n50948 , n50949 , n50950 , n50951 , n50952 , n398356 , n50954 , n50955 , 
 n398359 , n50957 , n398361 , n50959 , n50960 , n398364 , n50962 , n398366 , n398367 , n398368 , 
 n50966 , n398370 , n398371 , n50969 , n398373 , n50971 , n50972 , n398376 , n398377 , n50975 , 
 n398379 , n50977 , n398381 , n50979 , n50980 , n398384 , n398385 , n50983 , n50984 , n50985 , 
 n398389 , n398390 , n50988 , n398392 , n50990 , n50991 , n50992 , n398396 , n398397 , n50995 , 
 n398399 , n398400 , n398401 , n398402 , n51000 , n398404 , n51002 , n398406 , n51004 , n51005 , 
 n398409 , n398410 , n51008 , n398412 , n51010 , n51011 , n398415 , n51013 , n398417 , n51015 , 
 n51016 , n398420 , n398421 , n51019 , n398423 , n398424 , n51022 , n398426 , n398427 , n51025 , 
 n398429 , n51027 , n398431 , n398432 , n51030 , n51031 , n398435 , n398436 , n51034 , n398438 , 
 n398439 , n51037 , n398441 , n51039 , n51040 , n51041 , n398445 , n51043 , n398447 , n398448 , 
 n51046 , n398450 , n398451 , n51049 , n398453 , n398454 , n398455 , n398456 , n51054 , n398458 , 
 n398459 , n51057 , n398461 , n398462 , n51060 , n398464 , n398465 , n51063 , n398467 , n398468 , 
 n51066 , n398470 , n398471 , n398472 , n398473 , n51071 , n398475 , n51073 , n51074 , n51075 , 
 n51076 , n51077 , n398481 , n51079 , n51080 , n398484 , n398485 , n51083 , n398487 , n398488 , 
 n51086 , n51087 , n398491 , n51089 , n51090 , n398494 , n398495 , n51093 , n398497 , n51095 , 
 n398499 , n398500 , n51098 , n51099 , n398503 , n398504 , n51102 , n398506 , n398507 , n51105 , 
 n398509 , n398510 , n398511 , n51109 , n51110 , n398514 , n51112 , n51113 , n398517 , n51115 , 
 n51116 , n51117 , n51118 , n51119 , n51120 , n398524 , n51122 , n51123 , n51124 , n398528 , 
 n51126 , n51127 , n398531 , n51129 , n398533 , n398534 , n398535 , n51133 , n398537 , n51135 , 
 n51136 , n398540 , n51138 , n398542 , n398543 , n398544 , n51142 , n398546 , n398547 , n51145 , 
 n398549 , n398550 , n51148 , n398552 , n398553 , n51151 , n398555 , n398556 , n51154 , n51155 , 
 n51156 , n398560 , n51158 , n51159 , n51160 , n51161 , n51162 , n51163 , n51164 , n51165 , 
 n51166 , n51167 , n398571 , n398572 , n51170 , n398574 , n51172 , n51173 , n51174 , n51175 , 
 n51176 , n51177 , n51178 , n51179 , n51180 , n51181 , n51182 , n51183 , n51184 , n51185 , 
 n398589 , n398590 , n51188 , n51189 , n398593 , n51191 , n51192 , n398596 , n398597 , n398598 , 
 n51202 , n398600 , n398601 , n51205 , n398603 , n398604 , n398605 , n51209 , n398607 , n51211 , 
 n51212 , n51213 , n51214 , n51215 , n51216 , n51217 , n398615 , n398616 , n51220 , n398618 , 
 n398619 , n51223 , n398621 , n398622 , n51226 , n398624 , n51228 , n398626 , n398627 , n51231 , 
 n51232 , n398630 , n51234 , n51235 , n398633 , n398634 , n51238 , n51239 , n398637 , n398638 , 
 n51242 , n398640 , n398641 , n51245 , n398643 , n398644 , n398645 , n51249 , n398647 , n51251 , 
 n398649 , n51253 , n51254 , n398652 , n398653 , n51257 , n398655 , n398656 , n51260 , n398658 , 
 n398659 , n51263 , n51264 , n398662 , n398663 , n51267 , n398665 , n398666 , n51270 , n398668 , 
 n398669 , n51273 , n398671 , n398672 , n51276 , n398674 , n398675 , n51279 , n398677 , n51281 , 
 n398679 , n51283 , n398681 , n51285 , n51286 , n398684 , n398685 , n51289 , n398687 , n398688 , 
 n51292 , n398690 , n398691 , n51295 , n51296 , n51297 , n398695 , n51299 , n398697 , n398698 , 
 n51302 , n51303 , n51304 , n398702 , n398703 , n51307 , n51308 , n51309 , n398707 , n51311 , 
 n398709 , n51313 , n398711 , n51315 , n398713 , n398714 , n51318 , n51319 , n398717 , n398718 , 
 n51322 , n51323 , n398721 , n51325 , n398723 , n51327 , n51328 , n398726 , n398727 , n51331 , 
 n398729 , n51333 , n51334 , n51335 , n51336 , n51337 , n51338 , n398736 , n51340 , n398738 , 
 n51342 , n398740 , n398741 , n51345 , n51346 , n51347 , n398745 , n51349 , n398747 , n398748 , 
 n51352 , n398750 , n51354 , n51355 , n398753 , n398754 , n51358 , n398756 , n398757 , n51361 , 
 n398759 , n398760 , n51364 , n398762 , n398763 , n51367 , n51368 , n398766 , n51370 , n51371 , 
 n398769 , n51373 , n51374 , n398772 , n51376 , n398774 , n398775 , n51379 , n51380 , n51381 , 
 n51382 , n51383 , n51384 , n51385 , n398783 , n51387 , n398785 , n51389 , n398787 , n51391 , 
 n398789 , n51393 , n398791 , n398792 , n51396 , n398794 , n51398 , n51399 , n51400 , n51401 , 
 n51402 , n51403 , n51404 , n398802 , n51406 , n51407 , n398805 , n51409 , n398807 , n398808 , 
 n51412 , n398810 , n51414 , n398812 , n398813 , n51417 , n51418 , n51419 , n398817 , n51421 , 
 n398819 , n398820 , n51424 , n51425 , n398823 , n51427 , n51428 , n398826 , n398827 , n51431 , 
 n51432 , n398830 , n51434 , n398832 , n51436 , n398834 , n398835 , n51439 , n398837 , n51441 , 
 n398839 , n51443 , n398841 , n398842 , n51446 , n398844 , n398845 , n51449 , n398847 , n398848 , 
 n51452 , n398850 , n398851 , n51455 , n398853 , n398854 , n51458 , n398856 , n51460 , n51461 , 
 n398859 , n51463 , n398861 , n51465 , n51466 , n51467 , n51468 , n398866 , n398867 , n51471 , 
 n398869 , n51473 , n398871 , n51475 , n398873 , n398874 , n51478 , n398876 , n398877 , n51481 , 
 n398879 , n51483 , n51484 , n398882 , n398883 , n51487 , n398885 , n398886 , n51490 , n398888 , 
 n398889 , n51493 , n398891 , n51495 , n51496 , n51497 , n51498 , n398896 , n51500 , n398898 , 
 n51502 , n51503 , n51504 , n398902 , n51506 , n51507 , n51508 , n51509 , n51510 , n398908 , 
 n51512 , n398910 , n51514 , n51515 , n51516 , n51517 , n51518 , n51519 , n51520 , n51521 , 
 n51522 , n51523 , n51524 , n51525 , n398923 , n398924 , n51528 , n398926 , n51530 , n398928 , 
 n398929 , n51533 , n398931 , n51535 , n398933 , n51537 , n51538 , n398936 , n51540 , n398938 , 
 n398939 , n398940 , n51544 , n398942 , n398943 , n51547 , n398945 , n398946 , n51550 , n51551 , 
 n398949 , n51553 , n398951 , n51555 , n398953 , n398954 , n398955 , n398956 , n398957 , n51561 , 
 n398959 , n398960 , n51564 , n51565 , n51566 , n398964 , n51568 , n51569 , n51570 , n398968 , 
 n398969 , n51573 , n398971 , n398972 , n51576 , n398974 , n398975 , n51579 , n398977 , n51581 , 
 n398979 , n398980 , n51584 , n51585 , n398983 , n51587 , n398985 , n51589 , n398987 , n398988 , 
 n51592 , n51593 , n51594 , n51595 , n398993 , n51597 , n51598 , n51599 , n398997 , n51601 , 
 n398999 , n51603 , n51604 , n399002 , n399003 , n51607 , n399005 , n399006 , n51610 , n399008 , 
 n399009 , n399010 , n51614 , n399012 , n51616 , n51617 , n399015 , n51619 , n399017 , n51621 , 
 n51622 , n399020 , n399021 , n51625 , n399023 , n399024 , n51628 , n399026 , n399027 , n51631 , 
 n399029 , n51633 , n399031 , n399032 , n51636 , n51637 , n399035 , n399036 , n51640 , n399038 , 
 n399039 , n51643 , n399041 , n51645 , n399043 , n51647 , n51648 , n399046 , n51650 , n51651 , 
 n51652 , n399050 , n51654 , n399052 , n399053 , n51657 , n399055 , n51659 , n51660 , n399058 , 
 n399059 , n51663 , n399061 , n399062 , n51666 , n399064 , n399065 , n51669 , n399067 , n51671 , 
 n51672 , n399070 , n51674 , n399072 , n51676 , n51677 , n399075 , n399076 , n51680 , n399078 , 
 n399079 , n51683 , n399081 , n399082 , n51686 , n399084 , n51688 , n51689 , n399087 , n51691 , 
 n51692 , n399090 , n51694 , n399092 , n399093 , n51697 , n399095 , n51699 , n51700 , n399098 , 
 n399099 , n51703 , n399101 , n51705 , n399103 , n51707 , n399105 , n399106 , n51710 , n51711 , 
 n399109 , n51713 , n51714 , n399112 , n399113 , n51717 , n51718 , n399116 , n399117 , n51721 , 
 n399119 , n399120 , n51724 , n399122 , n51726 , n51727 , n51728 , n399126 , n51730 , n51731 , 
 n51732 , n399130 , n399131 , n51735 , n399133 , n51737 , n51738 , n399136 , n51740 , n399138 , 
 n51742 , n51743 , n399141 , n399142 , n51746 , n399144 , n399145 , n51749 , n399147 , n399148 , 
 n399149 , n51753 , n399151 , n399152 , n51756 , n399154 , n399155 , n51759 , n399157 , n51761 , 
 n399159 , n51763 , n51764 , n399162 , n51766 , n399164 , n399165 , n51769 , n399167 , n51771 , 
 n51772 , n51773 , n51774 , n51775 , n399173 , n399174 , n51778 , n399176 , n399177 , n51781 , 
 n399179 , n399180 , n399181 , n51785 , n399183 , n51787 , n51788 , n399186 , n399187 , n51791 , 
 n399189 , n399190 , n51794 , n399192 , n399193 , n51797 , n399195 , n51799 , n51800 , n399198 , 
 n399199 , n51803 , n399201 , n399202 , n51806 , n399204 , n399205 , n51809 , n399207 , n51811 , 
 n399209 , n51813 , n51814 , n399212 , n51816 , n399214 , n51818 , n51819 , n399217 , n51821 , 
 n51822 , n399220 , n51824 , n399222 , n399223 , n51827 , n399225 , n399226 , n399227 , n51831 , 
 n399229 , n399230 , n51834 , n399232 , n399233 , n51837 , n399235 , n399236 , n399237 , n399238 , 
 n51842 , n399240 , n399241 , n51845 , n399243 , n399244 , n51848 , n399246 , n51850 , n51851 , 
 n399249 , n399250 , n51854 , n399252 , n399253 , n51857 , n399255 , n399256 , n51860 , n399258 , 
 n51862 , n51863 , n399261 , n399262 , n51866 , n399264 , n399265 , n51869 , n399267 , n51871 , 
 n51872 , n51873 , n399271 , n399272 , n51876 , n399274 , n399275 , n51879 , n399277 , n51881 , 
 n51882 , n399280 , n399281 , n51885 , n399283 , n399284 , n51888 , n399286 , n399287 , n51891 , 
 n399289 , n399290 , n399291 , n51900 , n51901 , n399294 , n51903 , n51904 , n51905 , n399298 , 
 n51907 , n51908 , n51909 , n399302 , n51911 , n51912 , n51913 , n399306 , n51915 , n399308 , 
 n399309 , n51918 , n399311 , n51920 , n399313 , n399314 , n51923 , n399316 , n51925 , n399318 , 
 n51927 , n51928 , n51929 , n51930 , n51931 , n51932 , n399325 , n399326 , n51935 , n399328 , 
 n51937 , n399330 , n51939 , n51940 , n51941 , n399334 , n51943 , n51944 , n399337 , n51946 , 
 n399339 , n51948 , n399341 , n399342 , n51951 , n399344 , n51953 , n51954 , n399347 , n51956 , 
 n399349 , n51958 , n51959 , n51960 , n51961 , n51962 , n399355 , n399356 , n399357 , n51966 , 
 n399359 , n399360 , n51969 , n51970 , n399363 , n51972 , n51973 , n399366 , n51975 , n399368 , 
 n51977 , n399370 , n399371 , n51980 , n51981 , n51982 , n51983 , n399376 , n51985 , n51986 , 
 n399379 , n51988 , n399381 , n51990 , n51991 , n51992 , n51993 , n51994 , n399387 , n51996 , 
 n51997 , n399390 , n51999 , n52000 , n52001 , n399394 , n399395 , n399396 , n52005 , n399398 , 
 n52007 , n52008 , n399401 , n52010 , n399403 , n52012 , n52013 , n399406 , n399407 , n52016 , 
 n399409 , n399410 , n52019 , n399412 , n399413 , n399414 , n52023 , n399416 , n399417 , n52026 , 
 n399419 , n399420 , n52029 , n52030 , n52031 , n399424 , n399425 , n52034 , n52035 , n52036 , 
 n399429 , n399430 , n399431 , n52040 , n399433 , n52042 , n399435 , n52044 , n52045 , n399438 , 
 n399439 , n52048 , n399441 , n399442 , n52051 , n399444 , n399445 , n52054 , n52055 , n399448 , 
 n399449 , n52058 , n399451 , n399452 , n52061 , n399454 , n399455 , n52064 , n399457 , n399458 , 
 n52067 , n52068 , n399461 , n52070 , n52071 , n399464 , n399465 , n52074 , n399467 , n399468 , 
 n52077 , n399470 , n52079 , n52080 , n399473 , n399474 , n52083 , n399476 , n399477 , n52086 , 
 n399479 , n399480 , n52089 , n399482 , n399483 , n52092 , n52093 , n399486 , n52095 , n399488 , 
 n52097 , n52098 , n399491 , n399492 , n52101 , n399494 , n399495 , n52104 , n399497 , n52106 , 
 n52107 , n399500 , n399501 , n52110 , n399503 , n399504 , n52113 , n399506 , n52115 , n52116 , 
 n52117 , n52118 , n399511 , n399512 , n52121 , n399514 , n399515 , n399516 , n399517 , n52126 , 
 n399519 , n399520 , n52129 , n399522 , n399523 , n52132 , n52133 , n399526 , n52135 , n52136 , 
 n52137 , n52138 , n52139 , n399532 , n399533 , n52142 , n52143 , n399536 , n52145 , n399538 , 
 n399539 , n52148 , n52149 , n399542 , n52151 , n52152 , n399545 , n52154 , n52155 , n52156 , 
 n399549 , n399550 , n52159 , n52160 , n52161 , n399554 , n399555 , n52164 , n52165 , n52166 , 
 n399559 , n399560 , n52169 , n399562 , n399563 , n52172 , n399565 , n399566 , n52175 , n399568 , 
 n52177 , n52178 , n399571 , n399572 , n52181 , n399574 , n52183 , n399576 , n399577 , n52186 , 
 n52187 , n52188 , n52189 , n399582 , n399583 , n52192 , n399585 , n52194 , n52195 , n52196 , 
 n52197 , n399590 , n399591 , n52200 , n399593 , n52202 , n52203 , n52204 , n52205 , n399598 , 
 n399599 , n52208 , n399601 , n52210 , n52211 , n52212 , n52213 , n52214 , n52215 , n52216 , 
 n52217 , n52218 , n52219 , n52220 , n52221 , n52222 , n52223 , n399616 , n52225 , n52226 , 
 n52227 , n399620 , n52229 , n52230 , n52231 , n399624 , n52233 , n52234 , n52235 , n399628 , 
 n52237 , n52238 , n399631 , n52240 , n399633 , n52242 , n399635 , n52244 , n52245 , n52246 , 
 n52247 , n52248 , n399641 , n399642 , n52251 , n399644 , n52253 , n52254 , n399647 , n52256 , 
 n399649 , n52258 , n399651 , n52274 , n399653 , n399654 , n52339 , n52343 , n399657 , n52345 , 
 n52346 , n52347 , n52348 , n52349 , n52350 , n52351 , n52352 , n52353 , n52354 , n399668 , 
 n52356 , n399670 , n52358 , n52359 , n399673 , n399674 , n52362 , n399676 , n399677 , n52365 , 
 n399679 , n399680 , n399681 , n52369 , n399683 , n52371 , n399685 , n52373 , n399687 , n52375 , 
 n52376 , n52377 , n52378 , n52379 , n399693 , n52381 , n52382 , n52383 , n52384 , n52385 , 
 n52386 , n52387 , n52388 , n52389 , n52390 , n399704 , n399705 , n399706 , n52394 , n52395 , 
 n399709 , n399710 , n52398 , n399712 , n399713 , n52401 , n399715 , n52403 , n52404 , n399718 , 
 n52406 , n399720 , n52408 , n399722 , n399723 , n52411 , n399725 , n399726 , n52414 , n399728 , 
 n52416 , n399730 , n52418 , n52419 , n399733 , n399734 , n52422 , n399736 , n399737 , n52425 , 
 n399739 , n399740 , n52428 , n399742 , n52430 , n52431 , n52432 , n399746 , n52434 , n399748 , 
 n399749 , n399750 , n52438 , n399752 , n52440 , n52441 , n399755 , n52443 , n399757 , n52445 , 
 n52446 , n399760 , n399761 , n52449 , n52450 , n399764 , n399765 , n52453 , n399767 , n52455 , 
 n399769 , n399770 , n52458 , n399772 , n399773 , n52461 , n399775 , n52463 , n399777 , n52465 , 
 n52466 , n399780 , n399781 , n52469 , n399783 , n399784 , n52472 , n399786 , n399787 , n52475 , 
 n399789 , n52477 , n52478 , n52479 , n399793 , n52481 , n399795 , n399796 , n52484 , n52485 , 
 n52486 , n399800 , n399801 , n52489 , n52490 , n52491 , n399805 , n399806 , n52494 , n52495 , 
 n52496 , n399810 , n52498 , n52499 , n399813 , n52501 , n399815 , n399816 , n52504 , n52505 , 
 n399819 , n52507 , n52508 , n399822 , n52510 , n399824 , n52512 , n52513 , n52514 , n399828 , 
 n52516 , n52517 , n52518 , n52519 , n52520 , n52521 , n399835 , n52523 , n399837 , n52525 , 
 n52526 , n52527 , n399841 , n399842 , n52530 , n399844 , n52532 , n399846 , n399847 , n52535 , 
 n399849 , n399850 , n52538 , n399852 , n52540 , n52541 , n399855 , n52543 , n52544 , n399858 , 
 n399859 , n52547 , n52548 , n399862 , n399863 , n52551 , n52552 , n52553 , n399867 , n399868 , 
 n52556 , n399870 , n52558 , n52559 , n52560 , n52561 , n52562 , n52563 , n52564 , n52565 , 
 n52566 , n52567 , n52568 , n52569 , n52570 , n52571 , n52572 , n399886 , n399887 , n399888 , 
 n52576 , n399890 , n52578 , n399892 , n399893 , n399894 , n52582 , n399896 , n52584 , n52585 , 
 n399899 , n399900 , n52588 , n399902 , n52590 , n399904 , n399905 , n52593 , n399907 , n399908 , 
 n52596 , n399910 , n399911 , n52599 , n399913 , n399914 , n52602 , n52603 , n52604 , n399918 , 
 n399919 , n52607 , n399921 , n52609 , n52610 , n52611 , n52612 , n52613 , n52614 , n52615 , 
 n399929 , n52617 , n52618 , n52619 , n52620 , n399934 , n52622 , n52623 , n399937 , n52625 , 
 n399939 , n52627 , n52628 , n52629 , n52630 , n52631 , n52632 , n52633 , n399947 , n52635 , 
 n399949 , n52637 , n52638 , n399952 , n52640 , n52641 , n399955 , n52643 , n52644 , n52645 , 
 n52646 , n52647 , n52648 , n52649 , n52650 , n52651 , n52652 , n52653 , n52654 , n52655 , 
 n52656 , n399970 , n399971 , n52659 , n399973 , n399974 , n52662 , n52663 , n399977 , n52665 , 
 n399979 , n52667 , n399981 , n52669 , n52670 , n399984 , n52672 , n399986 , n399987 , n52675 , 
 n399989 , n52677 , n52678 , n399992 , n399993 , n52681 , n399995 , n399996 , n52684 , n399998 , 
 n399999 , n400000 , n52688 , n400002 , n400003 , n52691 , n400005 , n400006 , n52694 , n52695 , 
 n52696 , n400010 , n52698 , n400012 , n52700 , n52701 , n400015 , n400016 , n52704 , n400018 , 
 n400019 , n52707 , n400021 , n400022 , n400023 , n52711 , n400025 , n52713 , n52714 , n52715 , 
 n52716 , n400030 , n400031 , n52719 , n400033 , n400034 , n52722 , n400036 , n52724 , n52725 , 
 n400039 , n400040 , n52728 , n400042 , n400043 , n52731 , n400045 , n400046 , n52734 , n400048 , 
 n400049 , n400050 , n52741 , n400052 , n52743 , n52744 , n52745 , n52746 , n52747 , n52748 , 
 n52749 , n52750 , n52751 , n52752 , n52753 , n52754 , n52755 , n52756 , n52757 , n400068 , 
 n400069 , n52760 , n400071 , n52762 , n52763 , n400074 , n52765 , n52766 , n400077 , n400078 , 
 n52769 , n400080 , n400081 , n52772 , n400083 , n400084 , n52775 , n52776 , n400087 , n400088 , 
 n52779 , n400090 , n400091 , n52782 , n400093 , n400094 , n400095 , n52786 , n400097 , n52788 , 
 n52789 , n400100 , n400101 , n52792 , n400103 , n400104 , n52795 , n400106 , n400107 , n52798 , 
 n400109 , n52800 , n52801 , n400112 , n52803 , n400114 , n52805 , n400116 , n400117 , n52808 , 
 n400119 , n400120 , n52811 , n52812 , n400123 , n52814 , n400125 , n52816 , n400127 , n52818 , 
 n52819 , n400130 , n400131 , n52822 , n400133 , n400134 , n52825 , n400136 , n400137 , n52828 , 
 n52829 , n400140 , n400141 , n52832 , n400143 , n400144 , n52835 , n400146 , n400147 , n52838 , 
 n400149 , n400150 , n52841 , n400152 , n400153 , n400154 , n400155 , n52846 , n400157 , n400158 , 
 n52849 , n400160 , n400161 , n400162 , n52853 , n400164 , n52855 , n52856 , n52857 , n400168 , 
 n52859 , n400170 , n400171 , n52862 , n400173 , n52864 , n52865 , n400176 , n52867 , n400178 , 
 n52869 , n400180 , n400181 , n52872 , n400183 , n400184 , n52875 , n400186 , n52877 , n400188 , 
 n52879 , n52880 , n400191 , n400192 , n52883 , n400194 , n400195 , n52886 , n400197 , n400198 , 
 n52889 , n400200 , n52891 , n52892 , n400203 , n400204 , n52895 , n400206 , n400207 , n52898 , 
 n400209 , n400210 , n52901 , n52902 , n52903 , n400214 , n400215 , n52906 , n400217 , n52908 , 
 n400219 , n52910 , n400221 , n52912 , n52913 , n400224 , n400225 , n52916 , n400227 , n400228 , 
 n52919 , n400230 , n400231 , n52922 , n52923 , n400234 , n400235 , n52926 , n400237 , n400238 , 
 n52929 , n400240 , n400241 , n52932 , n52933 , n52934 , n400245 , n400246 , n52937 , n400248 , 
 n52939 , n400250 , n52941 , n52942 , n400253 , n52944 , n400255 , n52946 , n52947 , n400258 , 
 n52949 , n400260 , n52951 , n400262 , n400263 , n52954 , n400265 , n400266 , n400267 , n52958 , 
 n400269 , n400270 , n52961 , n400272 , n400273 , n52964 , n52965 , n52966 , n400277 , n400278 , 
 n52969 , n52970 , n52971 , n400282 , n400283 , n52974 , n52975 , n52976 , n400287 , n400288 , 
 n52979 , n52980 , n52981 , n52982 , n52983 , n400294 , n52985 , n400296 , n52987 , n52988 , 
 n400299 , n400300 , n52991 , n400302 , n400303 , n52994 , n400305 , n52996 , n400307 , n400308 , 
 n400309 , n53000 , n400311 , n53002 , n53003 , n400314 , n53005 , n400316 , n53007 , n400318 , 
 n400319 , n53010 , n400321 , n53012 , n400323 , n400324 , n53015 , n400326 , n53017 , n53018 , 
 n400329 , n53020 , n400331 , n53022 , n53023 , n53024 , n53025 , n53026 , n400337 , n53028 , 
 n400339 , n53030 , n53031 , n400342 , n400343 , n53034 , n400345 , n400346 , n53037 , n400348 , 
 n53039 , n53040 , n53041 , n53042 , n400353 , n53044 , n400355 , n53046 , n53047 , n53048 , 
 n53049 , n53050 , n53051 , n53052 , n400363 , n53054 , n400365 , n53056 , n400367 , n53058 , 
 n53059 , n53060 , n400371 , n53062 , n400373 , n53064 , n400375 , n400376 , n53067 , n53068 , 
 n53069 , n400380 , n53071 , n400382 , n53073 , n53074 , n400385 , n400386 , n53077 , n400388 , 
 n400389 , n53080 , n400391 , n53082 , n53083 , n400394 , n400395 , n53086 , n400397 , n53088 , 
 n400399 , n53090 , n400401 , n53092 , n400403 , n53094 , n400405 , n53096 , n53097 , n53098 , 
 n400409 , n53100 , n400411 , n53102 , n53103 , n53104 , n53105 , n53106 , n400417 , n53108 , 
 n400419 , n53110 , n53111 , n400422 , n400423 , n53114 , n400425 , n53116 , n53117 , n53118 , 
 n53119 , n400430 , n53121 , n53122 , n53123 , n400434 , n400435 , n400436 , n53127 , n400438 , 
 n53129 , n400440 , n53131 , n53132 , n400443 , n53134 , n53135 , n53136 , n400447 , n53138 , 
 n400449 , n400450 , n53141 , n400452 , n400453 , n53144 , n400455 , n53146 , n53147 , n400458 , 
 n400459 , n53150 , n400461 , n400462 , n53153 , n400464 , n400465 , n53156 , n400467 , n53158 , 
 n53159 , n400470 , n400471 , n53162 , n400473 , n400474 , n53165 , n400476 , n400477 , n53168 , 
 n53169 , n53170 , n53171 , n53172 , n53173 , n53174 , n53175 , n400486 , n400487 , n53178 , 
 n400489 , n53180 , n400491 , n53182 , n53183 , n400494 , n400495 , n53186 , n400497 , n53188 , 
 n400499 , n53190 , n53191 , n400502 , n400503 , n53194 , n400505 , n400506 , n53197 , n400508 , 
 n400509 , n53200 , n400511 , n400512 , n53203 , n400514 , n400515 , n53206 , n400517 , n400518 , 
 n53209 , n400520 , n400521 , n53212 , n400523 , n53214 , n400525 , n53216 , n53217 , n400528 , 
 n400529 , n53220 , n400531 , n400532 , n53223 , n400534 , n400535 , n53226 , n400537 , n53228 , 
 n53229 , n400540 , n400541 , n53232 , n400543 , n400544 , n53235 , n400546 , n400547 , n53238 , 
 n53239 , n400550 , n400551 , n53242 , n400553 , n53244 , n400555 , n53246 , n53247 , n53248 , 
 n53249 , n53250 , n53251 , n53252 , n53253 , n53254 , n53255 , n400566 , n53257 , n400568 , 
 n400569 , n53260 , n400571 , n400572 , n53263 , n400574 , n400575 , n53266 , n400577 , n400578 , 
 n53269 , n400580 , n53271 , n400582 , n400583 , n53274 , n400585 , n53276 , n400587 , n53278 , 
 n53279 , n53280 , n53281 , n400592 , n400593 , n53284 , n400595 , n53286 , n400597 , n53288 , 
 n400599 , n53290 , n53291 , n53292 , n53293 , n400604 , n53295 , n400606 , n400607 , n53298 , 
 n400609 , n53300 , n53301 , n53302 , n400613 , n400614 , n53305 , n400616 , n53307 , n400618 , 
 n53309 , n400620 , n400621 , n53312 , n53313 , n400624 , n53315 , n53316 , n400627 , n53318 , 
 n53319 , n53320 , n53321 , n53322 , n53323 , n53324 , n53325 , n53326 , n53327 , n53328 , 
 n53329 , n53330 , n53331 , n53332 , n53333 , n53334 , n53335 , n53336 , n53337 , n53338 , 
 n53339 , n53340 , n53341 , n53342 , n53343 , n53344 , n53345 , n53346 , n53347 , n53348 , 
 n53349 , n53350 , n53351 , n53352 , n53353 , n53354 , n53355 , n53356 , n53357 , n53358 , 
 n53359 , n53360 , n53361 , n53362 , n53363 , n53364 , n53365 , n53366 , n53367 , n53368 , 
 n53369 , n53370 , n53371 , n53372 , n53373 , n53374 , n53375 , n53376 , n53377 , n53378 , 
 n53379 , n53380 , n53381 , n53382 , n53383 , n53384 , n53385 , n53386 , n53387 , n53388 , 
 n53389 , n53390 , n53391 , n53392 , n53393 , n53394 , n53395 , n53396 , n53397 , n53398 , 
 n53399 , n53400 , n53401 , n53402 , n53403 , n53404 , n53405 , n53406 , n53407 , n53408 , 
 n53409 , n53410 , n53411 , n53412 , n53413 , n53414 , n53415 , n53416 , n53417 , n53418 , 
 n53419 , n53420 , n53421 , n53422 , n53423 , n53424 , n53425 , n53426 , n53427 , n53428 , 
 n53429 , n53430 , n53431 , n53432 , n53433 , n53434 , n53435 , n53436 , n53437 , n53438 , 
 n53439 , n53440 , n53441 , n53442 , n53443 , n53444 , n53445 , n53446 , n53447 , n53448 , 
 n53449 , n53450 , n53451 , n53452 , n53453 , n53454 , n53455 , n53456 , n53457 , n53458 , 
 n53459 , n53460 , n53461 , n53462 , n53463 , n53464 , n53465 , n53466 , n53467 , n53468 , 
 n53469 , n53470 , n53471 , n53472 , n53473 , n53474 , n53475 , n53476 , n53477 , n53478 , 
 n53479 , n53480 , n53481 , n53482 , n53483 , n53484 , n53485 , n53486 , n53487 , n53488 , 
 n53489 , n53490 , n53491 , n53492 , n53493 , n53494 , n53495 , n53496 , n53497 , n53498 , 
 n53499 , n53500 , n53501 , n53502 , n53503 , n53504 , n53505 , n53506 , n53507 , n53508 , 
 n53509 , n53510 , n53511 , n53512 , n53513 , n53514 , n53515 , n53516 , n53517 , n53518 , 
 n53519 , n53520 , n53521 , n53522 , n53523 , n53524 , n53525 , n53526 , n53527 , n53528 , 
 n53529 , n53530 , n53531 , n53532 , n53533 , n53534 , n53535 , n53536 , n53537 , n53538 , 
 n53539 , n53540 , n53541 , n53542 , n53543 , n53544 , n53545 , n53546 , n53547 , n53548 , 
 n53549 , n53550 , n53551 , n53552 , n53553 , n53554 , n53555 , n53556 , n53557 , n53558 , 
 n53559 , n53560 , n53561 , n53562 , n53563 , n53564 , n53565 , n53566 , n53567 , n53568 , 
 n53569 , n53570 , n53571 , n53572 , n53573 , n53574 , n53575 , n53576 , n53577 , n53578 , 
 n53579 , n53580 , n53581 , n53582 , n53583 , n53584 , n53585 , n53586 , n53587 , n53588 , 
 n53589 , n53590 , n53591 , n53592 , n53593 , n53594 , n53595 , n53596 , n53597 , n53598 , 
 n53599 , n53600 , n53601 , n53602 , n53603 , n53604 , n53605 , n53606 , n53607 , n53608 , 
 n53609 , n53610 , n53611 , n53612 , n53613 , n53614 , n53615 , n53616 , n53617 , n53618 , 
 n53619 , n53620 , n53621 , n53622 , n53623 , n53624 , n53625 , n53626 , n53627 , n53628 , 
 n53629 , n53630 , n53631 , n53632 , n53633 , n53634 , n53635 , n53636 , n53637 , n53638 , 
 n53639 , n53640 , n53641 , n53642 , n53643 , n53644 , n53645 , n53646 , n53647 , n53648 , 
 n53649 , n53650 , n53651 , n53652 , n53653 , n53654 , n53655 , n53656 , n53657 , n53658 , 
 n53659 , n53660 , n53661 , n53662 , n53663 , n53664 , n53665 , n53666 , n53667 , n53668 , 
 n53669 , n53670 , n53671 , n53672 , n53673 , n53674 , n53675 , n53676 , n53677 , n53678 , 
 n53679 , n53680 , n53681 , n53682 , n53683 , n53684 , n53685 , n53686 , n53687 , n53688 , 
 n53689 , n53690 , n53691 , n53692 , n53693 , n53694 , n53695 , n53696 , n53697 , n53698 , 
 n53699 , n53700 , n53701 , n53702 , n53703 , n53704 , n53705 , n53706 , n53707 , n53708 , 
 n53709 , n53710 , n53711 , n53712 , n53713 , n53714 , n53715 , n53716 , n53717 , n53718 , 
 n53719 , n53720 , n53721 , n53722 , n53723 , n53724 , n53725 , n53726 , n53727 , n53728 , 
 n53729 , n53730 , n53731 , n53732 , n53733 , n53734 , n53735 , n53736 , n53737 , n401048 , 
 n53739 , n53740 , n53741 , n53742 , n53743 , n53744 , n53745 , n53746 , n53747 , n53748 , 
 n53749 , n53750 , n53751 , n53752 , n53753 , n53754 , n53755 , n53756 , n53757 , n53758 , 
 n53759 , n53760 , n53761 , n53762 , n53763 , n53764 , n53765 , n53766 , n53767 , n53768 , 
 n53769 , n53770 , n53771 , n53772 , n53773 , n53774 , n53775 , n53776 , n53777 , n53778 , 
 n53779 , n53780 , n53781 , n53782 , n53783 , n53784 , n53785 , n53786 , n53787 , n53788 , 
 n53789 , n53790 , n53791 , n53792 , n53793 , n53794 , n53795 , n53796 , n53797 , n53798 , 
 n53799 , n53800 , n53801 , n53802 , n53803 , n53804 , n53805 , n53806 , n53807 , n53808 , 
 n53809 , n53810 , n53811 , n53812 , n53813 , n53814 , n53815 , n53816 , n53817 , n53818 , 
 n53819 , n53820 , n53821 , n53822 , n53823 , n53824 , n53825 , n53826 , n53827 , n53828 , 
 n53829 , n53830 , n53831 , n53832 , n53833 , n53834 , n53835 , n53836 , n53837 , n53838 , 
 n53839 , n53840 , n53841 , n53842 , n53843 , n53844 , n53845 , n53846 , n53847 , n53848 , 
 n53849 , n53850 , n53851 , n53852 , n53853 , n53854 , n53855 , n53856 , n53857 , n53858 , 
 n53859 , n53860 , n53861 , n53862 , n53863 , n53864 , n53865 , n53866 , n53867 , n53868 , 
 n53869 , n53870 , n53871 , n53872 , n53873 , n53874 , n53875 , n53876 , n53877 , n53878 , 
 n53879 , n53880 , n53881 , n53882 , n53883 , n53884 , n53885 , n53886 , n53887 , n53888 , 
 n53889 , n53890 , n53891 , n53892 , n53893 , n53894 , n53895 , n53896 , n53897 , n53898 , 
 n53899 , n53900 , n53901 , n53902 , n53903 , n53904 , n53905 , n53906 , n53907 , n53908 , 
 n53909 , n53910 , n53911 , n53912 , n53913 , n53914 , n53915 , n53916 , n53917 , n53918 , 
 n53919 , n53920 , n53921 , n53922 , n53923 , n53924 , n53925 , n53926 , n53927 , n53928 , 
 n53929 , n53930 , n53931 , n53932 , n53933 , n53934 , n53935 , n53936 , n53937 , n53938 , 
 n53939 , n53940 , n53941 , n53942 , n53943 , n53944 , n53945 , n53946 , n53947 , n53948 , 
 n53949 , n53950 , n53951 , n53952 , n53953 , n53954 , n53955 , n53956 , n53957 , n53958 , 
 n53959 , n53960 , n53961 , n53962 , n53963 , n53964 , n53965 , n53966 , n53967 , n53968 , 
 n53969 , n53970 , n53971 , n53972 , n53973 , n53974 , n53975 , n53976 , n53977 , n53978 , 
 n53979 , n53980 , n53981 , n53982 , n53983 , n53984 , n53985 , n53986 , n53987 , n53988 , 
 n53989 , n53990 , n53991 , n53992 , n53993 , n53994 , n53995 , n53996 , n53997 , n53998 , 
 n53999 , n54000 , n54001 , n54002 , n54003 , n54004 , n54005 , n54006 , n54007 , n54008 , 
 n54009 , n54010 , n54011 , n54012 , n54013 , n54014 , n54015 , n54016 , n54017 , n54018 , 
 n54019 , n54020 , n54021 , n54022 , n54023 , n54024 , n54025 , n54026 , n54027 , n54028 , 
 n54029 , n54030 , n54031 , n54032 , n54033 , n54034 , n54035 , n54036 , n54037 , n54038 , 
 n54039 , n54040 , n54041 , n54042 , n54043 , n54044 , n54045 , n54046 , n54047 , n54048 , 
 n54049 , n54050 , n54051 , n54052 , n54053 , n54054 , n54055 , n54056 , n54057 , n54058 , 
 n54059 , n54060 , n54061 , n54062 , n54063 , n54064 , n54065 , n54066 , n54067 , n54068 , 
 n54069 , n54070 , n54071 , n54072 , n54073 , n54074 , n54075 , n54076 , n54077 , n54078 , 
 n54079 , n54080 , n54081 , n54082 , n54083 , n54084 , n54085 , n54086 , n54087 , n54088 , 
 n54089 , n54090 , n54091 , n54092 , n54093 , n54094 , n54095 , n54096 , n54097 , n54098 , 
 n54099 , n54100 , n54101 , n54102 , n54103 , n54104 , n54105 , n54106 , n54107 , n54108 , 
 n54109 , n54110 , n54111 , n54112 , n54113 , n54114 , n54115 , n54116 , n54117 , n54118 , 
 n54119 , n54120 , n54121 , n54122 , n54123 , n54124 , n54125 , n54126 , n54127 , n54128 , 
 n54129 , n54130 , n54131 , n54132 , n54133 , n54134 , n54135 , n54136 , n54137 , n54138 , 
 n54139 , n54140 , n54141 , n54142 , n54143 , n54144 , n54145 , n54146 , n54147 , n54148 , 
 n54149 , n54150 , n54151 , n54152 , n54153 , n54154 , n54155 , n54156 , n54157 , n54158 , 
 n54159 , n54160 , n54161 , n54162 , n54163 , n54164 , n54165 , n54166 , n54167 , n54168 , 
 n54169 , n54170 , n54171 , n54172 , n54173 , n54174 , n54175 , n54176 , n54177 , n54178 , 
 n54179 , n54180 , n54181 , n54182 , n54183 , n54184 , n54185 , n54186 , n54187 , n54188 , 
 n54189 , n54190 , n54191 , n54192 , n54193 , n54194 , n54195 , n54196 , n54197 , n54198 , 
 n54199 , n54200 , n54201 , n54202 , n54203 , n54204 , n54205 , n54206 , n54207 , n54208 , 
 n54209 , n54210 , n54211 , n54212 , n54213 , n54214 , n54215 , n54216 , n54217 , n54218 , 
 n54219 , n54220 , n54221 , n54222 , n54223 , n54224 , n54225 , n54226 , n54227 , n54228 , 
 n54229 , n54230 , n54231 , n54232 , n54233 , n54234 , n54235 , n54236 , n54237 , n54238 , 
 n54239 , n54240 , n54241 , n54242 , n54243 , n54244 , n54245 , n54246 , n54247 , n54248 , 
 n54249 , n54250 , n54251 , n54252 , n54253 , n54254 , n54255 , n54256 , n54257 , n54258 , 
 n54259 , n54260 , n54261 , n54262 , n54263 , n54264 , n54265 , n54266 , n54267 , n401578 , 
 n54269 , n54270 , n54271 , n54272 , n54273 , n54274 , n54275 , n54276 , n54277 , n54278 , 
 n54279 , n54280 , n54281 , n54282 , n54283 , n54284 , n54285 , n54286 , n54287 , n54288 , 
 n54289 , n54290 , n54291 , n54292 , n54293 , n54294 , n54295 , n54296 , n54297 , n401608 , 
 n401609 , n401610 , n54301 , n401612 , n401613 , n54304 , n54305 , n401616 , n54307 , n54308 , 
 n401619 , n401620 , n401621 , n54312 , n401623 , n401624 , n54315 , n401626 , n401627 , n54318 , 
 n54319 , n54320 , n54321 , n54322 , n54323 , n54324 , n54325 , n54326 , n54327 , n54328 , 
 n54329 , n54330 , n54331 , n54332 , n54333 , n54334 , n54335 , n54336 , n401647 , n401648 , 
 n54339 , n401650 , n401651 , n54342 , n54343 , n401654 , n401655 , n54346 , n401657 , n401658 , 
 n54349 , n401660 , n401661 , n401662 , n54353 , n401664 , n401665 , n54356 , n401667 , n401668 , 
 n401669 , n54360 , n401671 , n401672 , n54363 , n401674 , n401675 , n401676 , n54367 , n401678 , 
 n401679 , n54370 , n401681 , n401682 , n54373 , n401684 , n401685 , n54376 , n401687 , n54378 , 
 n401689 , n401690 , n54381 , n401692 , n401693 , n54384 , n401695 , n401696 , n401697 , n54388 , 
 n401699 , n401700 , n54391 , n54392 , n401703 , n54394 , n54395 , n401706 , n401707 , n54398 , 
 n401709 , n401710 , n401711 , n54402 , n401713 , n54404 , n401715 , n401716 , n54407 , n54408 , 
 n54409 , n54410 , n54411 , n54412 , n54413 , n54414 , n54415 , n54416 , n54417 , n54418 , 
 n54419 , n54420 , n54421 , n54422 , n54423 , n54424 , n54425 , n54426 , n54427 , n54428 , 
 n54429 , n54430 , n54431 , n54432 , n54433 , n401744 , n401745 , n54436 , n401747 , n401748 , 
 n54439 , n54440 , n401751 , n401752 , n54443 , n401754 , n401755 , n54446 , n401757 , n401758 , 
 n54449 , n54450 , n54451 , n401762 , n401763 , n401764 , n401765 , n54456 , n401767 , n401768 , 
 n54459 , n401770 , n54461 , n54462 , n401773 , n54464 , n401775 , n401776 , n401777 , n54468 , 
 n54469 , n401780 , n54471 , n54472 , n401783 , n401784 , n54475 , n401786 , n54477 , n401788 , 
 n401789 , n401790 , n54481 , n54482 , n401793 , n401794 , n54485 , n54486 , n54487 , n401798 , 
 n401799 , n401800 , n54491 , n401802 , n54493 , n54494 , n401805 , n54496 , n401807 , n54498 , 
 n54499 , n401810 , n401811 , n54502 , n401813 , n401814 , n54505 , n401816 , n401817 , n401818 , 
 n54509 , n401820 , n401821 , n54512 , n401823 , n401824 , n54515 , n401826 , n401827 , n54518 , 
 n54519 , n401830 , n54521 , n54522 , n401833 , n401834 , n54525 , n401836 , n54527 , n54528 , 
 n401839 , n54530 , n401841 , n54532 , n401843 , n401844 , n54535 , n401846 , n401847 , n54538 , 
 n54539 , n54540 , n401851 , n54542 , n54543 , n401854 , n54545 , n54546 , n54547 , n401858 , 
 n401859 , n401860 , n54551 , n401862 , n54553 , n401864 , n54555 , n54556 , n401867 , n54558 , 
 n401869 , n54560 , n401871 , n401872 , n54563 , n401874 , n401875 , n54566 , n54567 , n401878 , 
 n401879 , n54570 , n401881 , n401882 , n54573 , n401884 , n401885 , n54576 , n54577 , n401888 , 
 n401889 , n54580 , n54581 , n401892 , n401893 , n54584 , n54585 , n401896 , n54587 , n54588 , 
 n401899 , n54590 , n54591 , n54592 , n54593 , n54594 , n401905 , n54596 , n401907 , n401908 , 
 n54599 , n54600 , n54601 , n54602 , n54603 , n54604 , n54605 , n54606 , n54607 , n401918 , 
 n401919 , n54610 , n401921 , n54612 , n401923 , n54614 , n54615 , n54616 , n54617 , n401928 , 
 n401929 , n54620 , n401931 , n54622 , n401933 , n401934 , n54625 , n401936 , n401937 , n54628 , 
 n401939 , n401940 , n54631 , n54632 , n54633 , n401944 , n401945 , n54636 , n54637 , n54638 , 
 n54639 , n54640 , n54641 , n54642 , n54643 , n54644 , n54645 , n54646 , n401957 , n54648 , 
 n54649 , n54650 , n401961 , n401962 , n54653 , n54654 , n54655 , n401966 , n401967 , n54658 , 
 n401969 , n401970 , n401971 , n401972 , n54663 , n54664 , n401975 , n54666 , n54667 , n401978 , 
 n54669 , n54670 , n54671 , n54672 , n54673 , n54674 , n401985 , n54676 , n54677 , n54678 , 
 n401989 , n54680 , n54681 , n54682 , n401993 , n54684 , n54685 , n54686 , n401997 , n401998 , 
 n54689 , n54690 , n402001 , n402002 , n54693 , n402004 , n402005 , n54696 , n402007 , n54698 , 
 n402009 , n54700 , n54701 , n402012 , n54703 , n54704 , n54705 , n402016 , n402017 , n402018 , 
 n54709 , n402020 , n54711 , n402022 , n54713 , n54714 , n402025 , n402026 , n54717 , n402028 , 
 n402029 , n54720 , n402031 , n402032 , n54723 , n54724 , n402035 , n402036 , n54727 , n402038 , 
 n402039 , n54730 , n402041 , n402042 , n402043 , n402044 , n54764 , n402046 , n54766 , n402048 , 
 n54768 , n54769 , n402051 , n54771 , n402053 , n54773 , n54774 , n402056 , n402057 , n54777 , 
 n402059 , n402060 , n54780 , n402062 , n402063 , n402064 , n54784 , n402066 , n402067 , n54787 , 
 n402069 , n402070 , n54790 , n402072 , n402073 , n402074 , n54795 , n54796 , n54797 , n402078 , 
 n54799 , n54800 , n54801 , n402082 , n54803 , n402084 , n402085 , n54806 , n402087 , n54808 , 
 n402089 , n54810 , n54811 , n54812 , n402093 , n402094 , n54815 , n54816 , n402097 , n402098 , 
 n54819 , n54820 , n54821 , n402102 , n402103 , n54824 , n54825 , n54826 , n54827 , n54828 , 
 n54829 , n54830 , n54831 , n54832 , n54833 , n54834 , n54835 , n54836 , n54837 , n402118 , 
 n54839 , n54840 , n54841 , n402122 , n54843 , n402124 , n54845 , n54846 , n54847 , n54848 , 
 n54849 , n402130 , n54851 , n402132 , n54853 , n54854 , n402135 , n402136 , n54857 , n402138 , 
 n402139 , n54860 , n402141 , n402142 , n402143 , n54864 , n402145 , n54866 , n402147 , n402148 , 
 n54869 , n402150 , n54871 , n54872 , n54873 , n402154 , n54875 , n402156 , n54877 , n402158 , 
 n402159 , n54880 , n402161 , n402162 , n54883 , n402164 , n402165 , n54886 , n402167 , n54888 , 
 n402169 , n54890 , n54891 , n54892 , n54893 , n54894 , n402175 , n54896 , n402177 , n54898 , 
 n54899 , n402180 , n402181 , n54902 , n402183 , n402184 , n54905 , n402186 , n402187 , n402188 , 
 n54909 , n402190 , n54911 , n54912 , n54913 , n54914 , n54915 , n54916 , n54917 , n54918 , 
 n54919 , n54920 , n402201 , n54922 , n54923 , n54924 , n54925 , n54926 , n54927 , n54928 , 
 n54929 , n54930 , n54931 , n54932 , n402213 , n54934 , n402215 , n402216 , n54937 , n402218 , 
 n54939 , n402220 , n54941 , n54942 , n54943 , n54944 , n54945 , n54946 , n402227 , n402228 , 
 n54949 , n402230 , n54951 , n54952 , n54953 , n54954 , n402235 , n54956 , n54957 , n402238 , 
 n54959 , n54960 , n402241 , n402242 , n54963 , n402244 , n402245 , n54966 , n402247 , n402248 , 
 n54969 , n402250 , n54971 , n54972 , n402253 , n402254 , n54975 , n402256 , n402257 , n54978 , 
 n402259 , n54980 , n54981 , n54982 , n402263 , n54984 , n54985 , n54986 , n402267 , n54988 , 
 n54989 , n402270 , n54991 , n54992 , n54993 , n402274 , n402275 , n54996 , n402277 , n54998 , 
 n402279 , n55000 , n55001 , n55002 , n402283 , n402284 , n55005 , n55006 , n55007 , n402288 , 
 n402289 , n55010 , n55011 , n402292 , n402293 , n55014 , n402295 , n55016 , n402297 , n55018 , 
 n55019 , n402300 , n55021 , n402302 , n55023 , n55024 , n402305 , n55026 , n402307 , n402308 , 
 n402309 , n55030 , n402311 , n402312 , n55033 , n402314 , n402315 , n402316 , n55037 , n402318 , 
 n402319 , n55040 , n402321 , n402322 , n55043 , n55044 , n402325 , n402326 , n55047 , n55048 , 
 n402329 , n402330 , n55051 , n402332 , n55053 , n55054 , n55055 , n402336 , n55057 , n402338 , 
 n55059 , n55060 , n402341 , n402342 , n55063 , n402344 , n402345 , n55066 , n402347 , n402348 , 
 n402349 , n55075 , n402351 , n402352 , n55078 , n402354 , n402355 , n55081 , n402357 , n55083 , 
 n402359 , n55085 , n402361 , n55087 , n55088 , n402364 , n402365 , n55091 , n402367 , n402368 , 
 n55094 , n402370 , n402371 , n55097 , n402373 , n55099 , n402375 , n402376 , n55102 , n55103 , 
 n402379 , n402380 , n55106 , n402382 , n402383 , n55109 , n402385 , n402386 , n55112 , n402388 , 
 n55114 , n55115 , n402391 , n402392 , n55118 , n402394 , n402395 , n55121 , n402397 , n55123 , 
 n55124 , n402400 , n402401 , n55127 , n402403 , n402404 , n55130 , n402406 , n55132 , n55133 , 
 n55134 , n402410 , n402411 , n55137 , n402413 , n55139 , n55140 , n55141 , n55142 , n402418 , 
 n55144 , n55145 , n55146 , n402422 , n402423 , n55149 , n402425 , n402426 , n55152 , n55153 , 
 n55154 , n55155 , n55156 , n55157 , n55158 , n55159 , n55160 , n55161 , n55162 , n55163 , 
 n402439 , n55165 , n402441 , n402442 , n55168 , n402444 , n402445 , n402446 , n55172 , n402448 , 
 n55174 , n402450 , n402451 , n55177 , n402453 , n402454 , n55180 , n402456 , n402457 , n55183 , 
 n402459 , n402460 , n55186 , n55187 , n55188 , n402464 , n402465 , n55191 , n55192 , n402468 , 
 n402469 , n55195 , n55196 , n55197 , n55198 , n55199 , n55200 , n55201 , n55202 , n55203 , 
 n55204 , n55205 , n402481 , n55207 , n402483 , n402484 , n55210 , n55211 , n55212 , n55213 , 
 n55214 , n402490 , n55216 , n55217 , n402493 , n55219 , n402495 , n55221 , n55222 , n402498 , 
 n55259 , n55260 , n55261 , n402502 , n402503 , n55264 , n402505 , n55266 , n402507 , n55268 , 
 n402509 , n55270 , n55271 , n55272 , n55273 , n55274 , n55275 , n55276 , n55277 , n402518 , 
 n402519 , n55280 , n402521 , n55282 , n55283 , n402524 , n402525 , n55286 , n402527 , n402528 , 
 n55289 , n402530 , n402531 , n55292 , n402533 , n55294 , n55295 , n402536 , n402537 , n55298 , 
 n402539 , n402540 , n55301 , n402542 , n55303 , n55304 , n55305 , n55306 , n55307 , n55308 , 
 n55309 , n402550 , n55311 , n402552 , n55313 , n402554 , n402555 , n55316 , n402557 , n402558 , 
 n55319 , n402560 , n402561 , n55322 , n402563 , n402564 , n55325 , n55326 , n55327 , n402568 , 
 n402569 , n55330 , n55331 , n55332 , n402573 , n402574 , n55335 , n55336 , n402577 , n55338 , 
 n402579 , n402580 , n55341 , n402582 , n55343 , n402584 , n402585 , n55346 , n55347 , n55348 , 
 n55349 , n402590 , n55351 , n55352 , n402593 , n55354 , n402595 , n402596 , n55357 , n55358 , 
 n55359 , n55360 , n55361 , n402602 , n402603 , n55364 , n402605 , n402606 , n55367 , n402608 , 
 n402609 , n402610 , n55371 , n402612 , n55373 , n55374 , n55375 , n55376 , n55377 , n55378 , 
 n55379 , n402620 , n402621 , n55382 , n402623 , n402624 , n55385 , n402626 , n402627 , n55388 , 
 n55389 , n55390 , n402631 , n402632 , n55393 , n55394 , n55395 , n55396 , n55397 , n402638 , 
 n55399 , n402640 , n402641 , n55402 , n402643 , n55404 , n402645 , n55406 , n55407 , n402648 , 
 n402649 , n55410 , n402651 , n402652 , n55413 , n402654 , n402655 , n55416 , n402657 , n55418 , 
 n55419 , n402660 , n402661 , n55422 , n402663 , n402664 , n55425 , n402666 , n402667 , n55428 , 
 n55429 , n55430 , n402671 , n55432 , n402673 , n55434 , n402675 , n55436 , n55437 , n402678 , 
 n55439 , n402680 , n55441 , n55442 , n402683 , n402684 , n55445 , n402686 , n402687 , n55448 , 
 n402689 , n402690 , n402691 , n55452 , n55453 , n402694 , n402695 , n55456 , n402697 , n55458 , 
 n55459 , n402700 , n402701 , n55462 , n402703 , n402704 , n55465 , n402706 , n402707 , n55468 , 
 n402709 , n55470 , n55471 , n402712 , n402713 , n55474 , n402715 , n402716 , n55477 , n402718 , 
 n55479 , n55480 , n55481 , n55482 , n402723 , n402724 , n55485 , n402726 , n402727 , n55488 , 
 n402729 , n55490 , n55491 , n402732 , n55493 , n402734 , n402735 , n55496 , n55497 , n402738 , 
 n402739 , n55500 , n402741 , n402742 , n55503 , n402744 , n402745 , n55506 , n402747 , n402748 , 
 n55509 , n402750 , n402751 , n55512 , n55513 , n402754 , n402755 , n55516 , n55517 , n402758 , 
 n55519 , n402760 , n402761 , n55522 , n402763 , n55524 , n55525 , n402766 , n402767 , n55528 , 
 n55529 , n402770 , n402771 , n55532 , n402773 , n55534 , n55535 , n402776 , n402777 , n55538 , 
 n55539 , n402780 , n402781 , n55542 , n55543 , n402784 , n55545 , n402786 , n55547 , n55548 , 
 n402789 , n402790 , n55551 , n402792 , n402793 , n55554 , n402795 , n402796 , n55557 , n402798 , 
 n55559 , n55560 , n402801 , n402802 , n55563 , n402804 , n402805 , n55566 , n402807 , n402808 , 
 n55569 , n402810 , n55571 , n55572 , n55573 , n55574 , n55575 , n55576 , n402817 , n55583 , 
 n402819 , n55590 , n55591 , n55592 , n55593 , n402824 , n402825 , n55596 , n402827 , n402828 , 
 n55599 , n402830 , n55601 , n55602 , n402833 , n402834 , n55605 , n402836 , n402837 , n55608 , 
 n402839 , n402840 , n55611 , n402842 , n402843 , n55614 , n402845 , n55616 , n55617 , n402848 , 
 n55619 , n402850 , n55621 , n402852 , n402853 , n55624 , n402855 , n402856 , n402857 , n55628 , 
 n402859 , n55630 , n55631 , n402862 , n402863 , n55634 , n402865 , n402866 , n55637 , n402868 , 
 n402869 , n55640 , n402871 , n55642 , n55643 , n402874 , n55645 , n402876 , n55647 , n402878 , 
 n402879 , n55650 , n402881 , n402882 , n55653 , n402884 , n55655 , n55656 , n55657 , n55658 , 
 n55659 , n55660 , n402891 , n55662 , n55663 , n402894 , n402895 , n55666 , n402897 , n402898 , 
 n55669 , n402900 , n402901 , n55672 , n55673 , n55674 , n402905 , n55676 , n55677 , n402908 , 
 n55679 , n55680 , n402911 , n55682 , n402913 , n55684 , n55685 , n402916 , n402917 , n55688 , 
 n402919 , n402920 , n55691 , n402922 , n402923 , n55694 , n402925 , n55696 , n55697 , n55698 , 
 n402929 , n55700 , n402931 , n55702 , n55703 , n55704 , n55705 , n55706 , n402937 , n55708 , 
 n402939 , n55710 , n55711 , n402942 , n402943 , n55714 , n402945 , n402946 , n55717 , n402948 , 
 n55719 , n55720 , n402951 , n402952 , n55723 , n402954 , n402955 , n55726 , n402957 , n55728 , 
 n55729 , n402960 , n55731 , n402962 , n55733 , n55734 , n402965 , n402966 , n55737 , n402968 , 
 n402969 , n55740 , n402971 , n402972 , n402973 , n55744 , n402975 , n402976 , n55747 , n402978 , 
 n402979 , n55750 , n402981 , n55752 , n55753 , n402984 , n55755 , n402986 , n402987 , n402988 , 
 n55759 , n402990 , n55761 , n402992 , n402993 , n55764 , n402995 , n402996 , n55767 , n402998 , 
 n402999 , n55770 , n403001 , n403002 , n55773 , n403004 , n55775 , n403006 , n403007 , n403008 , 
 n55779 , n403010 , n55781 , n55782 , n55783 , n55784 , n55785 , n55786 , n403017 , n403018 , 
 n55789 , n403020 , n403021 , n55792 , n403023 , n403024 , n55795 , n403026 , n403027 , n55798 , 
 n403029 , n403030 , n55801 , n55802 , n55803 , n403034 , n403035 , n55806 , n403037 , n55808 , 
 n403039 , n403040 , n55811 , n403042 , n403043 , n55814 , n403045 , n55816 , n55817 , n403048 , 
 n55819 , n403050 , n55821 , n403052 , n403053 , n55824 , n403055 , n403056 , n55827 , n403058 , 
 n55829 , n55830 , n55831 , n403062 , n403063 , n55834 , n403065 , n403066 , n55837 , n403068 , 
 n403069 , n55840 , n403071 , n403072 , n55843 , n55844 , n55845 , n55846 , n403077 , n55848 , 
 n403079 , n403080 , n403081 , n55852 , n403083 , n403084 , n55855 , n403086 , n55857 , n403088 , 
 n403089 , n403090 , n55861 , n403092 , n403093 , n55864 , n55865 , n403096 , n55867 , n55868 , 
 n55869 , n55870 , n55871 , n55872 , n55873 , n55874 , n55875 , n403106 , n55877 , n403108 , 
 n403109 , n403110 , n403111 , n55882 , n403113 , n403114 , n55885 , n55886 , n403117 , n403118 , 
 n55889 , n403120 , n403121 , n55892 , n403123 , n403124 , n55895 , n403126 , n55897 , n403128 , 
 n403129 , n55900 , n403131 , n55902 , n403133 , n403134 , n55905 , n403136 , n55907 , n403138 , 
 n403139 , n55910 , n403141 , n55912 , n403143 , n403144 , n55915 , n403146 , n403147 , n55918 , 
 n55919 , n403150 , n403151 , n55922 , n55923 , n403154 , n403155 , n403156 , n55927 , n403158 , 
 n403159 , n55930 , n403161 , n403162 , n55933 , n403164 , n403165 , n55936 , n403167 , n403168 , 
 n55939 , n55940 , n403171 , n55942 , n55943 , n55944 , n403175 , n403176 , n403177 , n55948 , 
 n403179 , n55950 , n403181 , n403182 , n55953 , n403184 , n403185 , n55956 , n55957 , n403188 , 
 n55959 , n55960 , n403191 , n403192 , n55963 , n403194 , n403195 , n403196 , n55967 , n403198 , 
 n55969 , n403200 , n403201 , n55972 , n55973 , n55974 , n55975 , n55976 , n55977 , n55978 , 
 n55979 , n55980 , n55981 , n55982 , n55983 , n55984 , n403215 , n403216 , n55987 , n403218 , 
 n403219 , n55990 , n55991 , n403222 , n403223 , n55994 , n403225 , n55996 , n55997 , n55998 , 
 n403229 , n403230 , n56001 , n403232 , n56003 , n403234 , n403235 , n403236 , n403237 , n56008 , 
 n56009 , n403240 , n56011 , n56012 , n403243 , n403244 , n403245 , n56016 , n403247 , n403248 , 
 n56019 , n56020 , n403251 , n403252 , n56023 , n403254 , n403255 , n56026 , n403257 , n403258 , 
 n56029 , n56030 , n403261 , n403262 , n403263 , n56034 , n403265 , n403266 , n56037 , n56038 , 
 n403269 , n403270 , n56041 , n56042 , n56043 , n56044 , n56045 , n56046 , n56047 , n403278 , 
 n403279 , n56050 , n403281 , n56052 , n403283 , n403284 , n56055 , n56056 , n403287 , n56058 , 
 n56059 , n403290 , n403291 , n56062 , n403293 , n56064 , n403295 , n403296 , n56067 , n403298 , 
 n403299 , n56070 , n403301 , n403302 , n403303 , n56074 , n403305 , n403306 , n403307 , n56078 , 
 n403309 , n403310 , n56081 , n403312 , n403313 , n56084 , n403315 , n403316 , n56087 , n403318 , 
 n403319 , n56090 , n56091 , n403322 , n403323 , n403324 , n56095 , n403326 , n403327 , n56098 , 
 n56099 , n403330 , n403331 , n56102 , n56103 , n56104 , n403335 , n403336 , n56107 , n56108 , 
 n56109 , n403340 , n56111 , n56112 , n56113 , n56114 , n56115 , n403346 , n56117 , n56118 , 
 n56119 , n403350 , n403351 , n56122 , n403353 , n403354 , n403355 , n56126 , n403357 , n56128 , 
 n403359 , n403360 , n56131 , n403362 , n403363 , n403364 , n56135 , n403366 , n56137 , n403368 , 
 n56139 , n56140 , n403371 , n403372 , n56143 , n403374 , n403375 , n56146 , n403377 , n403378 , 
 n56149 , n56150 , n403381 , n403382 , n56153 , n403384 , n403385 , n56156 , n403387 , n403388 , 
 n56159 , n403390 , n56161 , n403392 , n56163 , n56164 , n403395 , n403396 , n56167 , n403398 , 
 n403399 , n56170 , n403401 , n403402 , n56173 , n403404 , n56175 , n56176 , n56177 , n403408 , 
 n56179 , n56180 , n56181 , n403412 , n403413 , n56184 , n56185 , n403416 , n56187 , n403418 , 
 n403419 , n403420 , n56191 , n403422 , n403423 , n56194 , n403425 , n403426 , n403427 , n56198 , 
 n403429 , n56200 , n403431 , n56202 , n56203 , n403434 , n403435 , n56206 , n403437 , n403438 , 
 n56209 , n403440 , n403441 , n56212 , n56213 , n403444 , n56215 , n403446 , n56217 , n56218 , 
 n403449 , n403450 , n56221 , n403452 , n403453 , n56224 , n403455 , n403456 , n403457 , n56228 , 
 n403459 , n403460 , n56231 , n403462 , n403463 , n56234 , n403465 , n403466 , n56237 , n403468 , 
 n56239 , n403470 , n403471 , n56242 , n56243 , n56244 , n403475 , n403476 , n56247 , n56248 , 
 n56249 , n403480 , n403481 , n56252 , n56253 , n56254 , n403485 , n56256 , n56257 , n56258 , 
 n56259 , n56260 , n403491 , n56262 , n56263 , n56264 , n403495 , n403496 , n56267 , n403498 , 
 n56269 , n403500 , n56271 , n56272 , n56273 , n403504 , n56275 , n403506 , n403507 , n56278 , 
 n403509 , n403510 , n56281 , n403512 , n403513 , n56284 , n56285 , n56286 , n403517 , n403518 , 
 n56289 , n56290 , n56291 , n403522 , n56293 , n403524 , n56295 , n56296 , n403527 , n56298 , 
 n56299 , n56300 , n56301 , n56302 , n56303 , n403534 , n56305 , n403536 , n403537 , n56308 , 
 n56309 , n403540 , n403541 , n403542 , n403543 , n403544 , n56335 , n403546 , n56337 , n56338 , 
 n403549 , n403550 , n56341 , n403552 , n403553 , n56344 , n403555 , n403556 , n56347 , n403558 , 
 n56349 , n403560 , n56351 , n56352 , n403563 , n56354 , n403565 , n56356 , n403567 , n403568 , 
 n56359 , n56360 , n403571 , n403572 , n56363 , n403574 , n403575 , n56366 , n403577 , n403578 , 
 n403579 , n56370 , n403581 , n403582 , n56373 , n403584 , n403585 , n56376 , n56378 , n403588 , 
 n403589 , n56381 , n403591 , n56383 , n403593 , n56385 , n403595 , n403596 , n56388 , n56389 , 
 n403599 , n403600 , n56392 , n403602 , n403603 , n56395 , n403605 , n56397 , n403607 , n56399 , 
 n56400 , n56401 , n56402 , n56403 , n56404 , n403614 , n56406 , n56407 , n56408 , n403618 , 
 n403619 , n56411 , n56412 , n403622 , n403623 , n56415 , n56416 , n56417 , n56418 , n403628 , 
 n56420 , n403630 , n56422 , n56423 , n403633 , n403634 , n56426 , n403636 , n403637 , n56429 , 
 n403639 , n56431 , n56432 , n56449 , n56450 , n56451 , n56452 , n56453 , n56454 , n56455 , 
 n56456 , n403650 , n56458 , n403652 , n56460 , n56461 , n56462 , n56463 , n56464 , n403658 , 
 n56466 , n403660 , n56468 , n403662 , n56470 , n56471 , n403665 , n403666 , n56474 , n403668 , 
 n403669 , n56477 , n403671 , n403672 , n56480 , n403674 , n403675 , n56483 , n56484 , n403678 , 
 n403679 , n56487 , n403681 , n403682 , n56490 , n403684 , n403685 , n56493 , n403687 , n56495 , 
 n56496 , n403690 , n56498 , n403692 , n56500 , n56501 , n403695 , n403696 , n56504 , n403698 , 
 n403699 , n56507 , n403701 , n56509 , n56510 , n56511 , n56512 , n56513 , n56514 , n56515 , 
 n56516 , n403710 , n56518 , n403712 , n56520 , n403714 , n56522 , n403716 , n56524 , n403718 , 
 n403719 , n56527 , n403721 , n56529 , n403723 , n56531 , n403725 , n56533 , n56534 , n403728 , 
 n56536 , n403730 , n56538 , n403732 , n403733 , n56541 , n56542 , n56543 , n56544 , n403738 , 
 n403739 , n56547 , n403741 , n56549 , n56550 , n56551 , n56552 , n403746 , n403747 , n56555 , 
 n403749 , n403750 , n56558 , n403752 , n56560 , n56561 , n56562 , n403756 , n56564 , n403758 , 
 n403759 , n56567 , n56568 , n56569 , n56570 , n56571 , n403765 , n403766 , n56574 , n56575 , 
 n403769 , n56577 , n56578 , n403772 , n403773 , n56581 , n403775 , n403776 , n56584 , n403778 , 
 n403779 , n56587 , n56588 , n403782 , n56590 , n403784 , n56592 , n56593 , n56594 , n403788 , 
 n56596 , n403790 , n56598 , n56599 , n403793 , n403794 , n56602 , n403796 , n403797 , n56605 , 
 n403799 , n56607 , n56608 , n56609 , n56610 , n56611 , n403805 , n56613 , n403807 , n56615 , 
 n403809 , n56617 , n56618 , n403812 , n403813 , n56621 , n403815 , n403816 , n56624 , n403818 , 
 n56626 , n56627 , n56628 , n56629 , n56630 , n56631 , n403825 , n56633 , n56634 , n56635 , 
 n403829 , n56637 , n403831 , n56639 , n56640 , n403834 , n403835 , n56643 , n403837 , n403838 , 
 n56646 , n403840 , n403841 , n56649 , n403843 , n56651 , n56652 , n403846 , n403847 , n56655 , 
 n403849 , n403850 , n56658 , n403852 , n56660 , n56661 , n56662 , n56663 , n403857 , n56665 , 
 n403859 , n56667 , n56668 , n403862 , n403863 , n56671 , n56672 , n403866 , n56674 , n56675 , 
 n56676 , n56677 , n403871 , n403872 , n56680 , n56681 , n56682 , n403876 , n56684 , n403878 , 
 n56686 , n56687 , n403881 , n56689 , n403883 , n403884 , n56692 , n403886 , n403887 , n56695 , 
 n403889 , n56697 , n56698 , n56699 , n403893 , n56701 , n403895 , n403896 , n56704 , n403898 , 
 n403899 , n56707 , n403901 , n403902 , n56710 , n56711 , n56712 , n403906 , n403907 , n56715 , 
 n403909 , n403910 , n56718 , n56719 , n56720 , n403914 , n56722 , n403916 , n56724 , n56725 , 
 n403919 , n403920 , n56728 , n403922 , n56730 , n56731 , n56732 , n56733 , n56734 , n56735 , 
 n56736 , n56737 , n56738 , n56739 , n56740 , n56741 , n56742 , n56743 , n56744 , n403938 , 
 n56746 , n403940 , n56748 , n56749 , n56750 , n56751 , n56752 , n403946 , n403947 , n403948 , 
 n56756 , n56757 , n403951 , n56759 , n56760 , n403954 , n403955 , n56763 , n403957 , n56765 , 
 n56766 , n56767 , n56768 , n56769 , n403963 , n403964 , n56772 , n56773 , n403967 , n56775 , 
 n56776 , n403970 , n56778 , n56779 , n403973 , n403974 , n56782 , n403976 , n56784 , n56785 , 
 n56803 , n56804 , n56805 , n56808 , n56809 , n56810 , n403985 , n56812 , n403987 , n56814 , 
 n56815 , n56816 , n56817 , n56818 , n56819 , n403994 , n403995 , n56822 , n403997 , n56824 , 
 n403999 , n56826 , n404001 , n404002 , n56829 , n404004 , n56831 , n56832 , n404007 , n404008 , 
 n56835 , n56836 , n404011 , n404012 , n404013 , n56840 , n404015 , n56842 , n56843 , n404018 , 
 n404019 , n56846 , n56847 , n404022 , n56849 , n56850 , n404025 , n56852 , n56853 , n56854 , 
 n56855 , n56856 , n404031 , n56858 , n404033 , n56860 , n56861 , n404036 , n404037 , n56864 , 
 n404039 , n404040 , n56867 , n404042 , n404043 , n56870 , n404045 , n56872 , n56873 , n404048 , 
 n404049 , n56876 , n404051 , n404052 , n56879 , n404054 , n56881 , n404056 , n56883 , n404058 , 
 n56885 , n56886 , n404061 , n404062 , n56889 , n404064 , n404065 , n56892 , n404067 , n404068 , 
 n56895 , n404070 , n56897 , n56898 , n404073 , n56900 , n404075 , n56902 , n404077 , n404078 , 
 n56905 , n404080 , n56907 , n56908 , n56909 , n404084 , n404085 , n56912 , n404087 , n56914 , 
 n404089 , n56916 , n56917 , n404092 , n56919 , n404094 , n56921 , n404096 , n404097 , n56924 , 
 n404099 , n404100 , n404101 , n56928 , n404103 , n404104 , n56931 , n404106 , n404107 , n56934 , 
 n404109 , n56936 , n56937 , n56938 , n56939 , n56940 , n56941 , n56942 , n56943 , n56944 , 
 n56945 , n56946 , n56947 , n56948 , n404123 , n56950 , n56951 , n56952 , n56953 , n56954 , 
 n56955 , n404130 , n404131 , n56958 , n404133 , n56960 , n404135 , n56962 , n56963 , n404138 , 
 n404139 , n56966 , n404141 , n404142 , n56969 , n404144 , n404145 , n56972 , n56973 , n404148 , 
 n404149 , n56976 , n404151 , n404152 , n56979 , n404154 , n404155 , n56982 , n404157 , n56984 , 
 n404159 , n56986 , n56987 , n404162 , n404163 , n56990 , n404165 , n404166 , n56993 , n404168 , 
 n404169 , n56996 , n404171 , n56998 , n56999 , n404174 , n404175 , n57002 , n404177 , n404178 , 
 n57005 , n404180 , n404181 , n57008 , n57009 , n404184 , n404185 , n57012 , n57013 , n404188 , 
 n57015 , n404190 , n57017 , n57018 , n404193 , n404194 , n57021 , n404196 , n404197 , n57024 , 
 n404199 , n57026 , n57027 , n57028 , n57029 , n404204 , n57031 , n404206 , n57033 , n57034 , 
 n404209 , n404210 , n57037 , n404212 , n404213 , n57040 , n404215 , n57042 , n57043 , n57044 , 
 n404219 , n404220 , n57047 , n404222 , n57049 , n57050 , n404225 , n57052 , n404227 , n57054 , 
 n57055 , n404230 , n404231 , n57058 , n404233 , n404234 , n57061 , n404236 , n404237 , n57064 , 
 n404239 , n57066 , n57067 , n404242 , n404243 , n57070 , n404245 , n404246 , n57073 , n404248 , 
 n57075 , n404250 , n57077 , n404252 , n57079 , n404254 , n404255 , n57082 , n57083 , n57084 , 
 n404259 , n404260 , n57087 , n57088 , n57089 , n404264 , n57091 , n57092 , n57093 , n57094 , 
 n404269 , n57096 , n404271 , n57098 , n57099 , n57100 , n57101 , n57102 , n57103 , n404278 , 
 n57105 , n57106 , n404281 , n404282 , n57109 , n404284 , n57111 , n404286 , n57113 , n404288 , 
 n57115 , n57116 , n404291 , n404292 , n57119 , n404294 , n404295 , n57122 , n404297 , n404298 , 
 n57125 , n57126 , n404301 , n404302 , n57129 , n404304 , n404305 , n57132 , n404307 , n404308 , 
 n57135 , n404310 , n57137 , n57138 , n404313 , n404314 , n57141 , n57142 , n404317 , n57144 , 
 n57145 , n57146 , n57147 , n57148 , n57149 , n57150 , n404325 , n57152 , n404327 , n404328 , 
 n404329 , n57156 , n404331 , n57158 , n404333 , n57160 , n57161 , n404336 , n404337 , n57164 , 
 n404339 , n404340 , n57167 , n404342 , n404343 , n57170 , n404345 , n57172 , n404347 , n404348 , 
 n57175 , n404350 , n404351 , n57178 , n404353 , n57180 , n57181 , n57182 , n57183 , n57184 , 
 n57185 , n57186 , n57187 , n57188 , n57189 , n57190 , n57191 , n57192 , n57193 , n57194 , 
 n57195 , n57196 , n57197 , n57198 , n57199 , n404374 , n57201 , n404376 , n57203 , n404378 , 
 n57205 , n404380 , n404381 , n57208 , n57209 , n57210 , n404385 , n57212 , n57213 , n57214 , 
 n57215 , n57216 , n57217 , n57218 , n57219 , n57220 , n57221 , n404396 , n57223 , n404398 , 
 n404399 , n404400 , n404401 , n57228 , n404403 , n404404 , n57231 , n404406 , n404407 , n57234 , 
 n404409 , n57236 , n404411 , n57238 , n57239 , n404414 , n404415 , n57242 , n404417 , n404418 , 
 n57245 , n404420 , n404421 , n404422 , n57249 , n404424 , n404425 , n57252 , n57253 , n404428 , 
 n57255 , n57256 , n404431 , n404432 , n57259 , n57260 , n57261 , n404436 , n57263 , n57264 , 
 n57265 , n404440 , n57267 , n57268 , n57269 , n57270 , n404445 , n404446 , n57273 , n57274 , 
 n404449 , n404450 , n57277 , n57278 , n404453 , n404454 , n57281 , n404456 , n404457 , n57284 , 
 n404459 , n57286 , n404461 , n57288 , n57289 , n57290 , n404465 , n57292 , n57293 , n57294 , 
 n57295 , n57296 , n404471 , n57298 , n404473 , n57300 , n404475 , n57302 , n57303 , n404478 , 
 n404479 , n57306 , n404481 , n404482 , n57309 , n404484 , n404485 , n404486 , n57313 , n404488 , 
 n404489 , n57316 , n57317 , n404492 , n57319 , n57320 , n404495 , n404496 , n57323 , n404498 , 
 n404499 , n57326 , n57327 , n57328 , n57329 , n404504 , n57331 , n404506 , n57333 , n57334 , 
 n404509 , n404510 , n57337 , n404512 , n404513 , n57340 , n404515 , n404516 , n57343 , n404518 , 
 n57345 , n57346 , n404521 , n404522 , n57349 , n404524 , n404525 , n57352 , n404527 , n404528 , 
 n57355 , n57356 , n404531 , n404532 , n57359 , n404534 , n57361 , n404536 , n57363 , n404538 , 
 n57365 , n57366 , n404541 , n404542 , n57369 , n404544 , n404545 , n57372 , n404547 , n404548 , 
 n57375 , n57376 , n404551 , n404552 , n57379 , n404554 , n404555 , n57382 , n404557 , n404558 , 
 n57385 , n57386 , n57387 , n404562 , n57389 , n404564 , n57391 , n404566 , n57393 , n57394 , 
 n57395 , n57396 , n57397 , n57398 , n57399 , n57400 , n57401 , n404576 , n57403 , n404578 , 
 n57405 , n57406 , n404581 , n57408 , n404583 , n57410 , n57411 , n57412 , n57413 , n57414 , 
 n404589 , n57416 , n404591 , n57418 , n404593 , n57420 , n57421 , n57422 , n57423 , n404598 , 
 n404599 , n57426 , n404601 , n404602 , n57429 , n404604 , n57431 , n57432 , n57433 , n404608 , 
 n57435 , n404610 , n404611 , n57438 , n404613 , n57440 , n404615 , n57442 , n57443 , n404618 , 
 n404619 , n57446 , n404621 , n404622 , n57449 , n404624 , n57451 , n57452 , n57453 , n404628 , 
 n404629 , n57456 , n404631 , n57458 , n404633 , n57460 , n57461 , n404636 , n404637 , n57464 , 
 n404639 , n57466 , n404641 , n57468 , n57469 , n57470 , n57471 , n57472 , n404647 , n404648 , 
 n57475 , n404650 , n57477 , n404652 , n404653 , n57480 , n404655 , n404656 , n57483 , n404658 , 
 n404659 , n57486 , n404661 , n404662 , n57489 , n404664 , n57491 , n57492 , n57493 , n57494 , 
 n57495 , n404670 , n404671 , n404672 , n57499 , n404674 , n57501 , n57502 , n57503 , n57504 , 
 n57505 , n57506 , n57507 , n404682 , n404683 , n57510 , n404685 , n404686 , n57513 , n404688 , 
 n404689 , n57516 , n404691 , n57518 , n404693 , n57520 , n57521 , n404696 , n404697 , n57524 , 
 n404699 , n404700 , n57527 , n404702 , n404703 , n57530 , n404705 , n57532 , n57533 , n404708 , 
 n404709 , n57536 , n404711 , n404712 , n57539 , n404714 , n404715 , n57542 , n57543 , n57544 , 
 n404719 , n404720 , n57547 , n404722 , n57549 , n404724 , n57551 , n404726 , n404727 , n57554 , 
 n57555 , n404730 , n57557 , n404732 , n57559 , n57560 , n404735 , n404736 , n57563 , n404738 , 
 n404739 , n57566 , n404741 , n404742 , n57569 , n404744 , n57571 , n404746 , n404747 , n57574 , 
 n404749 , n404750 , n57577 , n57578 , n404753 , n404754 , n57581 , n404756 , n57583 , n404758 , 
 n57585 , n57586 , n404761 , n57588 , n404763 , n404764 , n57591 , n404766 , n57593 , n404768 , 
 n57595 , n57596 , n404771 , n404772 , n57599 , n57600 , n404775 , n404776 , n57603 , n57604 , 
 n404779 , n404780 , n57607 , n57608 , n404783 , n404784 , n57611 , n404786 , n404787 , n57614 , 
 n404789 , n404790 , n57617 , n404792 , n57619 , n57620 , n57621 , n57622 , n404797 , n404798 , 
 n57625 , n404800 , n57627 , n57628 , n57629 , n57630 , n57631 , n57632 , n404807 , n57634 , 
 n404809 , n57636 , n404811 , n404812 , n57639 , n404814 , n404815 , n57642 , n404817 , n57644 , 
 n404819 , n57646 , n57647 , n404822 , n404823 , n57650 , n404825 , n404826 , n57653 , n404828 , 
 n57655 , n57656 , n57657 , n404832 , n404833 , n57660 , n404835 , n57662 , n57663 , n57664 , 
 n57665 , n57666 , n57667 , n57668 , n57669 , n57670 , n57671 , n57672 , n404847 , n57674 , 
 n404849 , n57676 , n57677 , n404852 , n404853 , n57680 , n404855 , n404856 , n57683 , n404858 , 
 n404859 , n57686 , n404861 , n404862 , n57689 , n404864 , n57691 , n57692 , n404867 , n404868 , 
 n57695 , n404870 , n404871 , n57698 , n404873 , n57700 , n57701 , n404876 , n57703 , n57704 , 
 n57705 , n404880 , n57707 , n57708 , n57709 , n57710 , n404885 , n57712 , n57713 , n57714 , 
 n404889 , n404890 , n57717 , n57718 , n404893 , n404894 , n57721 , n57722 , n57723 , n57724 , 
 n404899 , n404900 , n57727 , n404902 , n57729 , n57730 , n57731 , n57732 , n57733 , n57734 , 
 n404909 , n57736 , n57737 , n57738 , n404913 , n57740 , n57741 , n57742 , n57743 , n404918 , 
 n57745 , n404920 , n404921 , n57748 , n57749 , n57750 , n57751 , n57752 , n57753 , n57754 , 
 n57755 , n57768 , n57769 , n57770 , n57771 , n57776 , n57777 , n57778 , n404937 , n57780 , 
 n404939 , n57782 , n57783 , n404942 , n57785 , n404944 , n57787 , n57788 , n57789 , n57790 , 
 n57791 , n57792 , n57793 , n404952 , n57797 , n57800 , n57801 , n57802 , n57803 , n404958 , 
 n57805 , n404960 , n404961 , n57808 , n57809 , n404964 , n57811 , n404966 , n57813 , n57814 , 
 n57816 , n57817 , n57820 , n57821 , n57822 , n57823 , n57824 , n57825 , n404977 , n57827 , 
 n404979 , n57829 , n57830 , n57831 , n404983 , n57833 , n57834 , n404986 , n57836 , n404988 , 
 n57838 , n57839 , n57840 , n404992 , n57842 , n404994 , n57844 , n57845 , n404997 , n57847 , 
 n404999 , n57849 , n57850 , n405002 , n405003 , n57853 , n405005 , n405006 , n57856 , n405008 , 
 n405009 , n405010 , n57860 , n405012 , n405013 , n57863 , n405015 , n405016 , n57866 , n57867 , 
 n57868 , n57869 , n57870 , n57871 , n57872 , n57873 , n57874 , n57875 , n57876 , n57877 , 
 n57878 , n57879 , n57880 , n57881 , n57882 , n57883 , n57884 , n57885 , n57886 , n57887 , 
 n57888 , n57889 , n57890 , n57891 , n405043 , n405044 , n405045 , n57895 , n405047 , n57897 , 
 n405049 , n405050 , n57900 , n405052 , n57902 , n57903 , n405055 , n57905 , n405057 , n405058 , 
 n57908 , n57909 , n57910 , n57911 , n57912 , n405064 , n57914 , n57915 , n405067 , n405068 , 
 n57918 , n57919 , n405071 , n57921 , n405073 , n57923 , n405075 , n57925 , n405077 , n405078 , 
 n57928 , n405080 , n57930 , n57931 , n405083 , n57933 , n405085 , n57935 , n57936 , n57937 , 
 n57938 , n57939 , n57940 , n57941 , n57942 , n57943 , n57944 , n405096 , n57946 , n405098 , 
 n57948 , n57949 , n405101 , n405102 , n57952 , n405104 , n405105 , n57955 , n405107 , n57957 , 
 n57958 , n57959 , n405111 , n405112 , n57962 , n405114 , n57964 , n57965 , n57966 , n405118 , 
 n57968 , n405120 , n57970 , n57971 , n405123 , n405124 , n57974 , n405126 , n405127 , n57977 , 
 n405129 , n405130 , n57980 , n405132 , n57982 , n57983 , n405135 , n405136 , n57986 , n405138 , 
 n57988 , n57989 , n57990 , n57991 , n57992 , n57993 , n57994 , n57995 , n57996 , n57997 , 
 n57998 , n57999 , n58000 , n58001 , n58002 , n58003 , n58004 , n405156 , n58006 , n405158 , 
 n58008 , n58009 , n405161 , n58011 , n405163 , n58013 , n58014 , n405166 , n405167 , n58017 , 
 n405169 , n405170 , n58020 , n405172 , n405173 , n405174 , n58024 , n405176 , n405177 , n58027 , 
 n405179 , n58029 , n58030 , n58031 , n58032 , n58033 , n58034 , n58035 , n58036 , n58037 , 
 n58038 , n405190 , n405191 , n58041 , n58042 , n405194 , n405195 , n58045 , n405197 , n405198 , 
 n58048 , n58049 , n405201 , n405202 , n405203 , n58053 , n405205 , n405206 , n58056 , n58057 , 
 n405209 , n405210 , n405211 , n58061 , n405213 , n58063 , n405215 , n405216 , n58066 , n405218 , 
 n405219 , n58069 , n58070 , n405222 , n405223 , n405224 , n58074 , n405226 , n58076 , n405228 , 
 n405229 , n58079 , n405231 , n405232 , n58082 , n58083 , n58084 , n58085 , n58086 , n58087 , 
 n58088 , n58089 , n58090 , n405242 , n405243 , n58093 , n405245 , n405246 , n58096 , n58097 , 
 n405249 , n405250 , n58100 , n405252 , n58102 , n405254 , n58104 , n58105 , n58106 , n58107 , 
 n405259 , n405260 , n58110 , n405262 , n405263 , n58113 , n405265 , n405266 , n58116 , n405268 , 
 n58118 , n405270 , n58120 , n58121 , n405273 , n405274 , n405275 , n58125 , n405277 , n405278 , 
 n58128 , n405280 , n405281 , n58131 , n405283 , n405284 , n58134 , n58135 , n405287 , n405288 , 
 n58138 , n58139 , n405291 , n405292 , n58142 , n405294 , n405295 , n405296 , n58146 , n405298 , 
 n58148 , n405300 , n405301 , n405302 , n58152 , n58153 , n405305 , n405306 , n58156 , n58157 , 
 n58158 , n58159 , n58160 , n58161 , n58162 , n58163 , n58164 , n58165 , n58166 , n405318 , 
 n405319 , n58169 , n405321 , n405322 , n58172 , n58173 , n405325 , n405326 , n58176 , n58177 , 
 n58178 , n405330 , n405331 , n58181 , n405333 , n58183 , n405335 , n405336 , n405337 , n58187 , 
 n58188 , n405340 , n405341 , n405342 , n58192 , n405344 , n405345 , n58195 , n58196 , n405348 , 
 n405349 , n58199 , n58200 , n58201 , n405353 , n405354 , n58204 , n58205 , n405357 , n405358 , 
 n58208 , n58209 , n405361 , n405362 , n58212 , n405364 , n58214 , n405366 , n58216 , n58217 , 
 n58218 , n405370 , n405371 , n58221 , n58222 , n58223 , n405375 , n58225 , n58226 , n405378 , 
 n405379 , n58229 , n405381 , n405382 , n58232 , n405384 , n405385 , n405386 , n58236 , n405388 , 
 n405389 , n58239 , n405391 , n405392 , n58242 , n405394 , n405395 , n58245 , n405397 , n405398 , 
 n58248 , n405400 , n405401 , n58251 , n405403 , n405404 , n405405 , n58255 , n405407 , n405408 , 
 n58258 , n405410 , n405411 , n405412 , n58262 , n405414 , n405415 , n58265 , n405417 , n405418 , 
 n58268 , n405420 , n405421 , n58271 , n405423 , n405424 , n58274 , n58275 , n58276 , n405428 , 
 n405429 , n58279 , n58280 , n405432 , n405433 , n58283 , n405435 , n405436 , n58286 , n405438 , 
 n58288 , n405440 , n405441 , n58291 , n405443 , n405444 , n405445 , n405446 , n58296 , n405448 , 
 n405449 , n58299 , n58300 , n405452 , n405453 , n405454 , n58304 , n405456 , n405457 , n58307 , 
 n58308 , n405460 , n405461 , n405462 , n405463 , n58313 , n405465 , n405466 , n58316 , n58317 , 
 n405469 , n405470 , n405471 , n58321 , n405473 , n405474 , n58324 , n405476 , n405477 , n58327 , 
 n58328 , n405480 , n405481 , n58331 , n405483 , n405484 , n58334 , n405486 , n405487 , n58337 , 
 n58338 , n405490 , n405491 , n58341 , n405493 , n405494 , n405495 , n58345 , n405497 , n58347 , 
 n405499 , n405500 , n58350 , n58351 , n58352 , n405504 , n405505 , n58355 , n405507 , n405508 , 
 n58358 , n58359 , n405511 , n405512 , n58362 , n405514 , n405515 , n58365 , n58366 , n58367 , 
 n405519 , n405520 , n58370 , n405522 , n58372 , n405524 , n58374 , n58375 , n58376 , n58377 , 
 n405529 , n405530 , n58380 , n405532 , n405533 , n58383 , n405535 , n405536 , n58386 , n405538 , 
 n405539 , n58389 , n405541 , n405542 , n58392 , n405544 , n405545 , n58395 , n405547 , n58397 , 
 n58398 , n58399 , n58400 , n58401 , n58402 , n58403 , n405555 , n58405 , n405557 , n58407 , 
 n405559 , n58409 , n58410 , n58411 , n405563 , n405564 , n58414 , n58415 , n58416 , n405568 , 
 n58418 , n58419 , n405571 , n58421 , n405573 , n405574 , n58424 , n405576 , n405577 , n58427 , 
 n405579 , n405580 , n405581 , n58431 , n405583 , n58433 , n405585 , n405586 , n58436 , n405588 , 
 n405589 , n58439 , n405591 , n405592 , n58442 , n58443 , n58444 , n405596 , n405597 , n58447 , 
 n405599 , n58449 , n58450 , n58451 , n58452 , n58453 , n58454 , n58455 , n58456 , n58457 , 
 n58458 , n58459 , n58460 , n58461 , n58462 , n58463 , n58464 , n58465 , n405617 , n58467 , 
 n405619 , n58469 , n58470 , n405622 , n58472 , n405624 , n405625 , n58475 , n405627 , n58477 , 
 n58478 , n58479 , n58480 , n58481 , n58482 , n58483 , n58484 , n58485 , n405637 , n58487 , 
 n405639 , n58489 , n58490 , n405642 , n405643 , n58493 , n58494 , n405646 , n58496 , n58497 , 
 n405649 , n58499 , n405651 , n405652 , n405653 , n58503 , n58504 , n405656 , n58506 , n58507 , 
 n405659 , n58509 , n405661 , n58511 , n58512 , n405664 , n405665 , n58515 , n405667 , n58517 , 
 n405669 , n58519 , n58520 , n405672 , n58522 , n405674 , n58524 , n58525 , n405677 , n405678 , 
 n58528 , n405680 , n405681 , n58531 , n405683 , n405684 , n405685 , n58535 , n405687 , n405688 , 
 n58538 , n405690 , n58540 , n58541 , n58542 , n58543 , n58544 , n58545 , n58546 , n405698 , 
 n405699 , n58549 , n405701 , n58551 , n58552 , n58553 , n58554 , n58555 , n58556 , n58557 , 
 n58558 , n58559 , n58560 , n58561 , n405713 , n58563 , n405715 , n58565 , n58566 , n58567 , 
 n58568 , n58569 , n58570 , n58571 , n58572 , n58573 , n405725 , n58575 , n58576 , n405728 , 
 n58578 , n58579 , n58580 , n58581 , n58582 , n405734 , n58584 , n405736 , n405737 , n58587 , 
 n405739 , n58589 , n58590 , n405742 , n405743 , n58593 , n405745 , n405746 , n58596 , n405748 , 
 n405749 , n405750 , n58600 , n405752 , n58602 , n58603 , n58604 , n58605 , n405757 , n405758 , 
 n58608 , n405760 , n58610 , n405762 , n58612 , n405764 , n58614 , n58615 , n405767 , n405768 , 
 n58618 , n405770 , n405771 , n58621 , n405773 , n58623 , n58624 , n58625 , n58626 , n405778 , 
 n58628 , n405780 , n58630 , n58631 , n405783 , n58633 , n405785 , n405786 , n405787 , n58637 , 
 n405789 , n405790 , n58640 , n405792 , n405793 , n405794 , n58644 , n405796 , n58646 , n58647 , 
 n58648 , n58649 , n58650 , n58651 , n405803 , n58653 , n58654 , n58655 , n405807 , n405808 , 
 n58658 , n405810 , n405811 , n58661 , n405813 , n58663 , n58664 , n405816 , n405817 , n58667 , 
 n405819 , n405820 , n58670 , n405822 , n58672 , n58673 , n58674 , n58675 , n58676 , n58677 , 
 n58678 , n58679 , n58680 , n58681 , n58682 , n58683 , n58684 , n58685 , n58686 , n58687 , 
 n405839 , n58689 , n405841 , n58691 , n58692 , n405844 , n405845 , n58695 , n405847 , n405848 , 
 n58698 , n405850 , n405851 , n58701 , n405853 , n58703 , n58704 , n405856 , n405857 , n58707 , 
 n405859 , n405860 , n58710 , n405862 , n405863 , n405864 , n58714 , n405866 , n58716 , n58717 , 
 n405869 , n405870 , n58720 , n405872 , n405873 , n58723 , n405875 , n405876 , n58726 , n405878 , 
 n58728 , n58729 , n405881 , n405882 , n58732 , n405884 , n405885 , n58735 , n405887 , n405888 , 
 n58738 , n405890 , n58740 , n405892 , n58742 , n58743 , n405895 , n58745 , n405897 , n405898 , 
 n58748 , n405900 , n58750 , n58751 , n405903 , n405904 , n58754 , n405906 , n405907 , n58757 , 
 n405909 , n405910 , n405911 , n58761 , n405913 , n405914 , n58764 , n405916 , n405917 , n58767 , 
 n405919 , n58769 , n405921 , n58771 , n58772 , n58773 , n58774 , n58775 , n58776 , n58777 , 
 n58778 , n58779 , n405931 , n58781 , n405933 , n58783 , n58784 , n58785 , n58786 , n58787 , 
 n58788 , n58789 , n58790 , n58791 , n58792 , n405944 , n58794 , n58795 , n58796 , n405948 , 
 n58798 , n58799 , n405951 , n405952 , n58802 , n405954 , n405955 , n58805 , n405957 , n58807 , 
 n405959 , n405960 , n58810 , n405962 , n58812 , n58813 , n405965 , n58815 , n405967 , n58817 , 
 n58818 , n405970 , n405971 , n58821 , n405973 , n405974 , n58824 , n405976 , n58826 , n58827 , 
 n405979 , n405980 , n58830 , n405982 , n58832 , n58833 , n58834 , n58835 , n58836 , n58837 , 
 n58838 , n405990 , n405991 , n58841 , n405993 , n405994 , n58844 , n405996 , n58846 , n58847 , 
 n405999 , n406000 , n58850 , n406002 , n406003 , n58853 , n406005 , n58855 , n58856 , n406008 , 
 n58858 , n406010 , n58860 , n58861 , n406013 , n406014 , n58864 , n406016 , n406017 , n58867 , 
 n406019 , n58869 , n58870 , n58871 , n406023 , n406024 , n58874 , n406026 , n58876 , n58877 , 
 n406029 , n406030 , n58880 , n406032 , n58882 , n406034 , n58884 , n58885 , n58886 , n58887 , 
 n58888 , n58889 , n58890 , n58891 , n406043 , n58893 , n406045 , n406046 , n58896 , n406048 , 
 n58898 , n58899 , n406051 , n406052 , n406053 , n406054 , n58927 , n406056 , n58929 , n58930 , 
 n406059 , n58932 , n406061 , n58934 , n58935 , n406064 , n58937 , n406066 , n58939 , n406068 , 
 n406069 , n58942 , n406071 , n406072 , n406073 , n58946 , n406075 , n406076 , n58949 , n406078 , 
 n406079 , n58952 , n58953 , n58954 , n58955 , n58956 , n58957 , n58958 , n406087 , n406088 , 
 n58961 , n406090 , n406091 , n58964 , n406093 , n406094 , n58967 , n58968 , n406097 , n58970 , 
 n58971 , n406100 , n406101 , n58974 , n58976 , n406104 , n406105 , n58979 , n58980 , n58981 , 
 n406109 , n58983 , n58984 , n58985 , n406113 , n406114 , n58988 , n406116 , n406117 , n58991 , 
 n58992 , n58993 , n406121 , n406122 , n58996 , n58997 , n406125 , n58999 , n406127 , n59001 , 
 n59002 , n406130 , n406131 , n59005 , n59006 , n406134 , n59008 , n59009 , n406137 , n406138 , 
 n59012 , n406140 , n59014 , n406142 , n406143 , n59017 , n406145 , n59019 , n406147 , n59021 , 
 n406149 , n59023 , n59024 , n406152 , n406153 , n59027 , n406155 , n406156 , n59030 , n406158 , 
 n406159 , n59033 , n406161 , n59035 , n59036 , n406164 , n406165 , n59039 , n406167 , n406168 , 
 n59042 , n406170 , n59044 , n59045 , n406173 , n406174 , n59048 , n406176 , n406177 , n406178 , 
 n59052 , n406180 , n59054 , n406182 , n59056 , n59057 , n406185 , n406186 , n59060 , n406188 , 
 n59062 , n406190 , n59064 , n59065 , n406193 , n406194 , n59068 , n406196 , n406197 , n59071 , 
 n406199 , n406200 , n59074 , n59075 , n406203 , n406204 , n59078 , n406206 , n406207 , n59081 , 
 n406209 , n406210 , n59084 , n59085 , n59086 , n406214 , n406215 , n59089 , n59090 , n59091 , 
 n406219 , n59093 , n406221 , n406222 , n59096 , n406224 , n59098 , n406226 , n59100 , n59101 , 
 n59102 , n59103 , n406231 , n59105 , n59106 , n406234 , n59108 , n406236 , n59110 , n59111 , 
 n59112 , n59113 , n59114 , n59115 , n59116 , n59117 , n59118 , n59119 , n59120 , n59121 , 
 n59122 , n59123 , n406251 , n59125 , n59126 , n59127 , n406255 , n59129 , n59130 , n59131 , 
 n59132 , n59133 , n406261 , n406262 , n59136 , n59137 , n406265 , n59139 , n59140 , n406268 , 
 n406269 , n59143 , n406271 , n406272 , n59146 , n59147 , n59148 , n59149 , n59150 , n59151 , 
 n59152 , n59153 , n59154 , n59155 , n59156 , n406284 , n59158 , n59159 , n406287 , n59161 , 
 n406289 , n59163 , n406291 , n59165 , n59166 , n406294 , n406295 , n59169 , n406297 , n406298 , 
 n59172 , n406300 , n406301 , n59175 , n59176 , n406304 , n59178 , n406306 , n59180 , n59181 , 
 n406309 , n406310 , n59184 , n406312 , n406313 , n59187 , n406315 , n406316 , n406317 , n59191 , 
 n406319 , n406320 , n59194 , n406322 , n59196 , n59197 , n59198 , n406326 , n406327 , n59201 , 
 n406329 , n59203 , n59204 , n59205 , n59206 , n406334 , n59208 , n406336 , n59210 , n59211 , 
 n406339 , n59213 , n406341 , n406342 , n59216 , n406344 , n59218 , n406346 , n59220 , n59221 , 
 n406349 , n59223 , n406351 , n406352 , n59226 , n406354 , n59228 , n59229 , n59230 , n406358 , 
 n406359 , n59233 , n406361 , n59235 , n59236 , n406364 , n406365 , n59239 , n406367 , n406368 , 
 n59242 , n406370 , n59244 , n59245 , n406373 , n406374 , n59248 , n59249 , n406377 , n406378 , 
 n406379 , n59253 , n406381 , n59255 , n59256 , n406384 , n406385 , n59259 , n406387 , n406388 , 
 n59262 , n406390 , n406391 , n59265 , n406393 , n59267 , n59268 , n406396 , n406397 , n59271 , 
 n406399 , n406400 , n59274 , n406402 , n406403 , n59277 , n406405 , n59279 , n406407 , n59281 , 
 n59282 , n59283 , n59284 , n59285 , n406413 , n59287 , n406415 , n59289 , n406417 , n59291 , 
 n406419 , n406420 , n59294 , n406422 , n406423 , n59297 , n406425 , n406426 , n59300 , n406428 , 
 n406429 , n59303 , n406431 , n59305 , n406433 , n59307 , n406435 , n406436 , n59310 , n406438 , 
 n406439 , n59313 , n59314 , n406442 , n406443 , n59317 , n59318 , n406446 , n406447 , n406448 , 
 n59322 , n406450 , n406451 , n59325 , n59326 , n406454 , n59328 , n59329 , n406457 , n406458 , 
 n59332 , n59333 , n406461 , n406462 , n59336 , n59337 , n406465 , n406466 , n406467 , n406468 , 
 n59342 , n406470 , n406471 , n59345 , n59346 , n406474 , n406475 , n406476 , n59350 , n406478 , 
 n406479 , n59353 , n59354 , n406482 , n406483 , n406484 , n406485 , n59359 , n406487 , n406488 , 
 n59362 , n59363 , n406491 , n406492 , n406493 , n59367 , n406495 , n406496 , n59370 , n59371 , 
 n406499 , n406500 , n59374 , n406502 , n406503 , n59377 , n406505 , n406506 , n59380 , n59381 , 
 n406509 , n406510 , n406511 , n59385 , n406513 , n406514 , n59388 , n59389 , n406517 , n406518 , 
 n59392 , n59393 , n59394 , n406522 , n406523 , n59397 , n406525 , n59399 , n406527 , n59401 , 
 n59402 , n406530 , n406531 , n59405 , n59406 , n406534 , n406535 , n59409 , n59410 , n406538 , 
 n406539 , n59413 , n59414 , n406542 , n59416 , n59417 , n59418 , n406546 , n59420 , n59421 , 
 n59422 , n406550 , n59424 , n59425 , n59426 , n59427 , n59428 , n59429 , n59430 , n59431 , 
 n59432 , n59433 , n59434 , n59435 , n406563 , n59437 , n406565 , n406566 , n406567 , n59441 , 
 n406569 , n59443 , n406571 , n406572 , n406573 , n59447 , n59448 , n406576 , n406577 , n59451 , 
 n406579 , n59453 , n406581 , n406582 , n59456 , n59457 , n406585 , n406586 , n59460 , n59461 , 
 n406589 , n59463 , n59464 , n59465 , n59466 , n59467 , n59468 , n59469 , n406597 , n59471 , 
 n406599 , n406600 , n59474 , n406602 , n406603 , n59477 , n406605 , n59479 , n406607 , n406608 , 
 n59482 , n406610 , n406611 , n59485 , n59486 , n406614 , n406615 , n406616 , n59490 , n406618 , 
 n406619 , n59493 , n59494 , n406622 , n59496 , n59497 , n59498 , n406626 , n406627 , n406628 , 
 n59502 , n406630 , n59504 , n406632 , n406633 , n59507 , n406635 , n406636 , n59510 , n406638 , 
 n406639 , n59513 , n59514 , n406642 , n406643 , n406644 , n59518 , n406646 , n406647 , n59521 , 
 n59522 , n406650 , n406651 , n406652 , n406653 , n59527 , n406655 , n406656 , n59530 , n59531 , 
 n406659 , n406660 , n406661 , n59535 , n406663 , n406664 , n59538 , n59539 , n406667 , n406668 , 
 n59542 , n406670 , n406671 , n59545 , n406673 , n406674 , n59548 , n59549 , n406677 , n406678 , 
 n406679 , n59553 , n406681 , n406682 , n59556 , n59557 , n406685 , n406686 , n59560 , n59561 , 
 n59562 , n406690 , n406691 , n59565 , n59566 , n59567 , n406695 , n59569 , n59570 , n59571 , 
 n406699 , n406700 , n59574 , n406702 , n406703 , n59577 , n59578 , n406706 , n406707 , n59581 , 
 n406709 , n406710 , n406711 , n59585 , n406713 , n59587 , n406715 , n406716 , n406717 , n59591 , 
 n59592 , n406720 , n406721 , n59595 , n59596 , n406724 , n406725 , n59599 , n406727 , n406728 , 
 n59602 , n59603 , n406731 , n406732 , n59606 , n406734 , n59608 , n59609 , n59610 , n406738 , 
 n406739 , n59613 , n406741 , n406742 , n59616 , n59617 , n406745 , n406746 , n406747 , n59621 , 
 n406749 , n406750 , n59624 , n59625 , n406753 , n406754 , n59628 , n406756 , n59630 , n406758 , 
 n406759 , n59633 , n59634 , n406762 , n406763 , n59637 , n406765 , n59639 , n406767 , n59641 , 
 n406769 , n59643 , n406771 , n406772 , n59646 , n406774 , n406775 , n59649 , n59650 , n406778 , 
 n406779 , n406780 , n59654 , n406782 , n406783 , n59657 , n59658 , n406786 , n59660 , n59661 , 
 n59662 , n59663 , n59664 , n59665 , n59666 , n59667 , n59668 , n59669 , n406797 , n59671 , 
 n59672 , n59673 , n406801 , n59675 , n59676 , n59677 , n59678 , n59679 , n59680 , n59681 , 
 n59682 , n406810 , n59684 , n59685 , n59686 , n406814 , n406815 , n59689 , n406817 , n59691 , 
 n406819 , n59693 , n406821 , n406822 , n59696 , n406824 , n406825 , n59699 , n59700 , n406828 , 
 n406829 , n59703 , n59704 , n406832 , n59706 , n406834 , n59708 , n406836 , n59710 , n59711 , 
 n406839 , n406840 , n59714 , n406842 , n406843 , n59717 , n406845 , n406846 , n59720 , n59721 , 
 n59722 , n406850 , n59724 , n59725 , n59726 , n406854 , n59728 , n406856 , n59730 , n406858 , 
 n59732 , n59733 , n406861 , n406862 , n59736 , n406864 , n406865 , n59739 , n406867 , n406868 , 
 n59742 , n59743 , n406871 , n59745 , n406873 , n59747 , n59748 , n406876 , n406877 , n59751 , 
 n406879 , n406880 , n59754 , n406882 , n406883 , n406884 , n59758 , n406886 , n406887 , n59761 , 
 n406889 , n59763 , n59764 , n59765 , n59766 , n59767 , n406895 , n406896 , n59770 , n406898 , 
 n59772 , n406900 , n406901 , n59775 , n406903 , n406904 , n59778 , n59779 , n406907 , n59781 , 
 n406909 , n59783 , n59784 , n59785 , n59786 , n406914 , n59788 , n406916 , n406917 , n59791 , 
 n406919 , n406920 , n406921 , n59795 , n59796 , n406924 , n59798 , n59799 , n406927 , n406928 , 
 n59802 , n59803 , n406931 , n406932 , n59806 , n59807 , n59808 , n406936 , n59810 , n59811 , 
 n59812 , n406940 , n59814 , n406942 , n406943 , n406944 , n59818 , n406946 , n406947 , n406948 , 
 n59822 , n406950 , n406951 , n59825 , n406953 , n59827 , n406955 , n406956 , n59830 , n406958 , 
 n59832 , n406960 , n59834 , n59835 , n59836 , n406964 , n59838 , n406966 , n406967 , n406968 , 
 n406969 , n59843 , n406971 , n406972 , n59846 , n406974 , n406975 , n59849 , n59850 , n59851 , 
 n406979 , n59853 , n59854 , n59855 , n59856 , n59857 , n406985 , n59859 , n59860 , n406988 , 
 n59862 , n59863 , n59864 , n59865 , n59866 , n59867 , n59868 , n59869 , n59870 , n59871 , 
 n59872 , n59873 , n59874 , n59875 , n59876 , n59877 , n59878 , n59879 , n59880 , n59881 , 
 n59882 , n59883 , n59885 , n59886 , n407013 , n59891 , n59892 , n59893 , n59894 , n59895 , 
 n59896 , n59897 , n59898 , n59899 , n407023 , n59901 , n407025 , n59903 , n59904 , n407028 , 
 n407029 , n59907 , n407031 , n407032 , n59910 , n407034 , n407035 , n407036 , n59914 , n407038 , 
 n59916 , n407040 , n59918 , n59919 , n407043 , n407044 , n59922 , n59945 , n407047 , n407048 , 
 n59948 , n407050 , n59950 , n407052 , n59952 , n59953 , n407055 , n407056 , n59956 , n407058 , 
 n407059 , n59959 , n407061 , n407062 , n59962 , n407064 , n59964 , n407066 , n407067 , n59967 , 
 n407069 , n59969 , n407071 , n59971 , n407073 , n407074 , n59974 , n59975 , n59976 , n407078 , 
 n59978 , n59979 , n407081 , n407082 , n59982 , n59983 , n407085 , n59985 , n407087 , n59987 , 
 n407089 , n407090 , n59990 , n407092 , n59992 , n59993 , n59994 , n59995 , n59996 , n407098 , 
 n407099 , n59999 , n407101 , n60001 , n407103 , n407104 , n60004 , n407106 , n407107 , n60007 , 
 n407109 , n407110 , n60010 , n407112 , n407113 , n407114 , n60015 , n407116 , n407117 , n407118 , 
 n60021 , n407120 , n60023 , n60024 , n407123 , n60026 , n407125 , n60028 , n60029 , n407128 , 
 n407129 , n60032 , n60033 , n407132 , n60035 , n407134 , n60037 , n60038 , n60039 , n60040 , 
 n60041 , n60042 , n60043 , n407142 , n60045 , n407144 , n60047 , n60048 , n407147 , n60050 , 
 n60051 , n407150 , n407151 , n60054 , n407153 , n60056 , n407155 , n407156 , n407157 , n60060 , 
 n60061 , n407160 , n407161 , n60064 , n60065 , n60066 , n60067 , n60068 , n60069 , n60070 , 
 n60071 , n60072 , n407171 , n60074 , n60075 , n60076 , n407175 , n60078 , n407177 , n60080 , 
 n60081 , n407180 , n407181 , n60084 , n60085 , n407184 , n407185 , n60088 , n407187 , n60090 , 
 n60091 , n407190 , n407191 , n60094 , n60095 , n407194 , n407195 , n60098 , n407197 , n60100 , 
 n407199 , n60102 , n60103 , n407202 , n407203 , n60106 , n407205 , n407206 , n60109 , n407208 , 
 n60111 , n60112 , n60113 , n60114 , n407213 , n60116 , n60117 , n60118 , n60119 , n60120 , 
 n60121 , n60122 , n60123 , n60124 , n60125 , n60126 , n407225 , n60128 , n60129 , n60130 , 
 n407229 , n407230 , n407231 , n407232 , n60135 , n407234 , n407235 , n60138 , n60139 , n407238 , 
 n60141 , n60142 , n407241 , n60144 , n407243 , n60146 , n407245 , n407246 , n60149 , n407248 , 
 n60151 , n407250 , n60153 , n60154 , n60155 , n407254 , n60157 , n407256 , n407257 , n407258 , 
 n407259 , n60162 , n60163 , n407262 , n407263 , n60166 , n407265 , n407266 , n60169 , n407268 , 
 n407269 , n60172 , n60173 , n60174 , n407273 , n60176 , n407275 , n60178 , n407277 , n407278 , 
 n60181 , n407280 , n60183 , n60184 , n407283 , n60186 , n407285 , n60188 , n407287 , n60190 , 
 n60191 , n60192 , n60193 , n60194 , n60195 , n407294 , n60197 , n407296 , n60199 , n60200 , 
 n407299 , n407300 , n60203 , n407302 , n407303 , n60206 , n407305 , n407306 , n407307 , n60210 , 
 n60211 , n407310 , n60213 , n407312 , n407313 , n60216 , n60217 , n407316 , n60219 , n60220 , 
 n60221 , n407320 , n60223 , n407322 , n60225 , n60226 , n60227 , n407326 , n60229 , n60230 , 
 n407329 , n60232 , n407331 , n60234 , n60235 , n60236 , n407335 , n407336 , n60258 , n407338 , 
 n60260 , n60261 , n407341 , n60263 , n60264 , n60265 , n60266 , n407346 , n60268 , n407348 , 
 n407349 , n60271 , n407351 , n407352 , n60274 , n60275 , n407355 , n60277 , n60278 , n60279 , 
 n407359 , n407360 , n60282 , n407362 , n60284 , n407364 , n60286 , n60287 , n407367 , n407368 , 
 n60290 , n407370 , n407371 , n60293 , n407373 , n407374 , n60296 , n60297 , n407377 , n407378 , 
 n60300 , n407380 , n407381 , n60303 , n407383 , n407384 , n60306 , n60307 , n60308 , n60309 , 
 n60310 , n60311 , n60312 , n407392 , n60314 , n60315 , n60316 , n407396 , n407397 , n60319 , 
 n60320 , n60321 , n407401 , n407402 , n60324 , n407404 , n60326 , n60327 , n407407 , n60329 , 
 n407409 , n60331 , n60332 , n407412 , n60334 , n407414 , n60336 , n60337 , n407417 , n407418 , 
 n60340 , n407420 , n407421 , n60343 , n407423 , n407424 , n407425 , n60347 , n60348 , n407428 , 
 n60350 , n60351 , n407431 , n60353 , n407433 , n60355 , n60356 , n60357 , n60358 , n60359 , 
 n60360 , n407440 , n407441 , n407442 , n60364 , n407444 , n60366 , n60367 , n407447 , n407448 , 
 n60370 , n407450 , n407451 , n60373 , n407453 , n407454 , n60376 , n407456 , n60378 , n60379 , 
 n407459 , n407460 , n60382 , n407462 , n407463 , n60385 , n407465 , n60387 , n60388 , n407468 , 
 n60390 , n407470 , n60392 , n60393 , n407473 , n407474 , n60396 , n407476 , n407477 , n60399 , 
 n407479 , n60401 , n60402 , n60403 , n60404 , n60405 , n60406 , n60407 , n60408 , n407488 , 
 n60410 , n407490 , n60412 , n60413 , n407493 , n407494 , n60416 , n407496 , n407497 , n60419 , 
 n407499 , n60421 , n60422 , n407502 , n407503 , n60425 , n407505 , n60427 , n60428 , n60429 , 
 n60430 , n60431 , n407511 , n60433 , n60434 , n60435 , n60436 , n60437 , n60438 , n60439 , 
 n60440 , n60441 , n60442 , n60443 , n407523 , n60445 , n60446 , n60447 , n407527 , n407528 , 
 n60450 , n407530 , n60452 , n407532 , n407533 , n60455 , n407535 , n60457 , n60458 , n407538 , 
 n60460 , n407540 , n60462 , n60463 , n407543 , n407544 , n60466 , n407546 , n407547 , n60469 , 
 n407549 , n407550 , n407551 , n60473 , n407553 , n407554 , n60476 , n407556 , n407557 , n60479 , 
 n60480 , n60481 , n60482 , n60483 , n407563 , n60485 , n407565 , n60487 , n60488 , n407568 , 
 n407569 , n60491 , n407571 , n407572 , n60494 , n407574 , n407575 , n60497 , n407577 , n60499 , 
 n60500 , n60501 , n60502 , n60503 , n60504 , n60505 , n407585 , n60507 , n60508 , n407588 , 
 n407589 , n60511 , n407591 , n407592 , n60514 , n407594 , n407595 , n60517 , n60518 , n407598 , 
 n60520 , n407600 , n407601 , n60523 , n407603 , n60525 , n407605 , n407606 , n60528 , n60529 , 
 n407609 , n60531 , n407611 , n60533 , n60534 , n407614 , n407615 , n60537 , n407617 , n407618 , 
 n60540 , n407620 , n407621 , n60543 , n407623 , n60545 , n60546 , n407626 , n407627 , n60549 , 
 n407629 , n407630 , n60552 , n407632 , n407633 , n60555 , n407635 , n60557 , n60558 , n407638 , 
 n407639 , n60561 , n407641 , n407642 , n60564 , n407644 , n60566 , n407646 , n60568 , n407648 , 
 n60570 , n60571 , n407651 , n60573 , n407653 , n60575 , n60576 , n407656 , n407657 , n60579 , 
 n407659 , n407660 , n60582 , n407662 , n407663 , n407664 , n60586 , n407666 , n407667 , n60589 , 
 n407669 , n60591 , n407671 , n407672 , n407673 , n60595 , n407675 , n407676 , n60598 , n407678 , 
 n407679 , n60601 , n407681 , n407682 , n60604 , n407684 , n407685 , n60607 , n60608 , n60609 , 
 n407689 , n60611 , n407691 , n407692 , n60617 , n60618 , n60619 , n60620 , n60621 , n60622 , 
 n60623 , n60624 , n60625 , n60626 , n60627 , n60628 , n60629 , n60630 , n60631 , n60632 , 
 n407709 , n60634 , n407711 , n60636 , n60637 , n60638 , n60639 , n60640 , n407717 , n407718 , 
 n407719 , n60644 , n407721 , n407722 , n60647 , n407724 , n60649 , n407726 , n407727 , n60652 , 
 n60653 , n407730 , n60655 , n407732 , n407733 , n407734 , n60659 , n407736 , n407737 , n60662 , 
 n407739 , n60664 , n60665 , n60666 , n60667 , n60668 , n407745 , n60670 , n60671 , n60672 , 
 n60673 , n60674 , n407751 , n407752 , n407753 , n60678 , n407755 , n60680 , n407757 , n60682 , 
 n407759 , n407760 , n60685 , n407762 , n60687 , n60688 , n407765 , n407766 , n407767 , n60692 , 
 n407769 , n60694 , n407771 , n60696 , n60697 , n407774 , n60699 , n407776 , n60701 , n407778 , 
 n407779 , n60704 , n407781 , n407782 , n60707 , n60708 , n407785 , n407786 , n60711 , n407788 , 
 n407789 , n60714 , n407791 , n407792 , n60717 , n407794 , n60719 , n407796 , n60721 , n60722 , 
 n407799 , n60724 , n407801 , n60726 , n60727 , n407804 , n407805 , n60730 , n407807 , n407808 , 
 n60733 , n407810 , n407811 , n407812 , n60737 , n407814 , n407815 , n60740 , n407817 , n407818 , 
 n60743 , n60744 , n60745 , n60746 , n407823 , n60748 , n407825 , n60750 , n60751 , n407828 , 
 n407829 , n60754 , n407831 , n407832 , n60757 , n407834 , n407835 , n60760 , n407837 , n60762 , 
 n407839 , n60764 , n60765 , n407842 , n407843 , n60768 , n407845 , n407846 , n60771 , n407848 , 
 n407849 , n60774 , n407851 , n60776 , n60777 , n407854 , n407855 , n60780 , n407857 , n407858 , 
 n60783 , n407860 , n407861 , n407862 , n60787 , n407864 , n60789 , n60790 , n407867 , n407868 , 
 n60793 , n407870 , n407871 , n60796 , n407873 , n407874 , n60799 , n407876 , n60801 , n60802 , 
 n407879 , n407880 , n60805 , n407882 , n407883 , n60808 , n407885 , n407886 , n60811 , n407888 , 
 n60813 , n407890 , n60815 , n60816 , n407893 , n60818 , n407895 , n60820 , n60821 , n407898 , 
 n407899 , n60824 , n407901 , n407902 , n60827 , n407904 , n407905 , n407906 , n60831 , n407908 , 
 n407909 , n60834 , n407911 , n407912 , n60837 , n60838 , n407915 , n407916 , n60841 , n60842 , 
 n60843 , n407920 , n60845 , n407922 , n60847 , n60848 , n60849 , n407926 , n60851 , n407928 , 
 n60853 , n60854 , n407931 , n60856 , n60857 , n407934 , n60859 , n407936 , n60861 , n407938 , 
 n60863 , n407940 , n60865 , n60866 , n407943 , n407944 , n60869 , n407946 , n60871 , n60872 , 
 n60873 , n407950 , n60875 , n407952 , n60877 , n60878 , n60879 , n60880 , n60881 , n60882 , 
 n60883 , n60884 , n407961 , n60886 , n407963 , n60888 , n60889 , n60890 , n60891 , n60892 , 
 n60893 , n60894 , n60895 , n407972 , n60897 , n407974 , n407975 , n60900 , n407977 , n407978 , 
 n60903 , n60904 , n407981 , n407982 , n60907 , n60908 , n407985 , n60910 , n60911 , n407988 , 
 n60913 , n60914 , n60915 , n60916 , n60917 , n407994 , n60919 , n60920 , n60921 , n407998 , 
 n407999 , n60924 , n60925 , n60926 , n408003 , n408004 , n60929 , n60930 , n60931 , n408008 , 
 n60933 , n60934 , n60935 , n60936 , n60937 , n60940 , n408015 , n408016 , n60943 , n408018 , 
 n60945 , n60946 , n60947 , n408022 , n408023 , n60950 , n408025 , n60952 , n408027 , n60954 , 
 n60955 , n408030 , n408031 , n60958 , n408033 , n408034 , n60961 , n408036 , n408037 , n60964 , 
 n408039 , n60966 , n408041 , n408042 , n60969 , n408044 , n408045 , n408046 , n408047 , n408048 , 
 n408049 , n408050 , n61007 , n61008 , n408053 , n61010 , n61011 , n61012 , n61013 , n408058 , 
 n61015 , n61016 , n61017 , n61018 , n61019 , n61020 , n61021 , n61022 , n61023 , n61024 , 
 n61025 , n61026 , n61027 , n61028 , n61029 , n61030 , n61031 , n61032 , n61033 , n61034 , 
 n61035 , n61036 , n408081 , n61038 , n408083 , n61040 , n61041 , n61042 , n61043 , n408088 , 
 n61045 , n61046 , n61047 , n408092 , n61049 , n61050 , n61051 , n408096 , n61053 , n61054 , 
 n408099 , n61056 , n61057 , n408102 , n61059 , n61060 , n61061 , n61062 , n61065 , n61066 , 
 n61067 , n61068 , n61069 , n61070 , n408113 , n61072 , n408115 , n61074 , n61075 , n408118 , 
 n408119 , n61078 , n408121 , n408122 , n61081 , n408124 , n408125 , n408126 , n61085 , n408128 , 
 n408129 , n61088 , n61089 , n408132 , n61091 , n61092 , n408135 , n61094 , n61095 , n61096 , 
 n61097 , n61098 , n61099 , n61100 , n61101 , n61102 , n408145 , n61104 , n408147 , n61106 , 
 n408149 , n61108 , n408151 , n61110 , n408153 , n61112 , n408155 , n61114 , n61115 , n408158 , 
 n408159 , n61118 , n408161 , n408162 , n61121 , n408164 , n408165 , n61124 , n408167 , n61126 , 
 n61127 , n408170 , n408171 , n61130 , n408173 , n408174 , n61133 , n408176 , n408177 , n61136 , 
 n408179 , n408180 , n61139 , n61140 , n61141 , n61142 , n408185 , n408186 , n61145 , n408188 , 
 n408189 , n408190 , n61149 , n408192 , n408193 , n408194 , n61153 , n408196 , n408197 , n61156 , 
 n408199 , n408200 , n408201 , n61160 , n408203 , n61162 , n408205 , n61164 , n61165 , n408208 , 
 n408209 , n61168 , n408211 , n408212 , n61171 , n408214 , n408215 , n61174 , n61175 , n408218 , 
 n408219 , n61178 , n408221 , n408222 , n61181 , n408224 , n408225 , n61184 , n61185 , n61186 , 
 n408229 , n408230 , n408231 , n61190 , n408233 , n408234 , n61193 , n408236 , n408237 , n61196 , 
 n61197 , n408240 , n61199 , n61200 , n408243 , n408244 , n61203 , n61204 , n408247 , n61206 , 
 n408249 , n61208 , n408251 , n408252 , n61211 , n408254 , n408255 , n61214 , n408257 , n61216 , 
 n61217 , n61218 , n408261 , n61220 , n408263 , n61222 , n61223 , n408266 , n408267 , n61226 , 
 n408269 , n61228 , n61229 , n61230 , n61231 , n61232 , n61233 , n61234 , n61235 , n61236 , 
 n61237 , n61238 , n61239 , n61240 , n61241 , n61242 , n61243 , n61244 , n61245 , n61246 , 
 n61247 , n61248 , n61249 , n61250 , n61251 , n408294 , n61253 , n408296 , n61255 , n408298 , 
 n61257 , n61258 , n408301 , n408302 , n61261 , n408304 , n408305 , n61264 , n408307 , n408308 , 
 n61267 , n408310 , n61269 , n61270 , n408313 , n408314 , n61273 , n408316 , n408317 , n61276 , 
 n408319 , n408320 , n61279 , n61280 , n61281 , n408324 , n408325 , n61284 , n61285 , n61286 , 
 n408329 , n408330 , n61289 , n61290 , n408333 , n408334 , n61293 , n408336 , n61295 , n408338 , 
 n61297 , n61298 , n61299 , n408342 , n61301 , n408344 , n408345 , n61304 , n408347 , n408348 , 
 n61307 , n408350 , n61309 , n61310 , n408353 , n408354 , n61313 , n408356 , n408357 , n61316 , 
 n408359 , n408360 , n408361 , n61320 , n408363 , n408364 , n61323 , n408366 , n61325 , n61326 , 
 n408369 , n61328 , n408371 , n61330 , n408373 , n61332 , n61333 , n408376 , n61335 , n408378 , 
 n61337 , n61338 , n61339 , n408382 , n61341 , n408384 , n408385 , n408386 , n61345 , n408388 , 
 n408389 , n61348 , n408391 , n408392 , n408393 , n61352 , n408395 , n61354 , n61355 , n408398 , 
 n408399 , n61358 , n408401 , n408402 , n61361 , n408404 , n408405 , n61364 , n408407 , n61366 , 
 n61367 , n408410 , n408411 , n61370 , n408413 , n408414 , n61373 , n408416 , n408417 , n61376 , 
 n408419 , n61378 , n408421 , n61380 , n61381 , n408424 , n408425 , n61384 , n408427 , n408428 , 
 n61387 , n408430 , n408431 , n408432 , n61391 , n408434 , n61393 , n61394 , n408437 , n408438 , 
 n61397 , n408440 , n408441 , n61400 , n408443 , n408444 , n61403 , n408446 , n61405 , n61406 , 
 n408449 , n408450 , n61409 , n408452 , n408453 , n61412 , n408455 , n408456 , n61415 , n61416 , 
 n61417 , n408460 , n408461 , n61420 , n61421 , n61422 , n408465 , n408466 , n61425 , n61426 , 
 n61427 , n61428 , n61429 , n61430 , n61431 , n408474 , n408475 , n61434 , n408477 , n61436 , 
 n408479 , n61438 , n408481 , n408482 , n61441 , n408484 , n408485 , n61444 , n61445 , n61446 , 
 n408489 , n408490 , n61449 , n61450 , n61451 , n408494 , n61453 , n61454 , n61455 , n408498 , 
 n61457 , n61458 , n61459 , n408502 , n408503 , n408504 , n61463 , n408506 , n61465 , n61466 , 
 n61467 , n61468 , n61469 , n408512 , n61471 , n408514 , n61473 , n61474 , n61475 , n61476 , 
 n408519 , n61478 , n408521 , n61480 , n408523 , n61482 , n408525 , n408526 , n61485 , n408528 , 
 n408529 , n61488 , n61489 , n61490 , n408533 , n408534 , n61493 , n61494 , n61495 , n408538 , 
 n408539 , n408540 , n408541 , n61500 , n408543 , n61502 , n61503 , n408546 , n408547 , n61506 , 
 n408549 , n61508 , n61509 , n61510 , n61511 , n61512 , n61513 , n61514 , n61515 , n61516 , 
 n61517 , n61518 , n61519 , n61520 , n61521 , n61522 , n408565 , n61524 , n408567 , n61526 , 
 n408569 , n408570 , n61529 , n61530 , n408573 , n61532 , n408575 , n408576 , n61535 , n61536 , 
 n408579 , n408580 , n408581 , n61540 , n61541 , n408584 , n61543 , n408586 , n408587 , n61546 , 
 n61547 , n408590 , n61549 , n61550 , n408593 , n61552 , n408595 , n61554 , n61555 , n61556 , 
 n61557 , n61558 , n408601 , n61560 , n408603 , n408604 , n61563 , n61564 , n61565 , n408608 , 
 n61567 , n408610 , n408611 , n61570 , n408613 , n61572 , n408615 , n408616 , n61575 , n408618 , 
 n61577 , n408620 , n61579 , n61580 , n61581 , n61582 , n61583 , n408626 , n408627 , n61586 , 
 n408629 , n408630 , n61589 , n408632 , n408633 , n61592 , n408635 , n408636 , n61595 , n408638 , 
 n61597 , n61598 , n61599 , n61600 , n61601 , n408644 , n61603 , n61604 , n408647 , n61606 , 
 n408649 , n408650 , n61609 , n408652 , n61611 , n61612 , n408655 , n408656 , n61615 , n408658 , 
 n408659 , n61618 , n408661 , n408662 , n408663 , n61622 , n408665 , n408666 , n61625 , n408668 , 
 n408669 , n61628 , n61629 , n408672 , n61631 , n408674 , n408675 , n61634 , n408677 , n61636 , 
 n61637 , n408680 , n61639 , n408682 , n61641 , n61642 , n408685 , n408686 , n61645 , n408688 , 
 n408689 , n61648 , n408691 , n408692 , n61651 , n408694 , n61653 , n61654 , n408697 , n408698 , 
 n61657 , n408700 , n408701 , n61660 , n408703 , n408704 , n408705 , n61664 , n408707 , n61666 , 
 n408709 , n61668 , n61669 , n61670 , n61671 , n61672 , n61673 , n408716 , n61675 , n408718 , 
 n408719 , n61678 , n61679 , n408722 , n61681 , n408724 , n61683 , n61684 , n408727 , n408728 , 
 n61687 , n408730 , n408731 , n61690 , n408733 , n408734 , n408735 , n61694 , n408737 , n408738 , 
 n61697 , n408740 , n408741 , n61700 , n408743 , n61702 , n408745 , n61704 , n61705 , n408748 , 
 n408749 , n61708 , n408751 , n408752 , n61711 , n408754 , n408755 , n61714 , n408757 , n61716 , 
 n61717 , n408760 , n408761 , n61720 , n408763 , n408764 , n61723 , n408766 , n408767 , n61726 , 
 n61727 , n61728 , n408771 , n408772 , n61731 , n408774 , n408775 , n61734 , n408777 , n408778 , 
 n61737 , n61738 , n408781 , n408782 , n61741 , n61742 , n61743 , n408786 , n408787 , n61746 , 
 n61747 , n61748 , n408791 , n408792 , n61751 , n408794 , n408795 , n61754 , n408797 , n61756 , 
 n61757 , n408800 , n61759 , n408802 , n61761 , n408804 , n61763 , n61764 , n61765 , n61767 , 
 n61768 , n61769 , n61770 , n61771 , n61773 , n61774 , n61775 , n61776 , n61777 , n61778 , 
 n61779 , n61780 , n61781 , n61782 , n61783 , n61784 , n61785 , n61786 , n61787 , n61788 , 
 n61789 , n61790 , n61791 , n61792 , n61793 , n61794 , n61795 , n61796 , n61797 , n61798 , 
 n61799 , n61800 , n61801 , n61802 , n61803 , n61804 , n408845 , n61806 , n61807 , n61808 , 
 n61809 , n408850 , n408851 , n61829 , n408853 , n61831 , n408855 , n408856 , n61834 , n61835 , 
 n61836 , n61837 , n408861 , n61839 , n408863 , n61841 , n61842 , n408866 , n408867 , n61845 , 
 n61846 , n408870 , n408871 , n61849 , n61850 , n61851 , n408875 , n408876 , n61854 , n61855 , 
 n408879 , n61857 , n61858 , n408882 , n61860 , n61861 , n61862 , n61863 , n61864 , n408888 , 
 n61866 , n408890 , n408891 , n61869 , n61870 , n408894 , n61872 , n61873 , n408897 , n408898 , 
 n61876 , n61877 , n408901 , n408902 , n61880 , n61881 , n408905 , n61883 , n61884 , n408908 , 
 n408909 , n408910 , n61888 , n408912 , n408913 , n61891 , n408915 , n61893 , n61894 , n61895 , 
 n61896 , n61897 , n408921 , n408922 , n61900 , n408924 , n61902 , n408926 , n408927 , n61905 , 
 n408929 , n408930 , n61908 , n408932 , n408933 , n61911 , n408935 , n408936 , n408937 , n61915 , 
 n408939 , n61917 , n408941 , n408942 , n61920 , n408944 , n408945 , n61923 , n408947 , n408948 , 
 n408949 , n61929 , n408951 , n408952 , n408953 , n408954 , n61934 , n408956 , n61936 , n408958 , 
 n408959 , n61939 , n408961 , n61941 , n61942 , n61943 , n61944 , n61945 , n61946 , n61947 , 
 n61948 , n61949 , n61950 , n61951 , n61952 , n61953 , n61954 , n61955 , n61956 , n61957 , 
 n61958 , n61959 , n61960 , n61961 , n408983 , n61963 , n408985 , n61965 , n61966 , n61967 , 
 n61968 , n408990 , n408991 , n408992 , n408993 , n61996 , n408995 , n408996 , n61999 , n408998 , 
 n62001 , n409000 , n62003 , n62004 , n409003 , n62006 , n409005 , n62008 , n409007 , n409008 , 
 n62011 , n409010 , n409011 , n62014 , n409013 , n62016 , n409015 , n409016 , n62019 , n409018 , 
 n409019 , n62022 , n409021 , n62024 , n409023 , n62026 , n62027 , n409026 , n409027 , n62030 , 
 n409029 , n409030 , n62033 , n409032 , n409033 , n62036 , n409035 , n62038 , n62039 , n409038 , 
 n409039 , n62042 , n409041 , n409042 , n62045 , n409044 , n409045 , n62048 , n409047 , n409048 , 
 n62051 , n62052 , n409051 , n62054 , n409053 , n62056 , n62057 , n62058 , n62059 , n62060 , 
 n62061 , n409060 , n409061 , n62064 , n409063 , n409064 , n62067 , n409066 , n409067 , n62070 , 
 n62071 , n62072 , n62073 , n409072 , n62075 , n409074 , n62077 , n409076 , n62079 , n62080 , 
 n62081 , n409080 , n62083 , n409082 , n409083 , n409084 , n62087 , n409086 , n62089 , n62090 , 
 n409089 , n409090 , n62093 , n409092 , n409093 , n62096 , n409095 , n409096 , n62099 , n409098 , 
 n409099 , n62102 , n409101 , n62104 , n409103 , n62106 , n409105 , n409106 , n62109 , n409108 , 
 n62111 , n409110 , n409111 , n409112 , n409113 , n62116 , n409115 , n409116 , n62119 , n62120 , 
 n409119 , n409120 , n409121 , n62124 , n409123 , n409124 , n62127 , n62128 , n409127 , n409128 , 
 n62131 , n62132 , n62133 , n62134 , n62135 , n62136 , n62137 , n62138 , n62139 , n409138 , 
 n62141 , n409140 , n409141 , n409142 , n62145 , n409144 , n62147 , n409146 , n409147 , n409148 , 
 n62151 , n62152 , n409151 , n409152 , n62155 , n409154 , n62157 , n409156 , n62159 , n62160 , 
 n62161 , n62162 , n409161 , n62164 , n409163 , n409164 , n62167 , n62168 , n409167 , n62170 , 
 n62171 , n409170 , n409171 , n62174 , n409173 , n409174 , n62177 , n409176 , n62179 , n409178 , 
 n409179 , n62182 , n409181 , n409182 , n409183 , n62186 , n409185 , n409186 , n409187 , n62190 , 
 n409189 , n409190 , n62193 , n409192 , n409193 , n62196 , n409195 , n409196 , n62199 , n409198 , 
 n409199 , n62202 , n62203 , n409202 , n409203 , n409204 , n62207 , n409206 , n409207 , n62210 , 
 n62211 , n409210 , n409211 , n62214 , n62215 , n62216 , n409215 , n409216 , n62219 , n62220 , 
 n62221 , n409220 , n62223 , n62224 , n409223 , n62226 , n62227 , n62228 , n62229 , n62230 , 
 n62231 , n62232 , n62233 , n62234 , n62235 , n62236 , n409235 , n409236 , n62239 , n409238 , 
 n409239 , n62242 , n62243 , n409242 , n409243 , n409244 , n62247 , n409246 , n409247 , n62250 , 
 n62251 , n409250 , n409251 , n409252 , n409253 , n62256 , n409255 , n409256 , n62259 , n62260 , 
 n409259 , n409260 , n62263 , n409262 , n409263 , n409264 , n62267 , n409266 , n62269 , n409268 , 
 n409269 , n409270 , n62273 , n62274 , n409273 , n409274 , n62277 , n62278 , n409277 , n409278 , 
 n62281 , n409280 , n409281 , n62284 , n62285 , n409284 , n409285 , n62288 , n409287 , n409288 , 
 n62291 , n409290 , n409291 , n62294 , n409293 , n409294 , n62297 , n62298 , n409297 , n409298 , 
 n409299 , n62302 , n409301 , n409302 , n62305 , n62306 , n409305 , n409306 , n62309 , n62310 , 
 n62311 , n409310 , n62313 , n62314 , n62315 , n409314 , n409315 , n62318 , n62319 , n409318 , 
 n62321 , n62322 , n409321 , n409322 , n409323 , n62326 , n409325 , n409326 , n62329 , n62330 , 
 n409329 , n409330 , n409331 , n409332 , n62335 , n409334 , n409335 , n62338 , n62339 , n409338 , 
 n409339 , n409340 , n62343 , n409342 , n409343 , n62346 , n62347 , n409346 , n409347 , n62350 , 
 n62351 , n62352 , n409351 , n409352 , n62355 , n62356 , n62357 , n409356 , n62359 , n409358 , 
 n62361 , n62362 , n62363 , n62364 , n62365 , n62366 , n409365 , n409366 , n62369 , n409368 , 
 n409369 , n62372 , n62373 , n409372 , n409373 , n409374 , n62377 , n409376 , n409377 , n62380 , 
 n62381 , n409380 , n409381 , n409382 , n62385 , n409384 , n409385 , n62388 , n62389 , n409388 , 
 n409389 , n409390 , n62393 , n409392 , n409393 , n62396 , n62397 , n409396 , n62399 , n409398 , 
 n409399 , n62402 , n409401 , n409402 , n62405 , n62406 , n409405 , n409406 , n409407 , n62410 , 
 n409409 , n409410 , n62413 , n62414 , n409413 , n62416 , n62417 , n62418 , n409417 , n409418 , 
 n409419 , n62422 , n409421 , n409422 , n62425 , n62426 , n409425 , n409426 , n409427 , n62430 , 
 n409429 , n409430 , n62433 , n409432 , n62435 , n409434 , n409435 , n409436 , n409437 , n62440 , 
 n409439 , n409440 , n62443 , n62444 , n409443 , n409444 , n409445 , n62448 , n409447 , n409448 , 
 n62451 , n62452 , n409451 , n409452 , n62455 , n62456 , n62457 , n62458 , n62459 , n62460 , 
 n62461 , n62462 , n62463 , n62464 , n62465 , n62466 , n62467 , n409466 , n62469 , n409468 , 
 n409469 , n409470 , n62473 , n409472 , n62475 , n409474 , n409475 , n409476 , n62479 , n62480 , 
 n409479 , n409480 , n409481 , n409482 , n62485 , n409484 , n409485 , n62488 , n62489 , n409488 , 
 n62491 , n62492 , n409491 , n409492 , n62495 , n62496 , n62497 , n409496 , n62499 , n409498 , 
 n409499 , n62502 , n409501 , n409502 , n62505 , n409504 , n409505 , n62508 , n409507 , n409508 , 
 n62511 , n409510 , n62513 , n409512 , n409513 , n409514 , n62517 , n409516 , n409517 , n409518 , 
 n62521 , n409520 , n409521 , n62524 , n409523 , n409524 , n62527 , n409526 , n409527 , n62530 , 
 n409529 , n409530 , n62533 , n62534 , n409533 , n409534 , n409535 , n62538 , n409537 , n409538 , 
 n62541 , n62542 , n409541 , n409542 , n62545 , n62546 , n62547 , n409546 , n409547 , n62550 , 
 n62551 , n62552 , n409551 , n409552 , n62555 , n62556 , n62557 , n409556 , n409557 , n62560 , 
 n62561 , n62562 , n409561 , n62564 , n62565 , n409564 , n62567 , n62568 , n62569 , n62570 , 
 n62571 , n62572 , n62573 , n62574 , n62575 , n62576 , n62577 , n62578 , n62579 , n62580 , 
 n62581 , n62582 , n62583 , n62584 , n409583 , n62586 , n409585 , n409586 , n409587 , n409588 , 
 n62591 , n409590 , n409591 , n62594 , n409593 , n409594 , n62597 , n62598 , n62599 , n409598 , 
 n62601 , n62602 , n62603 , n409602 , n409603 , n62606 , n409605 , n409606 , n409607 , n409608 , 
 n62611 , n409610 , n409611 , n62614 , n409613 , n409614 , n62617 , n409616 , n409617 , n409618 , 
 n62621 , n409620 , n62623 , n409622 , n62625 , n62626 , n409625 , n409626 , n62629 , n409628 , 
 n409629 , n62632 , n409631 , n409632 , n62635 , n62636 , n409635 , n409636 , n62639 , n409638 , 
 n409639 , n62642 , n409641 , n409642 , n62645 , n409644 , n409645 , n62648 , n409647 , n62650 , 
 n409649 , n62652 , n62653 , n409652 , n409653 , n62656 , n409655 , n409656 , n62659 , n409658 , 
 n409659 , n62662 , n409661 , n62664 , n409663 , n409664 , n62667 , n409666 , n409667 , n62670 , 
 n409669 , n62672 , n409671 , n62674 , n409673 , n62676 , n62677 , n409676 , n409677 , n62680 , 
 n62681 , n409680 , n409681 , n62684 , n62685 , n409684 , n409685 , n62688 , n409687 , n409688 , 
 n62691 , n409690 , n409691 , n62694 , n62695 , n409694 , n62697 , n409696 , n62699 , n62700 , 
 n409699 , n409700 , n62703 , n409702 , n409703 , n62706 , n409705 , n409706 , n62709 , n409708 , 
 n62711 , n62712 , n409711 , n409712 , n62715 , n409714 , n409715 , n62718 , n409717 , n409718 , 
 n62721 , n409720 , n62723 , n409722 , n62725 , n62726 , n409725 , n409726 , n62729 , n409728 , 
 n409729 , n62732 , n409731 , n409732 , n62735 , n409734 , n62737 , n62738 , n409737 , n409738 , 
 n62741 , n409740 , n409741 , n62744 , n409743 , n409744 , n62747 , n62748 , n409747 , n409748 , 
 n62751 , n409750 , n62753 , n409752 , n62755 , n409754 , n62757 , n62758 , n409757 , n409758 , 
 n62761 , n409760 , n409761 , n62764 , n409763 , n409764 , n62767 , n62768 , n409767 , n409768 , 
 n62771 , n409770 , n409771 , n62774 , n409773 , n409774 , n62777 , n409776 , n409777 , n62780 , 
 n409779 , n409780 , n62783 , n409782 , n409783 , n62786 , n409785 , n62788 , n409787 , n409788 , 
 n62791 , n62792 , n62793 , n409792 , n409793 , n62796 , n62797 , n409796 , n409797 , n62800 , 
 n62801 , n62802 , n409801 , n409802 , n62805 , n62806 , n409805 , n409806 , n62809 , n62810 , 
 n409809 , n62812 , n409811 , n62814 , n409813 , n62816 , n62817 , n409816 , n409817 , n62820 , 
 n409819 , n409820 , n62823 , n409822 , n409823 , n62826 , n409825 , n62828 , n62829 , n409828 , 
 n62831 , n409830 , n62833 , n409832 , n409833 , n62836 , n409835 , n409836 , n62839 , n62840 , 
 n62841 , n409840 , n409841 , n62844 , n62845 , n62846 , n409845 , n409846 , n62849 , n62850 , 
 n62851 , n409850 , n409851 , n62854 , n62855 , n62856 , n409855 , n409856 , n62859 , n409858 , 
 n62861 , n62862 , n62863 , n62864 , n409863 , n62866 , n409865 , n409866 , n62869 , n62870 , 
 n409869 , n62872 , n62873 , n409872 , n62875 , n62876 , n62877 , n62878 , n62879 , n409878 , 
 n62881 , n62882 , n409881 , n409882 , n62885 , n409884 , n62887 , n409886 , n62889 , n62890 , 
 n62891 , n409890 , n62893 , n409892 , n409893 , n62896 , n62897 , n62898 , n409897 , n62900 , 
 n409899 , n62902 , n409901 , n62904 , n62905 , n409904 , n409905 , n62908 , n409907 , n409908 , 
 n62911 , n409910 , n409911 , n409912 , n62915 , n62916 , n409915 , n62918 , n409917 , n409918 , 
 n62921 , n62922 , n409921 , n409922 , n62925 , n62926 , n62927 , n409926 , n409927 , n62930 , 
 n62931 , n62932 , n409931 , n409932 , n62935 , n62936 , n62937 , n62938 , n62939 , n62940 , 
 n62941 , n62942 , n62943 , n62944 , n409943 , n62946 , n409945 , n409946 , n62949 , n409948 , 
 n409949 , n62952 , n62953 , n409952 , n409953 , n62956 , n409955 , n409956 , n62959 , n409958 , 
 n409959 , n62962 , n409961 , n62964 , n62965 , n62966 , n62967 , n62968 , n62969 , n409968 , 
 n62971 , n409970 , n62973 , n62974 , n409973 , n62976 , n62977 , n62978 , n62979 , n409978 , 
 n62981 , n62982 , n62983 , n409982 , n409983 , n62986 , n409985 , n409986 , n62989 , n409988 , 
 n62991 , n62992 , n62993 , n62994 , n409993 , n62996 , n409995 , n62998 , n409997 , n63000 , 
 n409999 , n63002 , n63003 , n410002 , n63005 , n410004 , n410005 , n63008 , n63009 , n63010 , 
 n63011 , n410010 , n410011 , n63014 , n410013 , n410014 , n63017 , n410016 , n63019 , n63020 , 
 n63021 , n410020 , n63023 , n63024 , n410023 , n63026 , n63027 , n63028 , n410027 , n63030 , 
 n63031 , n410030 , n410031 , n63034 , n410033 , n410034 , n63037 , n410036 , n63039 , n410038 , 
 n410039 , n410040 , n63043 , n410042 , n63045 , n410044 , n63047 , n63048 , n410047 , n410048 , 
 n63051 , n410050 , n410051 , n63054 , n410053 , n410054 , n63057 , n63058 , n410057 , n63060 , 
 n410059 , n63062 , n410061 , n410062 , n63065 , n410064 , n410065 , n63068 , n410067 , n63070 , 
 n410069 , n63072 , n63073 , n410072 , n63075 , n410074 , n63077 , n63078 , n410077 , n410078 , 
 n63081 , n410080 , n410081 , n63084 , n410083 , n410084 , n410085 , n63088 , n410087 , n410088 , 
 n63091 , n410090 , n63093 , n410092 , n63095 , n410094 , n63097 , n410096 , n63099 , n410098 , 
 n63101 , n63102 , n410101 , n410102 , n63105 , n63106 , n410105 , n410106 , n63109 , n63110 , 
 n410109 , n410110 , n63113 , n410112 , n410113 , n63116 , n410115 , n410116 , n63119 , n63120 , 
 n410119 , n63122 , n410121 , n63124 , n63125 , n410124 , n410125 , n63128 , n410127 , n410128 , 
 n63131 , n410130 , n410131 , n63134 , n410133 , n410134 , n63137 , n410136 , n63139 , n63140 , 
 n410139 , n410140 , n63143 , n410142 , n410143 , n63146 , n410145 , n410146 , n410147 , n63150 , 
 n410149 , n63152 , n63153 , n63154 , n63155 , n63156 , n63157 , n410156 , n410157 , n63160 , 
 n410159 , n410160 , n63163 , n410162 , n410163 , n63166 , n410165 , n410166 , n63169 , n410168 , 
 n410169 , n63172 , n410171 , n63174 , n63175 , n410174 , n410175 , n63178 , n63179 , n410178 , 
 n410179 , n63182 , n63183 , n63184 , n410183 , n410184 , n410185 , n63188 , n410187 , n63190 , 
 n63191 , n410190 , n63193 , n410192 , n63195 , n63196 , n410195 , n410196 , n63199 , n410198 , 
 n410199 , n63202 , n410201 , n410202 , n410203 , n63206 , n410205 , n410206 , n63209 , n410208 , 
 n410209 , n63212 , n410211 , n63214 , n410213 , n63216 , n63217 , n410216 , n410217 , n63220 , 
 n63221 , n410220 , n410221 , n63224 , n410223 , n410224 , n63227 , n410226 , n63229 , n63230 , 
 n410229 , n410230 , n63233 , n410232 , n410233 , n63236 , n410235 , n410236 , n63239 , n63240 , 
 n63241 , n410240 , n410241 , n63244 , n410243 , n410244 , n410245 , n63248 , n410247 , n63250 , 
 n410249 , n410250 , n63253 , n410252 , n410253 , n63256 , n63257 , n63258 , n410257 , n410258 , 
 n63261 , n410260 , n63263 , n63264 , n63265 , n63266 , n63267 , n410266 , n63269 , n63270 , 
 n410269 , n410270 , n63273 , n63274 , n410273 , n410274 , n410275 , n410276 , n63279 , n63280 , 
 n410279 , n63282 , n63283 , n410282 , n410283 , n63286 , n410285 , n63288 , n63289 , n410288 , 
 n410289 , n63292 , n410291 , n410292 , n63295 , n410294 , n410295 , n63298 , n410297 , n63300 , 
 n410299 , n63302 , n63303 , n410302 , n410303 , n63306 , n410305 , n410306 , n63309 , n410308 , 
 n410309 , n63312 , n410311 , n63314 , n63315 , n410314 , n410315 , n63318 , n410317 , n410318 , 
 n63321 , n410320 , n410321 , n63324 , n63325 , n63326 , n63327 , n410326 , n63329 , n410328 , 
 n63331 , n63332 , n410331 , n410332 , n63335 , n410334 , n410335 , n63338 , n410337 , n63340 , 
 n63341 , n63342 , n410341 , n63344 , n63345 , n63346 , n63347 , n410346 , n63349 , n410348 , 
 n63351 , n63352 , n410351 , n410352 , n63355 , n410354 , n410355 , n63358 , n410357 , n63360 , 
 n63361 , n63362 , n410361 , n63364 , n63365 , n63366 , n63367 , n63368 , n63369 , n410368 , 
 n410369 , n410370 , n63373 , n63374 , n410373 , n63376 , n63377 , n410376 , n410377 , n63380 , 
 n410379 , n63382 , n63383 , n410382 , n410383 , n63386 , n410385 , n410386 , n63389 , n410388 , 
 n410389 , n63392 , n410391 , n63394 , n410393 , n63396 , n63397 , n410396 , n63399 , n410398 , 
 n63401 , n410400 , n410401 , n63404 , n63405 , n410404 , n410405 , n63408 , n410407 , n410408 , 
 n63411 , n410410 , n410411 , n63414 , n410413 , n63416 , n410415 , n63418 , n410417 , n410418 , 
 n63421 , n410420 , n63423 , n410422 , n63425 , n410424 , n63427 , n63428 , n410427 , n410428 , 
 n63431 , n410430 , n410431 , n63434 , n410433 , n410434 , n63437 , n410436 , n63439 , n63440 , 
 n410439 , n410440 , n63443 , n410442 , n410443 , n63446 , n410445 , n410446 , n63449 , n63450 , 
 n63451 , n63452 , n63453 , n410452 , n410453 , n410454 , n63457 , n410456 , n410457 , n63460 , 
 n63461 , n410460 , n410461 , n410462 , n63465 , n410464 , n410465 , n63468 , n63469 , n410468 , 
 n410469 , n410470 , n63473 , n410472 , n410473 , n63476 , n63477 , n410476 , n410477 , n410478 , 
 n63481 , n410480 , n410481 , n63484 , n63485 , n410484 , n63487 , n410486 , n410487 , n63490 , 
 n410489 , n410490 , n63493 , n63494 , n410493 , n410494 , n410495 , n63498 , n410497 , n410498 , 
 n63501 , n63502 , n410501 , n63504 , n63505 , n63506 , n410505 , n410506 , n410507 , n63510 , 
 n410509 , n63512 , n410511 , n410512 , n63515 , n410514 , n410515 , n63518 , n410517 , n410518 , 
 n63521 , n63522 , n410521 , n410522 , n410523 , n63526 , n410525 , n410526 , n63529 , n63530 , 
 n410529 , n410530 , n410531 , n410532 , n63535 , n410534 , n410535 , n63538 , n63539 , n410538 , 
 n410539 , n63542 , n410541 , n410542 , n410543 , n63546 , n410545 , n63548 , n410547 , n410548 , 
 n410549 , n63552 , n63553 , n410552 , n410553 , n63556 , n63557 , n63558 , n63559 , n63560 , 
 n63561 , n63562 , n63563 , n63564 , n410563 , n410564 , n63567 , n63568 , n410567 , n410568 , 
 n63571 , n63572 , n410571 , n410572 , n63575 , n410574 , n410575 , n63578 , n410577 , n410578 , 
 n63581 , n410580 , n410581 , n63584 , n63585 , n410584 , n410585 , n410586 , n63589 , n410588 , 
 n410589 , n63592 , n63593 , n410592 , n410593 , n63596 , n63597 , n63598 , n410597 , n410598 , 
 n63601 , n63602 , n63603 , n410602 , n63605 , n63606 , n410605 , n410606 , n63609 , n63610 , 
 n410609 , n63612 , n63613 , n63614 , n63615 , n63616 , n63617 , n63618 , n63619 , n410618 , 
 n63621 , n63622 , n63623 , n410622 , n63625 , n410624 , n63627 , n410626 , n63629 , n410628 , 
 n63631 , n63632 , n410631 , n410632 , n410633 , n63636 , n410635 , n410636 , n63639 , n410638 , 
 n63641 , n410640 , n410641 , n410642 , n410643 , n63646 , n410645 , n410646 , n63649 , n63650 , 
 n410649 , n410650 , n410651 , n63654 , n410653 , n410654 , n63657 , n63658 , n410657 , n410658 , 
 n63661 , n410660 , n410661 , n63664 , n410663 , n410664 , n63667 , n63668 , n410667 , n410668 , 
 n410669 , n63672 , n410671 , n410672 , n63675 , n63676 , n410675 , n410676 , n63679 , n63680 , 
 n63681 , n410680 , n410681 , n63684 , n63685 , n410684 , n410685 , n63688 , n410687 , n410688 , 
 n63691 , n410690 , n410691 , n63694 , n63695 , n410694 , n410695 , n410696 , n63699 , n410698 , 
 n410699 , n63702 , n63703 , n410702 , n410703 , n63706 , n63707 , n410706 , n410707 , n63710 , 
 n410709 , n410710 , n63713 , n63714 , n410713 , n410714 , n410715 , n63718 , n410717 , n410718 , 
 n410719 , n63722 , n410721 , n410722 , n63725 , n410724 , n410725 , n410726 , n410727 , n63730 , 
 n410729 , n410730 , n63733 , n410732 , n410733 , n63736 , n410735 , n410736 , n63739 , n410738 , 
 n410739 , n63742 , n63743 , n410742 , n63745 , n63746 , n410745 , n410746 , n410747 , n63750 , 
 n410749 , n410750 , n63753 , n63754 , n410753 , n410754 , n63757 , n63758 , n63759 , n410758 , 
 n410759 , n63762 , n63763 , n63764 , n410763 , n63766 , n63767 , n63768 , n63769 , n63770 , 
 n63771 , n63772 , n63773 , n63774 , n63775 , n410774 , n63777 , n63778 , n63779 , n410778 , 
 n410779 , n63782 , n410781 , n410782 , n63785 , n63786 , n410785 , n410786 , n410787 , n63790 , 
 n410789 , n410790 , n63793 , n63794 , n410793 , n410794 , n410795 , n63798 , n410797 , n63800 , 
 n410799 , n63802 , n410801 , n410802 , n63805 , n63806 , n410805 , n63808 , n63809 , n410808 , 
 n410809 , n410810 , n63813 , n410812 , n410813 , n63816 , n63817 , n410816 , n410817 , n410818 , 
 n410819 , n63822 , n410821 , n410822 , n63825 , n63826 , n410825 , n410826 , n410827 , n63830 , 
 n410829 , n410830 , n63833 , n63834 , n410833 , n410834 , n63837 , n410836 , n410837 , n63840 , 
 n410839 , n410840 , n63843 , n63844 , n410843 , n410844 , n410845 , n63848 , n410847 , n410848 , 
 n63851 , n63852 , n410851 , n410852 , n63855 , n63856 , n63857 , n410856 , n63859 , n63860 , 
 n63861 , n63862 , n63863 , n63864 , n63865 , n63866 , n63867 , n63868 , n410867 , n63870 , 
 n63871 , n63872 , n63873 , n63874 , n63875 , n63876 , n63877 , n63878 , n63879 , n63880 , 
 n63881 , n63882 , n63883 , n63884 , n63885 , n63886 , n63887 , n63888 , n63889 , n410888 , 
 n63891 , n410890 , n63893 , n410892 , n63895 , n63896 , n410895 , n410896 , n63899 , n410898 , 
 n410899 , n63902 , n410901 , n410902 , n63905 , n63906 , n410905 , n63908 , n410907 , n410908 , 
 n63911 , n63912 , n410911 , n410912 , n63915 , n410914 , n410915 , n63918 , n410917 , n410918 , 
 n63921 , n63922 , n63923 , n410922 , n410923 , n63926 , n410925 , n410926 , n63929 , n410928 , 
 n63931 , n63932 , n410931 , n410932 , n63935 , n410934 , n63937 , n410936 , n63939 , n410938 , 
 n410939 , n410940 , n63943 , n410942 , n63945 , n410944 , n410945 , n63948 , n410947 , n410948 , 
 n63951 , n410950 , n63953 , n410952 , n63955 , n63956 , n410955 , n410956 , n63959 , n63960 , 
 n410959 , n410960 , n63963 , n410962 , n410963 , n63966 , n410965 , n63968 , n63969 , n410968 , 
 n410969 , n63972 , n410971 , n63974 , n63975 , n410974 , n410975 , n63978 , n410977 , n410978 , 
 n63981 , n410980 , n410981 , n63984 , n410983 , n410984 , n63987 , n410986 , n410987 , n63990 , 
 n63991 , n63992 , n410991 , n410992 , n63995 , n63996 , n63997 , n410996 , n410997 , n64000 , 
 n64001 , n411000 , n64003 , n411002 , n64005 , n64006 , n64007 , n64008 , n411007 , n64010 , 
 n411009 , n411010 , n64013 , n411012 , n64015 , n411014 , n64017 , n64018 , n64019 , n64020 , 
 n411019 , n64022 , n411021 , n64024 , n411023 , n64026 , n64027 , n64028 , n64029 , n411028 , 
 n64031 , n411030 , n64033 , n64034 , n411033 , n411034 , n64037 , n64038 , n411037 , n64040 , 
 n64041 , n64042 , n64043 , n64044 , n411043 , n64046 , n64047 , n64048 , n64049 , n64050 , 
 n64051 , n64052 , n64053 , n64054 , n64055 , n64056 , n64057 , n64058 , n64059 , n64060 , 
 n411059 , n411060 , n64063 , n411062 , n64065 , n411064 , n64067 , n64068 , n411067 , n411068 , 
 n64071 , n64072 , n64073 , n411072 , n411073 , n64076 , n64077 , n64078 , n64079 , n64080 , 
 n64081 , n64082 , n64083 , n64084 , n64085 , n411084 , n64087 , n411086 , n411087 , n64090 , 
 n411089 , n411090 , n64093 , n64094 , n64095 , n411094 , n411095 , n64098 , n411097 , n411098 , 
 n64101 , n411100 , n411101 , n64104 , n64105 , n64106 , n411105 , n411106 , n411107 , n411108 , 
 n64135 , n64136 , n411111 , n64138 , n411113 , n64140 , n64141 , n411116 , n411117 , n64144 , 
 n411119 , n411120 , n64147 , n411122 , n64149 , n64150 , n64151 , n64152 , n64153 , n64154 , 
 n64155 , n64156 , n64157 , n411132 , n64159 , n411134 , n64161 , n411136 , n64163 , n411138 , 
 n64165 , n64166 , n411141 , n411142 , n64169 , n411144 , n411145 , n64172 , n411147 , n411148 , 
 n64175 , n64176 , n411151 , n64178 , n411153 , n64180 , n64181 , n411156 , n411157 , n64184 , 
 n411159 , n411160 , n64187 , n411162 , n411163 , n411164 , n64191 , n411166 , n411167 , n64194 , 
 n411169 , n411170 , n64197 , n64198 , n64199 , n64200 , n64201 , n64202 , n64203 , n64204 , 
 n64205 , n411180 , n64207 , n411182 , n64209 , n64210 , n411185 , n411186 , n64213 , n411188 , 
 n411189 , n64216 , n411191 , n411192 , n411193 , n64220 , n411195 , n64222 , n411197 , n64224 , 
 n411199 , n411200 , n64227 , n411202 , n64229 , n64230 , n411205 , n411206 , n64233 , n411208 , 
 n411209 , n64236 , n411211 , n411212 , n64239 , n411214 , n64241 , n64242 , n411217 , n411218 , 
 n64245 , n411220 , n64247 , n64248 , n411223 , n411224 , n64251 , n411226 , n411227 , n64254 , 
 n411229 , n411230 , n64257 , n411232 , n411233 , n64260 , n411235 , n64262 , n411237 , n64264 , 
 n411239 , n64266 , n64267 , n64268 , n64269 , n64270 , n64271 , n411246 , n64273 , n411248 , 
 n64275 , n411250 , n64277 , n64278 , n411253 , n64280 , n411255 , n64282 , n64283 , n64284 , 
 n64285 , n64286 , n64287 , n64288 , n64289 , n64290 , n64291 , n64292 , n64293 , n64294 , 
 n411269 , n64296 , n411271 , n64298 , n64299 , n411274 , n411275 , n64302 , n64303 , n411278 , 
 n64305 , n64306 , n411281 , n64308 , n64309 , n64310 , n64311 , n64312 , n411287 , n411288 , 
 n64315 , n411290 , n64317 , n411292 , n64319 , n64320 , n64321 , n64322 , n411297 , n64324 , 
 n411299 , n64326 , n411301 , n64328 , n64329 , n64330 , n64331 , n411306 , n411307 , n64334 , 
 n411309 , n64336 , n64337 , n64338 , n411313 , n64340 , n411315 , n64342 , n64343 , n64344 , 
 n411319 , n411320 , n411321 , n64348 , n411323 , n411324 , n411325 , n64352 , n411327 , n411328 , 
 n64355 , n64356 , n411331 , n411332 , n64359 , n411334 , n64361 , n64362 , n64363 , n64364 , 
 n411339 , n64366 , n411341 , n411342 , n64369 , n411344 , n411345 , n411346 , n64373 , n411348 , 
 n64375 , n411350 , n64377 , n411352 , n64379 , n411354 , n64381 , n64382 , n64383 , n64384 , 
 n64385 , n64386 , n411361 , n411362 , n64389 , n411364 , n411365 , n64392 , n411367 , n411368 , 
 n64395 , n64396 , n411371 , n64398 , n411373 , n64400 , n64401 , n64402 , n64403 , n64404 , 
 n64405 , n64406 , n64407 , n64408 , n64409 , n411384 , n64411 , n411386 , n64413 , n411388 , 
 n411389 , n64416 , n64417 , n64418 , n411393 , n411394 , n64421 , n64423 , n411397 , n411398 , 
 n64426 , n411400 , n411401 , n64429 , n411403 , n64431 , n411405 , n411406 , n64434 , n64435 , 
 n64436 , n411410 , n411411 , n64439 , n64440 , n64441 , n64442 , n64443 , n64444 , n64445 , 
 n64446 , n64447 , n411421 , n411422 , n411423 , n64474 , n64475 , n64476 , n64477 , n64478 , 
 n411429 , n64480 , n64481 , n64482 , n411433 , n64484 , n411435 , n64486 , n411437 , n64488 , 
 n64489 , n411440 , n411441 , n64492 , n411443 , n411444 , n64495 , n411446 , n411447 , n64498 , 
 n64499 , n64500 , n411451 , n411452 , n64503 , n411454 , n411455 , n64506 , n411457 , n64508 , 
 n411459 , n64510 , n64511 , n411462 , n411463 , n64514 , n411465 , n411466 , n64517 , n411468 , 
 n64519 , n64520 , n411471 , n411472 , n64523 , n411474 , n64525 , n411476 , n411477 , n64528 , 
 n411479 , n64530 , n411481 , n411482 , n64533 , n411484 , n64535 , n411486 , n64537 , n411488 , 
 n64539 , n64540 , n411491 , n411492 , n64543 , n411494 , n411495 , n64546 , n411497 , n411498 , 
 n64549 , n411500 , n64551 , n411502 , n64553 , n411504 , n411505 , n64556 , n411507 , n64558 , 
 n64559 , n411510 , n411511 , n64562 , n411513 , n411514 , n64565 , n411516 , n411517 , n64568 , 
 n64569 , n411520 , n64571 , n411522 , n64573 , n64574 , n411525 , n411526 , n64577 , n411528 , 
 n411529 , n64580 , n411531 , n411532 , n411533 , n64584 , n411535 , n411536 , n64587 , n411538 , 
 n411539 , n64590 , n411541 , n411542 , n64593 , n411544 , n64595 , n64596 , n64597 , n64598 , 
 n64599 , n64600 , n64601 , n64602 , n64603 , n411554 , n64605 , n64606 , n64607 , n64608 , 
 n411559 , n411560 , n64611 , n411562 , n64613 , n411564 , n411565 , n64616 , n64617 , n64618 , 
 n64619 , n64620 , n64621 , n64622 , n411573 , n64624 , n411575 , n411576 , n64627 , n64628 , 
 n411579 , n64630 , n411581 , n64632 , n64633 , n411584 , n411585 , n64636 , n64637 , n411588 , 
 n411589 , n411590 , n64641 , n64642 , n411593 , n64644 , n64645 , n411596 , n411597 , n64648 , 
 n411599 , n411600 , n64651 , n64652 , n64653 , n411604 , n64655 , n411606 , n64657 , n64658 , 
 n411609 , n411610 , n64661 , n411612 , n411613 , n64664 , n411615 , n411616 , n411617 , n64668 , 
 n411619 , n64670 , n411621 , n64672 , n411623 , n64674 , n411625 , n64676 , n64677 , n411628 , 
 n411629 , n64680 , n411631 , n411632 , n64683 , n411634 , n64685 , n64686 , n64687 , n411638 , 
 n411639 , n64690 , n411641 , n64692 , n411643 , n64694 , n64695 , n411646 , n411647 , n64698 , 
 n411649 , n411650 , n64701 , n411652 , n64703 , n411654 , n64705 , n411656 , n411657 , n64708 , 
 n411659 , n64710 , n64711 , n64712 , n64713 , n64714 , n411665 , n64716 , n64717 , n64718 , 
 n411669 , n64720 , n411671 , n64722 , n64723 , n411674 , n64725 , n411676 , n64727 , n64728 , 
 n411679 , n64730 , n411681 , n64732 , n411683 , n411684 , n64735 , n411686 , n64737 , n411688 , 
 n64739 , n411690 , n411691 , n64742 , n411693 , n411694 , n64745 , n411696 , n411697 , n64748 , 
 n411699 , n411700 , n64751 , n411702 , n64753 , n411704 , n64755 , n411706 , n64757 , n64758 , 
 n411709 , n411710 , n64761 , n411712 , n411713 , n64764 , n411715 , n411716 , n64767 , n64768 , 
 n64769 , n64770 , n64771 , n64772 , n411723 , n64774 , n411725 , n411726 , n64777 , n64778 , 
 n64779 , n64780 , n64781 , n64782 , n64783 , n64784 , n64785 , n64786 , n411737 , n64788 , 
 n64789 , n64790 , n64791 , n411742 , n64793 , n411744 , n64795 , n64796 , n411747 , n411748 , 
 n64799 , n411750 , n411751 , n411752 , n411753 , n411754 , n64805 , n64806 , n64807 , n64808 , 
 n64809 , n64810 , n64811 , n64812 , n411763 , n411764 , n64815 , n411766 , n64817 , n411768 , 
 n64819 , n64820 , n64821 , n411772 , n411773 , n64824 , n64825 , n64826 , n411777 , n64828 , 
 n411779 , n411780 , n411781 , n411782 , n64833 , n411784 , n411785 , n64836 , n411787 , n411788 , 
 n411789 , n64840 , n411791 , n64842 , n64843 , n411794 , n411795 , n64846 , n64847 , n411798 , 
 n64849 , n64850 , n64851 , n64852 , n64853 , n64854 , n64855 , n411806 , n64857 , n411808 , 
 n411809 , n411810 , n64861 , n64862 , n411813 , n64864 , n64865 , n411816 , n411817 , n64868 , 
 n411819 , n411820 , n64871 , n64872 , n411823 , n411824 , n64875 , n64876 , n64877 , n411828 , 
 n411829 , n64880 , n64881 , n411832 , n411833 , n64884 , n411835 , n411836 , n64887 , n411838 , 
 n411839 , n64890 , n411841 , n411842 , n64893 , n411844 , n64895 , n411846 , n411847 , n64898 , 
 n411849 , n64900 , n411851 , n64902 , n64903 , n64904 , n411855 , n411856 , n64907 , n64908 , 
 n64909 , n64910 , n411861 , n411862 , n64948 , n411864 , n64950 , n64951 , n411867 , n411868 , 
 n64954 , n411870 , n411871 , n64957 , n411873 , n64959 , n64960 , n64961 , n64962 , n64963 , 
 n64964 , n64965 , n64966 , n411882 , n64968 , n411884 , n411885 , n64971 , n411887 , n64973 , 
 n411889 , n64975 , n411891 , n411892 , n64978 , n64979 , n411895 , n411896 , n64982 , n411898 , 
 n411899 , n64985 , n411901 , n411902 , n64988 , n411904 , n411905 , n64991 , n64992 , n411908 , 
 n64994 , n411910 , n64996 , n64997 , n64998 , n64999 , n411915 , n411916 , n65002 , n411918 , 
 n411919 , n65005 , n411921 , n65007 , n411923 , n65009 , n411925 , n65011 , n411927 , n65013 , 
 n65014 , n65015 , n65016 , n65022 , n65024 , n411934 , n65026 , n411936 , n65028 , n65029 , 
 n411939 , n65031 , n411941 , n65033 , n65034 , n411944 , n411945 , n65037 , n411947 , n411948 , 
 n65040 , n411950 , n411951 , n411952 , n65044 , n411954 , n411955 , n65047 , n411957 , n411958 , 
 n411959 , n65051 , n411961 , n65053 , n65054 , n411964 , n411965 , n65057 , n411967 , n411968 , 
 n65060 , n411970 , n411971 , n65063 , n411973 , n65065 , n65066 , n411976 , n411977 , n65069 , 
 n411979 , n411980 , n65072 , n411982 , n411983 , n65075 , n411985 , n411986 , n65078 , n411988 , 
 n65080 , n411990 , n411991 , n65083 , n411993 , n411994 , n411995 , n411996 , n65088 , n411998 , 
 n411999 , n65091 , n412001 , n65093 , n65094 , n65095 , n412005 , n65097 , n412007 , n412008 , 
 n65100 , n65101 , n65102 , n412012 , n412013 , n65105 , n65106 , n65107 , n65108 , n65109 , 
 n65110 , n65111 , n412021 , n65113 , n65114 , n412024 , n65116 , n412026 , n65118 , n65119 , 
 n65120 , n65121 , n65122 , n65123 , n412033 , n65125 , n412035 , n412036 , n412037 , n412038 , 
 n65130 , n412040 , n412041 , n65133 , n412043 , n412044 , n65136 , n65137 , n65138 , n412048 , 
 n412049 , n65141 , n412051 , n65167 , n65171 , n412054 , n412055 , n65174 , n65175 , n65176 , 
 n65177 , n65178 , n412061 , n65180 , n412063 , n412064 , n65183 , n65184 , n412067 , n65186 , 
 n65187 , n412070 , n412071 , n65190 , n65191 , n65192 , n412075 , n412076 , n65195 , n412078 , 
 n412079 , n65198 , n65199 , n412082 , n412083 , n65202 , n65203 , n412086 , n412087 , n65206 , 
 n412089 , n412090 , n65209 , n412092 , n65211 , n412094 , n412095 , n412096 , n412097 , n65229 , 
 n412099 , n65231 , n65232 , n412102 , n412103 , n65235 , n412105 , n412106 , n65238 , n412108 , 
 n412109 , n412110 , n65245 , n65246 , n65247 , n412114 , n412115 , n65250 , n412117 , n412118 , 
 n65253 , n412120 , n412121 , n65256 , n412123 , n412124 , n65259 , n65260 , n412127 , n412128 , 
 n65263 , n412130 , n412131 , n65266 , n65267 , n412134 , n412135 , n412136 , n65271 , n412138 , 
 n412139 , n65274 , n65275 , n412142 , n65277 , n65278 , n412145 , n412146 , n65281 , n65282 , 
 n65283 , n412150 , n65285 , n412152 , n65287 , n412154 , n412155 , n65290 , n65291 , n412158 , 
 n65293 , n65294 , n412161 , n65296 , n65297 , n65298 , n65299 , n65300 , n412167 , n65302 , 
 n412169 , n65304 , n65305 , n412172 , n412173 , n65308 , n412175 , n412176 , n65311 , n412178 , 
 n65313 , n65314 , n412181 , n65316 , n412183 , n65318 , n65319 , n412186 , n412187 , n65322 , 
 n412189 , n412190 , n65325 , n412192 , n412193 , n412194 , n65329 , n412196 , n412197 , n65332 , 
 n412199 , n412200 , n65335 , n412202 , n65337 , n65338 , n65339 , n65340 , n65341 , n65342 , 
 n65343 , n65344 , n65345 , n65346 , n412213 , n412214 , n65349 , n412216 , n65351 , n65352 , 
 n65353 , n65354 , n412221 , n65356 , n65357 , n412224 , n412225 , n412226 , n412227 , n65382 , 
 n65383 , n412230 , n412231 , n65386 , n65387 , n65388 , n412235 , n412236 , n65391 , n65392 , 
 n65393 , n412240 , n412241 , n65396 , n412243 , n65398 , n412245 , n412246 , n65401 , n65402 , 
 n412249 , n65404 , n65405 , n412252 , n412253 , n65408 , n65409 , n412256 , n412257 , n65412 , 
 n65413 , n412260 , n412261 , n65416 , n65417 , n65418 , n412265 , n65420 , n412267 , n65435 , 
 n65436 , n412270 , n412271 , n65439 , n412273 , n65441 , n65442 , n412276 , n65448 , n65449 , 
 n65450 , n65451 , n65452 , n65453 , n65454 , n65455 , n65456 , n65457 , n65458 , n65459 , 
 n65460 , n65461 , n65462 , n65463 , n65464 , n65465 , n65466 , n65467 , n65468 , n65469 , 
 n65470 , n65471 , n412301 , n65473 , n412303 , n65475 , n65476 , n65477 , n65478 , n65479 , 
 n65480 , n65481 , n412311 , n65483 , n65484 , n65485 , n412315 , n412316 , n65488 , n412318 , 
 n412319 , n65491 , n65492 , n65493 , n412323 , n412324 , n65496 , n412326 , n412327 , n65499 , 
 n412329 , n65501 , n412331 , n412332 , n65504 , n412334 , n65506 , n65507 , n65508 , n65510 , 
 n412339 , n65512 , n65513 , n65514 , n65515 , n65516 , n412345 , n412346 , n65522 , n412348 , 
 n65524 , n65525 , n412351 , n65527 , n412353 , n412354 , n65530 , n412356 , n65532 , n65533 , 
 n65534 , n65535 , n65536 , n65537 , n65538 , n412364 , n65540 , n65541 , n65542 , n65543 , 
 n65544 , n412370 , n65546 , n65547 , n412373 , n412374 , n65550 , n412376 , n65552 , n412378 , 
 n412379 , n65555 , n412381 , n65557 , n65558 , n412384 , n412385 , n65561 , n412387 , n65563 , 
 n65564 , n65565 , n65566 , n65567 , n412393 , n65569 , n65570 , n65571 , n65572 , n412398 , 
 n65574 , n412400 , n65576 , n65577 , n65578 , n412404 , n65580 , n65581 , n65582 , n65583 , 
 n65584 , n65585 , n412411 , n412412 , n65588 , n65589 , n65590 , n65591 , n412417 , n65593 , 
 n65594 , n65595 , n412421 , n65597 , n65598 , n65599 , n65600 , n65601 , n65602 , n65603 , 
 n65604 , n65605 , n412431 , n65607 , n65608 , n412434 , n65610 , n412436 , n412437 , n65613 , 
 n65614 , n412440 , n412441 , n65617 , n412443 , n65619 , n65620 , n412446 , n65622 , n412448 , 
 n412449 , n65625 , n65626 , n412452 , n65628 , n412454 , n65630 , n65631 , n412457 , n412458 , 
 n65634 , n412460 , n65636 , n412462 , n65638 , n65639 , n412465 , n412466 , n412467 , n65643 , 
 n412469 , n65645 , n65646 , n412472 , n412473 , n65649 , n412475 , n65651 , n412477 , n412478 , 
 n65654 , n412480 , n412481 , n65657 , n65658 , n65659 , n412485 , n412486 , n65662 , n412488 , 
 n412489 , n65665 , n412491 , n65667 , n65668 , n65669 , n65670 , n65671 , n412497 , n65673 , 
 n412499 , n65675 , n65676 , n65677 , n65678 , n65679 , n65680 , n65681 , n65682 , n65683 , 
 n412509 , n412510 , n65686 , n412512 , n412513 , n65689 , n65690 , n65691 , n412517 , n65693 , 
 n65694 , n412520 , n412521 , n65697 , n65698 , n65699 , n65700 , n65701 , n412527 , n412528 , 
 n65704 , n412530 , n65706 , n65707 , n412533 , n65709 , n412535 , n65711 , n412537 , n65713 , 
 n412539 , n412540 , n65716 , n65717 , n412543 , n65719 , n412545 , n412546 , n412547 , n65723 , 
 n412549 , n65725 , n412551 , n412552 , n65728 , n412554 , n412555 , n65731 , n65732 , n65733 , 
 n65734 , n65735 , n412561 , n65737 , n65738 , n65739 , n412565 , n65741 , n412567 , n65743 , 
 n65744 , n65745 , n412571 , n65747 , n412573 , n65749 , n65750 , n412576 , n65752 , n412578 , 
 n412579 , n65755 , n412581 , n65757 , n65758 , n65759 , n65760 , n65761 , n412587 , n65763 , 
 n65764 , n65765 , n65766 , n65767 , n65768 , n65769 , n65770 , n65771 , n65772 , n65773 , 
 n65774 , n412600 , n65776 , n65777 , n65778 , n65779 , n412605 , n412606 , n65782 , n65783 , 
 n65784 , n412610 , n65786 , n412612 , n412613 , n65789 , n412615 , n65791 , n65792 , n65793 , 
 n65794 , n412620 , n412621 , n65797 , n412623 , n65799 , n65800 , n65801 , n412627 , n65803 , 
 n65804 , n65805 , n65806 , n65807 , n65808 , n65809 , n65810 , n65811 , n65812 , n65813 , 
 n65814 , n412640 , n412641 , n412642 , n65818 , n412644 , n412645 , n65821 , n65822 , n412648 , 
 n65824 , n412650 , n65826 , n65827 , n412653 , n412654 , n65830 , n412656 , n412657 , n65833 , 
 n412659 , n65835 , n65836 , n65837 , n65838 , n412664 , n65840 , n65841 , n65842 , n412668 , 
 n412669 , n412670 , n65846 , n412672 , n65848 , n65849 , n412675 , n412676 , n65852 , n412678 , 
 n412679 , n65855 , n412681 , n412682 , n65858 , n412684 , n65860 , n65861 , n412687 , n412688 , 
 n65864 , n412690 , n412691 , n65867 , n412693 , n412694 , n412695 , n65871 , n412697 , n65873 , 
 n412699 , n65875 , n65876 , n412702 , n65878 , n412704 , n65880 , n412706 , n412707 , n65883 , 
 n412709 , n412710 , n65886 , n65887 , n412713 , n412714 , n65890 , n412716 , n412717 , n65893 , 
 n412719 , n412720 , n65896 , n412722 , n65898 , n412724 , n65900 , n65901 , n412727 , n412728 , 
 n65904 , n412730 , n412731 , n65907 , n412733 , n412734 , n65910 , n412736 , n65912 , n65913 , 
 n412739 , n412740 , n65916 , n412742 , n412743 , n65919 , n412745 , n412746 , n412747 , n65923 , 
 n412749 , n65925 , n65926 , n412752 , n412753 , n65929 , n412755 , n412756 , n65932 , n412758 , 
 n412759 , n65935 , n412761 , n65937 , n65938 , n65939 , n412765 , n65941 , n412767 , n412768 , 
 n65944 , n412770 , n65946 , n412772 , n412773 , n412774 , n65950 , n412776 , n65952 , n412778 , 
 n65954 , n65955 , n412781 , n412782 , n65958 , n412784 , n412785 , n65961 , n412787 , n412788 , 
 n412789 , n65965 , n412791 , n412792 , n65968 , n412794 , n412795 , n65971 , n65972 , n65973 , 
 n412799 , n412800 , n65976 , n65977 , n65978 , n412804 , n412805 , n65981 , n412807 , n65983 , 
 n412809 , n65985 , n65986 , n412812 , n65988 , n412814 , n65990 , n65991 , n412817 , n412818 , 
 n65994 , n412820 , n412821 , n65997 , n412823 , n412824 , n412825 , n66001 , n412827 , n412828 , 
 n66004 , n412830 , n412831 , n66007 , n66008 , n66009 , n412835 , n66011 , n66012 , n66013 , 
 n66014 , n66015 , n66016 , n66017 , n66018 , n66019 , n66020 , n412846 , n66022 , n412848 , 
 n66024 , n66025 , n412851 , n412852 , n66028 , n412854 , n412855 , n66031 , n412857 , n412858 , 
 n66034 , n412860 , n66036 , n66037 , n412863 , n412864 , n66040 , n412866 , n412867 , n66043 , 
 n412869 , n412870 , n412871 , n412872 , n66048 , n412874 , n66050 , n412876 , n412877 , n66053 , 
 n66054 , n66055 , n412881 , n412882 , n66058 , n66059 , n66060 , n66061 , n66062 , n66063 , 
 n412889 , n412890 , n66066 , n412892 , n66068 , n66069 , n66070 , n66071 , n66072 , n412898 , 
 n66074 , n412900 , n66076 , n66077 , n412903 , n412904 , n66080 , n412906 , n412907 , n66083 , 
 n412909 , n412910 , n66086 , n412912 , n412913 , n66089 , n66090 , n412916 , n66092 , n412918 , 
 n66094 , n412920 , n412921 , n66097 , n66098 , n412924 , n412925 , n66101 , n412927 , n412928 , 
 n66104 , n412930 , n412931 , n66107 , n412933 , n66109 , n412935 , n66111 , n412937 , n66113 , 
 n66114 , n66115 , n412941 , n412942 , n66118 , n412944 , n412945 , n66121 , n66122 , n66123 , 
 n66124 , n66125 , n412951 , n66127 , n66128 , n412954 , n412955 , n66131 , n66132 , n412958 , 
 n66134 , n66135 , n412961 , n412962 , n66138 , n412964 , n412965 , n66141 , n412967 , n412968 , 
 n66144 , n412970 , n412971 , n66147 , n412973 , n412974 , n66150 , n412976 , n412977 , n66153 , 
 n66154 , n412980 , n412981 , n66157 , n412983 , n412984 , n412985 , n412986 , n66162 , n412988 , 
 n412989 , n66165 , n66166 , n412992 , n412993 , n412994 , n66170 , n412996 , n412997 , n66173 , 
 n66174 , n413000 , n413001 , n413002 , n66178 , n413004 , n66180 , n413006 , n66182 , n413008 , 
 n413009 , n66185 , n413011 , n413012 , n66188 , n66189 , n413015 , n413016 , n413017 , n66193 , 
 n413019 , n413020 , n66196 , n66197 , n413023 , n66199 , n66200 , n66201 , n413027 , n66203 , 
 n66204 , n413030 , n413031 , n66207 , n413033 , n413034 , n66210 , n413036 , n413037 , n66213 , 
 n66214 , n413040 , n413041 , n413042 , n66218 , n413044 , n413045 , n66221 , n66222 , n413048 , 
 n413049 , n413050 , n413051 , n66227 , n413053 , n413054 , n66230 , n66231 , n413057 , n413058 , 
 n413059 , n66235 , n413061 , n413062 , n66238 , n66239 , n413065 , n413066 , n66242 , n413068 , 
 n413069 , n66245 , n413071 , n66247 , n413073 , n413074 , n413075 , n66251 , n66252 , n413078 , 
 n413079 , n413080 , n66256 , n413082 , n413083 , n66259 , n66260 , n413086 , n413087 , n66263 , 
 n66264 , n66265 , n66266 , n66267 , n66268 , n66269 , n66270 , n413096 , n66272 , n413098 , 
 n413099 , n413100 , n66276 , n413102 , n66278 , n413104 , n413105 , n413106 , n66282 , n66283 , 
 n413109 , n413110 , n66286 , n413112 , n66288 , n413114 , n413115 , n66291 , n413117 , n413118 , 
 n66294 , n66295 , n413121 , n413122 , n66298 , n413124 , n413125 , n66301 , n66302 , n413128 , 
 n413129 , n66305 , n66306 , n413132 , n413133 , n66309 , n413135 , n66311 , n413137 , n413138 , 
 n66314 , n66315 , n66316 , n413142 , n413143 , n66319 , n66320 , n66321 , n413147 , n66323 , 
 n66324 , n413150 , n66326 , n66327 , n66328 , n66329 , n66330 , n66331 , n66332 , n66333 , 
 n66334 , n66335 , n66336 , n66337 , n66338 , n66339 , n66340 , n66341 , n66342 , n66343 , 
 n66344 , n66345 , n66346 , n66347 , n66348 , n66349 , n66350 , n413176 , n66352 , n66353 , 
 n66354 , n66355 , n66356 , n413182 , n66358 , n66359 , n413185 , n66361 , n413187 , n413188 , 
 n413189 , n66365 , n413191 , n413192 , n66368 , n66369 , n413195 , n413196 , n413197 , n413198 , 
 n66374 , n413200 , n413201 , n66377 , n66378 , n413204 , n413205 , n413206 , n66382 , n413208 , 
 n413209 , n66385 , n66386 , n413212 , n413213 , n66389 , n413215 , n413216 , n413217 , n413218 , 
 n66394 , n413220 , n413221 , n66397 , n66398 , n413224 , n413225 , n413226 , n66402 , n413228 , 
 n413229 , n66405 , n66406 , n413232 , n413233 , n66409 , n413235 , n66411 , n413237 , n66413 , 
 n413239 , n413240 , n66416 , n66417 , n413243 , n413244 , n413245 , n66421 , n413247 , n66423 , 
 n413249 , n413250 , n66426 , n66427 , n66428 , n413254 , n66430 , n413256 , n413257 , n66433 , 
 n413259 , n413260 , n66436 , n66437 , n413263 , n413264 , n413265 , n66441 , n413267 , n413268 , 
 n66444 , n66445 , n413271 , n413272 , n413273 , n413274 , n66450 , n413276 , n413277 , n66453 , 
 n66454 , n413280 , n413281 , n413282 , n66458 , n413284 , n413285 , n66461 , n66462 , n413288 , 
 n413289 , n66465 , n413291 , n66467 , n413293 , n413294 , n66470 , n413296 , n413297 , n66473 , 
 n66474 , n413300 , n413301 , n66477 , n413303 , n413304 , n66480 , n66481 , n413307 , n413308 , 
 n66484 , n66485 , n413311 , n413312 , n66488 , n66489 , n66490 , n413316 , n66492 , n66493 , 
 n66494 , n66495 , n66496 , n66497 , n66498 , n66499 , n66500 , n66501 , n66502 , n66503 , 
 n66504 , n413330 , n413331 , n66507 , n66508 , n413334 , n413335 , n413336 , n66512 , n413338 , 
 n413339 , n66515 , n66516 , n413342 , n413343 , n413344 , n66520 , n413346 , n413347 , n66523 , 
 n66524 , n413350 , n66526 , n413352 , n413353 , n66529 , n413355 , n413356 , n66532 , n66533 , 
 n413359 , n413360 , n413361 , n66537 , n413363 , n413364 , n66540 , n66541 , n413367 , n413368 , 
 n413369 , n66545 , n413371 , n413372 , n66548 , n66549 , n413375 , n413376 , n413377 , n66553 , 
 n413379 , n413380 , n66556 , n66557 , n413383 , n66559 , n66560 , n413386 , n66562 , n66563 , 
 n66564 , n66565 , n66566 , n66567 , n66568 , n66569 , n66570 , n66571 , n66572 , n413398 , 
 n66574 , n66575 , n66576 , n66577 , n66578 , n413404 , n66580 , n66581 , n66582 , n66583 , 
 n66584 , n413410 , n66586 , n66587 , n66588 , n413414 , n66590 , n66591 , n66592 , n66593 , 
 n66594 , n66595 , n66596 , n66597 , n413423 , n66599 , n413425 , n66601 , n413427 , n66603 , 
 n413429 , n413430 , n66606 , n413432 , n413433 , n66609 , n66610 , n66611 , n66612 , n413438 , 
 n413439 , n66615 , n413441 , n66617 , n66618 , n66619 , n66620 , n413446 , n66622 , n413448 , 
 n66624 , n413450 , n66626 , n66627 , n413453 , n413454 , n66630 , n413456 , n413457 , n66633 , 
 n413459 , n413460 , n66636 , n413462 , n66638 , n66639 , n66640 , n66641 , n66642 , n413468 , 
 n66644 , n66645 , n66646 , n413472 , n413473 , n66649 , n413475 , n413476 , n66652 , n66653 , 
 n413479 , n66655 , n413481 , n66657 , n413483 , n413484 , n66660 , n413486 , n413487 , n66663 , 
 n66664 , n413490 , n66666 , n413492 , n66668 , n413494 , n66670 , n66671 , n413497 , n413498 , 
 n66674 , n413500 , n413501 , n66677 , n413503 , n413504 , n66680 , n413506 , n66682 , n66683 , 
 n413509 , n413510 , n66686 , n413512 , n413513 , n66689 , n413515 , n413516 , n66692 , n66693 , 
 n66694 , n413520 , n413521 , n66697 , n66698 , n66699 , n413525 , n66701 , n66702 , n66703 , 
 n413529 , n413530 , n66706 , n413532 , n66708 , n413534 , n66710 , n413536 , n66712 , n413538 , 
 n66714 , n66715 , n413541 , n413542 , n66718 , n66719 , n413545 , n413546 , n413547 , n66723 , 
 n66724 , n413550 , n66726 , n66727 , n413553 , n66729 , n413555 , n413556 , n413557 , n66733 , 
 n413559 , n413560 , n66736 , n413562 , n66738 , n66739 , n66740 , n413566 , n413567 , n66743 , 
 n413569 , n413570 , n66746 , n413572 , n413573 , n66749 , n66750 , n413576 , n66752 , n413578 , 
 n413579 , n66755 , n66756 , n413582 , n413583 , n66759 , n413585 , n413586 , n66762 , n413588 , 
 n66764 , n66765 , n66766 , n66767 , n66768 , n66769 , n66770 , n66771 , n66772 , n413598 , 
 n413599 , n66775 , n413601 , n66777 , n66778 , n66779 , n66780 , n413606 , n66782 , n66783 , 
 n66784 , n413610 , n66786 , n66805 , n66806 , n413614 , n413615 , n413616 , n66810 , n413618 , 
 n66812 , n66813 , n413621 , n413622 , n66816 , n413624 , n413625 , n66819 , n413627 , n413628 , 
 n66822 , n413630 , n66824 , n66825 , n413633 , n413634 , n66828 , n413636 , n413637 , n66831 , 
 n413639 , n413640 , n413641 , n66835 , n413643 , n66837 , n413645 , n66839 , n413647 , n66841 , 
 n66842 , n413650 , n413651 , n66845 , n413653 , n413654 , n66848 , n413656 , n66850 , n66851 , 
 n66852 , n66853 , n66854 , n413662 , n413663 , n66857 , n413665 , n66859 , n66860 , n66861 , 
 n413669 , n66863 , n66864 , n66865 , n413673 , n413674 , n66868 , n66869 , n66870 , n413678 , 
 n413679 , n66873 , n413681 , n66875 , n413683 , n66877 , n413685 , n66879 , n66880 , n413688 , 
 n413689 , n66883 , n413691 , n413692 , n66886 , n413694 , n413695 , n66889 , n66890 , n413698 , 
 n66892 , n413700 , n66894 , n66895 , n413703 , n413704 , n66898 , n413706 , n413707 , n66901 , 
 n413709 , n413710 , n413711 , n66905 , n413713 , n413714 , n66908 , n413716 , n413717 , n66911 , 
 n66912 , n66913 , n413721 , n413722 , n66916 , n413724 , n66918 , n66919 , n66920 , n66921 , 
 n413729 , n66923 , n66925 , n66926 , n66927 , n413734 , n66929 , n413736 , n66931 , n66932 , 
 n413739 , n413740 , n66935 , n413742 , n413743 , n66938 , n413745 , n413746 , n413747 , n66942 , 
 n413749 , n413750 , n66945 , n66946 , n413753 , n66948 , n66949 , n413756 , n413757 , n66952 , 
 n413759 , n66954 , n66955 , n413762 , n413763 , n66958 , n413765 , n66960 , n66961 , n66962 , 
 n66963 , n66964 , n66965 , n413772 , n66967 , n413774 , n413775 , n66970 , n413777 , n66972 , 
 n413779 , n66974 , n413781 , n66976 , n66977 , n413784 , n413785 , n66980 , n66981 , n413788 , 
 n413789 , n66984 , n66985 , n413792 , n413793 , n66988 , n413795 , n413796 , n66991 , n413798 , 
 n413799 , n66994 , n413801 , n413802 , n66997 , n413804 , n66999 , n67000 , n67001 , n67002 , 
 n413809 , n67004 , n67005 , n413812 , n413813 , n67008 , n413815 , n413816 , n67011 , n413818 , 
 n413819 , n67014 , n413821 , n413822 , n67017 , n67018 , n413825 , n67020 , n413827 , n67022 , 
 n67023 , n413830 , n67025 , n413832 , n67027 , n413834 , n413835 , n67030 , n413837 , n67032 , 
 n67033 , n413840 , n413841 , n67036 , n413843 , n413844 , n67039 , n413846 , n413847 , n67042 , 
 n413849 , n67044 , n413851 , n413852 , n67047 , n413854 , n413855 , n67050 , n67051 , n413858 , 
 n67053 , n413860 , n67055 , n413862 , n67057 , n67058 , n413865 , n413866 , n67061 , n413868 , 
 n413869 , n67064 , n413871 , n67066 , n67067 , n67068 , n413875 , n67070 , n413877 , n67072 , 
 n67073 , n413880 , n67075 , n67076 , n67077 , n413884 , n413885 , n67080 , n413887 , n413888 , 
 n67083 , n413890 , n413891 , n67086 , n413893 , n413894 , n67089 , n67090 , n413897 , n67092 , 
 n413899 , n67094 , n413901 , n67096 , n67097 , n413904 , n413905 , n67100 , n413907 , n413908 , 
 n67103 , n413910 , n413911 , n67106 , n67107 , n413914 , n413915 , n67110 , n413917 , n413918 , 
 n67113 , n413920 , n413921 , n67116 , n67117 , n67118 , n67119 , n67120 , n67121 , n413928 , 
 n67123 , n413930 , n67125 , n67126 , n413933 , n413934 , n67129 , n67130 , n413937 , n67132 , 
 n67133 , n413940 , n413941 , n67136 , n67137 , n413944 , n67139 , n413946 , n67141 , n413948 , 
 n413949 , n67144 , n413951 , n413952 , n67147 , n67148 , n67149 , n413956 , n67151 , n413958 , 
 n67153 , n67154 , n413961 , n413962 , n67157 , n413964 , n413965 , n67160 , n413967 , n413968 , 
 n67163 , n413970 , n67165 , n67166 , n67167 , n67168 , n413975 , n67170 , n413977 , n67172 , 
 n413979 , n67174 , n413981 , n67176 , n67177 , n413984 , n413985 , n67180 , n413987 , n413988 , 
 n67183 , n413990 , n413991 , n67186 , n67187 , n413994 , n413995 , n67190 , n413997 , n413998 , 
 n67193 , n414000 , n67195 , n414002 , n67197 , n67198 , n67199 , n67200 , n414007 , n414008 , 
 n67203 , n414010 , n414011 , n67206 , n414013 , n414014 , n414015 , n67210 , n414017 , n67212 , 
 n414019 , n414020 , n67215 , n414022 , n414023 , n67218 , n414025 , n414026 , n414027 , n67222 , 
 n414029 , n67224 , n414031 , n414032 , n67227 , n414034 , n414035 , n67230 , n414037 , n414038 , 
 n67233 , n67234 , n67235 , n414042 , n414043 , n67238 , n67239 , n67240 , n414047 , n414048 , 
 n67243 , n414050 , n414051 , n414052 , n414053 , n67248 , n414055 , n414056 , n67251 , n414058 , 
 n67253 , n67254 , n414061 , n67256 , n414063 , n67258 , n67259 , n414066 , n67261 , n414068 , 
 n414069 , n67264 , n414071 , n67266 , n67267 , n414074 , n67283 , n67284 , n67285 , n67286 , 
 n67287 , n67288 , n67289 , n67290 , n414083 , n67292 , n414085 , n67294 , n67295 , n414088 , 
 n414089 , n67298 , n414091 , n414092 , n67301 , n414094 , n414095 , n414096 , n67305 , n414098 , 
 n67307 , n67308 , n67309 , n67310 , n67311 , n67312 , n67313 , n67314 , n67315 , n414108 , 
 n414109 , n67318 , n414111 , n67320 , n67321 , n67322 , n414115 , n67324 , n414117 , n67326 , 
 n67327 , n67328 , n67329 , n67330 , n414123 , n414124 , n67333 , n414126 , n414127 , n67336 , 
 n67337 , n67338 , n67339 , n67340 , n67341 , n67342 , n67343 , n67344 , n67345 , n67346 , 
 n414139 , n67348 , n414141 , n414142 , n67351 , n67352 , n414145 , n67354 , n414147 , n67356 , 
 n67357 , n67358 , n67359 , n67360 , n67361 , n414154 , n414155 , n67364 , n414157 , n414158 , 
 n67367 , n414160 , n414161 , n67370 , n414163 , n67372 , n67373 , n67374 , n414167 , n67376 , 
 n67377 , n414170 , n67379 , n414172 , n67381 , n67382 , n414175 , n414176 , n67385 , n414178 , 
 n414179 , n67388 , n414181 , n414182 , n67391 , n414184 , n67393 , n67394 , n414187 , n414188 , 
 n67397 , n414190 , n414191 , n67400 , n414193 , n67402 , n67403 , n67404 , n67405 , n67406 , 
 n67407 , n67408 , n414201 , n414202 , n67411 , n414204 , n67413 , n414206 , n414207 , n67416 , 
 n414209 , n67418 , n67419 , n67420 , n67421 , n67422 , n67423 , n67424 , n67425 , n67426 , 
 n414219 , n414220 , n67429 , n414222 , n67431 , n414224 , n414225 , n67434 , n414227 , n414228 , 
 n67437 , n414230 , n414231 , n414232 , n414233 , n67442 , n414235 , n414236 , n67445 , n414238 , 
 n67447 , n67448 , n67449 , n67450 , n67451 , n67452 , n67453 , n67454 , n67455 , n67456 , 
 n67457 , n67458 , n67460 , n414252 , n67462 , n414254 , n67464 , n67465 , n67466 , n67467 , 
 n67468 , n67469 , n67470 , n67471 , n67472 , n67473 , n67474 , n67475 , n67476 , n67477 , 
 n67478 , n67479 , n67480 , n67481 , n67482 , n67483 , n67484 , n67485 , n67486 , n67487 , 
 n67488 , n67489 , n67490 , n414282 , n414283 , n414284 , n414285 , n67495 , n414287 , n67497 , 
 n414289 , n414290 , n67500 , n67501 , n67502 , n414294 , n414295 , n67505 , n67506 , n67507 , 
 n414299 , n414300 , n67535 , n67536 , n67540 , n67541 , n414305 , n414306 , n67563 , n67564 , 
 n414309 , n67566 , n414311 , n67568 , n414313 , n67570 , n414315 , n67572 , n67573 , n414318 , 
 n414319 , n67576 , n414321 , n414322 , n67579 , n414324 , n414325 , n67582 , n67583 , n414328 , 
 n414329 , n67586 , n414331 , n414332 , n67589 , n414334 , n414335 , n67592 , n67594 , n414338 , 
 n67596 , n67597 , n414341 , n67599 , n67600 , n67601 , n414345 , n67603 , n67604 , n67605 , 
 n414349 , n67607 , n67608 , n67609 , n67610 , n67611 , n67612 , n67613 , n67614 , n67615 , 
 n67616 , n67617 , n67618 , n67619 , n67620 , n67621 , n67622 , n67623 , n414367 , n414368 , 
 n67626 , n414370 , n67628 , n67629 , n67630 , n414374 , n414375 , n67633 , n414377 , n67635 , 
 n414379 , n67637 , n67638 , n67639 , n67640 , n414384 , n67642 , n67643 , n414387 , n67645 , 
 n67646 , n67647 , n67648 , n67649 , n67650 , n414394 , n67652 , n67653 , n414397 , n414398 , 
 n67656 , n67657 , n414401 , n414402 , n67660 , n414404 , n67662 , n67663 , n414407 , n67665 , 
 n414409 , n67667 , n414411 , n414412 , n67670 , n414414 , n414415 , n414416 , n67674 , n67675 , 
 n414419 , n67677 , n67678 , n414422 , n414423 , n414424 , n414425 , n67683 , n414427 , n67685 , 
 n414429 , n414430 , n414431 , n414432 , n67690 , n414434 , n67692 , n414436 , n414437 , n67695 , 
 n67696 , n67697 , n414441 , n414442 , n67700 , n67701 , n414445 , n67703 , n414447 , n67724 , 
 n67725 , n67726 , n67727 , n414452 , n414453 , n67730 , n67731 , n414456 , n67733 , n414458 , 
 n67735 , n414460 , n67737 , n67738 , n414463 , n414464 , n67741 , n414466 , n414467 , n67744 , 
 n414469 , n414470 , n67747 , n414472 , n67749 , n67750 , n414475 , n414476 , n67753 , n414478 , 
 n414479 , n67756 , n414481 , n67758 , n414483 , n67760 , n414485 , n67762 , n67763 , n414488 , 
 n414489 , n67766 , n414491 , n414492 , n67769 , n414494 , n414495 , n67772 , n414497 , n67774 , 
 n67775 , n414500 , n414501 , n67778 , n414503 , n414504 , n67781 , n414506 , n414507 , n67784 , 
 n414509 , n67786 , n67787 , n414512 , n414513 , n67790 , n414515 , n414516 , n67793 , n414518 , 
 n67795 , n67796 , n67797 , n414522 , n414523 , n67800 , n414525 , n67802 , n67803 , n414528 , 
 n67805 , n414530 , n67807 , n67808 , n67809 , n414534 , n414535 , n67812 , n414537 , n414538 , 
 n67815 , n414540 , n414541 , n67818 , n414543 , n67820 , n67821 , n67822 , n67823 , n67824 , 
 n67825 , n67826 , n67827 , n67828 , n67829 , n67830 , n67831 , n67832 , n67833 , n67834 , 
 n67835 , n67836 , n67837 , n67838 , n67839 , n67840 , n67841 , n67842 , n414567 , n67844 , 
 n67845 , n414570 , n67847 , n67848 , n414573 , n67850 , n414575 , n414576 , n67853 , n414578 , 
 n67855 , n67856 , n414581 , n414582 , n67859 , n414584 , n67861 , n67862 , n414587 , n67864 , 
 n414589 , n67866 , n67867 , n414592 , n414593 , n67870 , n414595 , n414596 , n67873 , n414598 , 
 n414599 , n67876 , n414601 , n67878 , n67879 , n414604 , n414605 , n67882 , n414607 , n414608 , 
 n67885 , n414610 , n414611 , n67888 , n414613 , n67890 , n67891 , n67892 , n67893 , n67894 , 
 n67895 , n67896 , n414621 , n67898 , n414623 , n67900 , n67901 , n414626 , n67903 , n414628 , 
 n67905 , n414630 , n414631 , n67908 , n414633 , n414634 , n67911 , n414636 , n67913 , n67914 , 
 n67915 , n67916 , n67917 , n67918 , n67919 , n67920 , n67921 , n67922 , n414647 , n414648 , 
 n67925 , n414650 , n67927 , n67928 , n67929 , n67930 , n67931 , n67932 , n67933 , n414658 , 
 n414659 , n67936 , n414661 , n414662 , n67939 , n414664 , n414665 , n67942 , n67943 , n414668 , 
 n414669 , n414670 , n67947 , n414672 , n414673 , n67950 , n67951 , n414676 , n414677 , n414678 , 
 n414679 , n67956 , n67957 , n414682 , n67959 , n67960 , n414685 , n414686 , n67963 , n414688 , 
 n414689 , n414690 , n67967 , n414692 , n414693 , n67970 , n67971 , n414696 , n414697 , n67974 , 
 n67975 , n67976 , n67977 , n67978 , n67979 , n67980 , n67981 , n67982 , n67983 , n67984 , 
 n67985 , n67986 , n67987 , n414712 , n67989 , n414714 , n414715 , n414716 , n67993 , n414718 , 
 n414719 , n67996 , n67997 , n414722 , n414723 , n68000 , n68001 , n68002 , n414727 , n68004 , 
 n414729 , n414730 , n414731 , n68008 , n414733 , n414734 , n68011 , n68012 , n414737 , n414738 , 
 n414739 , n68016 , n414741 , n68018 , n68019 , n414744 , n414745 , n68022 , n68023 , n414748 , 
 n68025 , n68026 , n414751 , n414752 , n414753 , n68030 , n68031 , n414756 , n414757 , n68034 , 
 n414759 , n414760 , n68037 , n68038 , n68039 , n414764 , n414765 , n68042 , n68043 , n68044 , 
 n68045 , n68046 , n68047 , n68048 , n68049 , n68050 , n68051 , n68052 , n68053 , n414778 , 
 n68055 , n68056 , n68057 , n414782 , n414783 , n414784 , n68061 , n414786 , n414787 , n68064 , 
 n414789 , n414790 , n68067 , n414792 , n414793 , n68070 , n68071 , n414796 , n414797 , n414798 , 
 n68075 , n414800 , n414801 , n68078 , n68079 , n414804 , n414805 , n414806 , n414807 , n68084 , 
 n414809 , n414810 , n68087 , n68088 , n414813 , n414814 , n414815 , n68092 , n414817 , n414818 , 
 n68095 , n68096 , n414821 , n414822 , n68099 , n414824 , n414825 , n68102 , n414827 , n414828 , 
 n68105 , n68106 , n414831 , n414832 , n414833 , n68110 , n414835 , n414836 , n68113 , n68114 , 
 n414839 , n414840 , n414841 , n414842 , n68119 , n414844 , n414845 , n68122 , n68123 , n414848 , 
 n414849 , n414850 , n68127 , n414852 , n414853 , n68130 , n68131 , n414856 , n414857 , n68134 , 
 n414859 , n68136 , n414861 , n68138 , n414863 , n414864 , n68141 , n68142 , n414867 , n414868 , 
 n68145 , n414870 , n414871 , n68148 , n68149 , n414874 , n414875 , n68152 , n414877 , n414878 , 
 n414879 , n68156 , n68157 , n414882 , n414883 , n68160 , n68161 , n68162 , n414887 , n414888 , 
 n68165 , n68166 , n68167 , n414892 , n414893 , n68170 , n68171 , n68172 , n414897 , n68174 , 
 n68175 , n68176 , n68177 , n68178 , n68179 , n68180 , n68181 , n68182 , n68183 , n68184 , 
 n68185 , n68186 , n68187 , n68188 , n68189 , n68190 , n68191 , n414916 , n68193 , n68194 , 
 n414919 , n414920 , n68197 , n414922 , n414923 , n68200 , n68201 , n414926 , n414927 , n68204 , 
 n414929 , n68206 , n68207 , n68208 , n68209 , n68210 , n68211 , n68212 , n414937 , n68214 , 
 n68215 , n68216 , n68217 , n68218 , n68219 , n68220 , n414945 , n414946 , n414947 , n68224 , 
 n414949 , n414950 , n68227 , n68228 , n414953 , n68230 , n68231 , n68232 , n68233 , n414958 , 
 n68235 , n68236 , n414961 , n414962 , n414963 , n414964 , n68241 , n414966 , n414967 , n68244 , 
 n68245 , n414970 , n414971 , n414972 , n68249 , n414974 , n414975 , n68252 , n68253 , n414978 , 
 n414979 , n68256 , n414981 , n68258 , n414983 , n68260 , n68261 , n414986 , n414987 , n68264 , 
 n414989 , n414990 , n68267 , n68268 , n414993 , n414994 , n414995 , n68272 , n68273 , n414998 , 
 n414999 , n68276 , n68277 , n68278 , n415003 , n415004 , n68281 , n68282 , n68283 , n415008 , 
 n415009 , n68286 , n68287 , n68288 , n415013 , n415014 , n68291 , n68292 , n68293 , n415018 , 
 n415019 , n68296 , n68297 , n415022 , n415023 , n68300 , n68301 , n68302 , n68303 , n68304 , 
 n415029 , n68306 , n68307 , n68308 , n68309 , n68310 , n68311 , n68312 , n68313 , n415038 , 
 n68315 , n68316 , n68317 , n68318 , n68319 , n68320 , n68321 , n415046 , n68323 , n68324 , 
 n68325 , n415050 , n68327 , n68328 , n68329 , n68330 , n68331 , n68332 , n68333 , n68334 , 
 n68335 , n68336 , n68337 , n68338 , n68339 , n68340 , n68341 , n68342 , n68343 , n68344 , 
 n415069 , n68346 , n68347 , n68348 , n68349 , n68350 , n68351 , n68352 , n68353 , n68354 , 
 n68355 , n68356 , n68357 , n68358 , n68359 , n68360 , n68361 , n415086 , n68363 , n68364 , 
 n415089 , n68366 , n415091 , n68368 , n68369 , n415094 , n415095 , n68372 , n415097 , n68374 , 
 n68375 , n68376 , n415101 , n415102 , n68379 , n415104 , n415105 , n68382 , n415107 , n415108 , 
 n68385 , n415110 , n68387 , n68388 , n68389 , n68390 , n415115 , n415116 , n415117 , n68394 , 
 n68395 , n415120 , n415121 , n68398 , n68399 , n415124 , n68401 , n68402 , n68403 , n415128 , 
 n415129 , n68406 , n68407 , n415132 , n68409 , n68410 , n415135 , n68412 , n68413 , n68414 , 
 n68415 , n68416 , n68417 , n68418 , n68419 , n68420 , n415145 , n415146 , n68423 , n415148 , 
 n68425 , n415150 , n415151 , n68428 , n415153 , n415154 , n415155 , n68432 , n415157 , n68434 , 
 n68435 , n415160 , n415161 , n68438 , n415163 , n415164 , n68441 , n415166 , n415167 , n68444 , 
 n415169 , n68446 , n68447 , n415172 , n415173 , n68450 , n415175 , n415176 , n68453 , n415178 , 
 n415179 , n68456 , n415181 , n68458 , n415183 , n68460 , n415185 , n68462 , n68463 , n415188 , 
 n415189 , n68466 , n415191 , n415192 , n68469 , n415194 , n415195 , n68472 , n68473 , n415198 , 
 n68475 , n415200 , n68477 , n68478 , n415203 , n415204 , n68481 , n415206 , n415207 , n68484 , 
 n415209 , n415210 , n415211 , n68488 , n415213 , n415214 , n68491 , n415216 , n415217 , n68494 , 
 n68495 , n68496 , n415221 , n68498 , n68499 , n415224 , n415225 , n68502 , n415227 , n415228 , 
 n68505 , n415230 , n68507 , n415232 , n68509 , n68510 , n68511 , n415236 , n68513 , n68514 , 
 n415239 , n68520 , n415241 , n68522 , n68524 , n68525 , n68526 , n415246 , n415247 , n68529 , 
 n415249 , n415250 , n68532 , n68533 , n68534 , n415254 , n415255 , n68537 , n415257 , n68539 , 
 n68540 , n68541 , n68542 , n68543 , n68544 , n68545 , n68546 , n68547 , n415267 , n415268 , 
 n68550 , n415270 , n415271 , n68553 , n415273 , n68555 , n68556 , n415276 , n415277 , n68559 , 
 n415279 , n415280 , n68562 , n415282 , n68564 , n415284 , n68566 , n415286 , n415287 , n68569 , 
 n68570 , n68571 , n68572 , n68573 , n68574 , n68575 , n68576 , n68577 , n415297 , n415298 , 
 n68580 , n415300 , n68582 , n68583 , n415303 , n415304 , n68586 , n415306 , n68588 , n68589 , 
 n68590 , n415310 , n68592 , n415312 , n68594 , n68595 , n415315 , n415316 , n68598 , n415318 , 
 n415319 , n68601 , n415321 , n415322 , n415323 , n68605 , n415325 , n68607 , n68608 , n68609 , 
 n68610 , n68611 , n68612 , n68613 , n68614 , n68615 , n68616 , n68617 , n68618 , n68619 , 
 n415339 , n68621 , n415341 , n68623 , n68624 , n415344 , n415345 , n68627 , n415347 , n415348 , 
 n68630 , n415350 , n68632 , n68633 , n415353 , n415354 , n68636 , n415356 , n68638 , n68639 , 
 n68640 , n68641 , n68642 , n68643 , n68644 , n68645 , n68646 , n68647 , n68648 , n68649 , 
 n68650 , n68651 , n415371 , n68653 , n415373 , n68655 , n415375 , n68657 , n415377 , n68659 , 
 n68660 , n68661 , n68662 , n68663 , n415383 , n415384 , n68666 , n415386 , n68668 , n68669 , 
 n68670 , n68671 , n68672 , n68673 , n415393 , n68675 , n415395 , n68677 , n68678 , n415398 , 
 n415399 , n68681 , n415401 , n415402 , n68684 , n415404 , n68686 , n68687 , n68688 , n415408 , 
 n415409 , n68691 , n415411 , n68693 , n68694 , n68695 , n68696 , n68697 , n68698 , n68699 , 
 n68700 , n68701 , n68702 , n68703 , n68704 , n68705 , n415425 , n415426 , n68708 , n415428 , 
 n68710 , n68711 , n68712 , n68713 , n68714 , n68715 , n68716 , n68717 , n415437 , n68719 , 
 n68720 , n68721 , n68722 , n68723 , n68724 , n68725 , n68726 , n68727 , n68728 , n68729 , 
 n415449 , n68731 , n415451 , n68733 , n68734 , n415454 , n415455 , n68737 , n415457 , n415458 , 
 n68740 , n415460 , n68742 , n68743 , n68744 , n68745 , n68746 , n68747 , n68748 , n68749 , 
 n68750 , n68751 , n68752 , n415472 , n68754 , n415474 , n68756 , n68757 , n415477 , n68759 , 
 n415479 , n415480 , n68762 , n68763 , n415483 , n68765 , n415485 , n68767 , n68768 , n68769 , 
 n68770 , n415490 , n415491 , n68773 , n415493 , n415494 , n68776 , n415496 , n68778 , n415498 , 
 n68780 , n68781 , n415501 , n415502 , n68784 , n415504 , n68786 , n68787 , n415507 , n415508 , 
 n68790 , n415510 , n415511 , n68793 , n415513 , n415514 , n68796 , n68797 , n415517 , n68799 , 
 n415519 , n415520 , n68802 , n68803 , n415523 , n68805 , n68806 , n415526 , n415527 , n68809 , 
 n415529 , n68811 , n68812 , n415532 , n68814 , n415534 , n68816 , n415536 , n415537 , n68819 , 
 n415539 , n415540 , n68822 , n415542 , n68824 , n68825 , n415545 , n415546 , n68828 , n415548 , 
 n68830 , n68831 , n68832 , n68833 , n68834 , n415554 , n415555 , n68837 , n415557 , n68839 , 
 n68840 , n68841 , n415561 , n68843 , n68844 , n68845 , n68846 , n415566 , n68848 , n415568 , 
 n415569 , n68851 , n415571 , n68853 , n415573 , n68855 , n68856 , n415576 , n415577 , n68859 , 
 n415579 , n415580 , n68862 , n415582 , n415583 , n68865 , n68866 , n415586 , n68868 , n415588 , 
 n415589 , n68871 , n415591 , n68873 , n68874 , n415594 , n68876 , n415596 , n68878 , n68879 , 
 n415599 , n415600 , n68882 , n415602 , n415603 , n68885 , n415605 , n415606 , n68888 , n415608 , 
 n68890 , n68891 , n415611 , n415612 , n68894 , n415614 , n415615 , n68897 , n415617 , n68899 , 
 n415619 , n68901 , n415621 , n415622 , n68904 , n415624 , n68906 , n68907 , n415627 , n415628 , 
 n68910 , n415630 , n415631 , n68913 , n415633 , n68915 , n68916 , n68917 , n68918 , n68919 , 
 n68920 , n68921 , n415641 , n68923 , n415643 , n68925 , n68926 , n68927 , n68928 , n68929 , 
 n68930 , n415650 , n415651 , n68933 , n415653 , n415654 , n68936 , n415656 , n68938 , n68939 , 
 n68940 , n68941 , n68942 , n415662 , n68944 , n415664 , n68946 , n415666 , n68948 , n415668 , 
 n68950 , n68951 , n68952 , n68953 , n415673 , n68955 , n415675 , n68957 , n68958 , n415678 , 
 n415679 , n68961 , n415681 , n415682 , n68964 , n68965 , n415685 , n68967 , n68968 , n415688 , 
 n415689 , n68971 , n68972 , n68973 , n415693 , n68975 , n415695 , n415696 , n68978 , n415698 , 
 n415699 , n68981 , n415701 , n415702 , n68984 , n68985 , n68986 , n415706 , n415707 , n68989 , 
 n415709 , n415710 , n68992 , n415712 , n415713 , n68995 , n415715 , n415716 , n415717 , n68999 , 
 n415719 , n69001 , n415721 , n415722 , n69004 , n415724 , n415725 , n69007 , n415727 , n415728 , 
 n69010 , n415730 , n415731 , n69013 , n415733 , n415734 , n69016 , n415736 , n415737 , n69019 , 
 n415739 , n69021 , n69022 , n415742 , n69024 , n69025 , n69026 , n415746 , n415747 , n69029 , 
 n69030 , n415750 , n69032 , n415752 , n69034 , n69035 , n69036 , n69037 , n415757 , n69039 , 
 n415759 , n69041 , n69042 , n69043 , n415763 , n69045 , n415765 , n69047 , n69048 , n415768 , 
 n415769 , n69051 , n415771 , n69053 , n415773 , n69055 , n69056 , n69057 , n69058 , n415778 , 
 n415779 , n69061 , n415781 , n415782 , n69064 , n69065 , n415785 , n69067 , n69068 , n415788 , 
 n415789 , n415790 , n415791 , n69073 , n69074 , n415794 , n69076 , n69077 , n415797 , n415798 , 
 n415799 , n69081 , n69082 , n415802 , n69084 , n69085 , n415805 , n415806 , n69088 , n69089 , 
 n415809 , n69091 , n415811 , n415812 , n415813 , n69095 , n415815 , n69097 , n415817 , n415818 , 
 n69100 , n415820 , n415821 , n69103 , n415823 , n415824 , n415825 , n415826 , n69108 , n415828 , 
 n415829 , n69111 , n415831 , n415832 , n69114 , n69115 , n69116 , n415836 , n415837 , n69119 , 
 n69120 , n69121 , n415841 , n415842 , n69124 , n415844 , n415845 , n69127 , n69128 , n415848 , 
 n415849 , n69131 , n69132 , n415852 , n69134 , n415854 , n415855 , n69137 , n69138 , n69139 , 
 n69140 , n69144 , n69145 , n69146 , n415863 , n415864 , n415865 , n415866 , n69174 , n415868 , 
 n69176 , n415870 , n69178 , n69179 , n415873 , n415874 , n69182 , n415876 , n415877 , n69185 , 
 n415879 , n415880 , n69188 , n415882 , n69190 , n69191 , n415885 , n415886 , n69194 , n415888 , 
 n415889 , n69197 , n415891 , n415892 , n415893 , n69201 , n69202 , n69203 , n69204 , n69205 , 
 n415899 , n69207 , n69208 , n415902 , n415903 , n69211 , n415905 , n415906 , n69214 , n415908 , 
 n415909 , n69217 , n415911 , n69219 , n415913 , n69221 , n69222 , n415916 , n69224 , n415918 , 
 n415919 , n415920 , n415921 , n69229 , n415923 , n69231 , n415925 , n415926 , n69234 , n415928 , 
 n415929 , n69237 , n415931 , n415932 , n69240 , n415934 , n69242 , n415936 , n69244 , n69245 , 
 n69246 , n69247 , n69248 , n69249 , n69250 , n69251 , n69252 , n69253 , n69254 , n69255 , 
 n69256 , n69257 , n69258 , n69259 , n69260 , n69261 , n69262 , n69263 , n415957 , n69265 , 
 n415959 , n415960 , n69268 , n69269 , n415963 , n69271 , n415965 , n69273 , n415967 , n415968 , 
 n69276 , n69277 , n69278 , n69279 , n69280 , n69281 , n69282 , n69283 , n69284 , n69285 , 
 n69286 , n69287 , n69288 , n69289 , n69290 , n415984 , n69292 , n415986 , n69294 , n69295 , 
 n415989 , n415990 , n69298 , n415992 , n415993 , n69301 , n415995 , n415996 , n415997 , n69305 , 
 n415999 , n69307 , n69308 , n69309 , n69310 , n69311 , n416005 , n416006 , n416007 , n69315 , 
 n416009 , n416010 , n69318 , n416012 , n416013 , n69321 , n416015 , n416016 , n69324 , n416018 , 
 n416019 , n69327 , n416021 , n416022 , n69330 , n69331 , n69332 , n416026 , n416027 , n69335 , 
 n69337 , n416030 , n416031 , n69340 , n69341 , n69342 , n416035 , n416036 , n69345 , n416038 , 
 n416039 , n69348 , n69349 , n416042 , n416043 , n416044 , n416045 , n416046 , n69355 , n416048 , 
 n69357 , n416050 , n416051 , n69360 , n416053 , n416054 , n69363 , n416056 , n69365 , n416058 , 
 n69367 , n416060 , n69369 , n69370 , n69371 , n69372 , n69373 , n69374 , n69375 , n416068 , 
 n416069 , n69378 , n416071 , n416072 , n69381 , n416074 , n416075 , n416076 , n416077 , n69386 , 
 n416079 , n69388 , n416081 , n416082 , n69391 , n416084 , n69393 , n416086 , n69395 , n69396 , 
 n416089 , n416090 , n69399 , n416092 , n416093 , n69402 , n416095 , n416096 , n416097 , n69406 , 
 n416099 , n416100 , n69409 , n69410 , n416103 , n69412 , n69413 , n416106 , n416107 , n69416 , 
 n416109 , n69418 , n416111 , n416112 , n69421 , n69422 , n416115 , n69424 , n69425 , n416118 , 
 n69427 , n69428 , n69429 , n69430 , n69431 , n69432 , n416125 , n69434 , n416127 , n69436 , 
 n69437 , n69438 , n69439 , n69440 , n416133 , n69442 , n416135 , n69444 , n69445 , n416138 , 
 n416139 , n69448 , n416141 , n416142 , n69451 , n416144 , n69453 , n69454 , n69455 , n69456 , 
 n416149 , n69458 , n416151 , n69460 , n69461 , n416154 , n69463 , n416156 , n69465 , n69466 , 
 n416159 , n416160 , n69469 , n416162 , n416163 , n69472 , n416165 , n416166 , n69475 , n416168 , 
 n69477 , n69478 , n416171 , n416172 , n69481 , n416174 , n416175 , n69484 , n416177 , n69486 , 
 n416179 , n69488 , n416181 , n69490 , n69491 , n416184 , n416185 , n69494 , n416187 , n416188 , 
 n69497 , n416190 , n416191 , n69500 , n416193 , n69502 , n69503 , n416196 , n416197 , n69506 , 
 n416199 , n416200 , n69509 , n416202 , n69511 , n69512 , n416205 , n416206 , n69515 , n416208 , 
 n416209 , n69518 , n416211 , n69520 , n69521 , n416214 , n416215 , n69524 , n416217 , n416218 , 
 n69527 , n416220 , n416221 , n69530 , n416223 , n69532 , n69533 , n416226 , n416227 , n69536 , 
 n416229 , n416230 , n69539 , n416232 , n416233 , n416234 , n416235 , n69544 , n416237 , n69546 , 
 n416239 , n69548 , n69549 , n416242 , n416243 , n69552 , n416245 , n416246 , n69555 , n416248 , 
 n69557 , n416250 , n69559 , n416252 , n416253 , n69562 , n416255 , n416256 , n69565 , n69566 , 
 n69567 , n69568 , n69569 , n69570 , n69571 , n69572 , n69573 , n69574 , n69575 , n69576 , 
 n416269 , n69578 , n69579 , n69580 , n69581 , n416274 , n69583 , n416276 , n69585 , n69586 , 
 n416279 , n416280 , n69589 , n416282 , n416283 , n69592 , n416285 , n416286 , n69595 , n416288 , 
 n69597 , n416290 , n69599 , n416292 , n416293 , n69602 , n69603 , n416296 , n69605 , n416298 , 
 n416299 , n416300 , n69609 , n416302 , n416303 , n69612 , n416305 , n416306 , n69615 , n416308 , 
 n69617 , n69618 , n416311 , n416312 , n69621 , n416314 , n416315 , n69624 , n416317 , n416318 , 
 n69627 , n69628 , n69629 , n416322 , n416323 , n69632 , n416325 , n416326 , n416327 , n416328 , 
 n69637 , n416330 , n416331 , n69640 , n416333 , n69642 , n69643 , n416336 , n416337 , n69646 , 
 n416339 , n69648 , n69649 , n416342 , n416343 , n69652 , n416345 , n416346 , n69655 , n416348 , 
 n416349 , n69658 , n416351 , n416352 , n69661 , n416354 , n416355 , n69664 , n416357 , n416358 , 
 n69667 , n416360 , n416361 , n69670 , n416363 , n69672 , n416365 , n69674 , n69675 , n416368 , 
 n416369 , n69678 , n416371 , n416372 , n69681 , n416374 , n416375 , n69684 , n416377 , n69686 , 
 n69687 , n416380 , n416381 , n69690 , n416383 , n416384 , n69693 , n416386 , n416387 , n69696 , 
 n69697 , n69698 , n416391 , n69700 , n69701 , n69702 , n416395 , n69704 , n69705 , n69706 , 
 n416399 , n69708 , n69709 , n69710 , n416403 , n416404 , n69713 , n69714 , n416407 , n69716 , 
 n69717 , n69718 , n416411 , n69720 , n69721 , n69722 , n69723 , n69724 , n69725 , n69726 , 
 n69727 , n69728 , n69729 , n69730 , n69731 , n69732 , n69733 , n69734 , n69735 , n69736 , 
 n69737 , n69738 , n69739 , n69740 , n69741 , n69742 , n69743 , n69744 , n69745 , n69746 , 
 n69747 , n69748 , n69749 , n69750 , n69751 , n416444 , n69753 , n69754 , n69755 , n416448 , 
 n416449 , n69758 , n69759 , n69760 , n416453 , n416454 , n69763 , n69764 , n69765 , n416458 , 
 n69767 , n69768 , n69769 , n416462 , n416463 , n416464 , n69773 , n416466 , n69775 , n416468 , 
 n416469 , n69778 , n69779 , n416472 , n416473 , n69782 , n69783 , n69784 , n69785 , n69786 , 
 n69787 , n69788 , n69789 , n69790 , n69791 , n69792 , n416485 , n69799 , n416487 , n416488 , 
 n69815 , n416490 , n69834 , n416492 , n69836 , n69837 , n416495 , n416496 , n69840 , n69841 , 
 n416499 , n69843 , n69844 , n416502 , n69846 , n416504 , n69848 , n69849 , n69850 , n69851 , 
 n69852 , n69853 , n416511 , n416512 , n69856 , n416514 , n416515 , n69859 , n416517 , n416518 , 
 n69862 , n416520 , n416521 , n69865 , n416523 , n69867 , n416525 , n416526 , n69870 , n69871 , 
 n416529 , n69873 , n69874 , n416532 , n416533 , n69877 , n69878 , n69879 , n69880 , n416538 , 
 n69882 , n416540 , n416541 , n69885 , n69886 , n416544 , n416545 , n69889 , n416547 , n69891 , 
 n416549 , n69893 , n416551 , n69895 , n69896 , n416554 , n416555 , n69899 , n416557 , n416558 , 
 n69902 , n416560 , n416561 , n69905 , n416563 , n69907 , n69908 , n416566 , n416567 , n69911 , 
 n416569 , n416570 , n69914 , n416572 , n69916 , n69917 , n69918 , n69919 , n69920 , n69921 , 
 n69922 , n69923 , n69924 , n69925 , n69926 , n69927 , n69928 , n69929 , n69930 , n69931 , 
 n69932 , n69933 , n69934 , n416592 , n69936 , n416594 , n416595 , n416596 , n69940 , n416598 , 
 n416599 , n416600 , n69944 , n416602 , n416603 , n69947 , n416605 , n69949 , n69950 , n69952 , 
 n416609 , n69954 , n69956 , n416612 , n416613 , n69959 , n69960 , n69961 , n416617 , n69963 , 
 n69964 , n69965 , n416621 , n416622 , n416623 , n416624 , n69993 , n69994 , n416627 , n416628 , 
 n69997 , n69998 , n69999 , n416632 , n416633 , n70002 , n416635 , n70004 , n416637 , n70006 , 
 n70007 , n416640 , n416641 , n70010 , n416643 , n416644 , n70013 , n416646 , n416647 , n70016 , 
 n416649 , n70018 , n70019 , n416652 , n416653 , n70022 , n416655 , n416656 , n70025 , n416658 , 
 n416659 , n70028 , n416661 , n416662 , n70031 , n416664 , n70033 , n416666 , n70035 , n416668 , 
 n70037 , n70038 , n70039 , n70040 , n416673 , n70042 , n70043 , n416676 , n70045 , n416678 , 
 n70047 , n70048 , n416681 , n70050 , n416683 , n70052 , n70053 , n416686 , n416687 , n70056 , 
 n416689 , n416690 , n70059 , n416692 , n416693 , n416694 , n70063 , n416696 , n416697 , n70066 , 
 n416699 , n416700 , n70069 , n416702 , n416703 , n416704 , n70073 , n416706 , n70075 , n416708 , 
 n416709 , n70078 , n416711 , n416712 , n416713 , n416714 , n70083 , n416716 , n70085 , n416718 , 
 n416719 , n70088 , n70089 , n70090 , n70091 , n70092 , n70093 , n70094 , n70095 , n416728 , 
 n416729 , n70098 , n416731 , n70100 , n416733 , n70102 , n70103 , n70104 , n416737 , n416738 , 
 n70107 , n70108 , n416741 , n416742 , n70111 , n70112 , n70113 , n70114 , n416747 , n70116 , 
 n416749 , n70118 , n70119 , n416752 , n416753 , n70122 , n416755 , n416756 , n70125 , n416758 , 
 n70127 , n416760 , n70129 , n416762 , n70131 , n70132 , n416765 , n416766 , n70135 , n416768 , 
 n70137 , n70138 , n70139 , n70140 , n70141 , n70142 , n70143 , n70144 , n70145 , n70146 , 
 n416779 , n70148 , n70149 , n70150 , n70151 , n416784 , n416785 , n70154 , n416787 , n416788 , 
 n70157 , n70158 , n416791 , n416792 , n416793 , n70162 , n416795 , n416796 , n70165 , n70166 , 
 n416799 , n416800 , n416801 , n416802 , n70171 , n416804 , n416805 , n70174 , n70175 , n416808 , 
 n416809 , n70178 , n416811 , n416812 , n416813 , n70182 , n416815 , n416816 , n70185 , n70186 , 
 n416819 , n416820 , n70189 , n70190 , n70191 , n70192 , n70193 , n70194 , n70195 , n416828 , 
 n70197 , n416830 , n416831 , n416832 , n70201 , n416834 , n416835 , n70204 , n70205 , n416838 , 
 n416839 , n70208 , n70209 , n70210 , n416843 , n70212 , n416845 , n416846 , n416847 , n70216 , 
 n416849 , n416850 , n70219 , n70220 , n416853 , n416854 , n416855 , n70224 , n416857 , n70226 , 
 n70227 , n416860 , n416861 , n70230 , n70231 , n416864 , n70233 , n70234 , n416867 , n416868 , 
 n416869 , n70238 , n70239 , n416872 , n416873 , n70242 , n416875 , n416876 , n70245 , n70246 , 
 n70247 , n416880 , n416881 , n70250 , n416883 , n416884 , n70253 , n416886 , n416887 , n70256 , 
 n70257 , n416890 , n70259 , n70260 , n70261 , n416894 , n70263 , n70264 , n70265 , n416898 , 
 n416899 , n70268 , n70269 , n416902 , n416903 , n70272 , n70273 , n70274 , n416907 , n70276 , 
 n70277 , n70278 , n416911 , n70280 , n70281 , n70282 , n416915 , n70284 , n70285 , n70286 , 
 n70287 , n70288 , n70289 , n70290 , n416923 , n70292 , n70293 , n70294 , n416927 , n416928 , 
 n70297 , n416930 , n416931 , n70300 , n70301 , n416934 , n70303 , n70304 , n70305 , n70306 , 
 n416939 , n416940 , n70309 , n416942 , n416943 , n70312 , n70313 , n416946 , n416947 , n416948 , 
 n70317 , n416950 , n416951 , n70320 , n70321 , n416954 , n416955 , n416956 , n416957 , n70326 , 
 n416959 , n416960 , n70329 , n70330 , n416963 , n416964 , n416965 , n70334 , n416967 , n416968 , 
 n70337 , n70338 , n416971 , n416972 , n70341 , n70342 , n416975 , n416976 , n416977 , n416978 , 
 n70347 , n416980 , n416981 , n70350 , n70351 , n416984 , n416985 , n416986 , n70355 , n416988 , 
 n416989 , n70358 , n416991 , n416992 , n70361 , n70362 , n416995 , n416996 , n416997 , n70366 , 
 n70367 , n417000 , n417001 , n70370 , n417003 , n417004 , n70373 , n417006 , n417007 , n70376 , 
 n70377 , n417010 , n417011 , n417012 , n70381 , n417014 , n417015 , n70384 , n70385 , n417018 , 
 n417019 , n70388 , n70389 , n417022 , n70391 , n417024 , n417025 , n417026 , n70395 , n417028 , 
 n417029 , n70398 , n70399 , n417032 , n417033 , n70402 , n417035 , n70404 , n417037 , n417038 , 
 n70407 , n417040 , n417041 , n70410 , n70411 , n417044 , n417045 , n70414 , n417047 , n417048 , 
 n70417 , n70418 , n417051 , n417052 , n70421 , n70422 , n417055 , n417056 , n70425 , n70426 , 
 n70427 , n417060 , n417061 , n70430 , n70431 , n70432 , n417065 , n417066 , n70435 , n70436 , 
 n70437 , n417070 , n70439 , n70440 , n70441 , n417074 , n417075 , n417076 , n70445 , n417078 , 
 n417079 , n70448 , n70449 , n417082 , n417083 , n417084 , n70453 , n417086 , n417087 , n70456 , 
 n70457 , n417090 , n417091 , n417092 , n417093 , n70462 , n417095 , n417096 , n70465 , n70466 , 
 n417099 , n417100 , n417101 , n70470 , n417103 , n417104 , n70473 , n70474 , n417107 , n417108 , 
 n417109 , n417110 , n70479 , n417112 , n417113 , n70482 , n70483 , n417116 , n417117 , n70486 , 
 n70487 , n70488 , n417121 , n417122 , n70491 , n70492 , n70493 , n417126 , n417127 , n70496 , 
 n417129 , n70498 , n417131 , n417132 , n70501 , n417134 , n417135 , n70504 , n70505 , n417138 , 
 n417139 , n70508 , n417141 , n417142 , n70511 , n70512 , n417145 , n417146 , n70515 , n70516 , 
 n417149 , n417150 , n70519 , n70520 , n70521 , n417154 , n417155 , n70524 , n70525 , n70526 , 
 n417159 , n417160 , n70529 , n70530 , n70531 , n417164 , n70533 , n70534 , n70535 , n70536 , 
 n70537 , n70538 , n70539 , n70540 , n70541 , n70542 , n417175 , n417176 , n417177 , n70546 , 
 n417179 , n417180 , n70549 , n70550 , n417183 , n417184 , n417185 , n70554 , n417187 , n417188 , 
 n70557 , n70558 , n417191 , n417192 , n70561 , n70562 , n70563 , n417196 , n417197 , n70566 , 
 n70567 , n70568 , n417201 , n417202 , n70571 , n70572 , n417205 , n417206 , n70575 , n70576 , 
 n70577 , n417210 , n417211 , n70580 , n70581 , n70582 , n417215 , n70584 , n70585 , n417218 , 
 n70587 , n70588 , n70589 , n417222 , n70591 , n70592 , n70593 , n70594 , n70595 , n70596 , 
 n70597 , n70598 , n70599 , n70600 , n70601 , n70602 , n70603 , n70604 , n417237 , n417238 , 
 n70607 , n417240 , n70609 , n70610 , n70611 , n70612 , n70613 , n70614 , n417247 , n417248 , 
 n70617 , n417250 , n417251 , n70620 , n417253 , n417254 , n70623 , n70624 , n70625 , n70626 , 
 n417259 , n417260 , n70629 , n417262 , n70631 , n70632 , n70633 , n70634 , n417267 , n70636 , 
 n417269 , n70638 , n417271 , n70640 , n417273 , n70642 , n70643 , n70644 , n417277 , n417278 , 
 n417279 , n70648 , n417281 , n70650 , n70651 , n70652 , n70653 , n70654 , n70655 , n417288 , 
 n417289 , n70658 , n417291 , n417292 , n70661 , n417294 , n417295 , n70664 , n70665 , n70666 , 
 n417299 , n417300 , n417301 , n70670 , n417303 , n70672 , n70673 , n417306 , n70675 , n417308 , 
 n70677 , n70678 , n417311 , n417312 , n70681 , n417314 , n417315 , n70684 , n417317 , n417318 , 
 n417319 , n70688 , n417321 , n417322 , n70691 , n417324 , n417325 , n70694 , n70695 , n70696 , 
 n70697 , n70698 , n70699 , n70700 , n70701 , n417334 , n70703 , n417336 , n70705 , n70706 , 
 n417339 , n417340 , n70709 , n417342 , n70711 , n70712 , n417345 , n70714 , n417347 , n70716 , 
 n417349 , n417350 , n70719 , n70720 , n417353 , n417354 , n70723 , n417356 , n417357 , n70726 , 
 n417359 , n417360 , n417361 , n70730 , n417363 , n417364 , n70733 , n417366 , n417367 , n70736 , 
 n417369 , n70738 , n417371 , n70740 , n70741 , n417374 , n417375 , n70744 , n417377 , n417378 , 
 n70747 , n417380 , n417381 , n70750 , n417383 , n70752 , n70753 , n417386 , n417387 , n70756 , 
 n417389 , n417390 , n70759 , n417392 , n417393 , n70762 , n70763 , n70764 , n417397 , n417398 , 
 n70767 , n70768 , n70769 , n417402 , n417403 , n70772 , n70773 , n70774 , n417407 , n417408 , 
 n417409 , n70778 , n417411 , n70780 , n417413 , n70782 , n70783 , n417416 , n417417 , n70786 , 
 n417419 , n417420 , n70789 , n417422 , n417423 , n70792 , n70793 , n417426 , n417427 , n70796 , 
 n417429 , n417430 , n70799 , n417432 , n417433 , n70802 , n70803 , n417436 , n70805 , n417438 , 
 n70807 , n70808 , n417441 , n417442 , n70811 , n70812 , n417445 , n417446 , n70815 , n417448 , 
 n70817 , n70818 , n417451 , n417452 , n70821 , n417454 , n70823 , n417456 , n70825 , n70826 , 
 n70827 , n417460 , n417461 , n70830 , n417463 , n417464 , n70833 , n417466 , n417467 , n70836 , 
 n70838 , n417470 , n417471 , n70841 , n70842 , n70843 , n417475 , n417476 , n70846 , n70847 , 
 n70848 , n417480 , n417481 , n70851 , n70852 , n70853 , n417485 , n417486 , n70856 , n70857 , 
 n70858 , n417490 , n417491 , n70861 , n417493 , n417494 , n70864 , n417496 , n417497 , n70867 , 
 n417499 , n417500 , n70870 , n417502 , n417503 , n70873 , n417505 , n417506 , n70876 , n417508 , 
 n70878 , n417510 , n70880 , n417512 , n70882 , n417514 , n70884 , n70885 , n417517 , n417518 , 
 n70888 , n417520 , n417521 , n70891 , n417523 , n417524 , n70894 , n70895 , n417527 , n70897 , 
 n417529 , n70899 , n70900 , n417532 , n417533 , n70903 , n417535 , n417536 , n70906 , n417538 , 
 n417539 , n417540 , n70910 , n417542 , n417543 , n70913 , n417545 , n417546 , n70916 , n417548 , 
 n417549 , n417550 , n417551 , n70921 , n417553 , n70923 , n70924 , n417556 , n70926 , n417558 , 
 n417559 , n417560 , n70930 , n417562 , n70932 , n417564 , n417565 , n70935 , n417567 , n417568 , 
 n70938 , n417570 , n70940 , n417572 , n417573 , n70943 , n417575 , n70945 , n70946 , n417578 , 
 n417579 , n70949 , n417581 , n417582 , n70952 , n417584 , n417585 , n70955 , n417587 , n70957 , 
 n70958 , n417590 , n70960 , n417592 , n70962 , n70963 , n417595 , n417596 , n70966 , n417598 , 
 n417599 , n70969 , n417601 , n417602 , n417603 , n70973 , n417605 , n417606 , n70976 , n417608 , 
 n417609 , n417610 , n70980 , n417612 , n70982 , n70983 , n417615 , n70985 , n417617 , n417618 , 
 n417619 , n70989 , n417621 , n417622 , n70992 , n417624 , n417625 , n417626 , n70996 , n417628 , 
 n70998 , n417630 , n417631 , n71001 , n71002 , n417634 , n71004 , n71005 , n417637 , n71007 , 
 n71008 , n71009 , n417641 , n417642 , n71012 , n417644 , n417645 , n71015 , n71016 , n417648 , 
 n417649 , n417650 , n71020 , n417652 , n417653 , n71023 , n417655 , n417656 , n71026 , n71027 , 
 n417659 , n417660 , n417661 , n71031 , n71032 , n417664 , n417665 , n417666 , n417667 , n71037 , 
 n417669 , n417670 , n71040 , n71041 , n417673 , n417674 , n417675 , n71045 , n417677 , n417678 , 
 n71048 , n417680 , n417681 , n71051 , n71052 , n417684 , n417685 , n417686 , n71056 , n71057 , 
 n417689 , n417690 , n417691 , n417692 , n71062 , n417694 , n417695 , n71065 , n71066 , n417698 , 
 n417699 , n417700 , n71070 , n417702 , n417703 , n71073 , n417705 , n417706 , n71076 , n71077 , 
 n417709 , n417710 , n417711 , n71081 , n71082 , n417714 , n417715 , n417716 , n71086 , n71087 , 
 n71088 , n417720 , n71090 , n417722 , n417723 , n71093 , n71094 , n71095 , n417727 , n71097 , 
 n417729 , n417730 , n417731 , n71101 , n71102 , n417734 , n417735 , n71105 , n417737 , n71107 , 
 n417739 , n417740 , n417741 , n417742 , n417743 , n71113 , n71114 , n417746 , n417747 , n71117 , 
 n417749 , n417750 , n71120 , n71121 , n417753 , n417754 , n71124 , n417756 , n417757 , n71127 , 
 n71128 , n417760 , n417761 , n417762 , n71132 , n71133 , n417765 , n417766 , n71136 , n71137 , 
 n71138 , n417770 , n417771 , n71141 , n417773 , n417774 , n71144 , n417776 , n417777 , n71147 , 
 n71148 , n417780 , n417781 , n417782 , n71152 , n417784 , n417785 , n71155 , n417787 , n417788 , 
 n71158 , n71159 , n417791 , n417792 , n417793 , n71163 , n71164 , n417796 , n417797 , n417798 , 
 n71168 , n71169 , n71170 , n417802 , n71172 , n417804 , n417805 , n71175 , n417807 , n417808 , 
 n71178 , n71179 , n417811 , n417812 , n417813 , n71183 , n417815 , n71185 , n417817 , n417818 , 
 n71188 , n71189 , n417821 , n417822 , n71192 , n71193 , n417825 , n71195 , n71196 , n417828 , 
 n417829 , n417830 , n71200 , n71201 , n417833 , n417834 , n71204 , n417836 , n417837 , n71207 , 
 n71208 , n71209 , n417841 , n417842 , n71212 , n71213 , n71214 , n417846 , n417847 , n71217 , 
 n71218 , n71219 , n417851 , n417852 , n71222 , n417854 , n417855 , n71225 , n417857 , n417858 , 
 n71228 , n71229 , n417861 , n417862 , n417863 , n71233 , n417865 , n417866 , n71236 , n417868 , 
 n417869 , n71239 , n71240 , n417872 , n417873 , n417874 , n71244 , n71245 , n417877 , n417878 , 
 n417879 , n417880 , n71250 , n417882 , n417883 , n71253 , n71254 , n417886 , n417887 , n417888 , 
 n71258 , n417890 , n417891 , n71261 , n417893 , n417894 , n71264 , n71265 , n417897 , n417898 , 
 n417899 , n71269 , n71270 , n417902 , n417903 , n71273 , n417905 , n417906 , n71276 , n417908 , 
 n417909 , n71279 , n71280 , n417912 , n417913 , n417914 , n417915 , n71285 , n417917 , n417918 , 
 n71288 , n71289 , n417921 , n417922 , n71292 , n417924 , n417925 , n417926 , n417927 , n71297 , 
 n417929 , n417930 , n71300 , n71301 , n417933 , n417934 , n71304 , n417936 , n417937 , n71307 , 
 n417939 , n417940 , n71310 , n417942 , n417943 , n71313 , n71314 , n417946 , n417947 , n417948 , 
 n71318 , n71319 , n417951 , n417952 , n71322 , n417954 , n417955 , n71325 , n71326 , n71327 , 
 n417959 , n417960 , n71330 , n71331 , n71332 , n417964 , n417965 , n417966 , n71336 , n417968 , 
 n417969 , n71339 , n71340 , n417972 , n417973 , n417974 , n71344 , n417976 , n417977 , n71347 , 
 n417979 , n417980 , n71350 , n71351 , n417983 , n417984 , n417985 , n71355 , n71356 , n417988 , 
 n71358 , n71359 , n71360 , n71361 , n71362 , n71363 , n71364 , n71365 , n71366 , n417998 , 
 n417999 , n418000 , n418001 , n71371 , n418003 , n418004 , n71374 , n418006 , n418007 , n71377 , 
 n71378 , n418010 , n418011 , n418012 , n418013 , n71383 , n418015 , n418016 , n71386 , n418018 , 
 n418019 , n71389 , n418021 , n418022 , n71392 , n418024 , n418025 , n71395 , n71396 , n418028 , 
 n418029 , n418030 , n71400 , n71401 , n418033 , n418034 , n71404 , n71405 , n71406 , n418038 , 
 n71408 , n71409 , n418041 , n418042 , n71412 , n418044 , n418045 , n71415 , n418047 , n418048 , 
 n71418 , n71419 , n418051 , n418052 , n418053 , n71423 , n71424 , n418056 , n418057 , n71427 , 
 n418059 , n418060 , n71430 , n71431 , n71432 , n418064 , n418065 , n71435 , n418067 , n418068 , 
 n418069 , n71439 , n418071 , n418072 , n71442 , n418074 , n418075 , n71445 , n71446 , n418078 , 
 n418079 , n418080 , n71450 , n71451 , n418083 , n71453 , n418085 , n418086 , n71456 , n418088 , 
 n418089 , n71459 , n71460 , n418092 , n418093 , n418094 , n71464 , n418096 , n418097 , n71467 , 
 n71468 , n418100 , n71470 , n71471 , n71472 , n418104 , n418105 , n418106 , n71476 , n418108 , 
 n418109 , n71479 , n71480 , n418112 , n418113 , n418114 , n418115 , n71485 , n418117 , n418118 , 
 n71488 , n71489 , n418121 , n418122 , n71492 , n418124 , n418125 , n71495 , n418127 , n418128 , 
 n71498 , n71499 , n418131 , n418132 , n71502 , n418134 , n418135 , n71505 , n71506 , n71507 , 
 n418139 , n418140 , n71510 , n71511 , n71512 , n71513 , n418145 , n418146 , n71516 , n418148 , 
 n418149 , n71519 , n418151 , n418152 , n71522 , n71523 , n418155 , n418156 , n71526 , n418158 , 
 n418159 , n71529 , n418161 , n71531 , n71532 , n71533 , n71534 , n71535 , n71536 , n71537 , 
 n71538 , n71539 , n71540 , n418172 , n418173 , n71543 , n71544 , n71545 , n71546 , n418178 , 
 n418179 , n418180 , n418181 , n71551 , n418183 , n418184 , n71554 , n71555 , n418187 , n418188 , 
 n71558 , n71559 , n71560 , n418192 , n418193 , n71563 , n418195 , n418196 , n71566 , n71567 , 
 n71568 , n71569 , n71570 , n418202 , n71572 , n71573 , n71574 , n71575 , n418207 , n418208 , 
 n71578 , n71579 , n71580 , n418212 , n418213 , n71583 , n418215 , n418216 , n71586 , n418218 , 
 n71588 , n71589 , n71590 , n71591 , n71592 , n71593 , n71594 , n71595 , n71596 , n71597 , 
 n418229 , n71599 , n71600 , n418232 , n71602 , n71603 , n71604 , n418236 , n418237 , n71607 , 
 n418239 , n418240 , n71610 , n71611 , n418243 , n418244 , n418245 , n71615 , n418247 , n418248 , 
 n71618 , n71619 , n418251 , n418252 , n418253 , n418254 , n71624 , n418256 , n418257 , n71627 , 
 n71628 , n418260 , n418261 , n418262 , n71632 , n418264 , n418265 , n71635 , n71636 , n418268 , 
 n418269 , n418270 , n418271 , n418272 , n71642 , n418274 , n418275 , n71645 , n71646 , n418278 , 
 n418279 , n71649 , n418281 , n418282 , n71652 , n71653 , n418285 , n418286 , n71656 , n71657 , 
 n71658 , n71659 , n71660 , n71661 , n71662 , n71663 , n71664 , n418296 , n71666 , n418298 , 
 n418299 , n71669 , n418301 , n418302 , n71672 , n71673 , n418305 , n71675 , n418307 , n71677 , 
 n71678 , n71679 , n71680 , n71681 , n418313 , n71683 , n418315 , n418316 , n71686 , n418318 , 
 n418319 , n71689 , n71690 , n418322 , n418323 , n418324 , n418325 , n418326 , n71696 , n418328 , 
 n418329 , n71699 , n71700 , n418332 , n418333 , n71703 , n418335 , n418336 , n71706 , n71707 , 
 n418339 , n418340 , n71710 , n418342 , n71712 , n71713 , n71714 , n418346 , n71716 , n71717 , 
 n418349 , n418350 , n71720 , n71721 , n71722 , n418354 , n418355 , n418356 , n71726 , n418358 , 
 n418359 , n71729 , n71730 , n418362 , n418363 , n418364 , n71734 , n418366 , n418367 , n71737 , 
 n71738 , n418370 , n71740 , n418372 , n418373 , n71743 , n418375 , n418376 , n71746 , n71747 , 
 n418379 , n418380 , n418381 , n71751 , n418383 , n418384 , n71754 , n71755 , n418387 , n71757 , 
 n71758 , n71759 , n418391 , n71761 , n71762 , n71763 , n418395 , n418396 , n71766 , n71767 , 
 n71768 , n418400 , n71770 , n71771 , n71772 , n71773 , n71774 , n418406 , n71776 , n418408 , 
 n418409 , n71779 , n418411 , n418412 , n71782 , n71783 , n418415 , n418416 , n418417 , n71787 , 
 n418419 , n418420 , n71790 , n71791 , n418423 , n418424 , n71794 , n71795 , n418427 , n418428 , 
 n71798 , n418430 , n418431 , n71801 , n418433 , n418434 , n71804 , n71805 , n418437 , n418438 , 
 n418439 , n71809 , n418441 , n418442 , n71812 , n71813 , n418445 , n418446 , n418447 , n418448 , 
 n71818 , n418450 , n418451 , n71821 , n71822 , n418454 , n418455 , n71825 , n418457 , n418458 , 
 n418459 , n71829 , n418461 , n418462 , n71832 , n71833 , n418465 , n418466 , n71836 , n418468 , 
 n418469 , n71839 , n418471 , n418472 , n71842 , n71843 , n418475 , n418476 , n418477 , n71847 , 
 n418479 , n418480 , n71850 , n71851 , n418483 , n71853 , n71854 , n71855 , n418487 , n71857 , 
 n418489 , n71859 , n71860 , n418492 , n418493 , n71863 , n418495 , n418496 , n71866 , n71867 , 
 n418499 , n418500 , n418501 , n71871 , n71872 , n418504 , n71874 , n71875 , n71876 , n71877 , 
 n71878 , n418510 , n71880 , n71881 , n71882 , n418514 , n418515 , n71885 , n71886 , n71887 , 
 n418519 , n418520 , n418521 , n418522 , n71892 , n418524 , n418525 , n71895 , n71896 , n418528 , 
 n418529 , n418530 , n71900 , n418532 , n418533 , n71903 , n71904 , n418536 , n418537 , n71907 , 
 n418539 , n71909 , n418541 , n418542 , n71912 , n71913 , n71914 , n418546 , n71916 , n71917 , 
 n418549 , n71919 , n71920 , n71921 , n71922 , n71923 , n71924 , n71925 , n71926 , n418558 , 
 n71928 , n71929 , n71930 , n418562 , n71932 , n71933 , n71934 , n71935 , n71936 , n71937 , 
 n418569 , n71939 , n71940 , n71941 , n71942 , n71943 , n71944 , n418576 , n71946 , n71947 , 
 n418579 , n71949 , n71950 , n71951 , n71952 , n71953 , n71954 , n418586 , n71956 , n71957 , 
 n71958 , n71959 , n71960 , n71961 , n71962 , n71963 , n71964 , n71965 , n71966 , n71967 , 
 n71968 , n71969 , n71970 , n71971 , n71972 , n71973 , n71974 , n71975 , n71976 , n71977 , 
 n71978 , n418610 , n418611 , n71981 , n418613 , n71983 , n418615 , n71985 , n71986 , n418618 , 
 n418619 , n71989 , n418621 , n418622 , n71992 , n418624 , n418625 , n71995 , n71996 , n418628 , 
 n71998 , n418630 , n72000 , n72001 , n418633 , n418634 , n72004 , n418636 , n418637 , n72007 , 
 n418639 , n418640 , n418641 , n72011 , n418643 , n418644 , n72014 , n418646 , n418647 , n72017 , 
 n72018 , n72019 , n72020 , n72021 , n72022 , n72023 , n72024 , n72025 , n72026 , n72027 , 
 n72028 , n72029 , n418661 , n72031 , n72032 , n72033 , n418665 , n418666 , n72036 , n418668 , 
 n72038 , n418670 , n72040 , n72041 , n418673 , n72043 , n418675 , n72045 , n72046 , n418678 , 
 n418679 , n72049 , n418681 , n418682 , n72052 , n418684 , n418685 , n418686 , n72056 , n418688 , 
 n418689 , n72059 , n418691 , n418692 , n72062 , n72063 , n72064 , n418696 , n418697 , n72067 , 
 n418699 , n418700 , n72070 , n72071 , n418703 , n72073 , n418705 , n72075 , n72076 , n418708 , 
 n72078 , n72079 , n418711 , n418712 , n72082 , n418714 , n418715 , n72085 , n418717 , n418718 , 
 n72088 , n72089 , n418721 , n418722 , n72092 , n418724 , n72094 , n72095 , n418727 , n72097 , 
 n418729 , n418730 , n72100 , n418732 , n72102 , n418734 , n418735 , n72105 , n418737 , n418738 , 
 n72108 , n418740 , n418741 , n72111 , n418743 , n418744 , n72114 , n418746 , n72116 , n418748 , 
 n418749 , n72119 , n72120 , n418752 , n72122 , n72123 , n418755 , n418756 , n72126 , n418758 , 
 n72128 , n72129 , n418761 , n418762 , n72132 , n418764 , n418765 , n72135 , n418767 , n72137 , 
 n72138 , n72139 , n72140 , n418772 , n72142 , n418774 , n72144 , n72145 , n418777 , n418778 , 
 n72148 , n418780 , n418781 , n72151 , n418783 , n72153 , n72154 , n418786 , n418787 , n72157 , 
 n418789 , n72159 , n72160 , n72161 , n418793 , n72163 , n72164 , n418796 , n72166 , n418798 , 
 n72168 , n72169 , n418801 , n418802 , n72172 , n418804 , n418805 , n72175 , n418807 , n418808 , 
 n72178 , n418810 , n418811 , n72181 , n418813 , n72183 , n72184 , n418816 , n418817 , n72187 , 
 n418819 , n418820 , n72190 , n418822 , n418823 , n72193 , n72194 , n418826 , n418827 , n418828 , 
 n72198 , n418830 , n418831 , n72201 , n72202 , n418834 , n418835 , n418836 , n72206 , n418838 , 
 n418839 , n72209 , n72210 , n418842 , n72212 , n72213 , n72214 , n418846 , n418847 , n72217 , 
 n418849 , n418850 , n72220 , n72221 , n418853 , n418854 , n418855 , n72225 , n418857 , n418858 , 
 n72228 , n72229 , n418861 , n72231 , n72232 , n72233 , n72234 , n72235 , n72236 , n72237 , 
 n72238 , n418870 , n72240 , n72241 , n72242 , n72243 , n72244 , n72245 , n418877 , n418878 , 
 n72248 , n418880 , n418881 , n72251 , n72252 , n418884 , n418885 , n418886 , n72256 , n418888 , 
 n418889 , n72259 , n72260 , n418892 , n418893 , n418894 , n418895 , n72265 , n418897 , n418898 , 
 n72268 , n72269 , n418901 , n418902 , n72272 , n418904 , n418905 , n418906 , n72276 , n418908 , 
 n418909 , n72279 , n72280 , n418912 , n418913 , n72283 , n418915 , n418916 , n72286 , n418918 , 
 n418919 , n72289 , n418921 , n418922 , n418923 , n72293 , n418925 , n418926 , n72296 , n72297 , 
 n418929 , n418930 , n72300 , n418932 , n418933 , n72303 , n72304 , n418936 , n418937 , n418938 , 
 n72308 , n418940 , n72310 , n418942 , n418943 , n72313 , n418945 , n418946 , n72316 , n72317 , 
 n418949 , n418950 , n72320 , n418952 , n72322 , n418954 , n72324 , n72325 , n418957 , n418958 , 
 n418959 , n72329 , n418961 , n418962 , n72332 , n72333 , n418965 , n418966 , n72336 , n72337 , 
 n418969 , n418970 , n72340 , n72341 , n72342 , n418974 , n418975 , n72345 , n72346 , n72347 , 
 n418979 , n418980 , n72350 , n418982 , n72352 , n418984 , n418985 , n72355 , n418987 , n418988 , 
 n72358 , n72359 , n418991 , n418992 , n72362 , n418994 , n418995 , n72365 , n72366 , n418998 , 
 n418999 , n72369 , n419001 , n419002 , n72372 , n72373 , n419005 , n419006 , n419007 , n72377 , 
 n72378 , n419010 , n419011 , n72381 , n72382 , n72383 , n419015 , n419016 , n419017 , n419018 , 
 n72388 , n419020 , n419021 , n72391 , n72392 , n419024 , n419025 , n419026 , n72396 , n419028 , 
 n419029 , n72399 , n72400 , n419032 , n419033 , n72403 , n72404 , n72405 , n419037 , n419038 , 
 n72408 , n72409 , n419041 , n419042 , n419043 , n419044 , n419045 , n72415 , n419047 , n419048 , 
 n72418 , n72419 , n419051 , n419052 , n72422 , n72423 , n419055 , n419056 , n72426 , n419058 , 
 n72428 , n419060 , n419061 , n72431 , n419063 , n419064 , n72434 , n72435 , n419067 , n419068 , 
 n72438 , n419070 , n419071 , n72441 , n72442 , n419074 , n419075 , n72445 , n72446 , n419078 , 
 n419079 , n72449 , n72450 , n72451 , n419083 , n419084 , n72454 , n72455 , n72456 , n419088 , 
 n419089 , n72459 , n72460 , n72461 , n419093 , n72463 , n72464 , n72465 , n72466 , n72467 , 
 n72468 , n72469 , n419101 , n419102 , n72472 , n419104 , n419105 , n72475 , n72476 , n419108 , 
 n419109 , n419110 , n72480 , n419112 , n419113 , n72483 , n72484 , n419116 , n419117 , n419118 , 
 n419119 , n72489 , n419121 , n419122 , n72492 , n72493 , n419125 , n419126 , n419127 , n72497 , 
 n419129 , n419130 , n72500 , n72501 , n419133 , n419134 , n72504 , n72505 , n72506 , n419138 , 
 n419139 , n72509 , n72510 , n72511 , n419143 , n72513 , n72514 , n72515 , n72516 , n72517 , 
 n419149 , n72519 , n419151 , n419152 , n72522 , n419154 , n419155 , n72525 , n72526 , n419158 , 
 n419159 , n72529 , n419161 , n419162 , n72532 , n72533 , n419165 , n419166 , n72536 , n72537 , 
 n419169 , n72539 , n72540 , n72541 , n419173 , n419174 , n419175 , n72545 , n419177 , n419178 , 
 n72548 , n72549 , n419181 , n419182 , n419183 , n72553 , n419185 , n419186 , n72556 , n72557 , 
 n419189 , n419190 , n72560 , n72561 , n72562 , n419194 , n419195 , n72565 , n72566 , n72567 , 
 n419199 , n72569 , n72570 , n72571 , n419203 , n72573 , n72574 , n72575 , n72576 , n72577 , 
 n72578 , n72579 , n72580 , n72581 , n72582 , n72583 , n72584 , n72585 , n419217 , n72587 , 
 n72588 , n419220 , n419221 , n72591 , n72592 , n72593 , n72594 , n72595 , n419227 , n72597 , 
 n419229 , n72599 , n72600 , n419232 , n419233 , n72603 , n419235 , n419236 , n72606 , n419238 , 
 n419239 , n72609 , n419241 , n419242 , n72612 , n419244 , n72614 , n419246 , n72616 , n419248 , 
 n72618 , n419250 , n419251 , n72621 , n72622 , n419254 , n72624 , n419256 , n72626 , n419258 , 
 n419259 , n72629 , n419261 , n419262 , n72632 , n72633 , n419265 , n72635 , n419267 , n72637 , 
 n72638 , n72639 , n419271 , n419272 , n72642 , n419274 , n419275 , n72645 , n419277 , n419278 , 
 n419279 , n72649 , n419281 , n419282 , n419283 , n419284 , n419285 , n72655 , n72656 , n72657 , 
 n419289 , n72659 , n72660 , n72661 , n419293 , n72663 , n419295 , n419296 , n72666 , n419298 , 
 n72668 , n419300 , n72670 , n72671 , n419303 , n72673 , n419305 , n72675 , n72676 , n419308 , 
 n419309 , n72679 , n419311 , n419312 , n72682 , n419314 , n419315 , n419316 , n72686 , n419318 , 
 n419319 , n72689 , n419321 , n419322 , n72692 , n72693 , n419325 , n419326 , n72696 , n72697 , 
 n72698 , n419330 , n419331 , n72701 , n419333 , n419334 , n72704 , n419336 , n419337 , n419338 , 
 n419339 , n72709 , n72710 , n419342 , n72712 , n72713 , n419345 , n419346 , n72716 , n419348 , 
 n419349 , n72719 , n419351 , n72721 , n72722 , n419354 , n72724 , n419356 , n72726 , n72727 , 
 n419359 , n419360 , n72730 , n419362 , n419363 , n72733 , n419365 , n419366 , n419367 , n72737 , 
 n419369 , n419370 , n72740 , n419372 , n419373 , n72743 , n419375 , n72745 , n419377 , n72747 , 
 n419379 , n72749 , n72750 , n419382 , n419383 , n72753 , n419385 , n419386 , n72756 , n419388 , 
 n419389 , n72759 , n419391 , n419392 , n72762 , n72763 , n419395 , n72765 , n419397 , n72767 , 
 n72768 , n419400 , n419401 , n72771 , n419403 , n419404 , n72774 , n419406 , n419407 , n419408 , 
 n72778 , n419410 , n419411 , n72781 , n419413 , n419414 , n72784 , n72785 , n72786 , n419418 , 
 n419419 , n72789 , n419421 , n72791 , n419423 , n72793 , n72794 , n419426 , n72796 , n72797 , 
 n419429 , n419430 , n72800 , n72801 , n419433 , n419434 , n72804 , n419436 , n419437 , n72807 , 
 n72808 , n72809 , n72810 , n72811 , n72812 , n419444 , n419445 , n72815 , n419447 , n419448 , 
 n72818 , n419450 , n419451 , n72821 , n419453 , n419454 , n72824 , n72825 , n419457 , n419458 , 
 n419459 , n72829 , n419461 , n72831 , n72832 , n419464 , n419465 , n72835 , n419467 , n419468 , 
 n72838 , n419470 , n419471 , n72841 , n419473 , n72843 , n72844 , n419476 , n419477 , n72847 , 
 n72848 , n419480 , n72850 , n72851 , n419483 , n419484 , n419485 , n72855 , n419487 , n419488 , 
 n72858 , n419490 , n419491 , n72861 , n419493 , n72863 , n72864 , n72865 , n72866 , n72867 , 
 n419499 , n72869 , n72870 , n419502 , n72872 , n419504 , n72874 , n72875 , n72876 , n419508 , 
 n72878 , n419510 , n419511 , n419512 , n72882 , n419514 , n419515 , n72885 , n419517 , n419518 , 
 n419519 , n72889 , n72890 , n72891 , n72892 , n72893 , n72894 , n72895 , n419527 , n72897 , 
 n419529 , n72899 , n419531 , n419532 , n419533 , n72903 , n419535 , n419536 , n72906 , n419538 , 
 n419539 , n72909 , n419541 , n419542 , n419543 , n72913 , n72914 , n419546 , n419547 , n72917 , 
 n419549 , n419550 , n419551 , n72921 , n419553 , n72923 , n72924 , n419556 , n419557 , n72927 , 
 n419559 , n419560 , n72930 , n419562 , n419563 , n72933 , n419565 , n72935 , n72936 , n419568 , 
 n72938 , n419570 , n72940 , n72941 , n419573 , n419574 , n72944 , n419576 , n419577 , n72947 , 
 n419579 , n419580 , n419581 , n72951 , n419583 , n419584 , n72954 , n419586 , n419587 , n72957 , 
 n72958 , n72959 , n72960 , n72961 , n419593 , n419594 , n419595 , n72965 , n419597 , n72967 , 
 n72968 , n419600 , n419601 , n72971 , n419603 , n419604 , n72974 , n419606 , n419607 , n72977 , 
 n419609 , n72979 , n72980 , n72981 , n72982 , n72983 , n72984 , n419616 , n419617 , n72987 , 
 n419619 , n419620 , n72990 , n419622 , n419623 , n72993 , n419625 , n72995 , n419627 , n72997 , 
 n72998 , n419630 , n419631 , n73001 , n419633 , n419634 , n73004 , n419636 , n419637 , n73007 , 
 n73008 , n73009 , n419641 , n419642 , n419643 , n73013 , n419645 , n73015 , n73016 , n419648 , 
 n419649 , n73019 , n419651 , n419652 , n73022 , n419654 , n419655 , n73025 , n73026 , n419658 , 
 n73028 , n73029 , n419661 , n73031 , n419663 , n73033 , n73034 , n419666 , n419667 , n73037 , 
 n419669 , n419670 , n73040 , n419672 , n419673 , n419674 , n73044 , n419676 , n419677 , n73047 , 
 n419679 , n73049 , n73050 , n73051 , n73052 , n73053 , n73054 , n419686 , n73056 , n419688 , 
 n73058 , n419690 , n73060 , n73061 , n419693 , n419694 , n73064 , n419696 , n419697 , n73067 , 
 n419699 , n419700 , n73070 , n419702 , n73072 , n73073 , n419705 , n419706 , n73076 , n419708 , 
 n419709 , n73079 , n419711 , n419712 , n73082 , n73083 , n73084 , n419716 , n419717 , n73087 , 
 n419719 , n419720 , n73090 , n73091 , n73092 , n419724 , n419725 , n419726 , n73096 , n419728 , 
 n73098 , n73099 , n419731 , n73101 , n419733 , n73103 , n73104 , n419736 , n419737 , n73107 , 
 n419739 , n419740 , n73110 , n419742 , n419743 , n419744 , n73114 , n419746 , n419747 , n73117 , 
 n419749 , n73119 , n419751 , n73121 , n419753 , n73123 , n419755 , n73125 , n419757 , n419758 , 
 n73128 , n73129 , n419761 , n419762 , n73132 , n419764 , n419765 , n73135 , n419767 , n419768 , 
 n73138 , n73139 , n419771 , n419772 , n73142 , n73143 , n419775 , n73145 , n73146 , n419778 , 
 n419779 , n73149 , n419781 , n73151 , n419783 , n419784 , n73154 , n419786 , n73156 , n73157 , 
 n73158 , n73159 , n73160 , n73161 , n73162 , n73163 , n73164 , n73165 , n73166 , n73167 , 
 n419799 , n73169 , n419801 , n419802 , n73196 , n419804 , n419805 , n73199 , n419807 , n73201 , 
 n419809 , n73203 , n73204 , n419812 , n73206 , n419814 , n73208 , n419816 , n419817 , n73211 , 
 n419819 , n73213 , n73214 , n73215 , n73216 , n73217 , n73218 , n73219 , n419827 , n73221 , 
 n419829 , n419830 , n73224 , n419832 , n419833 , n73227 , n73228 , n73229 , n73230 , n73231 , 
 n73232 , n419840 , n73234 , n419842 , n73236 , n73237 , n73238 , n73239 , n73240 , n73241 , 
 n419849 , n419850 , n73244 , n419852 , n419853 , n73247 , n419855 , n419856 , n73250 , n419858 , 
 n419859 , n419860 , n73254 , n419862 , n73256 , n419864 , n419865 , n73259 , n419867 , n419868 , 
 n73262 , n419870 , n419871 , n73265 , n73266 , n73267 , n73268 , n73269 , n419877 , n73271 , 
 n73272 , n73273 , n73274 , n73275 , n419883 , n73277 , n419885 , n73279 , n73280 , n419888 , 
 n73282 , n419890 , n73284 , n73285 , n419893 , n419894 , n73288 , n419896 , n419897 , n73291 , 
 n419899 , n419900 , n419901 , n73295 , n419903 , n419904 , n73298 , n419906 , n419907 , n73301 , 
 n73302 , n73303 , n73304 , n419912 , n73306 , n73307 , n73308 , n73309 , n419917 , n73311 , 
 n419919 , n419920 , n73314 , n419922 , n73316 , n73317 , n419925 , n419926 , n73320 , n419928 , 
 n419929 , n73323 , n419931 , n419932 , n73326 , n419934 , n73328 , n419936 , n73330 , n73331 , 
 n419939 , n73333 , n419941 , n73335 , n73336 , n419944 , n419945 , n73339 , n419947 , n419948 , 
 n419949 , n419950 , n419951 , n419952 , n73346 , n419954 , n419955 , n73349 , n419957 , n419958 , 
 n73352 , n419960 , n419961 , n73355 , n419963 , n73357 , n73358 , n73359 , n73360 , n73361 , 
 n419969 , n73363 , n73364 , n73365 , n73366 , n73367 , n73368 , n419976 , n419977 , n73371 , 
 n419979 , n419980 , n73374 , n419982 , n419983 , n73377 , n73378 , n73379 , n419987 , n419988 , 
 n419989 , n73383 , n419991 , n73385 , n73386 , n419994 , n419995 , n73389 , n419997 , n419998 , 
 n73392 , n420000 , n420001 , n73395 , n420003 , n73397 , n73398 , n420006 , n73400 , n420008 , 
 n73402 , n73403 , n420011 , n420012 , n73406 , n420014 , n420015 , n73409 , n420017 , n420018 , 
 n420019 , n73413 , n420021 , n420022 , n73416 , n420024 , n420025 , n73419 , n73420 , n73421 , 
 n73422 , n73423 , n420031 , n420032 , n420033 , n73427 , n420035 , n73429 , n73430 , n420038 , 
 n420039 , n73433 , n420041 , n420042 , n73436 , n420044 , n420045 , n73439 , n73440 , n73441 , 
 n420049 , n420050 , n73444 , n420052 , n420053 , n73447 , n73448 , n73449 , n420057 , n420058 , 
 n420059 , n73453 , n420061 , n73455 , n420063 , n73457 , n73458 , n420066 , n420067 , n73461 , 
 n420069 , n420070 , n73464 , n420072 , n420073 , n73467 , n73468 , n420076 , n73470 , n420078 , 
 n73472 , n73473 , n420081 , n73475 , n420083 , n73477 , n420085 , n420086 , n73480 , n420088 , 
 n420089 , n420090 , n73484 , n420092 , n420093 , n73487 , n420095 , n420096 , n73490 , n73491 , 
 n73492 , n420100 , n420101 , n420102 , n73496 , n420104 , n73498 , n73499 , n420107 , n420108 , 
 n73502 , n420110 , n420111 , n73505 , n420113 , n420114 , n73508 , n420116 , n73510 , n420118 , 
 n73512 , n73513 , n420121 , n73515 , n420123 , n73517 , n420125 , n73519 , n73520 , n73521 , 
 n73522 , n73523 , n420131 , n73525 , n420133 , n420134 , n73528 , n420136 , n420137 , n73531 , 
 n73532 , n73533 , n420141 , n420142 , n73536 , n73537 , n73538 , n420146 , n420147 , n73541 , 
 n420149 , n73543 , n73544 , n73545 , n73546 , n420154 , n420155 , n73549 , n420157 , n73551 , 
 n420159 , n73553 , n73554 , n420162 , n420163 , n73557 , n420165 , n420166 , n420167 , n420168 , 
 n420169 , n73563 , n420171 , n73565 , n420173 , n73567 , n73568 , n420176 , n73570 , n420178 , 
 n420179 , n420180 , n420181 , n420182 , n73576 , n420184 , n420185 , n73579 , n420187 , n420188 , 
 n73582 , n420190 , n73584 , n420192 , n73586 , n420194 , n73588 , n73589 , n420197 , n420198 , 
 n73592 , n420200 , n420201 , n73595 , n420203 , n73597 , n73598 , n420206 , n73600 , n420208 , 
 n73602 , n420210 , n73604 , n420212 , n73606 , n73607 , n73608 , n73609 , n73610 , n73611 , 
 n73612 , n73613 , n73614 , n73615 , n73616 , n73617 , n73618 , n73619 , n73620 , n73621 , 
 n420229 , n420230 , n73624 , n420232 , n73626 , n73627 , n420235 , n420236 , n73630 , n73631 , 
 n420239 , n73633 , n73634 , n420242 , n420243 , n420244 , n73638 , n420246 , n420247 , n73641 , 
 n420249 , n420250 , n73644 , n420252 , n73646 , n420254 , n73648 , n73649 , n420257 , n73651 , 
 n420259 , n73653 , n73654 , n420262 , n420263 , n73657 , n420265 , n420266 , n73660 , n420268 , 
 n420269 , n420270 , n73664 , n420272 , n420273 , n73667 , n420275 , n420276 , n73670 , n420278 , 
 n420279 , n73673 , n73674 , n73675 , n73676 , n73677 , n73678 , n73679 , n73680 , n73681 , 
 n420289 , n73683 , n420291 , n73685 , n420293 , n73687 , n420295 , n73689 , n73690 , n420298 , 
 n420299 , n73693 , n420301 , n420302 , n73696 , n420304 , n420305 , n73699 , n73700 , n420308 , 
 n420309 , n73703 , n420311 , n420312 , n73706 , n420314 , n420315 , n73709 , n420317 , n420318 , 
 n420319 , n420320 , n73714 , n420322 , n420323 , n73717 , n420325 , n73719 , n420327 , n73721 , 
 n73722 , n420330 , n420331 , n73725 , n73726 , n420334 , n420335 , n73729 , n420337 , n420338 , 
 n73732 , n420340 , n73734 , n420342 , n420343 , n73737 , n73738 , n420346 , n73740 , n73741 , 
 n420349 , n420350 , n73744 , n73745 , n420353 , n420354 , n73748 , n420356 , n420357 , n73751 , 
 n420359 , n420360 , n73754 , n420362 , n420363 , n73757 , n73758 , n420366 , n420367 , n73761 , 
 n73762 , n73763 , n420371 , n73765 , n420373 , n73767 , n420375 , n73769 , n73770 , n420378 , 
 n420379 , n73773 , n73774 , n420382 , n73776 , n73777 , n420385 , n420386 , n420387 , n73781 , 
 n420389 , n420390 , n73784 , n420392 , n420393 , n73787 , n420395 , n420396 , n73790 , n73791 , 
 n73792 , n73793 , n73794 , n73795 , n420403 , n420404 , n73798 , n73799 , n420407 , n420408 , 
 n73802 , n73803 , n73804 , n73805 , n73806 , n420414 , n73808 , n73809 , n73810 , n73811 , 
 n73812 , n73813 , n73814 , n73815 , n73816 , n73817 , n420425 , n73819 , n420427 , n73821 , 
 n73822 , n420430 , n420431 , n73825 , n420433 , n420434 , n73828 , n420436 , n73830 , n73831 , 
 n73832 , n420440 , n420441 , n73835 , n420443 , n73837 , n73838 , n73839 , n73840 , n73841 , 
 n73842 , n420450 , n73844 , n73845 , n420453 , n420454 , n420455 , n420456 , n73850 , n420458 , 
 n420459 , n73853 , n73854 , n420462 , n420463 , n420464 , n73858 , n420466 , n420467 , n73861 , 
 n73862 , n420470 , n420471 , n73865 , n73866 , n420474 , n420475 , n73869 , n420477 , n73871 , 
 n420479 , n73873 , n420481 , n420482 , n73876 , n73877 , n420485 , n420486 , n73880 , n420488 , 
 n420489 , n73883 , n73884 , n420492 , n420493 , n420494 , n73888 , n73889 , n420497 , n420498 , 
 n73892 , n73893 , n73894 , n420502 , n420503 , n73897 , n420505 , n420506 , n73900 , n420508 , 
 n420509 , n73903 , n73904 , n420512 , n420513 , n420514 , n73908 , n420516 , n420517 , n73911 , 
 n73912 , n420520 , n420521 , n420522 , n420523 , n73917 , n420525 , n420526 , n73920 , n73921 , 
 n420529 , n420530 , n420531 , n73925 , n420533 , n420534 , n73928 , n73929 , n420537 , n420538 , 
 n420539 , n420540 , n420541 , n73935 , n420543 , n420544 , n73938 , n73939 , n420547 , n420548 , 
 n73942 , n420550 , n420551 , n73945 , n73946 , n420554 , n420555 , n420556 , n420557 , n73951 , 
 n420559 , n420560 , n73954 , n73955 , n420563 , n420564 , n73958 , n420566 , n420567 , n73961 , 
 n420569 , n73963 , n73964 , n420572 , n420573 , n73967 , n73968 , n420576 , n420577 , n73971 , 
 n420579 , n420580 , n73974 , n73975 , n73976 , n420584 , n420585 , n73979 , n73980 , n73981 , 
 n420589 , n420590 , n73984 , n420592 , n420593 , n73987 , n420595 , n420596 , n73990 , n73991 , 
 n420599 , n420600 , n420601 , n73995 , n420603 , n420604 , n73998 , n73999 , n420607 , n420608 , 
 n74002 , n420610 , n74004 , n420612 , n420613 , n74007 , n420615 , n420616 , n74010 , n74011 , 
 n420619 , n74013 , n74014 , n420622 , n74016 , n74017 , n74018 , n420626 , n420627 , n74021 , 
 n420629 , n420630 , n74024 , n74025 , n420633 , n420634 , n420635 , n74029 , n420637 , n420638 , 
 n74032 , n74033 , n420641 , n74035 , n420643 , n74037 , n420645 , n420646 , n74040 , n420648 , 
 n420649 , n74043 , n74044 , n420652 , n420653 , n74047 , n74048 , n420656 , n420657 , n74051 , 
 n74052 , n420660 , n74054 , n74055 , n74056 , n420664 , n74058 , n74059 , n74060 , n420668 , 
 n74062 , n74063 , n74064 , n74065 , n74066 , n420674 , n420675 , n420676 , n420677 , n74071 , 
 n420679 , n420680 , n74074 , n74075 , n420683 , n420684 , n420685 , n74079 , n420687 , n420688 , 
 n74082 , n74083 , n420691 , n420692 , n74086 , n420694 , n74088 , n420696 , n74090 , n420698 , 
 n420699 , n74093 , n74094 , n420702 , n420703 , n74097 , n420705 , n420706 , n74100 , n74101 , 
 n420709 , n420710 , n420711 , n74105 , n74106 , n420714 , n420715 , n74109 , n74110 , n74111 , 
 n420719 , n74113 , n74114 , n74115 , n74116 , n74117 , n420725 , n74119 , n74120 , n74121 , 
 n420729 , n74123 , n74124 , n74125 , n74126 , n74127 , n420735 , n420736 , n420737 , n74131 , 
 n420739 , n420740 , n74134 , n74135 , n420743 , n420744 , n420745 , n74139 , n420747 , n420748 , 
 n74142 , n74143 , n420751 , n420752 , n420753 , n420754 , n74148 , n420756 , n420757 , n74151 , 
 n74152 , n420760 , n420761 , n420762 , n74156 , n420764 , n420765 , n74159 , n74160 , n420768 , 
 n420769 , n74163 , n74164 , n420772 , n420773 , n74167 , n420775 , n420776 , n74170 , n420778 , 
 n420779 , n74173 , n74174 , n420782 , n420783 , n420784 , n420785 , n420786 , n420787 , n74181 , 
 n74182 , n420790 , n420791 , n420792 , n420793 , n420794 , n74188 , n420796 , n420797 , n74191 , 
 n74192 , n420800 , n420801 , n74195 , n420803 , n420804 , n74198 , n74199 , n420807 , n420808 , 
 n420809 , n420810 , n74204 , n420812 , n420813 , n74207 , n420815 , n420816 , n420817 , n74211 , 
 n420819 , n420820 , n74214 , n74215 , n420823 , n420824 , n74218 , n420826 , n420827 , n74221 , 
 n74222 , n420830 , n420831 , n74225 , n74226 , n74227 , n420835 , n420836 , n74230 , n420838 , 
 n74232 , n420840 , n74234 , n74235 , n420843 , n420844 , n74238 , n420846 , n420847 , n74241 , 
 n74242 , n420850 , n420851 , n420852 , n74246 , n74247 , n420855 , n420856 , n74250 , n74251 , 
 n74252 , n420860 , n420861 , n74255 , n74256 , n74257 , n420865 , n420866 , n74260 , n74261 , 
 n74262 , n420870 , n420871 , n74265 , n74266 , n74267 , n420875 , n74269 , n74270 , n74271 , 
 n74272 , n74273 , n74274 , n74275 , n74276 , n420884 , n74278 , n74279 , n420887 , n420888 , 
 n74282 , n74283 , n74284 , n420892 , n420893 , n74287 , n74288 , n74289 , n420897 , n74291 , 
 n74292 , n74293 , n74294 , n74295 , n420903 , n74297 , n420905 , n420906 , n74300 , n420908 , 
 n420909 , n74303 , n420911 , n420912 , n74306 , n420914 , n74308 , n74309 , n420917 , n74311 , 
 n420919 , n420920 , n420921 , n74315 , n420923 , n420924 , n74318 , n420926 , n420927 , n74321 , 
 n420929 , n420930 , n74324 , n420932 , n420933 , n74327 , n74328 , n420936 , n420937 , n74331 , 
 n74332 , n74333 , n420941 , n74335 , n74336 , n74337 , n420945 , n74339 , n420947 , n74341 , 
 n74342 , n420950 , n74344 , n420952 , n74346 , n420954 , n420955 , n74349 , n74350 , n420958 , 
 n420959 , n74353 , n420961 , n420962 , n74356 , n420964 , n420965 , n420966 , n74360 , n420968 , 
 n420969 , n74363 , n420971 , n420972 , n74366 , n420974 , n74368 , n420976 , n74370 , n74371 , 
 n420979 , n74373 , n74374 , n74375 , n420983 , n420984 , n74378 , n420986 , n420987 , n74381 , 
 n420989 , n74383 , n74384 , n420992 , n74386 , n420994 , n420995 , n74389 , n420997 , n420998 , 
 n420999 , n74393 , n421001 , n421002 , n74396 , n421004 , n421005 , n74399 , n421007 , n421008 , 
 n74402 , n421010 , n74404 , n74405 , n74406 , n74407 , n74408 , n74409 , n74410 , n74411 , 
 n74412 , n421020 , n74414 , n421022 , n74416 , n421024 , n421025 , n74419 , n74420 , n421028 , 
 n421029 , n74423 , n421031 , n421032 , n74426 , n421034 , n74428 , n74429 , n74430 , n421038 , 
 n421039 , n74433 , n421041 , n74435 , n74436 , n74437 , n74438 , n74439 , n421047 , n74441 , 
 n74442 , n421050 , n421051 , n74445 , n74446 , n74447 , n421055 , n421056 , n74450 , n421058 , 
 n421059 , n74453 , n421061 , n74455 , n74456 , n74457 , n74458 , n421066 , n74460 , n74461 , 
 n74462 , n74463 , n421071 , n421072 , n74466 , n421074 , n74468 , n421076 , n74470 , n421078 , 
 n74472 , n421080 , n74474 , n74475 , n421083 , n421084 , n74478 , n421086 , n421087 , n74481 , 
 n421089 , n421090 , n74484 , n421092 , n74486 , n74487 , n421095 , n421096 , n74490 , n421098 , 
 n421099 , n74493 , n421101 , n421102 , n74496 , n74497 , n74498 , n421106 , n74500 , n74501 , 
 n74502 , n421110 , n74504 , n421112 , n421113 , n74507 , n421115 , n421116 , n421117 , n74511 , 
 n421119 , n74513 , n421121 , n421122 , n74516 , n421124 , n421125 , n74519 , n421127 , n421128 , 
 n74522 , n421130 , n421131 , n74525 , n421133 , n421134 , n74528 , n421136 , n421137 , n74531 , 
 n74532 , n74533 , n74534 , n74535 , n421143 , n421144 , n74538 , n421146 , n421147 , n74541 , 
 n421149 , n421150 , n74544 , n421152 , n74546 , n421154 , n74548 , n74549 , n421157 , n421158 , 
 n74552 , n421160 , n421161 , n74555 , n421163 , n421164 , n74558 , n421166 , n421167 , n74561 , 
 n421169 , n74563 , n74564 , n421172 , n421173 , n74567 , n74568 , n74569 , n74570 , n421178 , 
 n74572 , n74573 , n74574 , n74575 , n74576 , n74577 , n74578 , n74579 , n421187 , n74581 , 
 n421189 , n74583 , n421191 , n74585 , n421193 , n74587 , n74588 , n421196 , n74590 , n421198 , 
 n74592 , n421200 , n421201 , n74595 , n421203 , n421204 , n74598 , n74599 , n421207 , n421208 , 
 n74602 , n421210 , n421211 , n74605 , n421213 , n421214 , n74608 , n421216 , n421217 , n74611 , 
 n421219 , n74613 , n421221 , n74615 , n74616 , n421224 , n74618 , n421226 , n74620 , n74621 , 
 n421229 , n421230 , n74624 , n421232 , n421233 , n74627 , n421235 , n421236 , n421237 , n74631 , 
 n421239 , n421240 , n74634 , n421242 , n421243 , n74637 , n421245 , n421246 , n74640 , n74641 , 
 n74642 , n74643 , n421251 , n74645 , n421253 , n74647 , n74648 , n421256 , n421257 , n74651 , 
 n421259 , n421260 , n74654 , n421262 , n421263 , n74657 , n421265 , n74659 , n74660 , n421268 , 
 n74662 , n421270 , n421271 , n74665 , n74666 , n74667 , n74668 , n421276 , n421277 , n74671 , 
 n421279 , n74673 , n421281 , n74675 , n74676 , n421284 , n74678 , n421286 , n74680 , n74681 , 
 n421289 , n421290 , n74684 , n421292 , n421293 , n74687 , n421295 , n421296 , n421297 , n74691 , 
 n421299 , n421300 , n74694 , n421302 , n421303 , n74697 , n421305 , n74699 , n74700 , n74701 , 
 n74702 , n421310 , n74704 , n421312 , n74706 , n421314 , n74708 , n74709 , n421317 , n74711 , 
 n421319 , n74713 , n74714 , n421322 , n421323 , n74717 , n421325 , n421326 , n74720 , n421328 , 
 n421329 , n421330 , n74724 , n421332 , n421333 , n74727 , n421335 , n74729 , n74730 , n74731 , 
 n421339 , n421340 , n74734 , n421342 , n74736 , n74737 , n421345 , n74739 , n74740 , n74741 , 
 n421349 , n74743 , n421351 , n421352 , n74746 , n421354 , n421355 , n74749 , n74750 , n421358 , 
 n421359 , n74753 , n74754 , n421362 , n74756 , n74757 , n421365 , n74759 , n421367 , n74761 , 
 n74762 , n74763 , n74764 , n421372 , n74766 , n421374 , n74768 , n74769 , n74770 , n74771 , 
 n421379 , n421380 , n74774 , n421382 , n74776 , n421384 , n74778 , n74779 , n421387 , n421388 , 
 n74782 , n421390 , n421391 , n74785 , n421393 , n421394 , n74788 , n74789 , n421397 , n421398 , 
 n74792 , n421400 , n421401 , n74795 , n421403 , n421404 , n74798 , n421406 , n74800 , n74801 , 
 n74802 , n74803 , n421411 , n421412 , n421413 , n74807 , n74808 , n421416 , n74810 , n74811 , 
 n421419 , n421420 , n74814 , n421422 , n74816 , n74817 , n421425 , n74819 , n421427 , n74821 , 
 n74822 , n421430 , n421431 , n74825 , n421433 , n421434 , n74828 , n421436 , n421437 , n421438 , 
 n74832 , n421440 , n421441 , n74835 , n421443 , n421444 , n74838 , n421446 , n421447 , n74841 , 
 n74842 , n421450 , n74844 , n74845 , n421453 , n421454 , n74848 , n421456 , n421457 , n74851 , 
 n74852 , n421460 , n74854 , n74855 , n421463 , n421464 , n74858 , n421466 , n421467 , n74861 , 
 n421469 , n74869 , n421471 , n74886 , n74887 , n74888 , n74889 , n421476 , n421477 , n421478 , 
 n74893 , n421480 , n421481 , n421482 , n421483 , n74898 , n74899 , n421486 , n74901 , n74902 , 
 n421489 , n421490 , n74905 , n421492 , n421493 , n74908 , n74909 , n421496 , n421497 , n421498 , 
 n421499 , n74914 , n421501 , n421502 , n74917 , n421504 , n421505 , n421506 , n74921 , n421508 , 
 n74923 , n74924 , n421511 , n421512 , n74927 , n421514 , n421515 , n74930 , n421517 , n421518 , 
 n74933 , n421520 , n74935 , n421522 , n421523 , n421524 , n74939 , n421526 , n421527 , n74942 , 
 n421529 , n421530 , n74945 , n421532 , n421533 , n74948 , n74949 , n74950 , n421537 , n421538 , 
 n74955 , n421540 , n421541 , n74973 , n74974 , n421544 , n421545 , n421546 , n421547 , n74987 , 
 n421549 , n421550 , n74990 , n421552 , n421553 , n421554 , n421555 , n75013 , n75014 , n421558 , 
 n421559 , n75017 , n75018 , n75019 , n421563 , n421564 , n75022 , n421566 , n421567 , n421568 , 
 n421569 , n75030 , n421571 , n421572 , n75033 , n75034 , n421575 , n75036 , n421577 , n421578 , 
 n75039 , n75040 , n421581 , n421582 , n75043 , n421584 , n421585 , n75046 , n75047 , n421588 , 
 n421589 , n75050 , n421591 , n421592 , n75053 , n421594 , n421595 , n75056 , n75057 , n421598 , 
 n421599 , n75060 , n75061 , n421602 , n421603 , n421604 , n421605 , n75084 , n75085 , n75086 , 
 n421609 , n421610 , n75089 , n75091 , n421613 , n421614 , n75094 , n75095 , n75096 , n421618 , 
 n75098 , n75099 , n75100 , n421622 , n75102 , n421624 , n75104 , n75105 , n421627 , n421628 , 
 n75108 , n421630 , n421631 , n75111 , n421633 , n421634 , n421635 , n75115 , n421637 , n75117 , 
 n421639 , n75119 , n421641 , n75121 , n75122 , n421644 , n75124 , n421646 , n421647 , n75127 , 
 n421649 , n75129 , n421651 , n421652 , n75132 , n421654 , n421655 , n75135 , n421657 , n75137 , 
 n75138 , n421660 , n421661 , n75141 , n421663 , n421664 , n75144 , n421666 , n421667 , n421668 , 
 n75148 , n421670 , n75150 , n75151 , n421673 , n421674 , n75154 , n75155 , n421677 , n75157 , 
 n75158 , n421680 , n421681 , n75161 , n421683 , n75163 , n421685 , n421686 , n75166 , n421688 , 
 n421689 , n75169 , n421691 , n75171 , n421693 , n75173 , n75174 , n421696 , n421697 , n75177 , 
 n421699 , n421700 , n75180 , n421702 , n421703 , n75183 , n421705 , n75185 , n75186 , n421708 , 
 n421709 , n75189 , n421711 , n421712 , n75192 , n421714 , n421715 , n75195 , n75196 , n75197 , 
 n421719 , n75199 , n75200 , n75201 , n75202 , n75203 , n75204 , n75205 , n75206 , n75207 , 
 n421729 , n75209 , n421731 , n75211 , n75212 , n421734 , n421735 , n75215 , n421737 , n421738 , 
 n75218 , n421740 , n421741 , n75221 , n421743 , n75223 , n75224 , n421746 , n421747 , n75227 , 
 n421749 , n421750 , n75230 , n421752 , n75232 , n75233 , n75234 , n75235 , n421757 , n421758 , 
 n75238 , n421760 , n421761 , n75241 , n421763 , n421764 , n421765 , n75245 , n421767 , n75247 , 
 n421769 , n75249 , n75250 , n75251 , n421773 , n421774 , n75254 , n421776 , n75256 , n421778 , 
 n75258 , n421780 , n75260 , n75261 , n421783 , n421784 , n75264 , n421786 , n421787 , n75267 , 
 n421789 , n421790 , n75270 , n75271 , n421793 , n421794 , n75274 , n421796 , n421797 , n75277 , 
 n421799 , n421800 , n75280 , n75281 , n75282 , n421804 , n421805 , n421806 , n421807 , n75287 , 
 n75288 , n421810 , n75290 , n75291 , n421813 , n421814 , n75294 , n421816 , n75296 , n75297 , 
 n421819 , n75299 , n421821 , n75301 , n421823 , n421824 , n75304 , n421826 , n421827 , n421828 , 
 n75308 , n421830 , n75310 , n75311 , n421833 , n421834 , n75314 , n421836 , n421837 , n75317 , 
 n421839 , n421840 , n75320 , n421842 , n75322 , n75323 , n421845 , n421846 , n75326 , n421848 , 
 n421849 , n75329 , n421851 , n421852 , n75332 , n75333 , n421855 , n421856 , n75336 , n421858 , 
 n75338 , n421860 , n75340 , n75341 , n421863 , n75343 , n421865 , n75345 , n75346 , n421868 , 
 n421869 , n75349 , n421871 , n421872 , n75352 , n421874 , n421875 , n75355 , n421877 , n421878 , 
 n421879 , n75359 , n421881 , n421882 , n75362 , n421884 , n421885 , n75365 , n75366 , n75367 , 
 n421889 , n421890 , n75370 , n421892 , n75372 , n421894 , n75374 , n75375 , n421897 , n421898 , 
 n75378 , n75379 , n421901 , n421902 , n421903 , n75383 , n75384 , n421906 , n75386 , n75387 , 
 n421909 , n421910 , n75390 , n75391 , n75392 , n421914 , n421915 , n421916 , n421917 , n75417 , 
 n75418 , n421920 , n421921 , n75421 , n75422 , n75423 , n421925 , n421926 , n75426 , n421928 , 
 n421929 , n75429 , n75430 , n421932 , n75432 , n75433 , n421935 , n421936 , n75436 , n75437 , 
 n75438 , n75439 , n421941 , n75441 , n421943 , n421944 , n75444 , n421946 , n75446 , n421948 , 
 n421949 , n75449 , n75450 , n421952 , n75452 , n421954 , n75454 , n75455 , n421957 , n75457 , 
 n421959 , n75459 , n75460 , n421962 , n421963 , n75463 , n421965 , n421966 , n75466 , n421968 , 
 n421969 , n421970 , n75470 , n421972 , n421973 , n75473 , n421975 , n421976 , n75476 , n421978 , 
 n421979 , n75479 , n75480 , n421982 , n75482 , n75483 , n421985 , n421986 , n75486 , n421988 , 
 n421989 , n75489 , n421991 , n75491 , n75492 , n421994 , n421995 , n75495 , n421997 , n421998 , 
 n75498 , n422000 , n422001 , n75501 , n75502 , n422004 , n422005 , n75505 , n75506 , n75507 , 
 n422009 , n422010 , n75510 , n422012 , n422013 , n75513 , n422015 , n422016 , n75516 , n75517 , 
 n422019 , n422020 , n75520 , n422022 , n75522 , n422024 , n75524 , n75525 , n422027 , n422028 , 
 n75528 , n422030 , n422031 , n75531 , n422033 , n422034 , n75534 , n422036 , n75536 , n75537 , 
 n422039 , n422040 , n75540 , n422042 , n422043 , n75543 , n422045 , n422046 , n422047 , n75547 , 
 n422049 , n75549 , n75550 , n422052 , n75552 , n422054 , n75554 , n75555 , n422057 , n422058 , 
 n75558 , n422060 , n422061 , n75561 , n422063 , n422064 , n422065 , n75565 , n422067 , n422068 , 
 n75568 , n422070 , n422071 , n75571 , n75572 , n75573 , n422075 , n422076 , n75576 , n75577 , 
 n75578 , n422080 , n422081 , n75581 , n422083 , n75583 , n422085 , n75585 , n422087 , n75587 , 
 n75588 , n422090 , n75590 , n422092 , n75592 , n75593 , n422095 , n422096 , n75596 , n422098 , 
 n422099 , n75599 , n422101 , n422102 , n422103 , n75603 , n422105 , n422106 , n75606 , n422108 , 
 n75608 , n422110 , n75610 , n422112 , n75612 , n75613 , n422115 , n75615 , n422117 , n75617 , 
 n422119 , n422120 , n75620 , n422122 , n422123 , n75623 , n422125 , n75625 , n75626 , n422128 , 
 n422129 , n75629 , n422131 , n422132 , n75632 , n422134 , n422135 , n75635 , n422137 , n422138 , 
 n75638 , n75639 , n75640 , n75641 , n75642 , n422144 , n75644 , n422146 , n75646 , n75647 , 
 n422149 , n422150 , n75650 , n422152 , n422153 , n75653 , n422155 , n422156 , n75656 , n422158 , 
 n422159 , n75659 , n75660 , n75661 , n75662 , n422164 , n75664 , n422166 , n422167 , n75667 , 
 n422169 , n422170 , n422171 , n422172 , n75672 , n422174 , n422175 , n75675 , n422177 , n422178 , 
 n75678 , n422180 , n75680 , n422182 , n422183 , n75683 , n422185 , n75685 , n422187 , n75687 , 
 n75688 , n422190 , n422191 , n75691 , n422193 , n75693 , n75694 , n422196 , n422197 , n75697 , 
 n422199 , n75699 , n75700 , n422202 , n422203 , n75703 , n422205 , n422206 , n75706 , n422208 , 
 n422209 , n75709 , n75710 , n422212 , n422213 , n75713 , n422215 , n75715 , n75716 , n75717 , 
 n75718 , n422220 , n422221 , n422222 , n75722 , n422224 , n422225 , n75725 , n75726 , n422228 , 
 n422229 , n422230 , n75730 , n422232 , n422233 , n75733 , n75734 , n422236 , n75736 , n75737 , 
 n75738 , n422240 , n75740 , n422242 , n75742 , n422244 , n422245 , n75745 , n75746 , n422248 , 
 n422249 , n75749 , n422251 , n422252 , n75752 , n75753 , n422255 , n422256 , n422257 , n75757 , 
 n75758 , n422260 , n75760 , n75761 , n75762 , n75763 , n75764 , n75765 , n75766 , n75767 , 
 n422269 , n422270 , n422271 , n75771 , n422273 , n422274 , n75774 , n75775 , n422277 , n422278 , 
 n422279 , n75779 , n422281 , n422282 , n75782 , n75783 , n422285 , n75785 , n422287 , n75787 , 
 n422289 , n422290 , n75790 , n422292 , n422293 , n75793 , n75794 , n422296 , n422297 , n75797 , 
 n422299 , n422300 , n75800 , n75801 , n422303 , n422304 , n75804 , n75805 , n422307 , n75807 , 
 n75808 , n75809 , n422311 , n422312 , n422313 , n75813 , n422315 , n422316 , n75816 , n422318 , 
 n422319 , n422320 , n422321 , n75821 , n422323 , n422324 , n75824 , n75825 , n422327 , n422328 , 
 n422329 , n75829 , n422331 , n422332 , n75832 , n422334 , n422335 , n75835 , n75836 , n422338 , 
 n422339 , n422340 , n75840 , n75841 , n422343 , n422344 , n75844 , n422346 , n422347 , n422348 , 
 n422349 , n75849 , n422351 , n422352 , n75852 , n75853 , n422355 , n422356 , n75856 , n422358 , 
 n75858 , n422360 , n75860 , n422362 , n422363 , n75863 , n75864 , n422366 , n422367 , n75867 , 
 n422369 , n422370 , n75870 , n75871 , n422373 , n422374 , n422375 , n75875 , n75876 , n422378 , 
 n422379 , n75879 , n75880 , n75881 , n422383 , n75883 , n75884 , n75885 , n422387 , n422388 , 
 n422389 , n75889 , n422391 , n422392 , n75892 , n75893 , n422395 , n422396 , n75896 , n422398 , 
 n422399 , n75899 , n75900 , n422402 , n422403 , n422404 , n422405 , n422406 , n75906 , n422408 , 
 n422409 , n75909 , n75910 , n422412 , n422413 , n75913 , n422415 , n422416 , n75916 , n75917 , 
 n422419 , n422420 , n75920 , n422422 , n422423 , n75923 , n422425 , n422426 , n422427 , n422428 , 
 n422429 , n75929 , n422431 , n422432 , n75932 , n75933 , n422435 , n422436 , n75936 , n422438 , 
 n422439 , n75939 , n75940 , n422442 , n422443 , n75943 , n422445 , n422446 , n75946 , n75947 , 
 n75948 , n422450 , n75950 , n75951 , n422453 , n75953 , n422455 , n75955 , n422457 , n75957 , 
 n422459 , n422460 , n75960 , n75961 , n422463 , n422464 , n75964 , n422466 , n422467 , n75967 , 
 n75968 , n422470 , n422471 , n422472 , n75972 , n75973 , n422475 , n75975 , n75976 , n75977 , 
 n75978 , n75979 , n75980 , n75981 , n422483 , n422484 , n75984 , n75985 , n75986 , n422488 , 
 n422489 , n75989 , n75990 , n75991 , n422493 , n75993 , n75994 , n75995 , n75996 , n75997 , 
 n75998 , n75999 , n76000 , n422502 , n76002 , n76003 , n76004 , n76005 , n76006 , n76007 , 
 n76008 , n422510 , n422511 , n76011 , n422513 , n422514 , n76014 , n76015 , n422517 , n422518 , 
 n422519 , n76019 , n422521 , n422522 , n76022 , n76023 , n422525 , n422526 , n76026 , n76027 , 
 n422529 , n422530 , n422531 , n422532 , n76032 , n76033 , n422535 , n76035 , n76036 , n422538 , 
 n422539 , n76039 , n422541 , n422542 , n422543 , n76043 , n422545 , n422546 , n76046 , n76047 , 
 n422549 , n422550 , n76050 , n422552 , n422553 , n76053 , n422555 , n422556 , n76056 , n422558 , 
 n76058 , n422560 , n422561 , n422562 , n422563 , n422564 , n76064 , n422566 , n422567 , n76067 , 
 n76068 , n422570 , n422571 , n76071 , n422573 , n422574 , n76074 , n76075 , n422577 , n422578 , 
 n76078 , n422580 , n76080 , n422582 , n76082 , n76083 , n422585 , n422586 , n422587 , n76087 , 
 n422589 , n422590 , n76090 , n76091 , n422593 , n422594 , n76094 , n76095 , n422597 , n422598 , 
 n76098 , n76099 , n76100 , n422602 , n422603 , n76103 , n76104 , n76105 , n422607 , n422608 , 
 n76108 , n422610 , n422611 , n422612 , n422613 , n76113 , n422615 , n422616 , n76116 , n76117 , 
 n422619 , n422620 , n76120 , n76121 , n422623 , n422624 , n76124 , n76125 , n422627 , n422628 , 
 n76128 , n76129 , n76130 , n422632 , n422633 , n76133 , n76134 , n76135 , n76136 , n76137 , 
 n422639 , n76139 , n76140 , n76141 , n422643 , n76143 , n76144 , n76145 , n422647 , n76147 , 
 n76148 , n76149 , n76150 , n76151 , n76152 , n76153 , n76154 , n76155 , n76156 , n76157 , 
 n76158 , n76159 , n76160 , n76161 , n76162 , n422664 , n422665 , n76165 , n422667 , n76167 , 
 n76168 , n422670 , n422671 , n76171 , n422673 , n422674 , n76174 , n422676 , n422677 , n76177 , 
 n422679 , n76179 , n76180 , n76181 , n76182 , n76183 , n422685 , n76185 , n422687 , n76187 , 
 n422689 , n76189 , n76190 , n422692 , n422693 , n76193 , n422695 , n422696 , n76196 , n422698 , 
 n422699 , n76199 , n422701 , n76201 , n76202 , n422704 , n422705 , n76205 , n422707 , n422708 , 
 n76208 , n422710 , n422711 , n76211 , n422713 , n422714 , n76214 , n422716 , n76216 , n76217 , 
 n76218 , n76219 , n422721 , n76221 , n422723 , n76223 , n422725 , n76225 , n76226 , n422728 , 
 n76228 , n422730 , n76230 , n76231 , n422733 , n422734 , n76234 , n422736 , n422737 , n76237 , 
 n422739 , n422740 , n422741 , n76241 , n422743 , n422744 , n76244 , n422746 , n422747 , n76247 , 
 n76248 , n76249 , n422751 , n422752 , n76252 , n76253 , n76254 , n422756 , n76256 , n76257 , 
 n76258 , n76259 , n76260 , n422762 , n76262 , n76263 , n76264 , n422766 , n76279 , n76280 , 
 n76281 , n422770 , n76283 , n76285 , n422773 , n422774 , n422775 , n422776 , n76310 , n422778 , 
 n76312 , n76313 , n422781 , n422782 , n76316 , n76317 , n422785 , n76319 , n76320 , n422788 , 
 n422789 , n422790 , n76324 , n422792 , n422793 , n76327 , n422795 , n422796 , n76330 , n76331 , 
 n422799 , n76333 , n422801 , n422802 , n76336 , n422804 , n422805 , n76339 , n422807 , n76341 , 
 n422809 , n76343 , n76344 , n422812 , n422813 , n76347 , n422815 , n422816 , n76350 , n422818 , 
 n422819 , n76353 , n422821 , n76355 , n76356 , n422824 , n422825 , n76359 , n422827 , n422828 , 
 n76362 , n422830 , n422831 , n76365 , n422833 , n422834 , n76368 , n76369 , n76370 , n76371 , 
 n422839 , n76373 , n422841 , n422842 , n422843 , n76377 , n422845 , n76379 , n422847 , n422848 , 
 n76382 , n422850 , n422851 , n76385 , n76386 , n76387 , n422855 , n422856 , n76390 , n76391 , 
 n76392 , n422860 , n422861 , n76395 , n76397 , n422864 , n422865 , n76400 , n76401 , n76402 , 
 n422869 , n76404 , n76405 , n76406 , n422873 , n422874 , n76409 , n422876 , n422877 , n76412 , 
 n422879 , n76414 , n422881 , n422882 , n422883 , n76418 , n422885 , n422886 , n76421 , n422888 , 
 n422889 , n76424 , n422891 , n422892 , n76427 , n422894 , n422895 , n76430 , n422897 , n422898 , 
 n422899 , n76434 , n422901 , n76436 , n422903 , n422904 , n76439 , n422906 , n422907 , n422908 , 
 n76443 , n422910 , n76445 , n422912 , n76447 , n76448 , n422915 , n422916 , n76451 , n422918 , 
 n422919 , n76454 , n422921 , n422922 , n76457 , n422924 , n422925 , n422926 , n76461 , n422928 , 
 n422929 , n76464 , n422931 , n422932 , n422933 , n76468 , n422935 , n76470 , n76471 , n422938 , 
 n76473 , n422940 , n76475 , n76476 , n422943 , n422944 , n76479 , n422946 , n422947 , n76482 , 
 n422949 , n422950 , n422951 , n76486 , n422953 , n422954 , n76489 , n422956 , n422957 , n76492 , 
 n422959 , n76494 , n422961 , n76496 , n76497 , n76498 , n76499 , n76500 , n76501 , n76502 , 
 n422969 , n76504 , n422971 , n422972 , n76507 , n422974 , n422975 , n422976 , n422977 , n76538 , 
 n422979 , n76540 , n422981 , n76542 , n76543 , n422984 , n76545 , n422986 , n76547 , n76548 , 
 n422989 , n76550 , n422991 , n422992 , n76553 , n422994 , n422995 , n76556 , n422997 , n422998 , 
 n422999 , n76560 , n423001 , n423002 , n423003 , n423004 , n423005 , n76566 , n423007 , n76568 , 
 n423009 , n76570 , n423011 , n423012 , n76573 , n423014 , n423015 , n76576 , n423017 , n423018 , 
 n76579 , n423020 , n76581 , n423022 , n76583 , n76584 , n423025 , n76586 , n423027 , n76588 , 
 n76589 , n423030 , n423031 , n76592 , n423033 , n423034 , n76595 , n423036 , n423037 , n423038 , 
 n76599 , n423040 , n423041 , n76602 , n423043 , n423044 , n76605 , n76606 , n76607 , n76608 , 
 n76609 , n423050 , n76611 , n76612 , n423053 , n423054 , n76615 , n423056 , n423057 , n76618 , 
 n423059 , n76620 , n76621 , n76622 , n76623 , n76624 , n423065 , n423066 , n423067 , n76628 , 
 n423069 , n76630 , n76631 , n423072 , n423073 , n76634 , n423075 , n423076 , n76637 , n423078 , 
 n423079 , n76640 , n76641 , n76642 , n76643 , n76644 , n76645 , n76646 , n76647 , n76648 , 
 n76649 , n76650 , n76651 , n423092 , n76653 , n423094 , n76655 , n76656 , n423097 , n423098 , 
 n76659 , n423100 , n423101 , n76662 , n423103 , n76664 , n423105 , n76666 , n423107 , n76668 , 
 n76669 , n423110 , n423111 , n76672 , n423113 , n423114 , n76675 , n423116 , n76677 , n423118 , 
 n76679 , n423120 , n76681 , n423122 , n423123 , n76684 , n423125 , n76686 , n76687 , n423128 , 
 n76689 , n423130 , n76691 , n76692 , n423133 , n423134 , n76695 , n423136 , n423137 , n76698 , 
 n423139 , n423140 , n423141 , n76702 , n423143 , n423144 , n76705 , n423146 , n423147 , n76708 , 
 n76709 , n76710 , n76711 , n76712 , n423153 , n423154 , n76715 , n423156 , n423157 , n423158 , 
 n76735 , n76736 , n76737 , n76738 , n76739 , n423164 , n423165 , n76742 , n423167 , n423168 , 
 n76745 , n423170 , n423171 , n423172 , n76749 , n423174 , n76751 , n423176 , n423177 , n76754 , 
 n423179 , n76756 , n76757 , n423182 , n76759 , n423184 , n423185 , n76762 , n423187 , n423188 , 
 n76765 , n423190 , n76774 , n76775 , n423193 , n76777 , n423195 , n423196 , n76780 , n423198 , 
 n423199 , n76783 , n76784 , n76785 , n76786 , n423204 , n423205 , n76789 , n423207 , n76791 , 
 n423209 , n76793 , n76794 , n423212 , n76796 , n423214 , n76798 , n76799 , n423217 , n423218 , 
 n76802 , n423220 , n423221 , n76805 , n423223 , n423224 , n423225 , n76809 , n423227 , n423228 , 
 n76812 , n423230 , n423231 , n423232 , n423233 , n76817 , n423235 , n76819 , n423237 , n423238 , 
 n423239 , n423240 , n76824 , n423242 , n423243 , n76827 , n423245 , n423246 , n423247 , n76831 , 
 n423249 , n76833 , n423251 , n76835 , n76836 , n423254 , n423255 , n76839 , n423257 , n423258 , 
 n76842 , n423260 , n423261 , n76845 , n76846 , n423264 , n76848 , n423266 , n76850 , n423268 , 
 n423269 , n76853 , n423271 , n423272 , n423273 , n76857 , n423275 , n76859 , n76860 , n423278 , 
 n423279 , n76863 , n76864 , n423282 , n76866 , n76867 , n423285 , n423286 , n423287 , n76871 , 
 n423289 , n423290 , n76874 , n423292 , n423293 , n76877 , n76878 , n76879 , n76880 , n76881 , 
 n423299 , n423300 , n76884 , n423302 , n423303 , n76887 , n76888 , n76889 , n76890 , n76891 , 
 n423309 , n423310 , n76894 , n423312 , n423313 , n76897 , n423315 , n423316 , n76900 , n423318 , 
 n423319 , n76903 , n76904 , n423322 , n76906 , n76907 , n423325 , n423326 , n423327 , n76911 , 
 n76912 , n423330 , n423331 , n76915 , n423333 , n423334 , n76920 , n76921 , n423337 , n423338 , 
 n76924 , n76925 , n76926 , n76927 , n76928 , n76929 , n76930 , n76931 , n423347 , n76933 , 
 n423349 , n76935 , n76936 , n76937 , n76938 , n423354 , n423355 , n76941 , n423357 , n76943 , 
 n76944 , n76945 , n423361 , n423362 , n76948 , n423364 , n76950 , n423366 , n76952 , n76953 , 
 n423369 , n423370 , n76956 , n423372 , n423373 , n76959 , n423375 , n423376 , n423377 , n76963 , 
 n76964 , n423380 , n76966 , n76967 , n76968 , n76969 , n76970 , n76971 , n76972 , n423388 , 
 n76974 , n423390 , n76976 , n423392 , n423393 , n76979 , n423395 , n423396 , n76982 , n423398 , 
 n423399 , n76985 , n423401 , n423402 , n76988 , n76989 , n423405 , n76991 , n423407 , n423408 , 
 n423409 , n76995 , n423411 , n76997 , n76998 , n423414 , n423415 , n77001 , n423417 , n423418 , 
 n77004 , n423420 , n423421 , n423422 , n423423 , n77035 , n77036 , n77037 , n423427 , n423428 , 
 n77040 , n77042 , n423431 , n423432 , n77045 , n77046 , n423435 , n423436 , n77049 , n77050 , 
 n423439 , n77052 , n423441 , n423442 , n77055 , n77056 , n423445 , n423446 , n423447 , n423448 , 
 n423449 , n77062 , n77063 , n77064 , n77065 , n77066 , n77067 , n423456 , n423457 , n77070 , 
 n423459 , n423460 , n77073 , n423462 , n77075 , n77076 , n77077 , n77078 , n77079 , n423468 , 
 n423469 , n77082 , n423471 , n423472 , n77085 , n423474 , n77087 , n423476 , n423477 , n423478 , 
 n77091 , n423480 , n423481 , n77094 , n77095 , n423484 , n423485 , n77098 , n423487 , n423488 , 
 n77101 , n77102 , n423491 , n77104 , n423493 , n423494 , n77107 , n77108 , n423497 , n77110 , 
 n77111 , n423500 , n423501 , n77114 , n77115 , n423504 , n423505 , n77118 , n423507 , n423508 , 
 n77121 , n423510 , n423511 , n77124 , n77125 , n423514 , n77127 , n423516 , n77129 , n77130 , 
 n77131 , n77132 , n77133 , n77134 , n423523 , n423524 , n77137 , n423526 , n423527 , n77140 , 
 n423529 , n423530 , n77143 , n77144 , n423533 , n423534 , n77147 , n77148 , n77149 , n77150 , 
 n77151 , n423540 , n423541 , n77154 , n423543 , n77156 , n77157 , n423546 , n423547 , n77160 , 
 n423549 , n423550 , n77163 , n423552 , n423553 , n77166 , n423555 , n77168 , n77169 , n423558 , 
 n423559 , n77172 , n423561 , n423562 , n77175 , n423564 , n423565 , n423566 , n423567 , n77180 , 
 n423569 , n77182 , n423571 , n423572 , n77185 , n77186 , n423575 , n77188 , n423577 , n77190 , 
 n423579 , n423580 , n77193 , n423582 , n423583 , n77196 , n423585 , n77198 , n77199 , n423588 , 
 n423589 , n77202 , n423591 , n423592 , n77205 , n423594 , n423595 , n77208 , n77209 , n77210 , 
 n423599 , n423600 , n77213 , n77214 , n77215 , n77216 , n423605 , n77218 , n423607 , n77220 , 
 n77221 , n423610 , n423611 , n77224 , n423613 , n423614 , n77227 , n423616 , n423617 , n77230 , 
 n423619 , n77232 , n423621 , n77234 , n77235 , n423624 , n77237 , n423626 , n77239 , n77240 , 
 n423629 , n423630 , n77243 , n423632 , n423633 , n77246 , n423635 , n423636 , n423637 , n77250 , 
 n423639 , n423640 , n77253 , n423642 , n423643 , n77256 , n77257 , n77258 , n423647 , n423648 , 
 n77261 , n77262 , n77263 , n423652 , n423653 , n77266 , n423655 , n423656 , n423657 , n77270 , 
 n423659 , n423660 , n423661 , n77274 , n423663 , n423664 , n77277 , n423666 , n423667 , n77280 , 
 n423669 , n423670 , n77283 , n423672 , n77285 , n77286 , n77287 , n77297 , n423677 , n77299 , 
 n423679 , n77301 , n77302 , n423682 , n423683 , n77305 , n77306 , n423686 , n423687 , n77309 , 
 n423689 , n77311 , n77312 , n423692 , n423693 , n77315 , n77316 , n423696 , n423697 , n77319 , 
 n423699 , n423700 , n423701 , n423702 , n77352 , n423704 , n77354 , n423706 , n77356 , n423708 , 
 n77358 , n77359 , n423711 , n423712 , n77362 , n77363 , n423715 , n423716 , n77366 , n77367 , 
 n423719 , n423720 , n77370 , n77371 , n423723 , n423724 , n423725 , n77375 , n423727 , n77377 , 
 n77378 , n423730 , n77380 , n423732 , n77382 , n77383 , n423735 , n423736 , n77386 , n423738 , 
 n423739 , n77389 , n423741 , n423742 , n423743 , n77393 , n423745 , n423746 , n77396 , n423748 , 
 n423749 , n77399 , n423751 , n77401 , n423753 , n77403 , n423755 , n77405 , n77406 , n423758 , 
 n423759 , n77409 , n423761 , n423762 , n423763 , n77413 , n77414 , n423766 , n423767 , n77417 , 
 n77418 , n423770 , n423771 , n423772 , n423773 , n423774 , n77424 , n423776 , n423777 , n423778 , 
 n77428 , n77429 , n423781 , n423782 , n77432 , n423784 , n423785 , n423786 , n423787 , n423788 , 
 n77438 , n423790 , n423791 , n423792 , n423793 , n77443 , n423795 , n423796 , n423797 , n423798 , 
 n77448 , n423800 , n423801 , n423802 , n77452 , n423804 , n423805 , n423806 , n423807 , n77457 , 
 n423809 , n423810 , n423811 , n423812 , n423813 , n77463 , n77464 , n423816 , n423817 , n423818 , 
 n77468 , n77469 , n423821 , n423822 , n77472 , n423824 , n423825 , n423826 , n423827 , n423828 , 
 n423829 , n77479 , n423831 , n423832 , n77482 , n423834 , n423835 , n423836 , n423837 , n77487 , 
 n423839 , n77489 , n423841 , n423842 , n77492 , n423844 , n77494 , n423846 , n423847 , n423848 , 
 n77498 , n423850 , n423851 , n423852 , n423853 , n423854 , n423855 , n423856 , n423857 , n423858 , 
 n77508 , n423860 , n423861 , n423862 , n77512 , n77513 , n77514 , n423866 , n423867 , n423868 , 
 n423869 , n77519 , n423871 , n423872 , n77522 , n77523 , n423875 , n423876 , n423877 , n77527 , 
 n423879 , n423880 , n423881 , n423882 , n423883 , n77533 , n77534 , n423886 , n423887 , n77537 , 
 n423889 , n423890 , n423891 , n423892 , n423893 , n423894 , n77544 , n423896 , n423897 , n423898 , 
 n423899 , n77549 , n423901 , n423902 , n77552 , n77553 , n423905 , n423906 , n423907 , n77557 , 
 n423909 , n77559 , n423911 , n423912 , n423913 , n77563 , n423915 , n423916 , n423917 , n77567 , 
 n423919 , n423920 , n423921 , n423922 , n423923 , n423924 , n77574 , n423926 , n423927 , n77577 , 
 n77578 , n77579 , n423931 , n423932 , n77582 , n77583 , n77584 , n423936 , n423937 , n77587 , 
 n77588 , n77589 , n423941 , n423942 , n423943 , n423944 , n77594 , n423946 , n423947 , n77597 , 
 n77598 , n423950 , n423951 , n423952 , n423953 , n423954 , n77604 , n423956 , n423957 , n423958 , 
 n423959 , n77609 , n423961 , n423962 , n423963 , n423964 , n423965 , n423966 , n423967 , n77617 , 
 n423969 , n423970 , n423971 , n423972 , n423973 , n77623 , n423975 , n423976 , n423977 , n77627 , 
 n423979 , n423980 , n423981 , n423982 , n423983 , n423984 , n77634 , n423986 , n423987 , n77637 , 
 n77638 , n423990 , n423991 , n423992 , n77642 , n423994 , n77644 , n423996 , n423997 , n77647 , 
 n423999 , n77649 , n424001 , n424002 , n77652 , n424004 , n424005 , n424006 , n424007 , n424008 , 
 n424009 , n77659 , n424011 , n424012 , n77662 , n77663 , n424015 , n424016 , n424017 , n77667 , 
 n424019 , n424020 , n424021 , n424022 , n77672 , n424024 , n77674 , n424026 , n424027 , n424028 , 
 n77678 , n424030 , n424031 , n424032 , n77682 , n424034 , n424035 , n424036 , n424037 , n424038 , 
 n77688 , n77689 , n424041 , n424042 , n424043 , n77693 , n77694 , n424046 , n424047 , n77697 , 
 n77698 , n424050 , n424051 , n424052 , n77702 , n424054 , n424055 , n424056 , n424057 , n424058 , 
 n424059 , n424060 , n424061 , n424062 , n424063 , n77713 , n77714 , n424066 , n424067 , n77717 , 
 n77718 , n77719 , n424071 , n424072 , n77722 , n77723 , n77724 , n424076 , n424077 , n77727 , 
 n77728 , n77729 , n424081 , n424082 , n77732 , n77733 , n77734 , n424086 , n424087 , n77737 , 
 n424089 , n424090 , n424091 , n424092 , n424093 , n424094 , n77744 , n424096 , n424097 , n424098 , 
 n424099 , n77749 , n424101 , n424102 , n424103 , n424104 , n77754 , n424106 , n424107 , n77757 , 
 n77758 , n424110 , n424111 , n424112 , n424113 , n424114 , n77764 , n424116 , n424117 , n77767 , 
 n424119 , n424120 , n424121 , n424122 , n424123 , n424124 , n424125 , n424126 , n424127 , n424128 , 
 n77778 , n77779 , n424131 , n424132 , n77782 , n424134 , n77784 , n424136 , n424137 , n424138 , 
 n77788 , n77789 , n424141 , n424142 , n77792 , n424144 , n77794 , n424146 , n424147 , n77797 , 
 n77798 , n424150 , n424151 , n424152 , n77802 , n424154 , n77804 , n424156 , n424157 , n424158 , 
 n77808 , n424160 , n424161 , n424162 , n77812 , n424164 , n424165 , n424166 , n424167 , n77817 , 
 n424169 , n77819 , n424171 , n424172 , n77822 , n77823 , n77824 , n424176 , n424177 , n424178 , 
 n77828 , n424180 , n424181 , n424182 , n77832 , n424184 , n424185 , n424186 , n424187 , n424188 , 
 n77838 , n77839 , n424191 , n424192 , n424193 , n77843 , n77844 , n424196 , n424197 , n77847 , 
 n77848 , n77849 , n424201 , n424202 , n77852 , n77853 , n424205 , n424206 , n424207 , n77857 , 
 n424209 , n77859 , n424211 , n424212 , n424213 , n77863 , n77864 , n424216 , n424217 , n77867 , 
 n424219 , n77869 , n424221 , n424222 , n424223 , n77873 , n77874 , n424226 , n424227 , n77877 , 
 n424229 , n77879 , n424231 , n424232 , n424233 , n424234 , n77884 , n424236 , n424237 , n77887 , 
 n424239 , n424240 , n424241 , n424242 , n424243 , n77893 , n77894 , n424246 , n424247 , n424248 , 
 n77898 , n77899 , n424251 , n424252 , n424253 , n77903 , n424255 , n424256 , n424257 , n424258 , 
 n424259 , n77909 , n424261 , n424262 , n424263 , n77913 , n77914 , n424266 , n424267 , n77917 , 
 n424269 , n424270 , n424271 , n424272 , n424273 , n77923 , n424275 , n424276 , n424277 , n424278 , 
 n424279 , n77929 , n424281 , n424282 , n77932 , n424284 , n424285 , n424286 , n424287 , n77937 , 
 n424289 , n424290 , n424291 , n424292 , n424293 , n77943 , n424295 , n424296 , n424297 , n77947 , 
 n77948 , n424300 , n424301 , n424302 , n424303 , n424304 , n77954 , n424306 , n424307 , n424308 , 
 n424309 , n424310 , n424311 , n424312 , n77963 , n424314 , n424315 , n424316 , n77967 , n424318 , 
 n77969 , n424320 , n424321 , n424322 , n424323 , n77974 , n424325 , n424326 , n77977 , n424328 , 
 n424329 , n424330 , n424331 , n424332 , n77983 , n424334 , n424335 , n424336 , n424337 , n77988 , 
 n77989 , n424340 , n424341 , n77992 , n424343 , n424344 , n424345 , n424346 , n424347 , n77998 , 
 n424349 , n424350 , n424351 , n78002 , n78003 , n424354 , n424355 , n424356 , n78007 , n78008 , 
 n424359 , n424360 , n424361 , n424362 , n424363 , n78014 , n424365 , n424366 , n424367 , n78018 , 
 n424369 , n424370 , n424371 , n424372 , n424373 , n78024 , n424375 , n424376 , n78027 , n424378 , 
 n78029 , n424380 , n424381 , n78032 , n78033 , n78034 , n424385 , n424386 , n424387 , n78038 , 
 n424389 , n424390 , n424391 , n424392 , n78043 , n424394 , n78059 , n78060 , n424397 , n424398 , 
 n424399 , n78064 , n78066 , n78067 , n78068 , n424404 , n78070 , n78071 , n78072 , n78073 , 
 n424409 , n78075 , n78076 , n424412 , n424413 , n78079 , n424415 , n78081 , n424417 , n78083 , 
 n424419 , n78085 , n424421 , n78087 , n78088 , n424424 , n424425 , n78091 , n424427 , n424428 , 
 n78094 , n424430 , n424431 , n424432 , n424433 , n78099 , n78100 , n424436 , n424437 , n78103 , 
 n424439 , n424440 , n78106 , n424442 , n424443 , n424444 , n424445 , n78111 , n78112 , n424448 , 
 n78114 , n424450 , n424451 , n424452 , n78118 , n424454 , n424455 , n78121 , n424457 , n424458 , 
 n78124 , n424460 , n424461 , n78127 , n424463 , n424464 , n424465 , n424466 , n78132 , n424468 , 
 n424469 , n78135 , n78136 , n424472 , n424473 , n424474 , n78140 , n424476 , n424477 , n78143 , 
 n78144 , n424480 , n78146 , n78147 , n78148 , n424484 , n424485 , n78151 , n424487 , n78153 , 
 n424489 , n424490 , n424491 , n424492 , n424493 , n78159 , n424495 , n424496 , n78162 , n78163 , 
 n424499 , n424500 , n424501 , n424502 , n424503 , n78169 , n78170 , n424506 , n424507 , n78173 , 
 n424509 , n424510 , n78176 , n424512 , n424513 , n78179 , n78180 , n424516 , n424517 , n78183 , 
 n424519 , n424520 , n78186 , n424522 , n78188 , n78189 , n424525 , n424526 , n78192 , n78193 , 
 n424529 , n424530 , n78196 , n78197 , n78198 , n424534 , n78200 , n78201 , n78202 , n78203 , 
 n78204 , n424540 , n424541 , n424542 , n78208 , n424544 , n424545 , n78211 , n78212 , n424548 , 
 n424549 , n424550 , n78216 , n424552 , n424553 , n78219 , n78220 , n424556 , n424557 , n78223 , 
 n78224 , n78225 , n424561 , n424562 , n78228 , n78229 , n78230 , n424566 , n78232 , n78233 , 
 n424569 , n424570 , n424571 , n78237 , n424573 , n424574 , n78240 , n78241 , n424577 , n424578 , 
 n424579 , n78245 , n424581 , n424582 , n78248 , n78249 , n424585 , n424586 , n78252 , n78253 , 
 n424589 , n424590 , n78256 , n424592 , n424593 , n78259 , n424595 , n424596 , n424597 , n424598 , 
 n78264 , n424600 , n424601 , n78267 , n78268 , n424604 , n78270 , n78271 , n78272 , n424608 , 
 n78274 , n424610 , n424611 , n78277 , n424613 , n424614 , n78280 , n78281 , n424617 , n78283 , 
 n424619 , n78285 , n78286 , n424622 , n424623 , n78289 , n78290 , n424626 , n78292 , n78293 , 
 n78294 , n78295 , n78296 , n78297 , n78298 , n78299 , n78300 , n78301 , n78302 , n78303 , 
 n78304 , n78305 , n78306 , n78307 , n78308 , n78309 , n78310 , n78311 , n424647 , n424648 , 
 n424649 , n78315 , n424651 , n424652 , n78318 , n78319 , n424655 , n424656 , n424657 , n78323 , 
 n424659 , n424660 , n78326 , n78327 , n424663 , n424664 , n424665 , n424666 , n424667 , n78333 , 
 n424669 , n424670 , n78336 , n78337 , n424673 , n424674 , n78340 , n424676 , n424677 , n78343 , 
 n424679 , n424680 , n424681 , n424682 , n78348 , n424684 , n424685 , n78351 , n424687 , n78353 , 
 n424689 , n424690 , n424691 , n78357 , n424693 , n78359 , n424695 , n424696 , n424697 , n78363 , 
 n424699 , n424700 , n78366 , n78367 , n424703 , n424704 , n78370 , n424706 , n424707 , n78373 , 
 n78374 , n424710 , n78376 , n78377 , n78378 , n424714 , n78380 , n424716 , n424717 , n78383 , 
 n424719 , n78385 , n424721 , n424722 , n78388 , n424724 , n424725 , n78391 , n78392 , n424728 , 
 n424729 , n78395 , n78396 , n424732 , n424733 , n78399 , n78400 , n424736 , n424737 , n78403 , 
 n78404 , n78405 , n424741 , n424742 , n78408 , n78409 , n78410 , n78411 , n78412 , n424748 , 
 n78414 , n78415 , n78416 , n424752 , n78418 , n78419 , n78420 , n78421 , n78422 , n78423 , 
 n78424 , n78425 , n424761 , n78427 , n78428 , n78429 , n78430 , n424766 , n78432 , n78433 , 
 n78434 , n78435 , n78436 , n424772 , n78438 , n424774 , n78440 , n424776 , n78442 , n78443 , 
 n78444 , n78445 , n78446 , n78447 , n424783 , n78449 , n424785 , n78451 , n78452 , n424788 , 
 n424789 , n78455 , n424791 , n424792 , n78458 , n424794 , n424795 , n78461 , n424797 , n78463 , 
 n78464 , n424800 , n78466 , n424802 , n78468 , n78469 , n424805 , n424806 , n78472 , n424808 , 
 n424809 , n78475 , n424811 , n424812 , n78478 , n424814 , n424815 , n424816 , n78482 , n424818 , 
 n424819 , n78485 , n424821 , n78487 , n78488 , n424824 , n424825 , n78491 , n78492 , n78493 , 
 n424829 , n424830 , n78496 , n424832 , n78498 , n78499 , n78500 , n78501 , n78502 , n78503 , 
 n424839 , n78505 , n424841 , n424842 , n424843 , n78509 , n424845 , n78511 , n424847 , n78513 , 
 n424849 , n424850 , n78516 , n424852 , n424853 , n78519 , n78520 , n424856 , n78522 , n424858 , 
 n78524 , n424860 , n78526 , n424862 , n78528 , n424864 , n78530 , n424866 , n78532 , n78533 , 
 n424869 , n424870 , n78536 , n424872 , n424873 , n78539 , n424875 , n424876 , n78542 , n424878 , 
 n78544 , n78545 , n424881 , n424882 , n78548 , n424884 , n424885 , n78551 , n424887 , n424888 , 
 n78554 , n78555 , n78556 , n424892 , n424893 , n78559 , n424895 , n78561 , n424897 , n78563 , 
 n78564 , n424900 , n424901 , n78567 , n78568 , n424904 , n78570 , n78571 , n424907 , n424908 , 
 n424909 , n78575 , n424911 , n424912 , n78578 , n424914 , n424915 , n78581 , n78582 , n78583 , 
 n424919 , n424920 , n424921 , n78587 , n424923 , n78589 , n78590 , n424926 , n78592 , n424928 , 
 n424929 , n424930 , n424931 , n424932 , n78598 , n424934 , n424935 , n78601 , n424937 , n424938 , 
 n78604 , n78605 , n78606 , n424942 , n424943 , n78609 , n78610 , n78611 , n424947 , n424948 , 
 n78614 , n78615 , n424951 , n424952 , n78618 , n424954 , n78620 , n424956 , n78622 , n78623 , 
 n424959 , n78625 , n424961 , n78627 , n424963 , n424964 , n424965 , n78631 , n424967 , n424968 , 
 n78634 , n424970 , n424971 , n424972 , n78638 , n424974 , n424975 , n78641 , n424977 , n424978 , 
 n78644 , n78645 , n78646 , n424982 , n424983 , n424984 , n424985 , n78651 , n78652 , n424988 , 
 n78654 , n78655 , n424991 , n78657 , n424993 , n78659 , n424995 , n424996 , n78662 , n424998 , 
 n424999 , n78665 , n425001 , n78667 , n78668 , n78669 , n78670 , n78671 , n78672 , n425008 , 
 n425009 , n78675 , n425011 , n425012 , n78678 , n425014 , n425015 , n78681 , n425017 , n425018 , 
 n425019 , n78685 , n78686 , n425022 , n78688 , n78689 , n425025 , n425026 , n78692 , n425028 , 
 n425029 , n78695 , n78696 , n425032 , n425033 , n78699 , n78700 , n78701 , n425037 , n425038 , 
 n78704 , n425040 , n425041 , n78707 , n425043 , n425044 , n78710 , n425046 , n425047 , n78713 , 
 n425049 , n425050 , n78716 , n425052 , n78718 , n78719 , n78720 , n78721 , n78722 , n78723 , 
 n78724 , n425060 , n425061 , n425062 , n78728 , n425064 , n425065 , n78731 , n425067 , n78733 , 
 n78734 , n425070 , n425071 , n78737 , n78738 , n425074 , n425075 , n425076 , n78742 , n425078 , 
 n78744 , n78745 , n425081 , n78747 , n425083 , n78749 , n78750 , n425086 , n425087 , n78753 , 
 n425089 , n425090 , n78756 , n425092 , n425093 , n425094 , n78760 , n425096 , n425097 , n78763 , 
 n425099 , n425100 , n78766 , n425102 , n78768 , n425104 , n78770 , n78771 , n425107 , n425108 , 
 n78774 , n425110 , n425111 , n78777 , n425113 , n425114 , n78780 , n425116 , n78782 , n78783 , 
 n425119 , n425120 , n78786 , n425122 , n425123 , n78789 , n425125 , n425126 , n425127 , n78793 , 
 n425129 , n78795 , n78796 , n425132 , n78798 , n425134 , n78800 , n78801 , n425137 , n425138 , 
 n78804 , n425140 , n425141 , n78807 , n425143 , n425144 , n425145 , n78811 , n425147 , n425148 , 
 n78814 , n425150 , n425151 , n78817 , n425153 , n78819 , n425155 , n78821 , n78822 , n425158 , 
 n425159 , n78825 , n425161 , n425162 , n78828 , n425164 , n425165 , n78831 , n425167 , n78833 , 
 n78834 , n425170 , n425171 , n78837 , n425173 , n425174 , n78840 , n425176 , n425177 , n78843 , 
 n78844 , n78845 , n425181 , n425182 , n78848 , n78849 , n78850 , n425186 , n425187 , n78853 , 
 n425189 , n425190 , n425191 , n78857 , n78858 , n425194 , n78860 , n78861 , n425197 , n425198 , 
 n78864 , n425200 , n78866 , n425202 , n425203 , n425204 , n78870 , n78871 , n425207 , n425208 , 
 n78874 , n78875 , n78876 , n425212 , n78878 , n425214 , n425215 , n78881 , n425217 , n78883 , 
 n425219 , n78885 , n78886 , n425222 , n425223 , n78889 , n425225 , n425226 , n78892 , n425228 , 
 n425229 , n78895 , n425231 , n78897 , n425233 , n425234 , n78900 , n425236 , n425237 , n425238 , 
 n78904 , n425240 , n78906 , n78907 , n425243 , n425244 , n425245 , n425246 , n425247 , n78913 , 
 n425249 , n78915 , n78916 , n78917 , n425253 , n425254 , n78920 , n425256 , n78922 , n78923 , 
 n425259 , n78925 , n425261 , n78927 , n78928 , n78929 , n78930 , n78931 , n78932 , n78933 , 
 n78934 , n78935 , n78936 , n78937 , n78938 , n425274 , n425275 , n425276 , n78942 , n425278 , 
 n78944 , n78945 , n425281 , n78947 , n425283 , n78949 , n425285 , n425286 , n78952 , n78953 , 
 n425289 , n425290 , n78956 , n425292 , n425293 , n78959 , n425295 , n425296 , n425297 , n78963 , 
 n425299 , n425300 , n78966 , n425302 , n425303 , n78969 , n425305 , n425306 , n78972 , n425308 , 
 n78974 , n425310 , n78976 , n425312 , n425313 , n78979 , n78980 , n78981 , n78982 , n425318 , 
 n425319 , n78985 , n425321 , n425322 , n425323 , n78989 , n425325 , n425326 , n425327 , n78993 , 
 n425329 , n425330 , n78996 , n425332 , n425333 , n78999 , n79000 , n79001 , n425337 , n425338 , 
 n79004 , n79005 , n79006 , n425342 , n79008 , n79009 , n425345 , n79011 , n79012 , n425348 , 
 n425349 , n425350 , n425351 , n79040 , n79041 , n425354 , n79043 , n425356 , n79045 , n425358 , 
 n425359 , n425360 , n79049 , n425362 , n425363 , n79052 , n425365 , n79054 , n425367 , n79056 , 
 n425369 , n425370 , n425371 , n79060 , n425373 , n79062 , n425375 , n79064 , n79065 , n79066 , 
 n425379 , n79068 , n79069 , n425382 , n425383 , n79072 , n79073 , n79074 , n425387 , n425388 , 
 n79077 , n79078 , n79079 , n425392 , n425393 , n79082 , n79083 , n79084 , n79085 , n425398 , 
 n425399 , n425400 , n79089 , n425402 , n79091 , n425404 , n425405 , n79094 , n425407 , n425408 , 
 n79097 , n425410 , n425411 , n79100 , n425413 , n425414 , n79103 , n425416 , n425417 , n79106 , 
 n425419 , n425420 , n425421 , n425422 , n425423 , n425424 , n79130 , n425426 , n79132 , n425428 , 
 n425429 , n79135 , n425431 , n425432 , n79138 , n79139 , n425435 , n425436 , n425437 , n425438 , 
 n79166 , n425440 , n425441 , n425442 , n79170 , n79171 , n425445 , n79173 , n79174 , n425448 , 
 n425449 , n79177 , n425451 , n425452 , n79180 , n79181 , n425455 , n425456 , n425457 , n79185 , 
 n425459 , n79187 , n79188 , n425462 , n79190 , n425464 , n79192 , n79193 , n425467 , n425468 , 
 n79196 , n425470 , n425471 , n79199 , n425473 , n425474 , n425475 , n79203 , n425477 , n425478 , 
 n79206 , n425480 , n425481 , n79209 , n79210 , n425484 , n425485 , n79213 , n79214 , n79215 , 
 n79216 , n79217 , n79218 , n79219 , n79220 , n425494 , n425495 , n79223 , n425497 , n79225 , 
 n79226 , n425500 , n79228 , n425502 , n79230 , n79231 , n425505 , n425506 , n79234 , n425508 , 
 n425509 , n79237 , n425511 , n425512 , n425513 , n79241 , n425515 , n425516 , n79244 , n425518 , 
 n425519 , n79247 , n425521 , n79249 , n425523 , n79251 , n425525 , n425526 , n79254 , n79255 , 
 n425529 , n425530 , n79258 , n425532 , n425533 , n79261 , n425535 , n425536 , n79264 , n425538 , 
 n79266 , n79267 , n425541 , n425542 , n79270 , n425544 , n425545 , n79273 , n425547 , n425548 , 
 n79276 , n79277 , n79278 , n425552 , n79280 , n425554 , n79282 , n425556 , n79284 , n79285 , 
 n425559 , n425560 , n79288 , n79289 , n425563 , n79291 , n79292 , n425566 , n425567 , n425568 , 
 n79296 , n425570 , n425571 , n79299 , n425573 , n79301 , n79302 , n79303 , n425577 , n79305 , 
 n79306 , n79307 , n425581 , n425582 , n79310 , n79311 , n425585 , n425586 , n425587 , n425588 , 
 n79316 , n79317 , n425591 , n79319 , n79320 , n425594 , n425595 , n79323 , n425597 , n79325 , 
 n79326 , n425600 , n425601 , n79329 , n425603 , n425604 , n79332 , n425606 , n425607 , n79335 , 
 n425609 , n79337 , n79338 , n79339 , n425613 , n425614 , n79342 , n425616 , n79344 , n79345 , 
 n425619 , n79347 , n425621 , n425622 , n79350 , n79351 , n79352 , n425626 , n425627 , n79355 , 
 n425629 , n425630 , n79358 , n425632 , n79360 , n79361 , n425635 , n425636 , n79364 , n425638 , 
 n425639 , n79367 , n425641 , n425642 , n79370 , n425644 , n425645 , n79373 , n425647 , n79375 , 
 n425649 , n425650 , n425651 , n79379 , n79380 , n425654 , n425655 , n79383 , n79384 , n79385 , 
 n425659 , n425660 , n79388 , n425662 , n79390 , n425664 , n79392 , n79393 , n425667 , n79395 , 
 n425669 , n79397 , n79398 , n425672 , n425673 , n79401 , n425675 , n425676 , n79404 , n425678 , 
 n425679 , n425680 , n79408 , n425682 , n425683 , n79411 , n425685 , n425686 , n79414 , n79415 , 
 n79416 , n425690 , n425691 , n79419 , n79421 , n425694 , n425695 , n79424 , n425697 , n425698 , 
 n79430 , n425700 , n79432 , n79433 , n79434 , n425704 , n79436 , n79437 , n79438 , n79439 , 
 n79440 , n79441 , n79442 , n79443 , n425713 , n425714 , n79446 , n79447 , n425717 , n79449 , 
 n79450 , n425720 , n79452 , n79453 , n79454 , n79455 , n79456 , n79457 , n79458 , n425728 , 
 n79460 , n425730 , n79462 , n79463 , n79464 , n425734 , n79466 , n425736 , n425737 , n425738 , 
 n79470 , n425740 , n79472 , n79473 , n425743 , n425744 , n79476 , n425746 , n425747 , n79479 , 
 n425749 , n425750 , n425751 , n79483 , n425753 , n425754 , n79486 , n425756 , n79488 , n79489 , 
 n79490 , n79491 , n79492 , n79493 , n79494 , n425764 , n425765 , n79497 , n425767 , n79499 , 
 n425769 , n79501 , n79502 , n79503 , n425773 , n425774 , n79506 , n79507 , n79508 , n79509 , 
 n79510 , n79511 , n79512 , n79513 , n79514 , n79515 , n425785 , n425786 , n425787 , n79533 , 
 n79534 , n425790 , n79536 , n79537 , n79538 , n79539 , n79540 , n79541 , n79542 , n79543 , 
 n79544 , n425800 , n79546 , n79547 , n79548 , n425804 , n425805 , n79551 , n425807 , n79553 , 
 n425809 , n425810 , n79556 , n425812 , n425813 , n79559 , n425815 , n425816 , n79562 , n425818 , 
 n425819 , n79565 , n79566 , n79567 , n79568 , n79569 , n79570 , n79571 , n79572 , n79573 , 
 n79574 , n79575 , n79576 , n79577 , n79578 , n79579 , n79580 , n79581 , n79582 , n425838 , 
 n425839 , n79585 , n79586 , n425842 , n79588 , n79589 , n425845 , n425846 , n79592 , n79593 , 
 n425849 , n425850 , n425851 , n79597 , n425853 , n79599 , n79600 , n425856 , n79602 , n425858 , 
 n79604 , n79605 , n425861 , n425862 , n79608 , n425864 , n425865 , n79611 , n425867 , n425868 , 
 n425869 , n79615 , n425871 , n425872 , n79618 , n425874 , n425875 , n79621 , n79622 , n79623 , 
 n425879 , n425880 , n425881 , n79627 , n425883 , n79629 , n79630 , n425886 , n425887 , n79633 , 
 n425889 , n425890 , n79636 , n425892 , n425893 , n79639 , n425895 , n79641 , n79642 , n425898 , 
 n425899 , n79645 , n425901 , n425902 , n79648 , n425904 , n425905 , n79651 , n79652 , n79653 , 
 n79654 , n79655 , n425911 , n425912 , n79658 , n425914 , n79660 , n79661 , n425917 , n425918 , 
 n79664 , n425920 , n425921 , n79667 , n425923 , n425924 , n79670 , n425926 , n79672 , n79673 , 
 n425929 , n425930 , n79676 , n425932 , n425933 , n79679 , n425935 , n425936 , n79682 , n425938 , 
 n79684 , n425940 , n79686 , n79687 , n425943 , n79689 , n425945 , n79691 , n79692 , n425948 , 
 n425949 , n79695 , n425951 , n425952 , n79698 , n425954 , n425955 , n425956 , n79702 , n425958 , 
 n425959 , n79705 , n425961 , n425962 , n79708 , n79709 , n79710 , n425966 , n425967 , n425968 , 
 n79714 , n425970 , n79716 , n79717 , n425973 , n425974 , n79720 , n425976 , n425977 , n79723 , 
 n425979 , n425980 , n79726 , n425982 , n79728 , n79729 , n425985 , n425986 , n79732 , n425988 , 
 n425989 , n79735 , n425991 , n425992 , n79738 , n79739 , n79740 , n425996 , n425997 , n79743 , 
 n79744 , n79745 , n426001 , n426002 , n79748 , n79749 , n79750 , n426006 , n426007 , n426008 , 
 n79754 , n426010 , n79756 , n79757 , n426013 , n426014 , n79760 , n426016 , n426017 , n79763 , 
 n426019 , n426020 , n79766 , n426022 , n79768 , n79769 , n426025 , n79771 , n426027 , n79773 , 
 n426029 , n426030 , n79776 , n426032 , n426033 , n79779 , n79780 , n79781 , n426037 , n426038 , 
 n79784 , n79785 , n79786 , n426042 , n426043 , n79789 , n79790 , n79791 , n426047 , n426048 , 
 n426049 , n426050 , n79821 , n79822 , n426053 , n79824 , n79825 , n79826 , n79827 , n79828 , 
 n426059 , n426060 , n79831 , n426062 , n426063 , n79834 , n79835 , n426066 , n79837 , n79838 , 
 n426069 , n426070 , n426071 , n426072 , n79862 , n426074 , n79864 , n426076 , n79866 , n426078 , 
 n426079 , n426080 , n79870 , n426082 , n79872 , n79873 , n426085 , n426086 , n79876 , n426088 , 
 n426089 , n79879 , n426091 , n426092 , n79882 , n426094 , n79884 , n79885 , n426097 , n426098 , 
 n79888 , n426100 , n426101 , n79891 , n426103 , n426104 , n79894 , n79895 , n79896 , n79897 , 
 n426109 , n79899 , n79900 , n79901 , n79902 , n79903 , n79904 , n79905 , n79906 , n79907 , 
 n79908 , n79909 , n426121 , n426122 , n79912 , n426124 , n426125 , n426126 , n426127 , n426128 , 
 n79918 , n426130 , n426131 , n79921 , n79922 , n426134 , n426135 , n79925 , n426137 , n426138 , 
 n79928 , n79929 , n426141 , n426142 , n79932 , n426144 , n426145 , n426146 , n426147 , n79937 , 
 n426149 , n426150 , n79940 , n79941 , n426153 , n426154 , n79944 , n426156 , n79946 , n426158 , 
 n426159 , n426160 , n79950 , n79951 , n426163 , n79953 , n426165 , n426166 , n79956 , n426168 , 
 n426169 , n426170 , n79960 , n426172 , n79962 , n426174 , n426175 , n79965 , n426177 , n79967 , 
 n79968 , n79969 , n79970 , n79971 , n79972 , n426184 , n79974 , n79975 , n79976 , n426188 , 
 n79978 , n426190 , n426191 , n79981 , n426193 , n426194 , n79984 , n79985 , n426197 , n426198 , 
 n426199 , n79989 , n426201 , n79991 , n426203 , n426204 , n426205 , n79995 , n79996 , n426208 , 
 n79998 , n79999 , n80000 , n426212 , n426213 , n80003 , n426215 , n426216 , n80006 , n80007 , 
 n426219 , n426220 , n426221 , n80011 , n426223 , n426224 , n80014 , n80015 , n426227 , n426228 , 
 n426229 , n426230 , n80020 , n426232 , n426233 , n80023 , n80024 , n426236 , n426237 , n426238 , 
 n80028 , n426240 , n426241 , n80031 , n80032 , n426244 , n426245 , n80035 , n426247 , n426248 , 
 n80038 , n426250 , n80040 , n426252 , n426253 , n80043 , n80044 , n80045 , n426257 , n80047 , 
 n80048 , n426260 , n426261 , n80051 , n426263 , n426264 , n426265 , n426266 , n426267 , n426268 , 
 n426269 , n426270 , n426271 , n426272 , n426273 , n80063 , n426275 , n426276 , n80066 , n426278 , 
 n426279 , n426280 , n426281 , n426282 , n80072 , n426284 , n426285 , n80075 , n426287 , n426288 , 
 n426289 , n426290 , n426291 , n80081 , n426293 , n426294 , n80084 , n426296 , n426297 , n426298 , 
 n426299 , n426300 , n426301 , n426302 , n426303 , n80093 , n426305 , n426306 , n80096 , n426308 , 
 n426309 , n80099 , n80100 , n426312 , n426313 , n80103 , n426315 , n426316 , n80106 , n80107 , 
 n426319 , n426320 , n426321 , n80111 , n426323 , n426324 , n80114 , n80115 , n426327 , n80117 , 
 n80118 , n80119 , n80120 , n80121 , n80122 , n80123 , n80124 , n80125 , n80126 , n426338 , 
 n80128 , n80129 , n80130 , n80131 , n80132 , n426344 , n80134 , n80135 , n426347 , n426348 , 
 n80138 , n80139 , n80140 , n426352 , n426353 , n80143 , n80144 , n426356 , n426357 , n80147 , 
 n80148 , n80149 , n426361 , n426362 , n426363 , n80153 , n80154 , n426366 , n426367 , n80157 , 
 n80158 , n426370 , n426371 , n80161 , n426373 , n426374 , n80164 , n426376 , n426377 , n80167 , 
 n426379 , n80169 , n80170 , n80171 , n80172 , n426384 , n426385 , n80175 , n426387 , n80177 , 
 n426389 , n426390 , n80180 , n80181 , n426393 , n426394 , n426395 , n80185 , n80186 , n426398 , 
 n426399 , n80189 , n426401 , n426402 , n426403 , n426404 , n80194 , n426406 , n426407 , n80197 , 
 n426409 , n426410 , n426411 , n80201 , n426413 , n80203 , n80204 , n426416 , n426417 , n80207 , 
 n426419 , n80209 , n426421 , n426422 , n426423 , n80213 , n426425 , n426426 , n80216 , n426428 , 
 n426429 , n80219 , n426431 , n426432 , n80222 , n426434 , n426435 , n80225 , n426437 , n80227 , 
 n80228 , n80229 , n80230 , n426442 , n426443 , n80233 , n426445 , n80235 , n80236 , n426448 , 
 n80238 , n426450 , n426451 , n80241 , n426453 , n426454 , n426455 , n426456 , n80246 , n80247 , 
 n80248 , n426460 , n80250 , n80251 , n80252 , n426464 , n426465 , n426466 , n426467 , n80257 , 
 n426469 , n426470 , n80260 , n80261 , n426473 , n426474 , n80264 , n426476 , n80266 , n80267 , 
 n426479 , n426480 , n80270 , n426482 , n426483 , n80273 , n426485 , n426486 , n80276 , n426488 , 
 n80278 , n426490 , n80280 , n80281 , n80282 , n80283 , n80284 , n80285 , n426497 , n426498 , 
 n80288 , n426500 , n426501 , n80291 , n426503 , n426504 , n80294 , n80295 , n80296 , n426508 , 
 n426509 , n80299 , n80301 , n426512 , n426513 , n426514 , n426515 , n80326 , n80327 , n426518 , 
 n426519 , n80330 , n80331 , n80332 , n426523 , n426524 , n80335 , n80336 , n426527 , n80338 , 
 n80339 , n80340 , n80341 , n80342 , n80343 , n80344 , n80345 , n426536 , n426537 , n80348 , 
 n80349 , n80350 , n426541 , n426542 , n80353 , n80354 , n80355 , n426546 , n80357 , n426548 , 
 n426549 , n80360 , n426551 , n426552 , n80363 , n426554 , n426555 , n80366 , n426557 , n80368 , 
 n80369 , n426560 , n80371 , n426562 , n426563 , n426564 , n80375 , n426566 , n426567 , n80378 , 
 n426569 , n80380 , n426571 , n426572 , n80383 , n426574 , n80385 , n80386 , n426577 , n426578 , 
 n80389 , n426580 , n80391 , n426582 , n426583 , n80394 , n426585 , n80396 , n80397 , n426588 , 
 n426589 , n80400 , n426591 , n80402 , n80403 , n80404 , n80405 , n426596 , n80407 , n80408 , 
 n426599 , n426600 , n80411 , n80412 , n426603 , n426604 , n80415 , n426606 , n80417 , n426608 , 
 n80419 , n80420 , n426611 , n80422 , n426613 , n80424 , n80425 , n426616 , n80427 , n426618 , 
 n426619 , n80430 , n426621 , n426622 , n80433 , n426624 , n426625 , n80436 , n426627 , n426628 , 
 n80439 , n80440 , n426631 , n80442 , n80443 , n426634 , n80445 , n80446 , n80447 , n80448 , 
 n426639 , n80450 , n80451 , n426642 , n426643 , n80454 , n426645 , n80456 , n426647 , n426648 , 
 n80459 , n80460 , n426651 , n80462 , n80463 , n80464 , n426655 , n426656 , n80467 , n80468 , 
 n426659 , n426660 , n426661 , n80472 , n426663 , n426664 , n426665 , n80476 , n426667 , n80478 , 
 n80479 , n426670 , n426671 , n80482 , n426673 , n426674 , n80485 , n426676 , n426677 , n80488 , 
 n426679 , n80490 , n80491 , n426682 , n426683 , n80494 , n426685 , n426686 , n80497 , n426688 , 
 n426689 , n426690 , n80501 , n426692 , n80503 , n80504 , n80505 , n80506 , n80507 , n80508 , 
 n426699 , n426700 , n80511 , n426702 , n426703 , n80514 , n426705 , n426706 , n80517 , n426708 , 
 n426709 , n80520 , n80521 , n426712 , n80523 , n426714 , n426715 , n426716 , n80527 , n426718 , 
 n80529 , n80530 , n426721 , n426722 , n80533 , n426724 , n426725 , n80536 , n426727 , n426728 , 
 n426729 , n80540 , n426731 , n80542 , n80543 , n426734 , n80545 , n426736 , n80547 , n80548 , 
 n426739 , n426740 , n80551 , n426742 , n426743 , n80554 , n426745 , n426746 , n426747 , n80558 , 
 n426749 , n426750 , n80561 , n426752 , n426753 , n426754 , n80565 , n426756 , n426757 , n426758 , 
 n80569 , n80570 , n426761 , n426762 , n426763 , n80574 , n80575 , n80576 , n426767 , n80578 , 
 n426769 , n426770 , n80581 , n80582 , n80583 , n80584 , n426775 , n426776 , n80587 , n80588 , 
 n80589 , n80590 , n80591 , n80592 , n80593 , n80594 , n80595 , n80596 , n80597 , n80598 , 
 n80599 , n426790 , n80601 , n80602 , n80603 , n80604 , n426795 , n426796 , n426797 , n426798 , 
 n80609 , n426800 , n426801 , n80612 , n80613 , n426804 , n426805 , n426806 , n426807 , n426808 , 
 n80619 , n80620 , n426811 , n426812 , n426813 , n80624 , n80625 , n426816 , n426817 , n80628 , 
 n426819 , n80630 , n426821 , n426822 , n426823 , n80634 , n426825 , n80636 , n426827 , n426828 , 
 n426829 , n80640 , n426831 , n426832 , n80643 , n80644 , n426835 , n426836 , n80647 , n426838 , 
 n426839 , n80650 , n80651 , n426842 , n80653 , n80654 , n80655 , n426846 , n80657 , n426848 , 
 n426849 , n80660 , n426851 , n426852 , n80663 , n426854 , n426855 , n80666 , n80667 , n426858 , 
 n426859 , n426860 , n80671 , n426862 , n426863 , n426864 , n426865 , n426866 , n426867 , n80678 , 
 n426869 , n426870 , n426871 , n426872 , n80683 , n80684 , n80685 , n426876 , n426877 , n426878 , 
 n426879 , n80690 , n426881 , n426882 , n426883 , n426884 , n426885 , n80696 , n426887 , n426888 , 
 n80699 , n80700 , n426891 , n426892 , n80703 , n426894 , n426895 , n80706 , n80707 , n426898 , 
 n426899 , n80710 , n426901 , n426902 , n426903 , n426904 , n80715 , n426906 , n426907 , n80718 , 
 n80719 , n426910 , n426911 , n80722 , n426913 , n426914 , n80725 , n80726 , n426917 , n80728 , 
 n426919 , n426920 , n80731 , n80732 , n80733 , n80734 , n426925 , n80736 , n426927 , n80738 , 
 n80739 , n80740 , n426931 , n80742 , n426933 , n426934 , n80745 , n426936 , n426937 , n80748 , 
 n80749 , n426940 , n426941 , n426942 , n80753 , n426944 , n426945 , n80756 , n80757 , n426948 , 
 n426949 , n80760 , n80761 , n80762 , n426953 , n426954 , n80765 , n80766 , n80767 , n426958 , 
 n426959 , n80770 , n80771 , n426962 , n426963 , n426964 , n426965 , n80776 , n426967 , n426968 , 
 n80779 , n80780 , n426971 , n426972 , n426973 , n80784 , n426975 , n426976 , n80787 , n80788 , 
 n426979 , n80790 , n80791 , n80792 , n426983 , n426984 , n80795 , n426986 , n80797 , n426988 , 
 n426989 , n426990 , n426991 , n80802 , n426993 , n426994 , n80805 , n80806 , n426997 , n426998 , 
 n426999 , n80810 , n427001 , n427002 , n80813 , n80814 , n427005 , n427006 , n80817 , n427008 , 
 n427009 , n80820 , n427011 , n427012 , n80823 , n427014 , n427015 , n427016 , n427017 , n80828 , 
 n427019 , n427020 , n80831 , n80832 , n427023 , n427024 , n80835 , n80836 , n80837 , n427028 , 
 n80839 , n80840 , n80841 , n80842 , n80843 , n80844 , n80845 , n80846 , n427037 , n80848 , 
 n80849 , n80850 , n427041 , n80852 , n80853 , n80854 , n80855 , n427046 , n80857 , n80858 , 
 n80859 , n427050 , n427051 , n80862 , n80863 , n80864 , n427055 , n427056 , n80867 , n80868 , 
 n80869 , n427060 , n427061 , n80872 , n80873 , n427064 , n427065 , n80876 , n427067 , n80878 , 
 n427069 , n80880 , n80881 , n427072 , n80883 , n427074 , n427075 , n427076 , n80887 , n427078 , 
 n80889 , n80890 , n427081 , n427082 , n80893 , n427084 , n427085 , n80896 , n427087 , n427088 , 
 n80899 , n427090 , n427091 , n80902 , n427093 , n427094 , n80905 , n80906 , n80907 , n427098 , 
 n80909 , n80910 , n80911 , n427102 , n80913 , n427104 , n80915 , n427106 , n80917 , n80918 , 
 n80919 , n80920 , n80921 , n80922 , n427113 , n427114 , n80925 , n427116 , n427117 , n427118 , 
 n427119 , n427120 , n80931 , n80932 , n80933 , n427124 , n427125 , n80936 , n427127 , n80938 , 
 n427129 , n80940 , n80941 , n427132 , n427133 , n80944 , n427135 , n427136 , n80947 , n427138 , 
 n427139 , n80950 , n427141 , n80952 , n80953 , n427144 , n427145 , n80956 , n427147 , n427148 , 
 n80959 , n427150 , n427151 , n80962 , n80963 , n80964 , n427155 , n427156 , n80967 , n80968 , 
 n80969 , n427160 , n427161 , n80972 , n80973 , n80974 , n427165 , n427166 , n80977 , n80978 , 
 n80979 , n427170 , n427171 , n80982 , n80983 , n80984 , n427175 , n427176 , n80987 , n80988 , 
 n80989 , n427180 , n427181 , n80992 , n80993 , n80994 , n427185 , n427186 , n427187 , n427188 , 
 n80999 , n427190 , n427191 , n81002 , n81003 , n81004 , n427195 , n427196 , n427197 , n81008 , 
 n81009 , n427200 , n81011 , n81012 , n81013 , n81014 , n81015 , n81016 , n81017 , n81018 , 
 n81019 , n81020 , n81021 , n81022 , n81023 , n81024 , n81025 , n81026 , n81027 , n81028 , 
 n81029 , n81030 , n81031 , n81032 , n81033 , n81034 , n81035 , n81036 , n81037 , n81038 , 
 n427229 , n427230 , n81056 , n81057 , n427233 , n427234 , n81060 , n81061 , n81062 , n427238 , 
 n427239 , n427240 , n81066 , n427242 , n81068 , n81069 , n427245 , n81071 , n427247 , n81073 , 
 n81074 , n427250 , n427251 , n81077 , n427253 , n427254 , n81080 , n427256 , n427257 , n427258 , 
 n81084 , n427260 , n427261 , n81087 , n427263 , n427264 , n427265 , n427266 , n81092 , n427268 , 
 n81094 , n427270 , n427271 , n81097 , n427273 , n81099 , n81100 , n81101 , n81102 , n81103 , 
 n81104 , n81105 , n81106 , n81107 , n81108 , n81109 , n81110 , n427286 , n81112 , n81113 , 
 n81114 , n81115 , n427291 , n81117 , n427293 , n81119 , n81120 , n427296 , n81122 , n427298 , 
 n81124 , n427300 , n427301 , n427302 , n427303 , n81129 , n81130 , n427306 , n427307 , n427308 , 
 n427309 , n81135 , n427311 , n81137 , n81138 , n427314 , n427315 , n81141 , n427317 , n427318 , 
 n81144 , n427320 , n81146 , n81147 , n81148 , n81149 , n427325 , n81151 , n427327 , n81153 , 
 n427329 , n81155 , n81156 , n427332 , n427333 , n81159 , n427335 , n81161 , n81162 , n427338 , 
 n427339 , n81165 , n427341 , n427342 , n81168 , n427344 , n427345 , n81171 , n427347 , n427348 , 
 n81174 , n427350 , n427351 , n81177 , n81178 , n427354 , n81180 , n427356 , n427357 , n81183 , 
 n427359 , n81185 , n427361 , n427362 , n81188 , n81189 , n81190 , n81191 , n427367 , n81193 , 
 n427369 , n427370 , n81196 , n427372 , n81198 , n81199 , n81200 , n81201 , n81202 , n427378 , 
 n81204 , n427380 , n81206 , n427382 , n81208 , n427384 , n81210 , n81211 , n427387 , n427388 , 
 n81214 , n427390 , n427391 , n81217 , n427393 , n427394 , n81220 , n81221 , n427397 , n427398 , 
 n81224 , n427400 , n427401 , n81227 , n427403 , n427404 , n81230 , n81231 , n81232 , n427408 , 
 n427409 , n81235 , n81236 , n81237 , n427413 , n427414 , n81240 , n81241 , n81242 , n427418 , 
 n427419 , n81245 , n81246 , n427422 , n427423 , n427424 , n427425 , n81276 , n81277 , n427428 , 
 n427429 , n81280 , n81282 , n427432 , n427433 , n81285 , n81286 , n427436 , n427437 , n81289 , 
 n81290 , n81291 , n427441 , n427442 , n81294 , n81295 , n81296 , n427446 , n427447 , n81299 , 
 n81300 , n427450 , n81302 , n81303 , n81304 , n427454 , n427455 , n427456 , n81308 , n427458 , 
 n81310 , n81311 , n427461 , n81313 , n427463 , n81315 , n81316 , n427466 , n427467 , n81319 , 
 n427469 , n427470 , n81322 , n427472 , n427473 , n427474 , n81326 , n427476 , n427477 , n81329 , 
 n427479 , n427480 , n427481 , n81333 , n427483 , n81335 , n81336 , n427486 , n427487 , n81339 , 
 n427489 , n427490 , n81342 , n427492 , n427493 , n81345 , n427495 , n81347 , n81348 , n427498 , 
 n81350 , n427500 , n81352 , n427502 , n427503 , n81355 , n427505 , n81357 , n427507 , n427508 , 
 n427509 , n81361 , n427511 , n427512 , n427513 , n427514 , n81366 , n81367 , n427517 , n81369 , 
 n427519 , n81371 , n81372 , n81373 , n81374 , n427524 , n81376 , n81377 , n427527 , n81379 , 
 n427529 , n427530 , n427531 , n81383 , n427533 , n81385 , n427535 , n81387 , n427537 , n81389 , 
 n427539 , n81391 , n81392 , n427542 , n427543 , n81395 , n427545 , n427546 , n81398 , n427548 , 
 n427549 , n81401 , n427551 , n81403 , n81404 , n427554 , n427555 , n81407 , n427557 , n427558 , 
 n81410 , n427560 , n427561 , n81413 , n81414 , n81415 , n427565 , n427566 , n81418 , n81419 , 
 n81420 , n427570 , n427571 , n81423 , n81424 , n81425 , n427575 , n427576 , n81428 , n81429 , 
 n427579 , n427580 , n427581 , n427582 , n81448 , n81449 , n427585 , n427586 , n81452 , n81453 , 
 n427589 , n427590 , n427591 , n427592 , n81470 , n81471 , n427595 , n427596 , n81474 , n81475 , 
 n427599 , n427600 , n81478 , n81479 , n81480 , n427604 , n427605 , n81483 , n81484 , n81485 , 
 n427609 , n427610 , n81488 , n81489 , n427613 , n427614 , n81492 , n427616 , n427617 , n81507 , 
 n81508 , n427620 , n427621 , n81511 , n81512 , n81513 , n427625 , n427626 , n81516 , n81517 , 
 n81518 , n81519 , n427631 , n81521 , n427633 , n81523 , n81524 , n427636 , n427637 , n81527 , 
 n427639 , n427640 , n81530 , n427642 , n427643 , n427644 , n81534 , n427646 , n81536 , n81537 , 
 n81538 , n81539 , n81540 , n81541 , n81542 , n81543 , n81544 , n81545 , n81546 , n81547 , 
 n81548 , n427660 , n427661 , n427662 , n81552 , n427664 , n81554 , n81555 , n427667 , n427668 , 
 n81558 , n427670 , n427671 , n81561 , n427673 , n427674 , n81564 , n427676 , n81566 , n81567 , 
 n427679 , n427680 , n81570 , n427682 , n427683 , n81573 , n427685 , n427686 , n81576 , n427688 , 
 n81578 , n81579 , n427691 , n81581 , n427693 , n81583 , n81584 , n427696 , n81586 , n427698 , 
 n427699 , n427700 , n81590 , n427702 , n427703 , n81593 , n427705 , n427706 , n81596 , n81597 , 
 n427709 , n427710 , n81600 , n81601 , n427713 , n81603 , n81604 , n427716 , n427717 , n427718 , 
 n81608 , n427720 , n427721 , n81611 , n427723 , n427724 , n81614 , n81615 , n81616 , n427728 , 
 n427729 , n427730 , n81620 , n427732 , n81622 , n427734 , n427735 , n427736 , n427737 , n427738 , 
 n81628 , n427740 , n427741 , n81631 , n427743 , n427744 , n81634 , n81635 , n427747 , n81637 , 
 n427749 , n427750 , n427751 , n427752 , n427753 , n81643 , n427755 , n427756 , n81646 , n427758 , 
 n427759 , n427760 , n81650 , n427762 , n427763 , n81653 , n427765 , n427766 , n81656 , n427768 , 
 n81658 , n427770 , n427771 , n427772 , n81662 , n427774 , n81664 , n427776 , n427777 , n427778 , 
 n427779 , n427780 , n81670 , n427782 , n427783 , n81673 , n427785 , n427786 , n81676 , n81677 , 
 n81678 , n427790 , n81680 , n81681 , n81682 , n427794 , n427795 , n427796 , n81686 , n427798 , 
 n81688 , n81689 , n427801 , n427802 , n81692 , n427804 , n427805 , n81695 , n427807 , n427808 , 
 n81698 , n427810 , n81700 , n427812 , n427813 , n81703 , n427815 , n427816 , n427817 , n427818 , 
 n427819 , n81709 , n427821 , n427822 , n81712 , n427824 , n81714 , n81715 , n427827 , n427828 , 
 n81718 , n427830 , n427831 , n81721 , n427833 , n427834 , n81724 , n81725 , n81726 , n427838 , 
 n81728 , n427840 , n427841 , n81731 , n81732 , n427844 , n81734 , n81735 , n427847 , n427848 , 
 n81738 , n427850 , n427851 , n81741 , n427853 , n81743 , n81744 , n427856 , n427857 , n81747 , 
 n427859 , n427860 , n81750 , n427862 , n81752 , n81753 , n81754 , n81755 , n81756 , n81757 , 
 n81758 , n81759 , n81760 , n427872 , n81762 , n81763 , n427875 , n427876 , n81766 , n81767 , 
 n81768 , n81769 , n81770 , n427882 , n427883 , n81773 , n81774 , n427886 , n81776 , n81777 , 
 n427889 , n427890 , n81780 , n427892 , n427893 , n81783 , n427895 , n427896 , n81786 , n427898 , 
 n427899 , n427900 , n427901 , n81794 , n427903 , n427904 , n81797 , n81798 , n427907 , n427908 , 
 n427909 , n427910 , n81823 , n81824 , n427913 , n427914 , n81827 , n81828 , n427917 , n427918 , 
 n81831 , n81832 , n81833 , n427922 , n427923 , n81836 , n81837 , n81838 , n427927 , n427928 , 
 n81841 , n81842 , n427931 , n427932 , n81845 , n81846 , n81847 , n427936 , n427937 , n81850 , 
 n81851 , n427940 , n427941 , n427942 , n81872 , n427944 , n81885 , n81886 , n427947 , n427948 , 
 n427949 , n81893 , n427951 , n427952 , n81896 , n427954 , n81898 , n427956 , n427957 , n427958 , 
 n81902 , n427960 , n81904 , n81905 , n427963 , n427964 , n81908 , n427966 , n427967 , n81911 , 
 n427969 , n427970 , n81914 , n427972 , n81916 , n81917 , n427975 , n427976 , n81920 , n427978 , 
 n427979 , n81923 , n427981 , n427982 , n81926 , n427984 , n427985 , n81929 , n427987 , n427988 , 
 n81932 , n81933 , n81934 , n427992 , n427993 , n427994 , n427995 , n81939 , n81940 , n427998 , 
 n81942 , n81943 , n428001 , n428002 , n81946 , n428004 , n81948 , n81949 , n428007 , n428008 , 
 n81952 , n428010 , n428011 , n81955 , n428013 , n428014 , n81958 , n428016 , n428017 , n81961 , 
 n428019 , n81963 , n428021 , n428022 , n81966 , n81967 , n81968 , n428026 , n428027 , n81971 , 
 n428029 , n428030 , n81974 , n428032 , n428033 , n81977 , n428035 , n428036 , n428037 , n428038 , 
 n81985 , n428040 , n428041 , n81988 , n81989 , n81990 , n428045 , n428046 , n81993 , n81994 , 
 n81995 , n428050 , n428051 , n81998 , n81999 , n428054 , n428055 , n82002 , n428057 , n428058 , 
 n82005 , n428060 , n82007 , n428062 , n428063 , n428064 , n428065 , n82012 , n428067 , n82014 , 
 n428069 , n428070 , n428071 , n428072 , n82040 , n82041 , n428075 , n82043 , n428077 , n82072 , 
 n82073 , n82074 , n82077 , n428082 , n82079 , n428084 , n428085 , n82082 , n82083 , n428088 , 
 n82085 , n82086 , n428091 , n428092 , n82089 , n82090 , n428095 , n428096 , n82093 , n428098 , 
 n428099 , n82096 , n428101 , n428102 , n82099 , n428104 , n82101 , n428106 , n428107 , n82104 , 
 n428109 , n428110 , n82107 , n82108 , n428113 , n428114 , n428115 , n82112 , n428117 , n428118 , 
 n82115 , n82116 , n428121 , n82118 , n82119 , n82120 , n428125 , n428126 , n428127 , n82124 , 
 n428129 , n428130 , n82127 , n82128 , n428133 , n428134 , n82131 , n428136 , n428137 , n82134 , 
 n82135 , n428140 , n428141 , n428142 , n428143 , n82140 , n428145 , n428146 , n82143 , n428148 , 
 n82145 , n428150 , n428151 , n428152 , n82149 , n428154 , n428155 , n82152 , n428157 , n428158 , 
 n428159 , n82156 , n428161 , n428162 , n82159 , n82160 , n428165 , n428166 , n82163 , n428168 , 
 n428169 , n82166 , n82167 , n428172 , n428173 , n82170 , n82171 , n82172 , n428177 , n428178 , 
 n82175 , n428180 , n428181 , n82178 , n428183 , n428184 , n82181 , n428186 , n428187 , n82184 , 
 n82185 , n428190 , n428191 , n428192 , n82189 , n428194 , n428195 , n428196 , n82193 , n428198 , 
 n428199 , n428200 , n428201 , n82198 , n428203 , n428204 , n428205 , n428206 , n82203 , n428208 , 
 n428209 , n82206 , n82207 , n428212 , n428213 , n428214 , n82211 , n428216 , n428217 , n82214 , 
 n82215 , n428220 , n428221 , n82218 , n428223 , n428224 , n82221 , n428226 , n428227 , n82224 , 
 n428229 , n428230 , n428231 , n82228 , n428233 , n82230 , n428235 , n428236 , n82233 , n428238 , 
 n428239 , n82236 , n82237 , n82238 , n428243 , n428244 , n82241 , n82242 , n82243 , n428248 , 
 n82245 , n82246 , n82247 , n82248 , n82249 , n82250 , n82251 , n82252 , n82253 , n82254 , 
 n428259 , n428260 , n428261 , n82258 , n428263 , n428264 , n82261 , n82262 , n428267 , n428268 , 
 n428269 , n82266 , n428271 , n428272 , n82269 , n82270 , n428275 , n82272 , n428277 , n428278 , 
 n82275 , n428280 , n428281 , n82278 , n82279 , n428284 , n428285 , n428286 , n82283 , n428288 , 
 n428289 , n82286 , n82287 , n428292 , n428293 , n82290 , n82291 , n428296 , n428297 , n82294 , 
 n428299 , n428300 , n82297 , n428302 , n82299 , n428304 , n428305 , n428306 , n428307 , n428308 , 
 n82305 , n428310 , n428311 , n82308 , n82309 , n428314 , n428315 , n82312 , n428317 , n428318 , 
 n82315 , n82316 , n428321 , n428322 , n82319 , n82320 , n428325 , n428326 , n82323 , n82324 , 
 n82325 , n428330 , n428331 , n82328 , n82329 , n82330 , n428335 , n82332 , n82333 , n82334 , 
 n428339 , n82336 , n82337 , n82338 , n82339 , n428344 , n82341 , n82342 , n82343 , n82344 , 
 n82345 , n428350 , n82347 , n82348 , n82349 , n428354 , n82351 , n82352 , n82353 , n82354 , 
 n82355 , n428360 , n82357 , n82358 , n428363 , n428364 , n82361 , n428366 , n82363 , n428368 , 
 n82365 , n82366 , n428371 , n428372 , n82369 , n428374 , n428375 , n82372 , n428377 , n428378 , 
 n82375 , n428380 , n82377 , n82378 , n428383 , n428384 , n82381 , n428386 , n428387 , n82384 , 
 n428389 , n428390 , n82387 , n82388 , n82389 , n428394 , n82391 , n428396 , n82393 , n428398 , 
 n82395 , n82396 , n428401 , n428402 , n82399 , n428404 , n82401 , n82402 , n428407 , n428408 , 
 n82405 , n428410 , n428411 , n82408 , n428413 , n428414 , n82411 , n428416 , n428417 , n82414 , 
 n428419 , n428420 , n82417 , n428422 , n82419 , n82420 , n82421 , n82422 , n428427 , n82424 , 
 n82425 , n428430 , n428431 , n82428 , n428433 , n82430 , n82431 , n82432 , n428437 , n82434 , 
 n428439 , n82436 , n82437 , n82438 , n82439 , n82440 , n428445 , n82442 , n82443 , n82444 , 
 n82445 , n428450 , n82447 , n82448 , n82449 , n428454 , n428455 , n82452 , n428457 , n428458 , 
 n82466 , n82467 , n82468 , n428462 , n428463 , n82471 , n428465 , n428466 , n82474 , n428468 , 
 n82476 , n428470 , n428471 , n428472 , n428473 , n82481 , n428475 , n428476 , n82484 , n82485 , 
 n428479 , n428480 , n82488 , n82489 , n428483 , n428484 , n82492 , n82493 , n82494 , n428488 , 
 n82496 , n82497 , n82498 , n428492 , n428493 , n82501 , n82502 , n428496 , n82518 , n82519 , 
 n82520 , n82521 , n82522 , n428502 , n428503 , n82525 , n428505 , n82527 , n82528 , n82529 , 
 n82530 , n428510 , n428511 , n82533 , n428513 , n82535 , n82536 , n428516 , n82538 , n428518 , 
 n82540 , n428520 , n428521 , n82543 , n82544 , n428524 , n428525 , n82547 , n428527 , n428528 , 
 n82550 , n428530 , n428531 , n428532 , n82554 , n428534 , n428535 , n82557 , n428537 , n428538 , 
 n82560 , n82561 , n82562 , n82563 , n428543 , n428544 , n82566 , n428546 , n82568 , n82569 , 
 n428549 , n428550 , n82572 , n428552 , n82574 , n82575 , n428555 , n428556 , n82578 , n428558 , 
 n428559 , n82581 , n428561 , n428562 , n82584 , n428564 , n428565 , n82587 , n428567 , n428568 , 
 n82590 , n82591 , n82592 , n428572 , n82594 , n82595 , n82596 , n428576 , n428577 , n82599 , 
 n428579 , n428580 , n82602 , n82603 , n428583 , n428584 , n428585 , n82607 , n428587 , n428588 , 
 n82610 , n82611 , n428591 , n428592 , n428593 , n82615 , n428595 , n428596 , n82618 , n428598 , 
 n82620 , n428600 , n428601 , n428602 , n82624 , n428604 , n428605 , n428606 , n428607 , n428608 , 
 n82630 , n428610 , n428611 , n82633 , n82634 , n428614 , n428615 , n82637 , n428617 , n428618 , 
 n82640 , n82641 , n428621 , n428622 , n82644 , n428624 , n428625 , n428626 , n82648 , n428628 , 
 n428629 , n82651 , n82652 , n428632 , n428633 , n82655 , n428635 , n428636 , n82658 , n82659 , 
 n428639 , n428640 , n428641 , n428642 , n82664 , n428644 , n428645 , n82667 , n428647 , n428648 , 
 n82670 , n82671 , n82672 , n428652 , n82674 , n82675 , n82676 , n428656 , n82678 , n82679 , 
 n82680 , n428660 , n82682 , n82683 , n428663 , n428664 , n82686 , n82687 , n82688 , n428668 , 
 n428669 , n82691 , n82692 , n82693 , n428673 , n82695 , n82696 , n82697 , n82698 , n82699 , 
 n428679 , n82701 , n82702 , n428682 , n428683 , n82705 , n428685 , n82707 , n82708 , n428688 , 
 n82710 , n428690 , n82712 , n82713 , n428693 , n428694 , n82716 , n428696 , n428697 , n82719 , 
 n428699 , n428700 , n82722 , n82723 , n428703 , n428704 , n82726 , n428706 , n428707 , n82729 , 
 n428709 , n428710 , n82732 , n82733 , n82734 , n428714 , n428715 , n82737 , n82738 , n82739 , 
 n428719 , n428720 , n82742 , n82743 , n82744 , n428724 , n428725 , n82747 , n82748 , n82749 , 
 n428729 , n428730 , n428731 , n82753 , n428733 , n82755 , n82756 , n428736 , n82758 , n428738 , 
 n82760 , n82761 , n428741 , n428742 , n82764 , n428744 , n428745 , n82767 , n428747 , n428748 , 
 n428749 , n82771 , n428751 , n428752 , n82774 , n428754 , n428755 , n82777 , n428757 , n428758 , 
 n82780 , n428760 , n428761 , n82783 , n82784 , n82785 , n428765 , n428766 , n82788 , n82789 , 
 n82790 , n82791 , n428771 , n428772 , n82794 , n428774 , n82796 , n82797 , n82798 , n82799 , 
 n428779 , n82801 , n428781 , n82803 , n428783 , n82805 , n428785 , n428786 , n82808 , n428788 , 
 n82810 , n82811 , n82812 , n82813 , n82814 , n82815 , n428795 , n428796 , n82818 , n428798 , 
 n428799 , n82821 , n428801 , n428802 , n428803 , n82825 , n428805 , n82827 , n82828 , n428808 , 
 n428809 , n82831 , n428811 , n428812 , n82834 , n428814 , n428815 , n82837 , n428817 , n82839 , 
 n82840 , n428820 , n428821 , n82843 , n428823 , n428824 , n82846 , n428826 , n428827 , n82849 , 
 n428829 , n82851 , n82852 , n428832 , n428833 , n82855 , n428835 , n82857 , n428837 , n82859 , 
 n428839 , n428840 , n82862 , n82863 , n82864 , n428844 , n428845 , n82867 , n82868 , n82869 , 
 n428849 , n82871 , n428851 , n428852 , n82874 , n428854 , n428855 , n428856 , n428857 , n82879 , 
 n428859 , n428860 , n82882 , n428862 , n428863 , n82885 , n82886 , n82887 , n428867 , n82889 , 
 n82890 , n82891 , n82892 , n82893 , n82894 , n82895 , n82896 , n82897 , n82898 , n82899 , 
 n82900 , n82901 , n82902 , n82903 , n82904 , n428884 , n82906 , n82907 , n82908 , n82909 , 
 n82910 , n428890 , n428891 , n82915 , n82916 , n82917 , n428895 , n428896 , n82920 , n428898 , 
 n82922 , n428900 , n82924 , n428902 , n428903 , n82927 , n428905 , n82929 , n428907 , n82931 , 
 n428909 , n82933 , n428911 , n428912 , n82936 , n428914 , n82938 , n82939 , n428917 , n428918 , 
 n82942 , n82943 , n428921 , n428922 , n82946 , n82947 , n428925 , n428926 , n82950 , n428928 , 
 n82952 , n428930 , n428931 , n82955 , n428933 , n82957 , n428935 , n428936 , n82960 , n82961 , 
 n428939 , n428940 , n82964 , n428942 , n428943 , n428944 , n82968 , n428946 , n82970 , n82971 , 
 n82972 , n82973 , n428951 , n428952 , n428953 , n428954 , n82990 , n428956 , n428957 , n82993 , 
 n428959 , n82995 , n428961 , n428962 , n82998 , n83000 , n428965 , n428966 , n83004 , n83005 , 
 n83006 , n83007 , n83008 , n83009 , n83010 , n83011 , n83012 , n83014 , n428977 , n428978 , 
 n428979 , n83030 , n83031 , n428982 , n428983 , n83034 , n428985 , n428986 , n83037 , n428988 , 
 n428989 , n83040 , n83041 , n83042 , n83043 , n83044 , n428995 , n83046 , n428997 , n83048 , 
 n83049 , n429000 , n429001 , n429002 , n83076 , n83077 , n429005 , n429006 , n83080 , n83081 , 
 n83082 , n83083 , n429011 , n83085 , n429013 , n83087 , n429015 , n83089 , n429017 , n83091 , 
 n83092 , n429020 , n83094 , n83095 , n429023 , n429024 , n83098 , n429026 , n83100 , n429028 , 
 n83102 , n83103 , n83104 , n83105 , n83106 , n83107 , n429035 , n429036 , n83110 , n429038 , 
 n429039 , n83113 , n429041 , n429042 , n83116 , n83117 , n83118 , n429046 , n429047 , n429048 , 
 n429049 , n83148 , n83149 , n429052 , n429053 , n83152 , n429055 , n429056 , n429057 , n429058 , 
 n429059 , n429060 , n429061 , n429062 , n429063 , n429064 , n429065 , n429066 , n429067 , n429068 , 
 n83188 , n429070 , n429071 , n429072 , n429073 , n429074 , n83194 , n429076 , n429077 , n83197 , 
 n429079 , n429080 , n429081 , n429082 , n429083 , n83203 , n429085 , n429086 , n83206 , n429088 , 
 n429089 , n83209 , n429091 , n429092 , n429093 , n429094 , n429095 , n429096 , n429097 , n429098 , 
 n429099 , n429100 , n429101 , n429102 , n429103 , n429104 , n429105 , n429106 , n429107 , n429108 , 
 n429109 , n429110 , n429111 , n429112 , n429113 , n429114 , n429115 , n429116 , n429117 , n429118 , 
 n429119 , n429120 , n429121 , n429122 , n429123 , n429124 , n429125 , n429126 , n429127 , n429128 , 
 n83248 , n429130 , n429131 , n429132 , n429133 , n429134 , n429135 , n429136 , n429137 , n429138 , 
 n429139 , n429140 , n429141 , n429142 , n429143 , n429144 , n429145 , n429146 , n83266 , n429148 , 
 n429149 , n83269 , n429151 , n429152 , n83272 , n429154 , n429155 , n429156 , n429157 , n429158 , 
 n429159 , n429160 , n429161 , n429162 , n429163 , n429164 , n429165 , n429166 , n429167 , n429168 , 
 n429169 , n429170 , n429171 , n429172 , n429173 , n429174 , n429175 , n429176 , n83296 , n429178 , 
 n429179 , n83299 , n83300 , n429182 , n429183 , n83303 , n429185 , n83305 , n429187 , n429188 , 
 n429189 , n83309 , n429191 , n429192 , n83312 , n83313 , n429195 , n429196 , n429197 , n83317 , 
 n429199 , n429200 , n83320 , n83321 , n429203 , n83323 , n83324 , n429206 , n83326 , n83327 , 
 n83328 , n429210 , n83330 , n83331 , n429213 , n429214 , n83334 , n83335 , n83336 , n429218 , 
 n429219 , n83339 , n83340 , n83341 , n429223 , n83343 , n83344 , n83345 , n83346 , n83347 , 
 n429229 , n83349 , n83350 , n429232 , n429233 , n83353 , n429235 , n83355 , n429237 , n83357 , 
 n429239 , n83359 , n83360 , n83361 , n83362 , n429244 , n83364 , n83365 , n429247 , n429248 , 
 n83368 , n83369 , n429251 , n83371 , n429253 , n429254 , n83374 , n83375 , n429257 , n429258 , 
 n429259 , n83379 , n429261 , n429262 , n83382 , n429264 , n429265 , n83385 , n83386 , n83387 , 
 n429269 , n429270 , n83390 , n429272 , n429273 , n429274 , n429275 , n83414 , n429277 , n83416 , 
 n429279 , n83418 , n429281 , n429282 , n83421 , n83422 , n429285 , n429286 , n83425 , n429288 , 
 n429289 , n83428 , n429291 , n429292 , n83431 , n429294 , n83433 , n83434 , n429297 , n83436 , 
 n429299 , n83438 , n83439 , n429302 , n429303 , n83442 , n429305 , n429306 , n83445 , n429308 , 
 n429309 , n429310 , n83449 , n429312 , n429313 , n83452 , n429315 , n429316 , n83455 , n83457 , 
 n429319 , n429320 , n429321 , n83461 , n429323 , n83463 , n83464 , n429326 , n83466 , n83467 , 
 n83468 , n83469 , n429331 , n83471 , n429333 , n429334 , n83474 , n429336 , n429337 , n429338 , 
 n429339 , n429340 , n83480 , n429342 , n429343 , n429344 , n83484 , n83485 , n429347 , n429348 , 
 n83488 , n429350 , n429351 , n83491 , n429353 , n429354 , n83494 , n429356 , n83496 , n429358 , 
 n83498 , n83499 , n429361 , n429362 , n83502 , n429364 , n429365 , n83505 , n429367 , n429368 , 
 n429369 , n429370 , n83510 , n429372 , n429373 , n83513 , n429375 , n429376 , n83516 , n429378 , 
 n83518 , n429380 , n83520 , n83521 , n429383 , n429384 , n83524 , n429386 , n429387 , n83527 , 
 n429389 , n429390 , n83530 , n429392 , n83532 , n83533 , n429395 , n429396 , n83536 , n429398 , 
 n429399 , n83539 , n429401 , n429402 , n83542 , n83543 , n429405 , n429406 , n83546 , n429408 , 
 n429409 , n429410 , n83550 , n429412 , n83552 , n429414 , n429415 , n429416 , n429417 , n83557 , 
 n429419 , n429420 , n83560 , n429422 , n429423 , n83563 , n83564 , n83565 , n429427 , n429428 , 
 n429429 , n83569 , n429431 , n429432 , n429433 , n83573 , n429435 , n429436 , n429437 , n429438 , 
 n429439 , n83591 , n429441 , n429442 , n429443 , n83595 , n429445 , n429446 , n429447 , n83599 , 
 n429449 , n83601 , n429451 , n429452 , n429453 , n429454 , n429455 , n429456 , n429457 , n83609 , 
 n429459 , n429460 , n429461 , n429462 , n429463 , n83615 , n429465 , n429466 , n429467 , n429468 , 
 n429469 , n429470 , n429471 , n429472 , n429473 , n429474 , n429475 , n429476 , n429477 , n429478 , 
 n83653 , n429480 , n429481 , n429482 , n429483 , n429484 , n83659 , n429486 , n429487 , n429488 , 
 n83663 , n429490 , n429491 , n429492 , n429493 , n429494 , n83669 , n429496 , n429497 , n429498 , 
 n429499 , n429500 , n83675 , n429502 , n429503 , n429504 , n429505 , n429506 , n83681 , n429508 , 
 n429509 , n429510 , n429511 , n429512 , n429513 , n83689 , n429515 , n83691 , n429517 , n83693 , 
 n429519 , n429520 , n429521 , n83697 , n429523 , n83699 , n429525 , n429526 , n429527 , n83703 , 
 n429529 , n429530 , n429531 , n429532 , n429533 , n83709 , n429535 , n429536 , n429537 , n429538 , 
 n429539 , n83715 , n429541 , n429542 , n429543 , n83719 , n429545 , n429546 , n429547 , n83723 , 
 n429549 , n83725 , n83726 , n429552 , n429553 , n83729 , n429555 , n429556 , n429557 , n429558 , 
 n429559 , n83735 , n429561 , n83737 , n83738 , n429564 , n429565 , n83741 , n429567 , n429568 , 
 n83744 , n429570 , n429571 , n83747 , n429573 , n83749 , n83750 , n429576 , n429577 , n83753 , 
 n429579 , n429580 , n83756 , n429582 , n429583 , n83759 , n429585 , n83761 , n83762 , n429588 , 
 n429589 , n429590 , n429591 , n83767 , n429593 , n429594 , n429595 , n429596 , n83785 , n83786 , 
 n429599 , n429600 , n83789 , n429602 , n429603 , n429604 , n429605 , n429606 , n83809 , n429608 , 
 n429609 , n83812 , n83813 , n429612 , n429613 , n429614 , n429615 , n83818 , n83819 , n429618 , 
 n83821 , n429620 , n429621 , n429622 , n83825 , n429624 , n429625 , n83828 , n429627 , n83830 , 
 n83831 , n429630 , n429631 , n83834 , n429633 , n429634 , n83837 , n429636 , n429637 , n429638 , 
 n429639 , n83842 , n429641 , n429642 , n429643 , n429644 , n429645 , n83848 , n429647 , n429648 , 
 n83851 , n429650 , n429651 , n83866 , n429653 , n429654 , n429655 , n429656 , n429657 , n429658 , 
 n429659 , n429660 , n429661 , n429662 , n429663 , n429664 , n429665 , n429666 , n429667 , n429668 , 
 n429669 , n429670 , n429671 , n429672 , n429673 , n429674 , n429675 , n429676 , n429677 , n429678 , 
 n429679 , n429680 , n429681 , n429682 , n429683 , n429684 , n429685 , n83899 , n429687 , n83901 , 
 n429689 , n429690 , n83904 , n429692 , n429693 , n429694 , n429695 , n83909 , n429697 , n429698 , 
 n429699 , n83913 , n429701 , n429702 , n429703 , n83917 , n429705 , n429706 , n83920 , n83921 , 
 n429709 , n429710 , n83924 , n429712 , n429713 , n429714 , n429715 , n429716 , n429717 , n83931 , 
 n83932 , n429720 , n429721 , n83935 , n429723 , n429724 , n83938 , n83939 , n429727 , n429728 , 
 n83942 , n83943 , n83944 , n429732 , n83946 , n83947 , n83948 , n429736 , n429737 , n83951 , 
 n429739 , n429740 , n429741 , n429742 , n429743 , n429744 , n83958 , n429746 , n429747 , n83961 , 
 n429749 , n429750 , n429751 , n429752 , n83966 , n429754 , n429755 , n429756 , n83970 , n429758 , 
 n83972 , n429760 , n429761 , n83975 , n429763 , n429764 , n83978 , n429766 , n429767 , n83981 , 
 n83982 , n83983 , n429771 , n429772 , n83986 , n429774 , n83988 , n429776 , n83990 , n83991 , 
 n83992 , n83993 , n83994 , n83995 , n83996 , n429784 , n429785 , n83999 , n84000 , n84001 , 
 n84002 , n84003 , n429791 , n429792 , n84006 , n429794 , n84008 , n84009 , n84010 , n429798 , 
 n429799 , n429800 , n84014 , n429802 , n84016 , n84017 , n429805 , n84019 , n84020 , n84021 , 
 n84022 , n84023 , n84024 , n84025 , n429813 , n84027 , n429815 , n84029 , n84030 , n84031 , 
 n429819 , n84033 , n429821 , n429822 , n84036 , n84037 , n84038 , n84039 , n429827 , n84041 , 
 n429829 , n84043 , n84044 , n429832 , n429833 , n84047 , n429835 , n84049 , n429837 , n84051 , 
 n429839 , n84053 , n429841 , n84055 , n84056 , n429844 , n429845 , n84059 , n429847 , n429848 , 
 n84062 , n429850 , n429851 , n84065 , n429853 , n84067 , n84068 , n429856 , n429857 , n84071 , 
 n429859 , n429860 , n84074 , n429862 , n429863 , n84077 , n84078 , n429866 , n429867 , n84081 , 
 n84082 , n429870 , n429871 , n84085 , n84086 , n429874 , n84088 , n84089 , n429877 , n84091 , 
 n84092 , n84093 , n84094 , n84095 , n84124 , n429884 , n429885 , n84129 , n429887 , n429888 , 
 n84132 , n429890 , n84134 , n429892 , n84136 , n429894 , n84138 , n84139 , n429897 , n84141 , 
 n84142 , n84143 , n84144 , n84145 , n84146 , n429904 , n429905 , n429906 , n84171 , n84172 , 
 n429909 , n429910 , n84175 , n429912 , n429913 , n84178 , n429915 , n429916 , n429917 , n429918 , 
 n429919 , n84184 , n429921 , n429922 , n84187 , n84188 , n84189 , n429926 , n429927 , n84192 , 
 n429929 , n429930 , n84195 , n429932 , n429933 , n84198 , n429935 , n84200 , n429937 , n84202 , 
 n429939 , n429940 , n84205 , n429942 , n429943 , n84208 , n84209 , n84210 , n429947 , n429948 , 
 n84213 , n429950 , n429951 , n84216 , n84217 , n84218 , n84219 , n429956 , n429957 , n84222 , 
 n429959 , n429960 , n429961 , n84226 , n429963 , n84228 , n429965 , n429966 , n84231 , n429968 , 
 n429969 , n429970 , n429971 , n84236 , n429973 , n84238 , n429975 , n429976 , n429977 , n429978 , 
 n84263 , n429980 , n429981 , n84277 , n84278 , n429984 , n429985 , n84281 , n429987 , n84283 , 
 n429989 , n84285 , n429991 , n429992 , n429993 , n429994 , n84290 , n429996 , n84292 , n429998 , 
 n429999 , n430000 , n430001 , n430002 , n84298 , n84299 , n84300 , n84301 , n84302 , n430008 , 
 n84304 , n430010 , n430011 , n84307 , n84308 , n430014 , n84310 , n430016 , n84312 , n84313 , 
 n430019 , n430020 , n84316 , n430022 , n430023 , n84319 , n430025 , n84321 , n84322 , n84323 , 
 n84324 , n430030 , n84326 , n430032 , n430033 , n84329 , n84330 , n430036 , n430037 , n84333 , 
 n430039 , n430040 , n430041 , n84337 , n430043 , n430044 , n84343 , n430046 , n84345 , n84346 , 
 n84347 , n84348 , n430051 , n430052 , n430053 , n430054 , n84353 , n430056 , n430057 , n84356 , 
 n84357 , n430060 , n430061 , n430062 , n84361 , n430064 , n430065 , n84364 , n84365 , n430068 , 
 n430069 , n84368 , n430071 , n430072 , n84371 , n430074 , n430075 , n84374 , n430077 , n430078 , 
 n430079 , n430080 , n84379 , n430082 , n430083 , n84382 , n84383 , n430086 , n430087 , n430088 , 
 n430089 , n84388 , n430091 , n430092 , n430093 , n84392 , n430095 , n84394 , n430097 , n430098 , 
 n84397 , n430100 , n430101 , n84400 , n430103 , n430104 , n84403 , n430106 , n430107 , n430108 , 
 n84407 , n430110 , n84409 , n430112 , n430113 , n84412 , n430115 , n430116 , n84415 , n430118 , 
 n430119 , n84418 , n84419 , n84420 , n430123 , n430124 , n84423 , n84424 , n84425 , n430128 , 
 n430129 , n84428 , n430131 , n84430 , n84431 , n430134 , n430135 , n84434 , n430137 , n84436 , 
 n84437 , n430140 , n84439 , n84440 , n430143 , n84442 , n430145 , n430146 , n84445 , n430148 , 
 n430149 , n430150 , n84449 , n430152 , n84451 , n430154 , n430155 , n84454 , n430157 , n84456 , 
 n84457 , n84458 , n430161 , n84460 , n430163 , n84462 , n430165 , n84464 , n84465 , n430168 , 
 n430169 , n84485 , n430171 , n84492 , n84493 , n84494 , n84495 , n430176 , n430177 , n84498 , 
 n430179 , n84500 , n84501 , n84502 , n84503 , n84504 , n84505 , n84506 , n430187 , n84508 , 
 n430189 , n430190 , n430191 , n430192 , n430193 , n430194 , n84517 , n430196 , n84519 , n84520 , 
 n84521 , n84522 , n430201 , n84524 , n84525 , n430204 , n84527 , n430206 , n430207 , n430208 , 
 n84531 , n430210 , n430211 , n84534 , n430213 , n430214 , n84537 , n430216 , n430217 , n84540 , 
 n430219 , n430220 , n84543 , n430222 , n430223 , n430224 , n84547 , n84550 , n430227 , n430228 , 
 n84556 , n430230 , n430231 , n430232 , n84560 , n430234 , n430235 , n430236 , n430237 , n84584 , 
 n84585 , n84586 , n430241 , n430242 , n84589 , n430244 , n430245 , n430246 , n84613 , n430248 , 
 n430249 , n84616 , n84617 , n430252 , n84619 , n430254 , n430255 , n84626 , n430257 , n430258 , 
 n84629 , n84630 , n84631 , n430262 , n430263 , n84634 , n430265 , n84636 , n84637 , n84638 , 
 n430269 , n430270 , n430271 , n430272 , n84643 , n430274 , n430275 , n84646 , n430277 , n430278 , 
 n84649 , n430280 , n84651 , n430282 , n430283 , n430284 , n430285 , n430286 , n84657 , n84674 , 
 n84675 , n84676 , n430291 , n430292 , n84679 , n430294 , n430295 , n430296 , n430297 , n84687 , 
 n430299 , n430300 , n84690 , n84693 , n84695 , n84696 , n84697 , n84698 , n84701 , n84703 , 
 n84704 , n84705 , n84706 , n84707 , n430313 , n84709 , n84710 , n84711 , n430317 , n430318 , 
 n430319 , n430320 , n84735 , n84736 , n84737 , n84738 , n84739 , n84740 , n84741 , n84742 , 
 n84743 , n84744 , n84745 , n430332 , n84747 , n84749 , n430335 , n430336 , n84752 , n84753 , 
 n84754 , n84755 , n84756 , n84757 , n84758 , n84759 , n84760 , n430346 , n430347 , n430348 , 
 n430349 , n84784 , n430351 , n84786 , n84787 , n430354 , n430355 , n84790 , n84791 , n430358 , 
 n430359 , n430360 , n430361 , n430362 , n84797 , n430364 , n430365 , n84800 , n430367 , n430368 , 
 n430369 , n430370 , n84805 , n430372 , n84807 , n430374 , n430375 , n430376 , n430377 , n430378 , 
 n84819 , n84820 , n430381 , n430382 , n430383 , n430384 , n84830 , n84831 , n430387 , n430388 , 
 n430389 , n84837 , n430391 , n84839 , n84840 , n430394 , n430395 , n84843 , n84844 , n430398 , 
 n430399 , n84847 , n84848 , n84852 , n430403 , n430404 , n430405 , n430406 , n84874 , n84875 , 
 n430409 , n430410 , n84878 , n84879 , n84880 , n430414 , n430415 , n84883 , n84885 , n430418 , 
 n430419 , n84888 , n84889 , n84890 , n430423 , n430424 , n84893 , n84894 , n84895 , n430428 , 
 n430429 , n84898 , n430431 , n84900 , n430433 , n84906 , n84907 , n430436 , n430437 , n84910 , 
 n430439 , n430440 , n84913 , n84914 , n430443 , n430444 , n84917 , n430446 , n430447 , n84920 , 
 n430449 , n430450 , n84923 , n84925 , n430453 , n430454 , n84966 , n84967 , n430457 , n430458 , 
 n84970 , n84971 , n430461 , n430462 , n430463 , n430464 , n84976 , n84977 , n430467 , n430468 , 
 n430469 , n430470 , n430471 , n430472 , n430473 , n430474 , n430475 , n430476 , n430477 , n430478 , 
 n430479 , n85039 , n85040 , n430482 , n430483 , n430484 , n430485 , n85060 , n430487 , n430488 , 
 n85073 , n85074 , n430491 , n430492 , n85083 , n85084 , n430495 , n430496 , n430497 , n430498 , 
 n85092 , n430500 , n430501 , n85095 , n430503 , n85097 , n430505 , n430506 , n85100 , n85102 , 
 n430509 , n85104 , n85105 , n85106 , n430513 , n430514 , n430515 , n85110 , n430517 , n85112 , 
 n85113 , n430520 , n430521 , n85116 , n430523 , n430524 , n85119 , n430526 , n85121 , n430528 , 
 n85123 , n430530 , n85125 , n85126 , n430533 , n430534 , n85129 , n430536 , n85131 , n430538 , 
 n430539 , n430540 , n85135 , n430542 , n430543 , n85138 , n430545 , n85140 , n85141 , n430548 , 
 n430549 , n85144 , n430551 , n85146 , n430553 , n430554 , n85149 , n430556 , n430557 , n85166 , 
 n430559 , n85168 , n430561 , n430562 , n430563 , n430564 , n85176 , n430566 , n85178 , n430568 , 
 n85180 , n85181 , n430571 , n430572 , n85184 , n85185 , n430575 , n85187 , n85188 , n85189 , 
 n85190 , n430580 , n85192 , n85193 , n430583 , n430584 , n430585 , n85197 , n430587 , n430588 , 
 n85200 , n430590 , n85202 , n430592 , n85204 , n430594 , n85206 , n85207 , n430597 , n430598 , 
 n85210 , n85211 , n430601 , n430602 , n85214 , n430604 , n85216 , n85217 , n430607 , n430608 , 
 n85220 , n85221 , n430611 , n430612 , n430613 , n430614 , n85226 , n430616 , n85228 , n430618 , 
 n430619 , n85231 , n430621 , n430622 , n430623 , n430624 , n85240 , n430626 , n430627 , n85243 , 
 n430629 , n85245 , n85246 , n430632 , n85248 , n430634 , n430635 , n430636 , n85252 , n430638 , 
 n430639 , n85255 , n430641 , n85257 , n430643 , n85259 , n430645 , n430646 , n85280 , n85281 , 
 n430649 , n430650 , n85284 , n85285 , n85286 , n430654 , n430655 , n85289 , n430657 , n430658 , 
 n85292 , n85293 , n85294 , n430662 , n430663 , n85297 , n430665 , n430666 , n85300 , n85301 , 
 n430669 , n430670 , n85304 , n85305 , n85307 , n430674 , n430675 , n85310 , n430677 , n430678 , 
 n85313 , n430680 , n430681 , n85316 , n430683 , n430684 , n85319 , n430686 , n85321 , n85322 , 
 n430689 , n85324 , n430691 , n85326 , n430693 , n85328 , n85329 , n430696 , n85331 , n430698 , 
 n85333 , n430700 , n430701 , n85336 , n430703 , n85338 , n85339 , n430706 , n430707 , n85342 , 
 n430709 , n430710 , n85345 , n430712 , n430713 , n85348 , n85351 , n85352 , n430717 , n430718 , 
 n85355 , n85356 , n430721 , n430722 , n85359 , n85360 , n430725 , n85362 , n430727 , n430728 , 
 n85365 , n85366 , n430731 , n430732 , n85369 , n85370 , n85371 , n430736 , n430737 , n85374 , 
 n85375 , n430740 , n430741 , n85378 , n85379 , n430744 , n430745 , n85382 , n430747 , n85384 , 
 n85385 , n430750 , n85387 , n430752 , n85389 , n430754 , n85391 , n430756 , n85393 , n430758 , 
 n85395 , n85396 , n430761 , n430762 , n85399 , n430764 , n85401 , n430766 , n430767 , n85404 , 
 n430769 , n430770 , n85407 , n430772 , n85409 , n85410 , n85411 , n430776 , n85413 , n85414 , 
 n85415 , n85416 , n85417 , n85418 , n430783 , n430784 , n85421 , n430786 , n85423 , n85424 , 
 n85425 , n430790 , n430791 , n85428 , n430793 , n85430 , n85431 , n85432 , n430797 , n85434 , 
 n430799 , n85436 , n430801 , n85438 , n430803 , n85440 , n85441 , n85442 , n430807 , n430808 , 
 n85445 , n85446 , n85447 , n430812 , n430813 , n85450 , n85451 , n85452 , n430817 , n430818 , 
 n85455 , n85456 , n85457 , n430822 , n430823 , n85460 , n85461 , n85462 , n430827 , n85464 , 
 n85465 , n85466 , n85467 , n85468 , n85469 , n85470 , n85471 , n85472 , n85473 , n430838 , 
 n430839 , n85476 , n85477 , n85478 , n85479 , n430844 , n430845 , n85482 , n85483 , n430848 , 
 n430849 , n430850 , n85487 , n85488 , n430853 , n85490 , n430855 , n430856 , n85493 , n85494 , 
 n430859 , n430860 , n85497 , n430862 , n430863 , n430864 , n85501 , n430866 , n85503 , n85504 , 
 n430869 , n85506 , n430871 , n430872 , n430873 , n430874 , n85511 , n430876 , n430877 , n85514 , 
 n430879 , n430880 , n85517 , n430882 , n85519 , n85520 , n430885 , n85522 , n85523 , n85524 , 
 n85525 , n430890 , n430891 , n85528 , n430893 , n85530 , n430895 , n85532 , n85533 , n430898 , 
 n430899 , n85536 , n85537 , n430902 , n85539 , n430904 , n85541 , n430906 , n430907 , n85544 , 
 n430909 , n430910 , n85547 , n430912 , n85549 , n85550 , n430915 , n85552 , n85553 , n85554 , 
 n430919 , n85556 , n430921 , n430922 , n85559 , n430924 , n430925 , n85562 , n85563 , n85564 , 
 n430929 , n430930 , n85567 , n85568 , n85569 , n85571 , n430935 , n430936 , n430937 , n85575 , 
 n430939 , n85577 , n85578 , n430942 , n430943 , n430944 , n85582 , n430946 , n85584 , n430948 , 
 n430949 , n430950 , n430951 , n430952 , n430953 , n430954 , n85592 , n430956 , n430957 , n430958 , 
 n85596 , n430960 , n85598 , n430962 , n85600 , n430964 , n430965 , n430966 , n85604 , n430968 , 
 n430969 , n430970 , n430971 , n430972 , n85610 , n430974 , n430975 , n430976 , n85614 , n430978 , 
 n430979 , n430980 , n430981 , n430982 , n85620 , n430984 , n85622 , n430986 , n85624 , n430988 , 
 n430989 , n430990 , n430991 , n430992 , n85630 , n430994 , n85632 , n430996 , n430997 , n430998 , 
 n430999 , n431000 , n431001 , n431002 , n431003 , n431004 , n431005 , n431006 , n431007 , n85674 , 
 n431009 , n431010 , n85677 , n85678 , n85679 , n85680 , n85681 , n431016 , n431017 , n85684 , 
 n431019 , n431020 , n431021 , n431022 , n85689 , n431024 , n431025 , n431026 , n431027 , n431028 , 
 n85695 , n85696 , n85698 , n431032 , n85700 , n85701 , n85702 , n85703 , n85704 , n85705 , 
 n85706 , n85707 , n431041 , n85709 , n431043 , n85711 , n431045 , n85713 , n431047 , n85715 , 
 n85716 , n431050 , n431051 , n85719 , n431053 , n431054 , n85722 , n431056 , n431057 , n85725 , 
 n85726 , n431060 , n431061 , n85729 , n431063 , n431064 , n85732 , n431066 , n85734 , n85735 , 
 n85736 , n85737 , n85738 , n431072 , n431073 , n85741 , n431075 , n85743 , n85744 , n85745 , 
 n431079 , n85747 , n431081 , n85749 , n85750 , n431084 , n85752 , n431086 , n85754 , n431088 , 
 n431089 , n431090 , n85758 , n431092 , n431093 , n85761 , n431095 , n431096 , n431097 , n85765 , 
 n431099 , n431100 , n85768 , n431102 , n85770 , n85771 , n85772 , n85773 , n85774 , n85775 , 
 n85776 , n85777 , n85778 , n85779 , n85780 , n431114 , n85782 , n85783 , n85784 , n85785 , 
 n85786 , n85787 , n85788 , n431122 , n85790 , n85791 , n431125 , n85793 , n431127 , n85795 , 
 n85796 , n85797 , n431131 , n85799 , n85800 , n85801 , n85802 , n431136 , n431137 , n431138 , 
 n85806 , n431140 , n85808 , n85809 , n431143 , n431144 , n85812 , n431146 , n431147 , n85815 , 
 n431149 , n431150 , n431151 , n431152 , n431153 , n431154 , n85822 , n431156 , n431157 , n85825 , 
 n431159 , n431160 , n85828 , n431162 , n431163 , n85831 , n85832 , n85833 , n85834 , n431168 , 
 n85836 , n431170 , n85838 , n85839 , n431173 , n431174 , n85842 , n431176 , n431177 , n85845 , 
 n431179 , n431180 , n85848 , n431182 , n85850 , n85851 , n431185 , n431186 , n85854 , n431188 , 
 n431189 , n85857 , n431191 , n85859 , n85860 , n85861 , n85862 , n85863 , n85864 , n85865 , 
 n85866 , n85867 , n431201 , n431202 , n85870 , n431204 , n85872 , n85873 , n431207 , n431208 , 
 n85876 , n431210 , n431211 , n431212 , n85880 , n85881 , n431215 , n431216 , n85884 , n431218 , 
 n85886 , n431220 , n85888 , n85889 , n431223 , n85891 , n431225 , n85893 , n85894 , n431228 , 
 n431229 , n85897 , n431231 , n431232 , n85900 , n431234 , n431235 , n431236 , n85904 , n431238 , 
 n431239 , n85907 , n431241 , n431242 , n85910 , n431244 , n85912 , n85913 , n85914 , n85915 , 
 n85916 , n85917 , n85918 , n85919 , n85920 , n85921 , n85922 , n85923 , n85924 , n85925 , 
 n85926 , n85927 , n431261 , n85929 , n431263 , n431264 , n85932 , n85933 , n431267 , n431268 , 
 n431269 , n431270 , n85938 , n85939 , n431273 , n85941 , n431275 , n431276 , n85960 , n85961 , 
 n431279 , n85963 , n85964 , n431282 , n85966 , n85967 , n85968 , n431286 , n85970 , n431288 , 
 n85972 , n85973 , n431291 , n431292 , n85976 , n431294 , n431295 , n85979 , n431297 , n431298 , 
 n431299 , n85983 , n431301 , n85985 , n431303 , n431304 , n85988 , n431306 , n85990 , n431308 , 
 n85992 , n85993 , n431311 , n431312 , n85996 , n431314 , n431315 , n85999 , n431317 , n431318 , 
 n86002 , n86003 , n431321 , n431322 , n86006 , n431324 , n431325 , n86009 , n431327 , n431328 , 
 n86012 , n86013 , n86014 , n86015 , n431333 , n431334 , n86018 , n86019 , n86020 , n86021 , 
 n86022 , n431340 , n431341 , n86025 , n431343 , n86027 , n86028 , n86029 , n431347 , n86031 , 
 n431349 , n431350 , n86034 , n431352 , n86036 , n431354 , n86038 , n86039 , n431357 , n431358 , 
 n86042 , n431360 , n431361 , n86045 , n431363 , n431364 , n86048 , n431366 , n431367 , n86051 , 
 n431369 , n431370 , n86054 , n431372 , n86056 , n431374 , n86058 , n431376 , n86060 , n86061 , 
 n431379 , n431380 , n431381 , n431382 , n431383 , n86067 , n431385 , n431386 , n86070 , n86071 , 
 n431389 , n431390 , n86074 , n431392 , n431393 , n86077 , n431395 , n431396 , n86080 , n431398 , 
 n431399 , n86083 , n431401 , n431402 , n86086 , n431404 , n86088 , n86089 , n431407 , n86097 , 
 n431409 , n86099 , n431411 , n86101 , n431413 , n431414 , n86104 , n86105 , n431417 , n86107 , 
 n431419 , n86109 , n86110 , n431422 , n86112 , n431424 , n431425 , n86115 , n431427 , n86117 , 
 n86118 , n86119 , n86120 , n86121 , n86122 , n86123 , n86124 , n431436 , n86126 , n431438 , 
 n86128 , n431440 , n431441 , n431442 , n431443 , n86133 , n86134 , n431446 , n431447 , n86137 , 
 n431449 , n431450 , n86140 , n431452 , n86142 , n431454 , n86144 , n431456 , n431457 , n431458 , 
 n86148 , n431460 , n86150 , n431462 , n431463 , n86153 , n86154 , n86155 , n86156 , n431468 , 
 n431469 , n86159 , n431471 , n86161 , n86162 , n431474 , n86164 , n431476 , n86166 , n431478 , 
 n86168 , n431480 , n431481 , n86171 , n86172 , n431484 , n86174 , n431486 , n86176 , n431488 , 
 n431489 , n86179 , n431491 , n431492 , n431493 , n86183 , n431495 , n431496 , n86186 , n86189 , 
 n431499 , n86191 , n431501 , n431502 , n431503 , n431504 , n86199 , n431506 , n431507 , n86202 , 
 n431509 , n86206 , n86207 , n431512 , n86209 , n431514 , n431515 , n431516 , n431517 , n86217 , 
 n431519 , n431520 , n86220 , n431522 , n86222 , n86223 , n86224 , n86225 , n86226 , n431528 , 
 n431529 , n431530 , n86230 , n431532 , n86232 , n431534 , n86234 , n86235 , n431537 , n431538 , 
 n86238 , n431540 , n431541 , n86241 , n431543 , n431544 , n86244 , n86245 , n431547 , n431548 , 
 n86248 , n431550 , n431551 , n86251 , n431553 , n86253 , n431555 , n86255 , n431557 , n86257 , 
 n86258 , n431560 , n431561 , n86261 , n86262 , n431564 , n86264 , n86265 , n431567 , n431568 , 
 n86268 , n431570 , n86270 , n431572 , n431573 , n86273 , n431575 , n86275 , n86276 , n86277 , 
 n86278 , n86279 , n86280 , n431582 , n431583 , n86283 , n431585 , n431586 , n86286 , n431588 , 
 n431589 , n86289 , n86290 , n431592 , n86292 , n86293 , n431595 , n431596 , n431597 , n86297 , 
 n86298 , n431600 , n86300 , n86301 , n86302 , n86303 , n86304 , n86305 , n431607 , n86307 , 
 n431609 , n431610 , n86333 , n431612 , n431613 , n86336 , n86337 , n86338 , n86339 , n86340 , 
 n86341 , n431620 , n86343 , n431622 , n86345 , n431624 , n86347 , n86348 , n431627 , n431628 , 
 n86351 , n431630 , n431631 , n86354 , n431633 , n431634 , n86357 , n86358 , n431637 , n431638 , 
 n86361 , n86362 , n86363 , n86364 , n86365 , n431644 , n431645 , n86368 , n431647 , n86370 , 
 n431649 , n431650 , n431651 , n86384 , n431653 , n86386 , n431655 , n86388 , n86389 , n431658 , 
 n86391 , n431660 , n431661 , n86394 , n431663 , n86396 , n86397 , n431666 , n431667 , n431668 , 
 n431669 , n86402 , n431671 , n431672 , n86405 , n431674 , n431675 , n86408 , n86409 , n86410 , 
 n86411 , n431680 , n86413 , n431682 , n86415 , n86416 , n431685 , n431686 , n86419 , n431688 , 
 n431689 , n86422 , n431691 , n431692 , n431693 , n86426 , n431695 , n86428 , n86429 , n86430 , 
 n86431 , n86432 , n86433 , n86434 , n86435 , n86436 , n86437 , n86438 , n86439 , n86440 , 
 n86441 , n86442 , n86443 , n86444 , n86445 , n86446 , n86447 , n431716 , n431717 , n86450 , 
 n431719 , n86452 , n86453 , n431722 , n86455 , n431724 , n86457 , n86458 , n431727 , n86460 , 
 n431729 , n86462 , n86463 , n431732 , n431733 , n86466 , n431735 , n431736 , n86469 , n431738 , 
 n431739 , n431740 , n86473 , n431742 , n431743 , n86476 , n431745 , n86478 , n86479 , n86480 , 
 n431749 , n431750 , n86483 , n431752 , n86485 , n86486 , n431755 , n86488 , n431757 , n86490 , 
 n431759 , n86492 , n86493 , n431762 , n431763 , n86496 , n431765 , n431766 , n86499 , n431768 , 
 n431769 , n86502 , n86503 , n431772 , n431773 , n86506 , n431775 , n431776 , n86509 , n431778 , 
 n86511 , n431780 , n86513 , n431782 , n86515 , n86516 , n431785 , n431786 , n86519 , n431788 , 
 n431789 , n86522 , n431791 , n431792 , n86525 , n86526 , n431795 , n431796 , n86529 , n86530 , 
 n86531 , n86532 , n86533 , n431802 , n431803 , n86536 , n431805 , n86538 , n86539 , n86540 , 
 n86541 , n86542 , n431811 , n86544 , n431813 , n86546 , n431815 , n86548 , n86549 , n86550 , 
 n86551 , n86552 , n86553 , n86554 , n86555 , n86556 , n86557 , n86558 , n431827 , n86560 , 
 n431829 , n86562 , n431831 , n86564 , n431833 , n431834 , n86567 , n86568 , n431837 , n86570 , 
 n86571 , n86572 , n86573 , n431842 , n431843 , n86576 , n86577 , n86578 , n431847 , n86580 , 
 n86581 , n86582 , n431851 , n431852 , n86585 , n431854 , n431855 , n86588 , n431857 , n431858 , 
 n86591 , n86592 , n86593 , n431862 , n431863 , n86596 , n431865 , n431866 , n86599 , n86600 , 
 n86601 , n86602 , n431871 , n431872 , n86605 , n431874 , n431875 , n86608 , n431877 , n431878 , 
 n431879 , n86612 , n431881 , n86614 , n86615 , n431884 , n431885 , n86618 , n431887 , n431888 , 
 n86621 , n431890 , n86623 , n86624 , n86625 , n86626 , n86627 , n431896 , n86629 , n86630 , 
 n86631 , n86632 , n86633 , n86634 , n86635 , n86636 , n431905 , n86638 , n86639 , n86640 , 
 n86641 , n86642 , n431911 , n86644 , n86645 , n86646 , n86647 , n431916 , n86649 , n86650 , 
 n86651 , n86652 , n86653 , n86654 , n86655 , n431924 , n86657 , n431926 , n431927 , n431928 , 
 n86661 , n431930 , n86663 , n86664 , n431933 , n431934 , n86667 , n431936 , n431937 , n86670 , 
 n431939 , n86672 , n86673 , n86674 , n86675 , n86676 , n86677 , n86678 , n86679 , n86680 , 
 n86681 , n86682 , n431951 , n86684 , n86685 , n86686 , n86687 , n86688 , n431957 , n431958 , 
 n431959 , n86714 , n86715 , n86716 , n86717 , n86718 , n86719 , n86720 , n86721 , n86722 , 
 n86723 , n86724 , n86725 , n431972 , n86727 , n431974 , n86729 , n86730 , n86731 , n86732 , 
 n431979 , n86734 , n431981 , n86736 , n431983 , n86738 , n86739 , n86740 , n431987 , n86742 , 
 n431989 , n431990 , n86745 , n86746 , n86747 , n86748 , n86749 , n431996 , n431997 , n86752 , 
 n431999 , n432000 , n432001 , n86756 , n432003 , n86758 , n432005 , n432006 , n86761 , n432008 , 
 n86763 , n86764 , n432011 , n86766 , n432013 , n86768 , n432015 , n432016 , n86771 , n432018 , 
 n432019 , n86774 , n86775 , n86776 , n432023 , n432024 , n86779 , n432026 , n86781 , n86782 , 
 n432029 , n432030 , n86785 , n432032 , n432033 , n86788 , n432035 , n432036 , n86791 , n432038 , 
 n432039 , n86794 , n432041 , n86796 , n432043 , n432044 , n86799 , n432046 , n432047 , n432048 , 
 n86803 , n432050 , n86805 , n86806 , n432053 , n432054 , n86809 , n86810 , n432057 , n86812 , 
 n432059 , n86814 , n432061 , n432062 , n432063 , n86818 , n86819 , n432066 , n86821 , n86822 , 
 n432069 , n432070 , n86825 , n432072 , n432073 , n86828 , n86829 , n432076 , n86831 , n86832 , 
 n432079 , n432080 , n432081 , n86836 , n86837 , n432084 , n432085 , n86840 , n432087 , n432088 , 
 n432089 , n432090 , n86863 , n86866 , n86867 , n432094 , n432095 , n86870 , n432097 , n432098 , 
 n86873 , n86874 , n86875 , n86876 , n86877 , n86878 , n86879 , n86880 , n86881 , n86882 , 
 n86883 , n86884 , n86885 , n86886 , n86887 , n432114 , n86889 , n432116 , n86891 , n86892 , 
 n86893 , n86894 , n432121 , n86896 , n432123 , n86898 , n86899 , n86900 , n86901 , n86902 , 
 n432129 , n86904 , n86905 , n86907 , n432133 , n432134 , n86910 , n86911 , n86912 , n86913 , 
 n86914 , n432140 , n86916 , n432142 , n432143 , n86919 , n86920 , n86921 , n86922 , n86923 , 
 n432149 , n432150 , n86926 , n432152 , n432153 , n86929 , n432155 , n432156 , n86932 , n86933 , 
 n86934 , n86935 , n432161 , n432162 , n86938 , n432164 , n432165 , n86941 , n432167 , n432168 , 
 n86944 , n86945 , n86946 , n86947 , n86948 , n86949 , n432175 , n432176 , n86952 , n432178 , 
 n86954 , n86955 , n86956 , n86957 , n432183 , n432184 , n86960 , n432186 , n86962 , n432188 , 
 n86964 , n432190 , n432191 , n86967 , n432193 , n432194 , n432195 , n432196 , n86972 , n432198 , 
 n86974 , n432200 , n432201 , n86977 , n86978 , n86979 , n86980 , n86981 , n86982 , n432208 , 
 n86984 , n432210 , n86986 , n432212 , n86988 , n432214 , n432215 , n86991 , n86992 , n432218 , 
 n86994 , n432220 , n86996 , n86997 , n432223 , n86999 , n432225 , n432226 , n87002 , n432228 , 
 n432229 , n87005 , n87006 , n87007 , n432233 , n432234 , n87010 , n87011 , n87012 , n87013 , 
 n87014 , n87015 , n87016 , n87017 , n87018 , n87019 , n87020 , n432246 , n432247 , n432248 , 
 n87047 , n87048 , n87049 , n87050 , n87051 , n432254 , n432255 , n87054 , n432257 , n432258 , 
 n432259 , n432260 , n87062 , n432262 , n432263 , n87065 , n432265 , n432266 , n87068 , n432268 , 
 n432269 , n87071 , n432271 , n87073 , n432273 , n432274 , n87076 , n432276 , n432277 , n87079 , 
 n432279 , n432280 , n87082 , n432282 , n432283 , n87085 , n432285 , n432286 , n87088 , n432288 , 
 n87090 , n432290 , n432291 , n87093 , n432293 , n432294 , n87096 , n432296 , n432297 , n87099 , 
 n432299 , n87101 , n432301 , n87103 , n87104 , n432304 , n432305 , n87107 , n432307 , n432308 , 
 n87110 , n432310 , n432311 , n87113 , n432313 , n87115 , n432315 , n432316 , n87118 , n432318 , 
 n432319 , n87121 , n87122 , n432322 , n87124 , n432324 , n432325 , n432326 , n87128 , n432328 , 
 n432329 , n87131 , n432331 , n87133 , n87134 , n432334 , n87136 , n432336 , n432337 , n87150 , 
 n87151 , n87152 , n87153 , n432342 , n432343 , n432344 , n87157 , n432346 , n87159 , n87160 , 
 n432349 , n87162 , n432351 , n87164 , n432353 , n432354 , n87167 , n432356 , n432357 , n87170 , 
 n432359 , n87172 , n432361 , n432362 , n87175 , n432364 , n87177 , n87178 , n432367 , n432368 , 
 n87181 , n432370 , n432371 , n87184 , n432373 , n432374 , n87187 , n87188 , n87189 , n432378 , 
 n87191 , n87192 , n87193 , n87194 , n87195 , n87196 , n87197 , n87198 , n87199 , n87200 , 
 n87201 , n87202 , n87203 , n432392 , n87205 , n87206 , n87207 , n432396 , n432397 , n432398 , 
 n432399 , n87237 , n87238 , n87239 , n432403 , n432404 , n87242 , n432406 , n432407 , n87245 , 
 n432409 , n432410 , n87248 , n432412 , n432413 , n87251 , n87252 , n432416 , n432417 , n87255 , 
 n432419 , n432420 , n87258 , n87261 , n432423 , n432424 , n87264 , n432426 , n87266 , n87267 , 
 n87268 , n87270 , n432431 , n87272 , n87273 , n432434 , n87275 , n432436 , n87277 , n87278 , 
 n87279 , n87280 , n87281 , n87282 , n87283 , n87284 , n87285 , n432446 , n87287 , n87288 , 
 n432449 , n432450 , n87291 , n432452 , n432453 , n432454 , n87295 , n87296 , n87297 , n87298 , 
 n87299 , n87300 , n87301 , n87302 , n87303 , n87304 , n87305 , n432466 , n87307 , n87308 , 
 n432469 , n432470 , n87311 , n87312 , n432473 , n432474 , n432475 , n87316 , n432477 , n87318 , 
 n87319 , n432480 , n432481 , n87322 , n432483 , n432484 , n87325 , n432486 , n432487 , n87328 , 
 n87329 , n87330 , n432491 , n432492 , n87333 , n432494 , n432495 , n87336 , n87337 , n432498 , 
 n87339 , n432500 , n432501 , n87342 , n87343 , n432504 , n87345 , n87346 , n432507 , n87348 , 
 n432509 , n432510 , n87351 , n432512 , n432513 , n87354 , n87355 , n432516 , n432517 , n432518 , 
 n87359 , n432520 , n87364 , n87365 , n87366 , n87368 , n87369 , n87370 , n87371 , n87372 , 
 n87373 , n432530 , n87375 , n87376 , n87377 , n87378 , n87379 , n432536 , n432537 , n87382 , 
 n432539 , n432540 , n87385 , n87386 , n432543 , n87388 , n432545 , n432546 , n87391 , n87392 , 
 n432549 , n432550 , n432551 , n87396 , n432553 , n87398 , n87399 , n432556 , n87401 , n432558 , 
 n87403 , n87404 , n432561 , n87406 , n432563 , n432564 , n87409 , n432566 , n432567 , n87412 , 
 n87413 , n432570 , n87415 , n87416 , n87417 , n432574 , n87419 , n432576 , n432577 , n87422 , 
 n87423 , n87424 , n87425 , n87426 , n87427 , n87428 , n87429 , n87430 , n87431 , n87435 , 
 n87437 , n87438 , n87439 , n87440 , n87441 , n87442 , n432595 , n87458 , n432597 , n87460 , 
 n87461 , n432600 , n87463 , n432602 , n87465 , n432604 , n432605 , n87468 , n432607 , n432608 , 
 n432609 , n87472 , n87473 , n432612 , n87475 , n87476 , n432615 , n432616 , n87479 , n87480 , 
 n87481 , n87482 , n87483 , n87484 , n432623 , n432624 , n87487 , n432626 , n432627 , n87490 , 
 n432629 , n432630 , n87499 , n87500 , n87501 , n87502 , n87503 , n87504 , n87505 , n87506 , 
 n87507 , n87508 , n87509 , n432642 , n87511 , n432644 , n432645 , n87514 , n432647 , n432648 , 
 n432649 , n87518 , n87519 , n432652 , n432653 , n87522 , n432655 , n432656 , n87525 , n432658 , 
 n432659 , n432660 , n87531 , n432662 , n432663 , n432664 , n87535 , n432666 , n87537 , n432668 , 
 n432669 , n432670 , n87541 , n432672 , n87543 , n432674 , n432675 , n432676 , n87547 , n432678 , 
 n432679 , n432680 , n87551 , n432682 , n432683 , n432684 , n87555 , n432686 , n87557 , n432688 , 
 n432689 , n432690 , n432691 , n432692 , n87563 , n432694 , n432695 , n432696 , n432697 , n432698 , 
 n87569 , n432700 , n432701 , n432702 , n87573 , n432704 , n432705 , n432706 , n87577 , n432708 , 
 n87579 , n432710 , n87581 , n432712 , n432713 , n432714 , n87585 , n432716 , n87587 , n432718 , 
 n432719 , n432720 , n432721 , n432722 , n432723 , n432724 , n432725 , n432726 , n432727 , n432728 , 
 n432729 , n432730 , n432731 , n432732 , n432733 , n432734 , n432735 , n432736 , n432737 , n432738 , 
 n432739 , n432740 , n432741 , n432742 , n432743 , n432744 , n432745 , n432746 , n432747 , n432748 , 
 n432749 , n432750 , n432751 , n432752 , n432753 , n432754 , n432755 , n432756 , n432757 , n432758 , 
 n432759 , n432760 , n432761 , n432762 , n432763 , n432764 , n432765 , n432766 , n432767 , n432768 , 
 n432769 , n432770 , n432771 , n432772 , n432773 , n432774 , n432775 , n432776 , n432777 , n432778 , 
 n432779 , n432780 , n432781 , n432782 , n432783 , n432784 , n432785 , n432786 , n432787 , n432788 , 
 n432789 , n432790 , n432791 , n432792 , n432793 , n432794 , n432795 , n432796 , n432797 , n432798 , 
 n432799 , n432800 , n432801 , n432802 , n432803 , n432804 , n432805 , n432806 , n432807 , n432808 , 
 n432809 , n432810 , n432811 , n432812 , n432813 , n432814 , n432815 , n432816 , n432817 , n432818 , 
 n432819 , n432820 , n432821 , n432822 , n432823 , n432824 , n432825 , n432826 , n432827 , n432828 , 
 n432829 , n432830 , n432831 , n432832 , n432833 , n432834 , n432835 , n432836 , n432837 , n432838 , 
 n432839 , n432840 , n432841 , n432842 , n432843 , n432844 , n432845 , n432846 , n432847 , n432848 , 
 n432849 , n432850 , n432851 , n432852 , n432853 , n432854 , n432855 , n432856 , n432857 , n432858 , 
 n432859 , n432860 , n432861 , n432862 , n432863 , n432864 , n432865 , n432866 , n432867 , n432868 , 
 n432869 , n432870 , n432871 , n432872 , n432873 , n432874 , n432875 , n432876 , n432877 , n432878 , 
 n432879 , n432880 , n432881 , n432882 , n432883 , n432884 , n432885 , n432886 , n432887 , n432888 , 
 n432889 , n432890 , n432891 , n432892 , n432893 , n432894 , n432895 , n432896 , n432897 , n432898 , 
 n432899 , n432900 , n432901 , n432902 , n432903 , n432904 , n432905 , n432906 , n432907 , n432908 , 
 n432909 , n432910 , n432911 , n432912 , n432913 , n432914 , n432915 , n432916 , n432917 , n432918 , 
 n432919 , n432920 , n432921 , n432922 , n432923 , n432924 , n432925 , n432926 , n432927 , n432928 , 
 n432929 , n432930 , n432931 , n432932 , n432933 , n432934 , n432935 , n432936 , n432937 , n432938 , 
 n432939 , n432940 , n432941 , n432942 , n432943 , n432944 , n432945 , n432946 , n432947 , n432948 , 
 n432949 , n432950 , n432951 , n432952 , n432953 , n432954 , n432955 , n432956 , n432957 , n432958 , 
 n432959 , n432960 , n432961 , n432962 , n432963 , n432964 , n432965 , n432966 , n432967 , n432968 , 
 n432969 , n432970 , n432971 , n432972 , n432973 , n432974 , n432975 , n432976 , n432977 , n432978 , 
 n432979 , n432980 , n432981 , n432982 , n432983 , n432984 , n432985 , n432986 , n432987 , n432988 , 
 n432989 , n432990 , n432991 , n432992 , n432993 , n432994 , n432995 , n432996 , n432997 , n432998 , 
 n432999 , n433000 , n433001 , n433002 , n433003 , n433004 , n433005 , n433006 , n433007 , n433008 , 
 n433009 , n433010 , n433011 , n433012 , n433013 , n433014 , n433015 , n433016 , n433017 , n433018 , 
 n433019 , n433020 , n433021 , n433022 , n433023 , n433024 , n433025 , n433026 , n433027 , n433028 , 
 n433029 , n433030 , n433031 , n433032 , n433033 , n433034 , n433035 , n433036 , n433037 , n433038 , 
 n433039 , n433040 , n433041 , n433042 , n433043 , n433044 , n433045 , n433046 , n433047 , n433048 , 
 n433049 , n433050 , n433051 , n433052 , n433053 , n433054 , n433055 , n433056 , n433057 , n433058 , 
 n433059 , n433060 , n433061 , n433062 , n433063 , n433064 , n433065 , n433066 , n433067 , n433068 , 
 n433069 , n433070 , n433071 , n433072 , n433073 , n433074 , n433075 , n433076 , n433077 , n433078 , 
 n433079 , n433080 , n433081 , n433082 , n433083 , n433084 , n433085 , n433086 , n433087 , n433088 , 
 n433089 , n433090 , n433091 , n433092 , n433093 , n433094 , n433095 , n433096 , n433097 , n433098 , 
 n433099 , n433100 , n433101 , n433102 , n433103 , n433104 , n433105 , n433106 , n433107 , n433108 , 
 n433109 , n433110 , n433111 , n433112 , n433113 , n433114 , n433115 , n433116 , n433117 , n433118 , 
 n433119 , n433120 , n433121 , n433122 , n433123 , n433124 , n433125 , n433126 , n433127 , n433128 , 
 n433129 , n433130 , n433131 , n433132 , n433133 , n433134 , n433135 , n433136 , n433137 , n433138 , 
 n433139 , n433140 , n433141 , n433142 , n433143 , n433144 , n433145 , n433146 , n433147 , n433148 , 
 n433149 , n433150 , n433151 , n433152 , n433153 , n433154 , n433155 , n433156 , n433157 , n433158 , 
 n433159 , n433160 , n433161 , n433162 , n433163 , n433164 , n433165 , n433166 , n433167 , n433168 , 
 n433169 , n433170 , n433171 , n433172 , n433173 , n433174 , n433175 , n433176 , n433177 , n433178 , 
 n433179 , n433180 , n433181 , n433182 , n433183 , n433184 , n433185 , n433186 , n433187 , n433188 , 
 n433189 , n433190 , n433191 , n433192 , n433193 , n433194 , n433195 , n433196 , n433197 , n433198 , 
 n433199 , n433200 , n433201 , n433202 , n433203 , n433204 , n433205 , n433206 , n433207 , n433208 , 
 n433209 , n433210 , n433211 , n433212 , n433213 , n433214 , n433215 , n433216 , n433217 , n433218 , 
 n433219 , n433220 , n433221 , n433222 , n433223 , n433224 , n433225 , n433226 , n433227 , n433228 , 
 n433229 , n433230 , n433231 , n433232 , n433233 , n433234 , n433235 , n433236 , n433237 , n433238 , 
 n433239 , n433240 , n433241 , n433242 , n433243 , n433244 , n433245 , n433246 , n433247 , n433248 , 
 n433249 , n433250 , n433251 , n433252 , n433253 , n433254 , n433255 , n433256 , n433257 , n433258 , 
 n433259 , n433260 , n433261 , n433262 , n433263 , n433264 , n433265 , n433266 , n433267 , n433268 , 
 n433269 , n433270 , n433271 , n433272 , n433273 , n433274 , n433275 , n433276 , n433277 , n433278 , 
 n433279 , n433280 , n433281 , n433282 , n433283 , n433284 , n433285 , n433286 , n433287 , n433288 , 
 n433289 , n433290 , n433291 , n433292 , n433293 , n433294 , n433295 , n433296 , n433297 , n433298 , 
 n433299 , n433300 , n433301 , n433302 , n433303 , n433304 , n433305 , n433306 , n433307 , n433308 , 
 n433309 , n433310 , n433311 , n433312 , n433313 , n433314 , n433315 , n433316 , n433317 , n433318 , 
 n433319 , n433320 , n433321 , n433322 , n433323 , n433324 , n433325 , n433326 , n433327 , n433328 , 
 n433329 , n433330 , n433331 , n433332 , n433333 , n433334 , n433335 , n433336 , n433337 , n433338 , 
 n433339 , n433340 , n433341 , n433342 , n433343 , n433344 , n433345 , n433346 , n433347 , n433348 , 
 n433349 , n433350 , n433351 , n433352 , n433353 , n433354 , n433355 , n433356 , n433357 , n433358 , 
 n433359 , n433360 , n433361 , n433362 , n433363 , n433364 , n433365 , n433366 , n433367 , n433368 , 
 n433369 , n433370 , n433371 , n433372 , n433373 , n433374 , n433375 , n433376 , n433377 , n433378 , 
 n433379 , n433380 , n433381 , n433382 , n433383 , n433384 , n433385 , n433386 , n433387 , n433388 , 
 n433389 , n433390 , n433391 , n433392 , n433393 , n433394 , n433395 , n433396 , n433397 , n433398 , 
 n433399 , n433400 , n433401 , n433402 , n433403 , n433404 , n433405 , n433406 , n433407 , n433408 , 
 n433409 , n433410 , n433411 , n433412 , n433413 , n433414 , n433415 , n433416 , n433417 , n433418 , 
 n433419 , n433420 , n433421 , n433422 , n433423 , n433424 , n433425 , n433426 , n433427 , n433428 , 
 n433429 , n433430 , n433431 , n433432 , n433433 , n433434 , n433435 , n433436 , n433437 , n433438 , 
 n433439 , n433440 , n433441 , n433442 , n433443 , n433444 , n433445 , n433446 , n433447 , n433448 , 
 n433449 , n433450 , n433451 , n433452 , n433453 , n433454 , n433455 , n433456 , n433457 , n433458 , 
 n433459 , n433460 , n433461 , n433462 , n433463 , n433464 , n433465 , n433466 , n433467 , n433468 , 
 n433469 , n433470 , n433471 , n433472 , n433473 , n433474 , n433475 , n433476 , n433477 , n433478 , 
 n433479 , n433480 , n433481 , n433482 , n433483 , n433484 , n433485 , n433486 , n433487 , n433488 , 
 n433489 , n433490 , n433491 , n433492 , n433493 , n433494 , n433495 , n433496 , n433497 , n433498 , 
 n433499 , n433500 , n433501 , n433502 , n433503 , n433504 , n433505 , n433506 , n433507 , n433508 , 
 n433509 , n433510 , n433511 , n433512 , n433513 , n433514 , n433515 , n433516 , n433517 , n433518 , 
 n433519 , n433520 , n433521 , n433522 , n433523 , n433524 , n433525 , n433526 , n433527 , n433528 , 
 n433529 , n433530 , n433531 , n433532 , n433533 , n433534 , n433535 , n433536 , n433537 , n433538 , 
 n433539 , n433540 , n433541 , n433542 , n433543 , n433544 , n433545 , n433546 , n433547 , n433548 , 
 n433549 , n433550 , n433551 , n433552 , n433553 , n433554 , n433555 , n433556 , n433557 , n433558 , 
 n433559 , n433560 , n433561 , n433562 , n433563 , n433564 , n433565 , n433566 , n433567 , n433568 , 
 n433569 , n433570 , n433571 , n433572 , n433573 , n433574 , n433575 , n433576 , n433577 , n433578 , 
 n433579 , n433580 , n433581 , n433582 , n433583 , n433584 , n433585 , n433586 , n433587 , n433588 , 
 n433589 , n433590 , n433591 , n433592 , n433593 , n433594 , n433595 , n433596 , n433597 , n433598 , 
 n433599 , n433600 , n433601 , n433602 , n433603 , n433604 , n433605 , n433606 , n433607 , n433608 , 
 n433609 , n433610 , n433611 , n433612 , n433613 , n433614 , n433615 , n433616 , n433617 , n433618 , 
 n433619 , n433620 , n433621 , n433622 , n433623 , n433624 , n433625 , n433626 , n433627 , n433628 , 
 n433629 , n433630 , n433631 , n433632 , n433633 , n433634 , n433635 , n433636 , n433637 , n433638 , 
 n433639 , n433640 , n433641 , n433642 , n433643 , n433644 , n433645 , n433646 , n433647 , n433648 , 
 n433649 , n433650 , n433651 , n433652 , n433653 , n433654 , n433655 , n433656 , n433657 , n433658 , 
 n433659 , n433660 , n433661 , n433662 , n433663 , n433664 , n433665 , n433666 , n433667 , n433668 , 
 n433669 , n433670 , n433671 , n433672 , n433673 , n433674 , n433675 , n433676 , n433677 , n433678 , 
 n433679 , n433680 , n433681 , n433682 , n433683 , n433684 , n433685 , n433686 , n433687 , n433688 , 
 n433689 , n433690 , n433691 , n433692 , n433693 , n433694 , n433695 , n433696 , n433697 , n433698 , 
 n433699 , n433700 , n433701 , n433702 , n433703 , n433704 , n433705 , n433706 , n433707 , n433708 , 
 n433709 , n433710 , n433711 , n433712 , n433713 , n433714 , n433715 , n433716 , n433717 , n433718 , 
 n433719 , n433720 , n433721 , n433722 , n433723 , n433724 , n433725 , n433726 , n433727 , n433728 , 
 n433729 , n433730 , n433731 , n433732 , n433733 , n433734 , n433735 , n433736 , n433737 , n433738 , 
 n433739 , n433740 , n433741 , n433742 , n433743 , n433744 , n433745 , n433746 , n433747 , n433748 , 
 n433749 , n433750 , n433751 , n433752 , n433753 , n433754 , n433755 , n433756 , n433757 , n433758 , 
 n433759 , n433760 , n433761 , n433762 , n433763 , n433764 , n433765 , n433766 , n433767 , n433768 , 
 n433769 , n433770 , n433771 , n433772 , n433773 , n433774 , n433775 , n433776 , n433777 , n433778 , 
 n433779 , n433780 , n433781 , n433782 , n433783 , n433784 , n433785 , n433786 , n433787 , n433788 , 
 n433789 , n433790 , n433791 , n433792 , n433793 , n433794 , n433795 , n433796 , n433797 , n433798 , 
 n433799 , n433800 , n433801 , n433802 , n433803 , n433804 , n433805 , n433806 , n433807 , n433808 , 
 n433809 , n433810 , n433811 , n433812 , n433813 , n433814 , n433815 , n433816 , n433817 , n433818 , 
 n433819 , n433820 , n433821 , n433822 , n433823 , n433824 , n433825 , n433826 , n433827 , n433828 , 
 n433829 , n433830 , n433831 , n433832 , n433833 , n433834 , n433835 , n433836 , n433837 , n433838 , 
 n433839 , n433840 , n433841 , n433842 , n433843 , n433844 , n433845 , n433846 , n433847 , n433848 , 
 n433849 , n433850 , n433851 , n433852 , n433853 , n433854 , n433855 , n433856 , n433857 , n433858 , 
 n433859 , n433860 , n433861 , n433862 , n433863 , n433864 , n433865 , n433866 , n433867 , n433868 , 
 n433869 , n433870 , n433871 , n433872 , n433873 , n433874 , n433875 , n433876 , n433877 , n433878 , 
 n433879 , n433880 , n433881 , n433882 , n433883 , n433884 , n433885 , n433886 , n433887 , n433888 , 
 n433889 , n433890 , n433891 , n433892 , n433893 , n433894 , n433895 , n433896 , n433897 , n433898 , 
 n433899 , n433900 , n433901 , n433902 , n433903 , n433904 , n433905 , n433906 , n433907 , n433908 , 
 n433909 , n433910 , n433911 , n433912 , n433913 , n433914 , n433915 , n433916 , n433917 , n433918 , 
 n433919 , n433920 , n433921 , n433922 , n433923 , n433924 , n433925 , n433926 , n433927 , n433928 , 
 n433929 , n433930 , n433931 , n433932 , n433933 , n433934 , n433935 , n433936 , n433937 , n433938 , 
 n433939 , n433940 , n433941 , n433942 , n433943 , n433944 , n433945 , n433946 , n433947 , n433948 , 
 n433949 , n433950 , n433951 , n433952 , n433953 , n433954 , n433955 , n433956 , n433957 , n433958 , 
 n433959 , n433960 , n433961 , n433962 , n433963 , n433964 , n433965 , n433966 , n433967 , n433968 , 
 n433969 , n433970 , n433971 , n433972 , n433973 , n433974 , n433975 , n433976 , n433977 , n433978 , 
 n433979 , n433980 , n433981 , n433982 , n433983 , n433984 , n433985 , n433986 , n433987 , n433988 , 
 n433989 , n433990 , n433991 , n433992 , n433993 , n433994 , n433995 , n433996 , n433997 , n433998 , 
 n433999 , n434000 , n434001 , n434002 , n434003 , n434004 , n434005 , n434006 , n434007 , n434008 , 
 n434009 , n434010 , n434011 , n434012 , n434013 , n434014 , n434015 , n434016 , n434017 , n434018 , 
 n434019 , n434020 , n434021 , n434022 , n434023 , n434024 , n434025 , n434026 , n434027 , n434028 , 
 n434029 , n434030 , n434031 , n434032 , n434033 , n434034 , n434035 , n434036 , n434037 , n434038 , 
 n434039 , n434040 , n434041 , n434042 , n434043 , n434044 , n434045 , n434046 , n434047 , n434048 , 
 n434049 , n434050 , n434051 , n434052 , n434053 , n434054 , n434055 , n434056 , n434057 , n434058 , 
 n434059 , n434060 , n434061 , n434062 , n434063 , n434064 , n434065 , n434066 , n434067 , n434068 , 
 n434069 , n434070 , n434071 , n434072 , n434073 , n434074 , n434075 , n434076 , n434077 , n434078 , 
 n434079 , n434080 , n434081 , n434082 , n434083 , n434084 , n434085 , n434086 , n434087 , n434088 , 
 n434089 , n434090 , n434091 , n434092 , n434093 , n434094 , n434095 , n434096 , n434097 , n434098 , 
 n434099 , n434100 , n434101 , n434102 , n434103 , n434104 , n434105 , n434106 , n434107 , n434108 , 
 n434109 , n434110 , n434111 , n434112 , n434113 , n434114 , n434115 , n434116 , n434117 , n434118 , 
 n434119 , n434120 , n434121 , n434122 , n434123 , n434124 , n434125 , n434126 , n434127 , n434128 , 
 n434129 , n434130 , n434131 , n434132 , n434133 , n434134 , n434135 , n434136 , n434137 , n434138 , 
 n434139 , n434140 , n434141 , n434142 , n434143 , n434144 , n434145 , n434146 , n434147 , n434148 , 
 n434149 , n434150 , n434151 , n434152 , n434153 , n434154 , n434155 , n434156 , n434157 , n434158 , 
 n434159 , n434160 , n434161 , n434162 , n434163 , n434164 , n434165 , n434166 , n434167 , n434168 , 
 n434169 , n434170 , n434171 , n434172 , n434173 , n434174 , n434175 , n434176 , n434177 , n434178 , 
 n434179 , n434180 , n434181 , n434182 , n434183 , n434184 , n434185 , n434186 , n434187 , n434188 , 
 n434189 , n434190 , n434191 , n434192 , n434193 , n434194 , n434195 , n434196 , n434197 , n434198 , 
 n434199 , n434200 , n434201 , n434202 , n434203 , n434204 , n434205 , n434206 , n434207 , n434208 , 
 n434209 , n434210 , n434211 , n434212 , n434213 , n434214 , n434215 , n434216 , n434217 , n434218 , 
 n434219 , n434220 , n434221 , n434222 , n434223 , n434224 , n434225 , n434226 , n434227 , n434228 , 
 n434229 , n434230 , n434231 , n434232 , n434233 , n434234 , n434235 , n434236 , n434237 , n434238 , 
 n434239 , n434240 , n434241 , n434242 , n434243 , n434244 , n434245 , n434246 , n434247 , n434248 , 
 n434249 , n434250 , n434251 , n434252 , n434253 , n434254 , n434255 , n434256 , n434257 , n434258 , 
 n434259 , n434260 , n434261 , n434262 , n434263 , n434264 , n434265 , n434266 , n434267 , n434268 , 
 n434269 , n434270 , n434271 , n434272 , n434273 , n434274 , n434275 , n434276 , n434277 , n434278 , 
 n434279 , n434280 , n434281 , n434282 , n434283 , n434284 , n434285 , n434286 , n434287 , n434288 , 
 n434289 , n434290 , n434291 , n434292 , n434293 , n434294 , n434295 , n434296 , n434297 , n434298 , 
 n434299 , n434300 , n434301 , n434302 , n434303 , n434304 , n434305 , n434306 , n434307 , n434308 , 
 n434309 , n434310 , n434311 , n434312 , n434313 , n434314 , n434315 , n434316 , n434317 , n434318 , 
 n434319 , n434320 , n434321 , n434322 , n434323 , n434324 , n434325 , n434326 , n434327 , n434328 , 
 n434329 , n434330 , n434331 , n434332 , n434333 , n434334 , n434335 , n434336 , n434337 , n434338 , 
 n434339 , n434340 , n434341 , n434342 , n434343 , n434344 , n434345 , n434346 , n434347 , n434348 , 
 n434349 , n434350 , n434351 , n434352 , n434353 , n434354 , n434355 , n434356 , n434357 , n434358 , 
 n434359 , n434360 , n434361 , n434362 , n434363 , n434364 , n434365 , n434366 , n434367 , n434368 , 
 n434369 , n434370 , n434371 , n434372 , n434373 , n434374 , n434375 , n434376 , n434377 , n434378 , 
 n434379 , n434380 , n434381 , n434382 , n434383 , n434384 , n434385 , n434386 , n434387 , n434388 , 
 n434389 , n434390 , n434391 , n434392 , n434393 , n434394 , n434395 , n434396 , n434397 , n434398 , 
 n434399 , n434400 , n434401 , n434402 , n434403 , n434404 , n434405 , n434406 , n434407 , n434408 , 
 n434409 , n434410 , n434411 , n434412 , n434413 , n434414 , n434415 , n434416 , n434417 , n434418 , 
 n434419 , n434420 , n434421 , n434422 , n434423 , n434424 , n434425 , n434426 , n434427 , n434428 , 
 n434429 , n434430 , n434431 , n434432 , n434433 , n434434 , n434435 , n434436 , n434437 , n434438 , 
 n434439 , n434440 , n434441 , n434442 , n434443 , n434444 , n434445 , n434446 , n434447 , n434448 , 
 n434449 , n434450 , n434451 , n434452 , n434453 , n434454 , n434455 , n434456 , n434457 , n434458 , 
 n434459 , n434460 , n434461 , n434462 , n434463 , n434464 , n434465 , n434466 , n434467 , n434468 , 
 n434469 , n434470 , n434471 , n434472 , n434473 , n434474 , n434475 , n434476 , n434477 , n434478 , 
 n434479 , n434480 , n434481 , n434482 , n434483 , n434484 , n434485 , n434486 , n434487 , n434488 , 
 n434489 , n434490 , n434491 , n434492 , n434493 , n434494 , n434495 , n434496 , n434497 , n434498 , 
 n434499 , n434500 , n434501 , n434502 , n434503 , n434504 , n434505 , n434506 , n434507 , n434508 , 
 n434509 , n434510 , n434511 , n434512 , n434513 , n434514 , n434515 , n434516 , n434517 , n434518 , 
 n434519 , n434520 , n434521 , n434522 , n434523 , n434524 , n434525 , n434526 , n434527 , n434528 , 
 n434529 , n434530 , n434531 , n434532 , n434533 , n434534 , n434535 , n434536 , n434537 , n434538 , 
 n434539 , n434540 , n434541 , n434542 , n434543 , n434544 , n434545 , n434546 , n434547 , n434548 , 
 n434549 , n434550 , n434551 , n434552 , n434553 , n434554 , n434555 , n434556 , n434557 , n434558 , 
 n434559 , n434560 , n434561 , n434562 , n434563 , n434564 , n434565 , n434566 , n434567 , n434568 , 
 n434569 , n434570 , n434571 , n434572 , n434573 , n434574 , n434575 , n434576 , n434577 , n434578 , 
 n434579 , n434580 , n434581 , n434582 , n434583 , n434584 , n434585 , n434586 , n434587 , n434588 , 
 n434589 , n434590 , n434591 , n434592 , n434593 , n434594 , n434595 , n434596 , n434597 , n434598 , 
 n434599 , n434600 , n434601 , n434602 , n434603 , n434604 , n434605 , n434606 , n434607 , n434608 , 
 n434609 , n434610 , n434611 , n434612 , n434613 , n434614 , n434615 , n434616 , n434617 , n434618 , 
 n434619 , n434620 , n434621 , n434622 , n434623 , n434624 , n434625 , n434626 , n434627 , n434628 , 
 n434629 , n434630 , n434631 , n434632 , n434633 , n434634 , n434635 , n434636 , n434637 , n434638 , 
 n434639 , n434640 , n434641 , n434642 , n434643 , n434644 , n434645 , n434646 , n434647 , n434648 , 
 n434649 , n434650 , n434651 , n434652 , n434653 , n434654 , n434655 , n434656 , n434657 , n434658 , 
 n434659 , n434660 , n434661 , n434662 , n434663 , n434664 , n434665 , n434666 , n434667 , n434668 , 
 n434669 , n434670 , n434671 , n434672 , n434673 , n434674 , n434675 , n434676 , n434677 , n434678 , 
 n434679 , n434680 , n434681 , n434682 , n434683 , n434684 , n434685 , n434686 , n434687 , n434688 , 
 n434689 , n434690 , n434691 , n434692 , n434693 , n434694 , n434695 , n434696 , n434697 , n434698 , 
 n434699 , n434700 , n434701 , n434702 , n434703 , n434704 , n434705 , n434706 , n434707 , n434708 , 
 n434709 , n434710 , n434711 , n434712 , n434713 , n434714 , n434715 , n434716 , n434717 , n434718 , 
 n434719 , n434720 , n434721 , n434722 , n434723 , n434724 , n434725 , n434726 , n434727 , n434728 , 
 n434729 , n434730 , n434731 , n434732 , n434733 , n434734 , n434735 , n434736 , n434737 , n434738 , 
 n434739 , n434740 , n434741 , n434742 , n434743 , n434744 , n434745 , n434746 , n434747 , n434748 , 
 n434749 , n434750 , n434751 , n434752 , n434753 , n434754 , n434755 , n434756 , n434757 , n434758 , 
 n434759 , n434760 , n434761 , n434762 , n434763 , n434764 , n434765 , n434766 , n434767 , n434768 , 
 n434769 , n434770 , n434771 , n434772 , n434773 , n434774 , n434775 , n434776 , n434777 , n434778 , 
 n434779 , n434780 , n434781 , n434782 , n434783 , n434784 , n434785 , n434786 , n434787 , n434788 , 
 n434789 , n434790 , n434791 , n434792 , n434793 , n434794 , n434795 , n434796 , n434797 , n434798 , 
 n434799 , n434800 , n434801 , n434802 , n434803 , n434804 , n434805 , n434806 , n434807 , n434808 , 
 n434809 , n434810 , n434811 , n434812 , n434813 , n434814 , n434815 , n434816 , n434817 , n434818 , 
 n434819 , n434820 , n434821 , n434822 , n434823 , n434824 , n434825 , n434826 , n434827 , n434828 , 
 n434829 , n434830 , n434831 , n434832 , n434833 , n434834 , n434835 , n434836 , n434837 , n434838 , 
 n434839 , n434840 , n434841 , n434842 , n434843 , n434844 , n434845 , n434846 , n434847 , n434848 , 
 n434849 , n434850 , n434851 , n434852 , n434853 , n434854 , n434855 , n434856 , n434857 , n434858 , 
 n434859 , n434860 , n434861 , n434862 , n434863 , n434864 , n434865 , n434866 , n434867 , n434868 , 
 n434869 , n434870 , n434871 , n434872 , n434873 , n434874 , n434875 , n434876 , n434877 , n434878 , 
 n434879 , n434880 , n434881 , n434882 , n434883 , n434884 , n434885 , n434886 , n434887 , n434888 , 
 n434889 , n434890 , n434891 , n434892 , n434893 , n434894 , n434895 , n434896 , n434897 , n434898 , 
 n434899 , n434900 , n434901 , n434902 , n434903 , n434904 , n434905 , n434906 , n434907 , n434908 , 
 n434909 , n434910 , n434911 , n434912 , n434913 , n434914 , n434915 , n434916 , n434917 , n434918 , 
 n434919 , n434920 , n434921 , n434922 , n434923 , n434924 , n434925 , n434926 , n434927 , n434928 , 
 n434929 , n434930 , n434931 , n434932 , n434933 , n434934 , n434935 , n434936 , n434937 , n434938 , 
 n434939 , n434940 , n434941 , n434942 , n434943 , n434944 , n434945 , n434946 , n434947 , n434948 , 
 n434949 , n434950 , n434951 , n434952 , n434953 , n434954 , n434955 , n434956 , n434957 , n434958 , 
 n434959 , n434960 , n434961 , n434962 , n434963 , n434964 , n434965 , n434966 , n434967 , n434968 , 
 n434969 , n434970 , n434971 , n434972 , n434973 , n434974 , n434975 , n434976 , n434977 , n434978 , 
 n434979 , n434980 , n434981 , n434982 , n434983 , n434984 , n434985 , n434986 , n434987 , n434988 , 
 n434989 , n434990 , n434991 , n434992 , n434993 , n434994 , n434995 , n434996 , n434997 , n434998 , 
 n434999 , n435000 , n435001 , n435002 , n435003 , n435004 , n435005 , n435006 , n435007 , n435008 , 
 n435009 , n435010 , n435011 , n435012 , n435013 , n435014 , n435015 , n435016 , n435017 , n435018 , 
 n435019 , n435020 , n435021 , n435022 , n435023 , n435024 , n435025 , n435026 , n435027 , n435028 , 
 n435029 , n435030 , n435031 , n435032 , n435033 , n435034 , n435035 , n435036 , n435037 , n435038 , 
 n435039 , n435040 , n435041 , n435042 , n435043 , n435044 , n435045 , n435046 , n435047 , n435048 , 
 n435049 , n435050 , n435051 , n435052 , n435053 , n435054 , n435055 , n435056 , n435057 , n435058 , 
 n435059 , n435060 , n435061 , n435062 , n435063 , n435064 , n435065 , n435066 , n435067 , n435068 , 
 n435069 , n435070 , n435071 , n435072 , n435073 , n435074 , n435075 , n435076 , n435077 , n435078 , 
 n435079 , n435080 , n435081 , n435082 , n435083 , n435084 , n435085 , n435086 , n435087 , n435088 , 
 n435089 , n435090 , n435091 , n435092 , n435093 , n435094 , n435095 , n435096 , n435097 , n435098 , 
 n435099 , n435100 , n435101 , n435102 , n435103 , n435104 , n435105 , n435106 , n435107 , n435108 , 
 n435109 , n435110 , n435111 , n435112 , n435113 , n435114 , n435115 , n435116 , n435117 , n435118 , 
 n435119 , n435120 , n435121 , n435122 , n435123 , n435124 , n435125 , n435126 , n435127 , n435128 , 
 n435129 , n435130 , n435131 , n435132 , n435133 , n435134 , n435135 , n435136 , n435137 , n435138 , 
 n435139 , n435140 , n435141 , n435142 , n435143 , n435144 , n435145 , n435146 , n435147 , n435148 , 
 n435149 , n435150 , n435151 , n435152 , n435153 , n435154 , n435155 , n435156 , n435157 , n435158 , 
 n435159 , n435160 , n435161 , n435162 , n435163 , n435164 , n435165 , n435166 , n435167 , n435168 , 
 n435169 , n435170 , n435171 , n435172 , n435173 , n435174 , n435175 , n435176 , n435177 , n435178 , 
 n435179 , n435180 , n435181 , n435182 , n435183 , n435184 , n435185 , n435186 , n435187 , n435188 , 
 n435189 , n435190 , n435191 , n435192 , n435193 , n435194 , n435195 , n435196 , n435197 , n435198 , 
 n435199 , n435200 , n435201 , n435202 , n435203 , n435204 , n435205 , n435206 , n435207 , n435208 , 
 n435209 , n435210 , n435211 , n435212 , n435213 , n435214 , n435215 , n435216 , n435217 , n435218 , 
 n435219 , n435220 , n435221 , n435222 , n435223 , n435224 , n435225 , n435226 , n435227 , n435228 , 
 n435229 , n435230 , n435231 , n435232 , n435233 , n435234 , n435235 , n435236 , n435237 , n435238 , 
 n435239 , n435240 , n435241 , n435242 , n435243 , n435244 , n435245 , n435246 , n435247 , n435248 , 
 n435249 , n435250 , n435251 , n435252 , n435253 , n435254 , n435255 , n435256 , n435257 , n435258 , 
 n435259 , n435260 , n435261 , n435262 , n435263 , n435264 , n435265 , n435266 , n435267 , n435268 , 
 n435269 , n435270 , n435271 , n435272 , n435273 , n435274 , n435275 , n435276 , n435277 , n435278 , 
 n435279 , n435280 , n435281 , n435282 , n435283 , n435284 , n435285 , n435286 , n435287 , n435288 , 
 n435289 , n435290 , n435291 , n435292 , n435293 , n435294 , n435295 , n435296 , n435297 , n435298 , 
 n435299 , n435300 , n435301 , n435302 , n435303 , n435304 , n435305 , n435306 , n435307 , n435308 , 
 n435309 , n435310 , n435311 , n435312 , n435313 , n435314 , n435315 , n435316 , n435317 , n435318 , 
 n435319 , n435320 , n435321 , n435322 , n435323 , n435324 , n435325 , n435326 , n435327 , n435328 , 
 n435329 , n435330 , n435331 , n435332 , n435333 , n435334 , n435335 , n435336 , n435337 , n435338 , 
 n435339 , n435340 , n435341 , n435342 , n435343 , n435344 , n435345 , n435346 , n435347 , n435348 , 
 n435349 , n435350 , n435351 , n435352 , n435353 , n435354 , n435355 , n435356 , n435357 , n435358 , 
 n435359 , n435360 , n435361 , n435362 , n435363 , n435364 , n435365 , n435366 , n435367 , n435368 , 
 n435369 , n435370 , n435371 , n435372 , n435373 , n435374 , n435375 , n435376 , n435377 , n435378 , 
 n435379 , n435380 , n435381 , n435382 , n435383 , n435384 , n435385 , n435386 , n435387 , n435388 , 
 n435389 , n435390 , n435391 , n435392 , n435393 , n435394 , n435395 , n435396 , n435397 , n435398 , 
 n435399 , n435400 , n435401 , n435402 , n435403 , n435404 , n435405 , n435406 , n435407 , n435408 , 
 n435409 , n435410 , n435411 , n435412 , n435413 , n435414 , n435415 , n435416 , n435417 , n435418 , 
 n435419 , n435420 , n435421 , n435422 , n435423 , n435424 , n435425 , n435426 , n435427 , n435428 , 
 n435429 , n435430 , n435431 , n435432 , n435433 , n435434 , n435435 , n435436 , n435437 , n435438 , 
 n435439 , n435440 , n435441 , n435442 , n435443 , n435444 , n435445 , n435446 , n435447 , n435448 , 
 n435449 , n435450 , n435451 , n435452 , n435453 , n435454 , n435455 , n435456 , n435457 , n435458 , 
 n435459 , n435460 , n435461 , n435462 , n435463 , n435464 , n435465 , n435466 , n435467 , n435468 , 
 n435469 , n435470 , n435471 , n435472 , n435473 , n435474 , n435475 , n435476 , n435477 , n435478 , 
 n435479 , n435480 , n435481 , n435482 , n435483 , n435484 , n435485 , n435486 , n435487 , n435488 , 
 n435489 , n435490 , n435491 , n435492 , n435493 , n435494 , n435495 , n435496 , n435497 , n435498 , 
 n435499 , n435500 , n435501 , n435502 , n435503 , n435504 , n435505 , n435506 , n435507 , n435508 , 
 n435509 , n435510 , n435511 , n435512 , n435513 , n435514 , n435515 , n435516 , n435517 , n435518 , 
 n435519 , n435520 , n435521 , n435522 , n435523 , n435524 , n435525 , n435526 , n435527 , n435528 , 
 n435529 , n435530 , n435531 , n435532 , n435533 , n435534 , n435535 , n435536 , n435537 , n435538 , 
 n435539 , n435540 , n435541 , n435542 , n435543 , n435544 , n435545 , n435546 , n435547 , n435548 , 
 n435549 , n435550 , n435551 , n435552 , n435553 , n435554 , n435555 , n435556 , n435557 , n435558 , 
 n435559 , n435560 , n435561 , n435562 , n435563 , n435564 , n435565 , n435566 , n435567 , n435568 , 
 n435569 , n435570 , n435571 , n435572 , n435573 , n435574 , n435575 , n435576 , n435577 , n435578 , 
 n435579 , n435580 , n435581 , n435582 , n435583 , n435584 , n435585 , n435586 , n435587 , n435588 , 
 n435589 , n435590 , n435591 , n435592 , n435593 , n435594 , n435595 , n435596 , n435597 , n435598 , 
 n435599 , n435600 , n435601 , n435602 , n435603 , n435604 , n435605 , n435606 , n435607 , n435608 , 
 n435609 , n435610 , n435611 , n435612 , n435613 , n435614 , n435615 , n435616 , n435617 , n435618 , 
 n435619 , n435620 , n435621 , n435622 , n435623 , n435624 , n435625 , n435626 , n435627 , n435628 , 
 n435629 , n435630 , n435631 , n435632 , n435633 , n435634 , n435635 , n435636 , n435637 , n435638 , 
 n435639 , n435640 , n435641 , n435642 , n435643 , n435644 , n435645 , n435646 , n435647 , n435648 , 
 n435649 , n435650 , n435651 , n435652 , n435653 , n435654 , n435655 , n435656 , n435657 , n435658 , 
 n435659 , n435660 , n435661 , n435662 , n435663 , n435664 , n435665 , n435666 , n435667 , n435668 , 
 n435669 , n435670 , n435671 , n435672 , n435673 , n435674 , n435675 , n435676 , n435677 , n435678 , 
 n435679 , n435680 , n435681 , n435682 , n435683 , n435684 , n435685 , n435686 , n435687 , n435688 , 
 n435689 , n435690 , n435691 , n435692 , n435693 , n435694 , n435695 , n435696 , n435697 , n435698 , 
 n435699 , n435700 , n435701 , n435702 , n435703 , n435704 , n435705 , n435706 , n435707 , n435708 , 
 n435709 , n435710 , n435711 , n435712 , n435713 , n435714 , n435715 , n435716 , n435717 , n435718 , 
 n435719 , n435720 , n435721 , n435722 , n435723 , n435724 , n435725 , n435726 , n435727 , n435728 , 
 n435729 , n435730 , n435731 , n435732 , n435733 , n435734 , n435735 , n435736 , n435737 , n435738 , 
 n435739 , n435740 , n435741 , n435742 , n435743 , n435744 , n435745 , n435746 , n435747 , n435748 , 
 n435749 , n435750 , n435751 , n435752 , n435753 , n435754 , n435755 , n435756 , n435757 , n435758 , 
 n435759 , n435760 , n435761 , n435762 , n435763 , n435764 , n435765 , n435766 , n435767 , n435768 , 
 n435769 , n435770 , n435771 , n435772 , n435773 , n435774 , n435775 , n435776 , n435777 , n435778 , 
 n435779 , n435780 , n435781 , n435782 , n435783 , n435784 , n435785 , n435786 , n435787 , n435788 , 
 n435789 , n435790 , n435791 , n435792 , n435793 , n435794 , n435795 , n435796 , n435797 , n435798 , 
 n435799 , n435800 , n435801 , n435802 , n435803 , n435804 , n435805 , n435806 , n435807 , n435808 , 
 n435809 , n435810 , n435811 , n435812 , n435813 , n435814 , n435815 , n435816 , n435817 , n435818 , 
 n435819 , n435820 , n435821 , n435822 , n435823 , n435824 , n435825 , n435826 , n435827 , n435828 , 
 n435829 , n435830 , n435831 , n435832 , n435833 , n435834 , n435835 , n435836 , n435837 , n435838 , 
 n435839 , n435840 , n435841 , n435842 , n435843 , n435844 , n435845 , n435846 , n435847 , n435848 , 
 n435849 , n435850 , n435851 , n435852 , n435853 , n435854 , n435855 , n435856 , n435857 , n435858 , 
 n435859 , n435860 , n435861 , n435862 , n435863 , n435864 , n435865 , n435866 , n435867 , n435868 , 
 n435869 , n435870 , n435871 , n435872 , n435873 , n435874 , n435875 , n435876 , n435877 , n435878 , 
 n435879 , n435880 , n435881 , n435882 , n435883 , n435884 , n435885 , n435886 , n435887 , n435888 , 
 n435889 , n435890 , n435891 , n435892 , n435893 , n435894 , n435895 , n435896 , n435897 , n435898 , 
 n435899 , n435900 , n435901 , n435902 , n435903 , n435904 , n435905 , n435906 , n435907 , n435908 , 
 n435909 , n435910 , n435911 , n435912 , n435913 , n435914 , n435915 , n435916 , n435917 , n435918 , 
 n435919 , n435920 , n435921 , n435922 , n435923 , n435924 , n435925 , n435926 , n435927 , n435928 , 
 n435929 , n435930 , n435931 , n435932 , n435933 , n435934 , n435935 , n435936 , n435937 , n435938 , 
 n435939 , n435940 , n435941 , n435942 , n435943 , n435944 , n435945 , n435946 , n435947 , n435948 , 
 n435949 , n435950 , n435951 , n435952 , n435953 , n435954 , n435955 , n435956 , n435957 , n435958 , 
 n435959 , n435960 , n435961 , n435962 , n435963 , n435964 , n435965 , n435966 , n435967 , n435968 , 
 n435969 , n435970 , n435971 , n435972 , n435973 , n435974 , n435975 , n435976 , n435977 , n435978 , 
 n435979 , n435980 , n435981 , n435982 , n435983 , n435984 , n435985 , n435986 , n435987 , n435988 , 
 n435989 , n435990 , n435991 , n435992 , n435993 , n435994 , n435995 , n435996 , n435997 , n435998 , 
 n435999 , n436000 , n436001 , n436002 , n436003 , n436004 , n436005 , n436006 , n436007 , n436008 , 
 n436009 , n436010 , n436011 , n436012 , n436013 , n436014 , n436015 , n436016 , n436017 , n436018 , 
 n436019 , n436020 , n436021 , n436022 , n436023 , n436024 , n436025 , n436026 , n436027 , n436028 , 
 n436029 , n436030 , n436031 , n436032 , n436033 , n436034 , n436035 , n436036 , n436037 , n436038 , 
 n436039 , n436040 , n436041 , n436042 , n436043 , n436044 , n436045 , n436046 , n436047 , n436048 , 
 n436049 , n436050 , n436051 , n436052 , n436053 , n436054 , n436055 , n436056 , n436057 , n436058 , 
 n436059 , n436060 , n436061 , n436062 , n436063 , n436064 , n436065 , n436066 , n436067 , n436068 , 
 n436069 , n436070 , n436071 , n436072 , n436073 , n436074 , n436075 , n436076 , n436077 , n436078 , 
 n436079 , n436080 , n436081 , n436082 , n436083 , n436084 , n436085 , n436086 , n436087 , n436088 , 
 n436089 , n436090 , n436091 , n436092 , n436093 , n436094 , n436095 , n436096 , n436097 , n436098 , 
 n436099 , n436100 , n436101 , n436102 , n436103 , n436104 , n436105 , n436106 , n436107 , n436108 , 
 n436109 , n436110 , n436111 , n436112 , n436113 , n436114 , n436115 , n436116 , n436117 , n436118 , 
 n436119 , n436120 , n436121 , n436122 , n436123 , n436124 , n436125 , n436126 , n436127 , n436128 , 
 n436129 , n436130 , n436131 , n436132 , n436133 , n436134 , n436135 , n436136 , n436137 , n436138 , 
 n436139 , n436140 , n436141 , n436142 , n436143 , n436144 , n436145 , n436146 , n436147 , n436148 , 
 n436149 , n436150 , n436151 , n436152 , n436153 , n436154 , n436155 , n436156 , n436157 , n436158 , 
 n436159 , n436160 , n436161 , n436162 , n436163 , n436164 , n436165 , n436166 , n436167 , n436168 , 
 n436169 , n436170 , n436171 , n436172 , n436173 , n436174 , n436175 , n436176 , n436177 , n436178 , 
 n436179 , n436180 , n436181 , n436182 , n436183 , n436184 , n436185 , n436186 , n436187 , n436188 , 
 n436189 , n436190 , n436191 , n436192 , n436193 , n436194 , n436195 , n436196 , n436197 , n436198 , 
 n436199 , n436200 , n436201 , n436202 , n436203 , n436204 , n436205 , n436206 , n436207 , n436208 , 
 n436209 , n436210 , n436211 , n436212 , n436213 , n436214 , n436215 , n436216 , n436217 , n436218 , 
 n436219 , n436220 , n436221 , n436222 , n436223 , n436224 , n436225 , n436226 , n436227 , n436228 , 
 n436229 , n436230 , n436231 , n436232 , n436233 , n436234 , n436235 , n436236 , n436237 , n436238 , 
 n436239 , n436240 , n436241 , n436242 , n436243 , n436244 , n436245 , n436246 , n436247 , n436248 , 
 n436249 , n436250 , n436251 , n436252 , n436253 , n436254 , n436255 , n436256 , n436257 , n436258 , 
 n436259 , n436260 , n436261 , n436262 , n436263 , n436264 , n436265 , n436266 , n436267 , n436268 , 
 n436269 , n436270 , n436271 , n436272 , n436273 , n436274 , n436275 , n436276 , n436277 , n436278 , 
 n436279 , n436280 , n436281 , n436282 , n436283 , n436284 , n436285 , n436286 , n436287 , n436288 , 
 n436289 , n436290 , n436291 , n436292 , n436293 , n436294 , n436295 , n436296 , n436297 , n436298 , 
 n436299 , n436300 , n436301 , n436302 , n436303 , n436304 , n436305 , n436306 , n436307 , n436308 , 
 n436309 , n436310 , n436311 , n436312 , n436313 , n436314 , n436315 , n436316 , n436317 , n436318 , 
 n436319 , n436320 , n436321 , n436322 , n436323 , n436324 , n436325 , n436326 , n436327 , n436328 , 
 n436329 , n436330 , n436331 , n436332 , n436333 , n436334 , n436335 , n436336 , n436337 , n436338 , 
 n436339 , n436340 , n436341 , n436342 , n436343 , n436344 , n436345 , n436346 , n436347 , n436348 , 
 n436349 , n436350 , n436351 , n436352 , n436353 , n436354 , n436355 , n436356 , n436357 , n436358 , 
 n436359 , n436360 , n436361 , n436362 , n436363 , n436364 , n436365 , n436366 , n436367 , n436368 , 
 n436369 , n436370 , n436371 , n436372 , n436373 , n436374 , n436375 , n436376 , n436377 , n436378 , 
 n436379 , n436380 , n436381 , n436382 , n436383 , n436384 , n436385 , n436386 , n436387 , n436388 , 
 n436389 , n436390 , n436391 , n436392 , n436393 , n436394 , n436395 , n436396 , n436397 , n436398 , 
 n436399 , n436400 , n436401 , n436402 , n436403 , n436404 , n436405 , n436406 , n436407 , n436408 , 
 n436409 , n436410 , n436411 , n436412 , n436413 , n436414 , n436415 , n436416 , n436417 , n436418 , 
 n436419 , n436420 , n436421 , n436422 , n436423 , n436424 , n436425 , n436426 , n436427 , n436428 , 
 n436429 , n436430 , n436431 , n436432 , n436433 , n436434 , n436435 , n436436 , n436437 , n436438 , 
 n436439 , n436440 , n436441 , n436442 , n436443 , n436444 , n436445 , n436446 , n436447 , n436448 , 
 n436449 , n436450 , n436451 , n436452 , n436453 , n436454 , n436455 , n436456 , n436457 , n436458 , 
 n436459 , n436460 , n436461 , n436462 , n436463 , n436464 , n436465 , n436466 , n436467 , n436468 , 
 n436469 , n436470 , n436471 , n436472 , n436473 , n436474 , n436475 , n436476 , n436477 , n436478 , 
 n436479 , n436480 , n436481 , n436482 , n436483 , n436484 , n436485 , n436486 , n436487 , n436488 , 
 n436489 , n436490 , n436491 , n436492 , n436493 , n436494 , n436495 , n436496 , n436497 , n436498 , 
 n436499 , n436500 , n436501 , n436502 , n436503 , n436504 , n436505 , n436506 , n436507 , n436508 , 
 n436509 , n436510 , n436511 , n436512 , n436513 , n436514 , n436515 , n436516 , n436517 , n436518 , 
 n436519 , n436520 , n436521 , n436522 , n436523 , n436524 , n436525 , n436526 , n436527 , n436528 , 
 n436529 , n436530 , n436531 , n436532 , n436533 , n436534 , n436535 , n436536 , n436537 , n436538 , 
 n436539 , n436540 , n436541 , n436542 , n436543 , n436544 , n436545 , n436546 , n436547 , n436548 , 
 n436549 , n436550 , n436551 , n436552 , n436553 , n436554 , n436555 , n436556 , n436557 , n436558 , 
 n436559 , n436560 , n436561 , n436562 , n436563 , n436564 , n436565 , n436566 , n436567 , n436568 , 
 n436569 , n436570 , n436571 , n436572 , n436573 , n436574 , n436575 , n436576 , n436577 , n436578 , 
 n436579 , n436580 , n436581 , n436582 , n436583 , n436584 , n436585 , n436586 , n436587 , n436588 , 
 n436589 , n436590 , n436591 , n436592 , n436593 , n436594 , n436595 , n436596 , n436597 , n436598 , 
 n436599 , n436600 , n436601 , n436602 , n436603 , n436604 , n436605 , n436606 , n436607 , n436608 , 
 n436609 , n436610 , n436611 , n436612 , n436613 , n436614 , n436615 , n436616 , n436617 , n436618 , 
 n436619 , n436620 , n436621 , n436622 , n436623 , n436624 , n436625 , n436626 , n436627 , n436628 , 
 n436629 , n436630 , n436631 , n436632 , n436633 , n436634 , n436635 , n436636 , n436637 , n436638 , 
 n436639 , n436640 , n436641 , n436642 , n436643 , n436644 , n436645 , n436646 , n436647 , n436648 , 
 n436649 , n436650 , n436651 , n436652 , n436653 , n436654 , n436655 , n436656 , n436657 , n436658 , 
 n436659 , n436660 , n436661 , n436662 , n436663 , n436664 , n436665 , n436666 , n436667 , n436668 , 
 n436669 , n436670 , n436671 , n436672 , n436673 , n436674 , n436675 , n436676 , n436677 , n436678 , 
 n436679 , n436680 , n436681 , n436682 , n436683 , n436684 , n436685 , n436686 , n436687 , n436688 , 
 n436689 , n436690 , n436691 , n436692 , n436693 , n436694 , n436695 , n436696 , n436697 , n436698 , 
 n436699 , n436700 , n436701 , n436702 , n436703 , n436704 , n436705 , n436706 , n436707 , n436708 , 
 n436709 , n436710 , n436711 , n436712 , n436713 , n436714 , n436715 , n436716 , n436717 , n436718 , 
 n436719 , n436720 , n436721 , n436722 , n436723 , n436724 , n436725 , n436726 , n436727 , n436728 , 
 n436729 , n436730 , n436731 , n436732 , n436733 , n436734 , n436735 , n436736 , n436737 , n436738 , 
 n436739 , n436740 , n436741 , n436742 , n436743 , n436744 , n436745 , n436746 , n436747 , n436748 , 
 n436749 , n436750 , n436751 , n436752 , n436753 , n436754 , n436755 , n436756 , n436757 , n436758 , 
 n436759 , n436760 , n436761 , n436762 , n436763 , n436764 , n436765 , n436766 , n436767 , n436768 , 
 n436769 , n436770 , n436771 , n436772 , n436773 , n436774 , n436775 , n436776 , n436777 , n436778 , 
 n436779 , n436780 , n436781 , n436782 , n436783 , n436784 , n436785 , n436786 , n436787 , n436788 , 
 n436789 , n436790 , n436791 , n436792 , n436793 , n436794 , n436795 , n436796 , n436797 , n436798 , 
 n436799 , n436800 , n436801 , n436802 , n436803 , n436804 , n436805 , n436806 , n436807 , n436808 , 
 n436809 , n436810 , n436811 , n436812 , n436813 , n436814 , n436815 , n436816 , n436817 , n436818 , 
 n436819 , n436820 , n436821 , n436822 , n436823 , n436824 , n436825 , n436826 , n436827 , n436828 , 
 n436829 , n436830 , n436831 , n436832 , n436833 , n436834 , n436835 , n436836 , n436837 , n436838 , 
 n436839 , n436840 , n436841 , n436842 , n436843 , n436844 , n436845 , n436846 , n436847 , n436848 , 
 n436849 , n436850 , n436851 , n436852 , n436853 , n436854 , n436855 , n436856 , n436857 , n436858 , 
 n436859 , n436860 , n436861 , n436862 , n436863 , n436864 , n436865 , n436866 , n436867 , n436868 , 
 n436869 , n436870 , n436871 , n436872 , n436873 , n436874 , n436875 , n436876 , n436877 , n436878 , 
 n436879 , n436880 , n436881 , n436882 , n436883 , n436884 , n436885 , n436886 , n436887 , n436888 , 
 n436889 , n436890 , n436891 , n436892 , n436893 , n436894 , n436895 , n436896 , n436897 , n436898 , 
 n436899 , n436900 , n436901 , n436902 , n436903 , n436904 , n436905 , n436906 , n436907 , n436908 , 
 n436909 , n436910 , n436911 , n436912 , n436913 , n436914 , n436915 , n436916 , n436917 , n436918 , 
 n436919 , n436920 , n436921 , n436922 , n436923 , n436924 , n436925 , n436926 , n436927 , n436928 , 
 n436929 , n436930 , n436931 , n436932 , n436933 , n436934 , n436935 , n436936 , n436937 , n436938 , 
 n436939 , n436940 , n436941 , n436942 , n436943 , n436944 , n436945 , n436946 , n436947 , n436948 , 
 n436949 , n436950 , n436951 , n436952 , n436953 , n436954 , n436955 , n436956 , n436957 , n436958 , 
 n436959 , n436960 , n436961 , n436962 , n436963 , n436964 , n436965 , n436966 , n436967 , n436968 , 
 n436969 , n436970 , n436971 , n436972 , n436973 , n436974 , n436975 , n436976 , n436977 , n436978 , 
 n436979 , n436980 , n436981 , n436982 , n436983 , n436984 , n436985 , n436986 , n436987 , n436988 , 
 n436989 , n436990 , n436991 , n436992 , n436993 , n436994 , n436995 , n436996 , n436997 , n436998 , 
 n436999 , n437000 , n437001 , n437002 , n437003 , n437004 , n437005 , n437006 , n437007 , n437008 , 
 n437009 , n437010 , n437011 , n437012 , n437013 , n437014 , n437015 , n437016 , n437017 , n437018 , 
 n437019 , n437020 , n437021 , n437022 , n437023 , n437024 , n437025 , n437026 , n437027 , n437028 , 
 n437029 , n437030 , n437031 , n437032 , n437033 , n437034 , n437035 , n437036 , n437037 , n437038 , 
 n437039 , n437040 , n437041 , n437042 , n437043 , n437044 , n437045 , n437046 , n437047 , n437048 , 
 n437049 , n437050 , n437051 , n437052 , n437053 , n437054 , n437055 , n437056 , n437057 , n437058 , 
 n437059 , n437060 , n437061 , n437062 , n437063 , n437064 , n437065 , n437066 , n437067 , n437068 , 
 n437069 , n437070 , n437071 , n437072 , n437073 , n437074 , n437075 , n437076 , n437077 , n437078 , 
 n437079 , n437080 , n437081 , n437082 , n437083 , n437084 , n437085 , n437086 , n437087 , n437088 , 
 n437089 , n437090 , n437091 , n437092 , n437093 , n437094 , n437095 , n437096 , n437097 , n437098 , 
 n437099 , n437100 , n437101 , n437102 , n437103 , n437104 , n437105 , n437106 , n437107 , n437108 , 
 n437109 , n437110 , n437111 , n437112 , n437113 , n437114 , n437115 , n437116 , n437117 , n437118 , 
 n437119 , n437120 , n437121 , n437122 , n437123 , n437124 , n437125 , n437126 , n437127 , n437128 , 
 n437129 , n437130 , n437131 , n437132 , n437133 , n437134 , n437135 , n437136 , n437137 , n437138 , 
 n437139 , n437140 , n437141 , n437142 , n437143 , n437144 , n437145 , n437146 , n437147 , n437148 , 
 n437149 , n437150 , n437151 , n437152 , n437153 , n437154 , n437155 , n437156 , n437157 , n437158 , 
 n437159 , n437160 , n437161 , n437162 , n437163 , n437164 , n437165 , n437166 , n437167 , n437168 , 
 n437169 , n437170 , n437171 , n437172 , n437173 , n437174 , n437175 , n437176 , n437177 , n437178 , 
 n437179 , n437180 , n437181 , n437182 , n437183 , n437184 , n437185 , n437186 , n437187 , n437188 , 
 n437189 , n437190 , n437191 , n437192 , n437193 , n437194 , n437195 , n437196 , n437197 , n437198 , 
 n437199 , n437200 , n437201 , n437202 , n437203 , n437204 , n437205 , n437206 , n437207 , n437208 , 
 n437209 , n437210 , n437211 , n437212 , n437213 , n437214 , n437215 , n437216 , n437217 , n437218 , 
 n437219 , n437220 , n437221 , n437222 , n437223 , n437224 , n437225 , n437226 , n437227 , n437228 , 
 n437229 , n437230 , n437231 , n437232 , n437233 , n437234 , n437235 , n437236 , n437237 , n437238 , 
 n437239 , n437240 , n437241 , n437242 , n437243 , n437244 , n437245 , n437246 , n437247 , n437248 , 
 n437249 , n437250 , n437251 , n437252 , n437253 , n437254 , n437255 , n437256 , n437257 , n437258 , 
 n437259 , n437260 , n437261 , n437262 , n437263 , n437264 , n437265 , n437266 , n437267 , n437268 , 
 n437269 , n437270 , n437271 , n437272 , n437273 , n437274 , n437275 , n437276 , n437277 , n437278 , 
 n437279 , n437280 , n437281 , n437282 , n437283 , n437284 , n437285 , n437286 , n437287 , n437288 , 
 n437289 , n437290 , n437291 , n437292 , n437293 , n437294 , n437295 , n437296 , n437297 , n437298 , 
 n437299 , n437300 , n437301 , n437302 , n437303 , n437304 , n437305 , n437306 , n437307 , n437308 , 
 n437309 , n437310 , n437311 , n437312 , n437313 , n437314 , n437315 , n437316 , n437317 , n437318 , 
 n437319 , n437320 , n437321 , n437322 , n437323 , n437324 , n437325 , n437326 , n437327 , n437328 , 
 n437329 , n437330 , n437331 , n437332 , n437333 , n437334 , n437335 , n437336 , n437337 , n437338 , 
 n437339 , n437340 , n437341 , n437342 , n437343 , n437344 , n437345 , n437346 , n437347 , n437348 , 
 n437349 , n437350 , n437351 , n437352 , n437353 , n437354 , n437355 , n437356 , n437357 , n437358 , 
 n437359 , n437360 , n437361 , n437362 , n437363 , n437364 , n437365 , n437366 , n437367 , n437368 , 
 n437369 , n437370 , n437371 , n437372 , n437373 , n437374 , n437375 , n437376 , n437377 , n437378 , 
 n437379 , n437380 , n437381 , n437382 , n437383 , n437384 , n437385 , n437386 , n437387 , n437388 , 
 n437389 , n437390 , n437391 , n437392 , n437393 , n437394 , n437395 , n437396 , n437397 , n437398 , 
 n437399 , n437400 , n437401 , n437402 , n437403 , n437404 , n437405 , n437406 , n437407 , n437408 , 
 n437409 , n437410 , n437411 , n437412 , n437413 , n437414 , n437415 , n437416 , n437417 , n437418 , 
 n437419 , n437420 , n437421 , n437422 , n437423 , n437424 , n437425 , n437426 , n437427 , n437428 , 
 n437429 , n437430 , n437431 , n437432 , n437433 , n437434 , n437435 , n437436 , n437437 , n437438 , 
 n437439 , n437440 , n437441 , n437442 , n437443 , n437444 , n437445 , n437446 , n437447 , n437448 , 
 n437449 , n437450 , n437451 , n437452 , n437453 , n437454 , n437455 , n437456 , n437457 , n437458 , 
 n437459 , n437460 , n437461 , n437462 , n437463 , n437464 , n437465 , n437466 , n437467 , n437468 , 
 n437469 , n437470 , n437471 , n437472 , n437473 , n437474 , n437475 , n437476 , n437477 , n437478 , 
 n437479 , n437480 , n437481 , n437482 , n437483 , n437484 , n437485 , n437486 , n437487 , n437488 , 
 n437489 , n437490 , n437491 , n437492 , n437493 , n437494 , n437495 , n437496 , n437497 , n437498 , 
 n437499 , n437500 , n437501 , n437502 , n437503 , n437504 , n437505 , n437506 , n437507 , n437508 , 
 n437509 , n437510 , n437511 , n437512 , n437513 , n437514 , n437515 , n437516 , n437517 , n437518 , 
 n437519 , n437520 , n437521 , n437522 , n437523 , n437524 , n437525 , n437526 , n437527 , n437528 , 
 n437529 , n437530 , n437531 , n437532 , n437533 , n437534 , n437535 , n437536 , n437537 , n437538 , 
 n437539 , n437540 , n437541 , n437542 , n437543 , n437544 , n437545 , n437546 , n437547 , n437548 , 
 n437549 , n437550 , n437551 , n437552 , n437553 , n437554 , n437555 , n437556 , n437557 , n437558 , 
 n437559 , n437560 , n437561 , n437562 , n437563 , n437564 , n437565 , n437566 , n437567 , n437568 , 
 n437569 , n437570 , n437571 , n437572 , n437573 , n437574 , n437575 , n437576 , n437577 , n437578 , 
 n437579 , n437580 , n437581 , n437582 , n437583 , n437584 , n437585 , n437586 , n437587 , n437588 , 
 n437589 , n437590 , n437591 , n437592 , n437593 , n437594 , n437595 , n437596 , n437597 , n437598 , 
 n437599 , n437600 , n437601 , n437602 , n437603 , n437604 , n437605 , n437606 , n437607 , n437608 , 
 n437609 , n437610 , n437611 , n437612 , n437613 , n437614 , n437615 , n437616 , n437617 , n437618 , 
 n437619 , n437620 , n437621 , n437622 , n437623 , n437624 , n437625 , n437626 , n437627 , n437628 , 
 n437629 , n437630 , n437631 , n437632 , n437633 , n437634 , n437635 , n437636 , n437637 , n437638 , 
 n437639 , n437640 , n437641 , n437642 , n437643 , n437644 , n437645 , n437646 , n437647 , n437648 , 
 n437649 , n437650 , n437651 , n437652 , n437653 , n437654 , n437655 , n437656 , n437657 , n437658 , 
 n437659 , n437660 , n437661 , n437662 , n437663 , n437664 , n437665 , n437666 , n437667 , n437668 , 
 n437669 , n437670 , n437671 , n437672 , n437673 , n437674 , n437675 , n437676 , n437677 , n437678 , 
 n437679 , n437680 , n437681 , n437682 , n437683 , n437684 , n437685 , n437686 , n437687 , n437688 , 
 n437689 , n437690 , n437691 , n437692 , n437693 , n437694 , n437695 , n437696 , n437697 , n437698 , 
 n437699 , n437700 , n437701 , n437702 , n437703 , n437704 , n437705 , n437706 , n437707 , n437708 , 
 n437709 , n437710 , n437711 , n437712 , n437713 , n437714 , n437715 , n437716 , n437717 , n437718 , 
 n437719 , n437720 , n437721 , n437722 , n437723 , n437724 , n437725 , n437726 , n437727 , n437728 , 
 n437729 , n437730 , n437731 , n437732 , n437733 , n437734 , n437735 , n437736 , n437737 , n437738 , 
 n437739 , n437740 , n437741 , n437742 , n437743 , n437744 , n437745 , n437746 , n437747 , n437748 , 
 n437749 , n437750 , n437751 , n437752 , n437753 , n437754 , n437755 , n437756 , n437757 , n437758 , 
 n437759 , n437760 , n437761 , n437762 , n437763 , n437764 , n437765 , n437766 , n437767 , n437768 , 
 n437769 , n437770 , n437771 , n437772 , n437773 , n437774 , n437775 , n437776 , n437777 , n437778 , 
 n437779 , n437780 , n437781 , n437782 , n437783 , n437784 , n437785 , n437786 , n437787 , n437788 , 
 n437789 , n437790 , n437791 , n437792 , n437793 , n437794 , n437795 , n437796 , n437797 , n437798 , 
 n437799 , n437800 , n437801 , n437802 , n437803 , n437804 , n437805 , n437806 , n437807 , n437808 , 
 n437809 , n437810 , n437811 , n437812 , n437813 , n437814 , n437815 , n437816 , n437817 , n437818 , 
 n437819 , n437820 , n437821 , n437822 , n437823 , n437824 , n437825 , n437826 , n437827 , n437828 , 
 n437829 , n437830 , n437831 , n437832 , n437833 , n437834 , n437835 , n437836 , n437837 , n437838 , 
 n437839 , n437840 , n437841 , n437842 , n437843 , n437844 , n437845 , n437846 , n437847 , n437848 , 
 n437849 , n437850 , n437851 , n437852 , n437853 , n437854 , n437855 , n437856 , n437857 , n437858 , 
 n437859 , n437860 , n437861 , n437862 , n437863 , n437864 , n437865 , n437866 , n437867 , n437868 , 
 n437869 , n437870 , n437871 , n437872 , n437873 , n437874 , n437875 , n437876 , n437877 , n437878 , 
 n437879 , n437880 , n437881 , n437882 , n437883 , n437884 , n437885 , n437886 , n437887 , n437888 , 
 n437889 , n437890 , n437891 , n437892 , n437893 , n437894 , n437895 , n437896 , n437897 , n437898 , 
 n437899 , n437900 , n437901 , n437902 , n437903 , n437904 , n437905 , n437906 , n437907 , n437908 , 
 n437909 , n437910 , n437911 , n437912 , n437913 , n437914 , n437915 , n437916 , n437917 , n437918 , 
 n437919 , n437920 , n437921 , n437922 , n437923 , n437924 , n437925 , n437926 , n437927 , n437928 , 
 n437929 , n437930 , n437931 , n437932 , n437933 , n437934 , n437935 , n437936 , n437937 , n437938 , 
 n437939 , n437940 , n437941 , n437942 , n437943 , n437944 , n437945 , n437946 , n437947 , n437948 , 
 n437949 , n437950 , n437951 , n437952 , n437953 , n437954 , n437955 , n437956 , n437957 , n437958 , 
 n437959 , n437960 , n437961 , n437962 , n437963 , n437964 , n437965 , n437966 , n437967 , n437968 , 
 n437969 , n437970 , n437971 , n437972 , n437973 , n437974 , n437975 , n437976 , n437977 , n437978 , 
 n437979 , n437980 , n437981 , n437982 , n437983 , n437984 , n437985 , n437986 , n437987 , n437988 , 
 n437989 , n437990 , n437991 , n437992 , n437993 , n437994 , n437995 , n437996 , n437997 , n437998 , 
 n437999 , n438000 , n438001 , n438002 , n438003 , n438004 , n438005 , n438006 , n438007 , n438008 , 
 n438009 , n438010 , n438011 , n438012 , n438013 , n438014 , n438015 , n438016 , n438017 , n438018 , 
 n438019 , n438020 , n438021 , n438022 , n438023 , n438024 , n438025 , n438026 , n438027 , n438028 , 
 n438029 , n438030 , n438031 , n438032 , n438033 , n438034 , n438035 , n438036 , n438037 , n438038 , 
 n438039 , n438040 , n438041 , n438042 , n438043 , n438044 , n438045 , n438046 , n438047 , n438048 , 
 n438049 , n438050 , n438051 , n438052 , n438053 , n438054 , n438055 , n438056 , n438057 , n438058 , 
 n438059 , n438060 , n438061 , n438062 , n438063 , n438064 , n438065 , n438066 , n438067 , n438068 , 
 n438069 , n438070 , n438071 , n438072 , n438073 , n438074 , n438075 , n438076 , n438077 , n438078 , 
 n438079 , n438080 , n438081 , n438082 , n438083 , n438084 , n438085 , n438086 , n438087 , n438088 , 
 n438089 , n438090 , n438091 , n438092 , n438093 , n438094 , n438095 , n438096 , n438097 , n438098 , 
 n438099 , n438100 , n438101 , n438102 , n438103 , n438104 , n438105 , n438106 , n438107 , n438108 , 
 n438109 , n438110 , n438111 , n438112 , n438113 , n438114 , n438115 , n438116 , n438117 , n438118 , 
 n438119 , n438120 , n438121 , n438122 , n438123 , n438124 , n438125 , n438126 , n438127 , n438128 , 
 n438129 , n438130 , n438131 , n438132 , n438133 , n438134 , n438135 , n438136 , n438137 , n438138 , 
 n438139 , n438140 , n438141 , n438142 , n438143 , n438144 , n438145 , n438146 , n438147 , n438148 , 
 n438149 , n438150 , n438151 , n438152 , n438153 , n438154 , n438155 , n438156 , n438157 , n438158 , 
 n438159 , n438160 , n438161 , n438162 , n438163 , n438164 , n438165 , n438166 , n438167 , n438168 , 
 n438169 , n438170 , n438171 , n438172 , n438173 , n438174 , n438175 , n438176 , n438177 , n438178 , 
 n438179 , n438180 , n438181 , n438182 , n438183 , n438184 , n438185 , n438186 , n438187 , n438188 , 
 n438189 , n438190 , n438191 , n438192 , n438193 , n438194 , n438195 , n438196 , n438197 , n438198 , 
 n438199 , n438200 , n438201 , n438202 , n438203 , n438204 , n438205 , n438206 , n438207 , n438208 , 
 n438209 , n438210 , n438211 , n438212 , n438213 , n438214 , n438215 , n438216 , n438217 , n438218 , 
 n438219 , n438220 , n438221 , n438222 , n438223 , n438224 , n438225 , n438226 , n438227 , n438228 , 
 n438229 , n438230 , n438231 , n438232 , n438233 , n438234 , n438235 , n438236 , n438237 , n438238 , 
 n438239 , n438240 , n438241 , n438242 , n438243 , n438244 , n438245 , n438246 , n438247 , n438248 , 
 n438249 , n438250 , n438251 , n438252 , n438253 , n438254 , n438255 , n438256 , n438257 , n438258 , 
 n438259 , n438260 , n438261 , n438262 , n438263 , n438264 , n438265 , n438266 , n438267 , n438268 , 
 n438269 , n438270 , n438271 , n438272 , n438273 , n438274 , n438275 , n438276 , n438277 , n438278 , 
 n438279 , n438280 , n438281 , n438282 , n438283 , n438284 , n438285 , n438286 , n438287 , n438288 , 
 n438289 , n438290 , n438291 , n438292 , n438293 , n438294 , n438295 , n438296 , n438297 , n438298 , 
 n438299 , n438300 , n438301 , n438302 , n438303 , n438304 , n438305 , n438306 , n438307 , n438308 , 
 n438309 , n438310 , n438311 , n438312 , n438313 , n438314 , n438315 , n438316 , n438317 , n438318 , 
 n438319 , n438320 , n438321 , n438322 , n438323 , n438324 , n438325 , n438326 , n438327 , n438328 , 
 n438329 , n438330 , n438331 , n438332 , n438333 , n438334 , n438335 , n438336 , n438337 , n438338 , 
 n438339 , n438340 , n438341 , n438342 , n438343 , n438344 , n438345 , n438346 , n438347 , n438348 , 
 n438349 , n438350 , n438351 , n438352 , n438353 , n438354 , n438355 , n438356 , n438357 , n438358 , 
 n438359 , n438360 , n438361 , n438362 , n438363 , n438364 , n438365 , n438366 , n438367 , n438368 , 
 n438369 , n438370 , n438371 , n438372 , n438373 , n438374 , n438375 , n438376 , n438377 , n438378 , 
 n438379 , n438380 , n438381 , n438382 , n438383 , n438384 , n438385 , n438386 , n438387 , n438388 , 
 n438389 , n438390 , n438391 , n438392 , n438393 , n438394 , n438395 , n438396 , n438397 , n438398 , 
 n438399 , n438400 , n438401 , n438402 , n438403 , n438404 , n438405 , n438406 , n438407 , n438408 , 
 n438409 , n438410 , n438411 , n438412 , n438413 , n438414 , n438415 , n438416 , n438417 , n438418 , 
 n438419 , n438420 , n438421 , n438422 , n438423 , n438424 , n438425 , n438426 , n438427 , n438428 , 
 n438429 , n438430 , n438431 , n438432 , n438433 , n438434 , n438435 , n438436 , n438437 , n438438 , 
 n438439 , n438440 , n438441 , n438442 , n438443 , n438444 , n438445 , n438446 , n438447 , n438448 , 
 n438449 , n438450 , n438451 , n438452 , n438453 , n438454 , n438455 , n438456 , n438457 , n438458 , 
 n438459 , n438460 , n438461 , n438462 , n438463 , n438464 , n438465 , n438466 , n438467 , n438468 , 
 n438469 , n438470 , n438471 , n438472 , n438473 , n438474 , n438475 , n438476 , n438477 , n438478 , 
 n438479 , n438480 , n438481 , n438482 , n438483 , n438484 , n438485 , n438486 , n438487 , n438488 , 
 n438489 , n438490 , n438491 , n438492 , n438493 , n438494 , n438495 , n438496 , n438497 , n438498 , 
 n438499 , n438500 , n438501 , n438502 , n438503 , n438504 , n438505 , n438506 , n438507 , n438508 , 
 n438509 , n438510 , n438511 , n438512 , n438513 , n438514 , n438515 , n438516 , n438517 , n438518 , 
 n438519 , n438520 , n438521 , n438522 , n438523 , n438524 , n438525 , n438526 , n438527 , n438528 , 
 n438529 , n438530 , n438531 , n438532 , n438533 , n438534 , n438535 , n438536 , n438537 , n438538 , 
 n438539 , n438540 , n438541 , n438542 , n438543 , n438544 , n438545 , n438546 , n438547 , n438548 , 
 n438549 , n438550 , n438551 , n438552 , n438553 , n438554 , n438555 , n438556 , n438557 , n438558 , 
 n438559 , n438560 , n438561 , n438562 , n438563 , n438564 , n438565 , n438566 , n438567 , n438568 , 
 n438569 , n438570 , n438571 , n438572 , n438573 , n438574 , n438575 , n438576 , n438577 , n438578 , 
 n438579 , n438580 , n438581 , n438582 , n438583 , n438584 , n438585 , n438586 , n438587 , n438588 , 
 n438589 , n438590 , n438591 , n438592 , n438593 , n438594 , n438595 , n438596 , n438597 , n438598 , 
 n438599 , n438600 , n438601 , n438602 , n438603 , n438604 , n438605 , n438606 , n438607 , n438608 , 
 n438609 , n438610 , n438611 , n438612 , n438613 , n438614 , n438615 , n438616 , n438617 , n438618 , 
 n438619 , n438620 , n438621 , n438622 , n438623 , n438624 , n438625 , n438626 , n438627 , n438628 , 
 n438629 , n438630 , n438631 , n438632 , n438633 , n438634 , n438635 , n438636 , n438637 , n438638 , 
 n438639 , n438640 , n438641 , n438642 , n438643 , n438644 , n438645 , n438646 , n438647 , n438648 , 
 n438649 , n438650 , n438651 , n438652 , n438653 , n438654 , n438655 , n438656 , n438657 , n438658 , 
 n438659 , n438660 , n438661 , n438662 , n438663 , n438664 , n438665 , n438666 , n438667 , n438668 , 
 n438669 , n438670 , n438671 , n438672 , n438673 , n438674 , n438675 , n438676 , n438677 , n438678 , 
 n438679 , n438680 , n438681 , n438682 , n438683 , n438684 , n438685 , n438686 , n438687 , n438688 , 
 n438689 , n438690 , n438691 , n438692 , n438693 , n438694 , n438695 , n438696 , n438697 , n438698 , 
 n438699 , n438700 , n438701 , n438702 , n438703 , n438704 , n438705 , n438706 , n438707 , n438708 , 
 n438709 , n438710 , n438711 , n438712 , n438713 , n438714 , n438715 , n438716 , n438717 , n438718 , 
 n438719 , n438720 , n438721 , n438722 , n438723 , n438724 , n438725 , n438726 , n438727 , n438728 , 
 n438729 , n438730 , n438731 , n438732 , n438733 , n438734 , n438735 , n438736 , n438737 , n438738 , 
 n438739 , n438740 , n438741 , n438742 , n438743 , n438744 , n438745 , n438746 , n438747 , n438748 , 
 n438749 , n438750 , n438751 , n438752 , n438753 , n438754 , n438755 , n438756 , n438757 , n438758 , 
 n438759 , n438760 , n438761 , n438762 , n438763 , n438764 , n438765 , n438766 , n438767 , n438768 , 
 n438769 , n438770 , n438771 , n438772 , n438773 , n438774 , n438775 , n438776 , n438777 , n438778 , 
 n438779 , n438780 , n438781 , n438782 , n438783 , n438784 , n438785 , n438786 , n438787 , n438788 , 
 n438789 , n438790 , n438791 , n438792 , n438793 , n438794 , n438795 , n438796 , n438797 , n438798 , 
 n438799 , n438800 , n438801 , n438802 , n438803 , n438804 , n438805 , n438806 , n438807 , n438808 , 
 n438809 , n438810 , n438811 , n438812 , n438813 , n438814 , n438815 , n438816 , n438817 , n438818 , 
 n438819 , n438820 , n438821 , n438822 , n438823 , n438824 , n438825 , n438826 , n438827 , n438828 , 
 n438829 , n438830 , n438831 , n438832 , n438833 , n438834 , n438835 , n438836 , n438837 , n438838 , 
 n438839 , n438840 , n438841 , n438842 , n438843 , n438844 , n438845 , n438846 , n438847 , n438848 , 
 n438849 , n438850 , n438851 , n438852 , n438853 , n438854 , n438855 , n438856 , n438857 , n438858 , 
 n438859 , n438860 , n438861 , n438862 , n438863 , n438864 , n438865 , n438866 , n438867 , n438868 , 
 n438869 , n438870 , n438871 , n438872 , n438873 , n438874 , n438875 , n438876 , n438877 , n438878 , 
 n438879 , n438880 , n438881 , n438882 , n438883 , n438884 , n438885 , n438886 , n438887 , n438888 , 
 n438889 , n438890 , n438891 , n438892 , n438893 , n438894 , n438895 , n438896 , n438897 , n438898 , 
 n438899 , n438900 , n438901 , n438902 , n438903 , n438904 , n438905 , n438906 , n438907 , n438908 , 
 n438909 , n438910 , n438911 , n438912 , n438913 , n438914 , n438915 , n438916 , n438917 , n438918 , 
 n438919 , n438920 , n438921 , n438922 , n438923 , n438924 , n438925 , n438926 , n438927 , n438928 , 
 n438929 , n438930 , n438931 , n438932 , n438933 , n438934 , n438935 , n438936 , n438937 , n438938 , 
 n438939 , n438940 , n438941 , n438942 , n438943 , n438944 , n438945 , n438946 , n438947 , n438948 , 
 n438949 , n438950 , n438951 , n438952 , n438953 , n438954 , n438955 , n438956 , n438957 , n438958 , 
 n438959 , n438960 , n438961 , n438962 , n438963 , n438964 , n438965 , n438966 , n438967 , n438968 , 
 n438969 , n438970 , n438971 , n438972 , n438973 , n438974 , n438975 , n438976 , n438977 , n438978 , 
 n438979 , n438980 , n438981 , n438982 , n438983 , n438984 , n438985 , n438986 , n438987 , n438988 , 
 n438989 , n438990 , n438991 , n438992 , n438993 , n438994 , n438995 , n438996 , n438997 , n438998 , 
 n438999 , n439000 , n439001 , n439002 , n439003 , n439004 , n439005 , n439006 , n439007 , n439008 , 
 n439009 , n439010 , n439011 , n439012 , n439013 , n439014 , n439015 , n439016 , n439017 , n439018 , 
 n439019 , n439020 , n439021 , n439022 , n439023 , n439024 , n439025 , n439026 , n439027 , n439028 , 
 n439029 , n439030 , n439031 , n439032 , n439033 , n439034 , n439035 , n439036 , n439037 , n439038 , 
 n439039 , n439040 , n439041 , n439042 , n439043 , n439044 , n439045 , n439046 , n439047 , n439048 , 
 n439049 , n439050 , n439051 , n439052 , n439053 , n439054 , n439055 , n439056 , n439057 , n439058 , 
 n439059 , n439060 , n439061 , n439062 , n439063 , n439064 , n439065 , n439066 , n439067 , n439068 , 
 n439069 , n439070 , n439071 , n439072 , n439073 , n439074 , n439075 , n439076 , n439077 , n439078 , 
 n439079 , n439080 , n439081 , n439082 , n439083 , n439084 , n439085 , n439086 , n439087 , n439088 , 
 n439089 , n439090 , n439091 , n439092 , n439093 , n439094 , n439095 , n439096 , n439097 , n439098 , 
 n439099 , n439100 , n439101 , n439102 , n439103 , n439104 , n439105 , n439106 , n439107 , n439108 , 
 n439109 , n439110 , n439111 , n439112 , n439113 , n439114 , n439115 , n439116 , n439117 , n439118 , 
 n439119 , n439120 , n439121 , n439122 , n439123 , n439124 , n439125 , n439126 , n439127 , n439128 , 
 n439129 , n439130 , n439131 , n439132 , n439133 , n439134 , n439135 , n439136 , n439137 , n439138 , 
 n439139 , n439140 , n439141 , n439142 , n439143 , n439144 , n439145 , n439146 , n439147 , n439148 , 
 n439149 , n439150 , n439151 , n439152 , n439153 , n439154 , n439155 , n439156 , n439157 , n439158 , 
 n439159 , n439160 , n439161 , n439162 , n439163 , n439164 , n439165 , n439166 , n439167 , n439168 , 
 n439169 , n439170 , n439171 , n439172 , n439173 , n439174 , n439175 , n439176 , n439177 , n439178 , 
 n439179 , n439180 , n439181 , n439182 , n439183 , n439184 , n439185 , n439186 , n439187 , n439188 , 
 n439189 , n439190 , n439191 , n439192 , n439193 , n439194 , n439195 , n439196 , n439197 , n439198 , 
 n439199 , n439200 , n439201 , n439202 , n439203 , n439204 , n439205 , n439206 , n439207 , n439208 , 
 n439209 , n439210 , n439211 , n439212 , n439213 , n439214 , n439215 , n439216 , n439217 , n439218 , 
 n439219 , n439220 , n439221 , n439222 , n439223 , n439224 , n439225 , n439226 , n439227 , n439228 , 
 n439229 , n439230 , n439231 , n439232 , n439233 , n439234 , n439235 , n439236 , n439237 , n439238 , 
 n439239 , n439240 , n439241 , n439242 , n439243 , n439244 , n439245 , n439246 , n439247 , n439248 , 
 n439249 , n439250 , n439251 , n439252 , n439253 , n439254 , n439255 , n439256 , n439257 , n439258 , 
 n439259 , n439260 , n439261 , n439262 , n439263 , n439264 , n439265 , n439266 , n439267 , n439268 , 
 n439269 , n439270 , n439271 , n439272 , n439273 , n439274 , n439275 , n439276 , n439277 , n439278 , 
 n439279 , n439280 , n439281 , n439282 , n439283 , n439284 , n439285 , n439286 , n439287 , n439288 , 
 n439289 , n439290 , n439291 , n439292 , n439293 , n439294 , n439295 , n439296 , n439297 , n439298 , 
 n439299 , n439300 , n439301 , n439302 , n439303 , n439304 , n439305 , n439306 , n439307 , n439308 , 
 n439309 , n439310 , n439311 , n439312 , n439313 , n439314 , n439315 , n439316 , n439317 , n439318 , 
 n439319 , n439320 , n439321 , n439322 , n439323 , n439324 , n439325 , n439326 , n439327 , n439328 , 
 n439329 , n439330 , n439331 , n439332 , n439333 , n439334 , n439335 , n439336 , n439337 , n439338 , 
 n439339 , n439340 , n439341 , n439342 , n439343 , n439344 , n439345 , n439346 , n439347 , n439348 , 
 n439349 , n439350 , n439351 , n439352 , n439353 , n439354 , n439355 , n439356 , n439357 , n439358 , 
 n439359 , n439360 , n439361 , n439362 , n439363 , n439364 , n439365 , n439366 , n439367 , n439368 , 
 n439369 , n439370 , n439371 , n439372 , n439373 , n439374 , n439375 , n439376 , n439377 , n439378 , 
 n439379 , n439380 , n439381 , n439382 , n439383 , n439384 , n439385 , n439386 , n439387 , n439388 , 
 n439389 , n439390 , n439391 , n439392 , n439393 , n439394 , n439395 , n439396 , n439397 , n439398 , 
 n439399 , n439400 , n439401 , n439402 , n439403 , n439404 , n439405 , n439406 , n439407 , n439408 , 
 n439409 , n439410 , n439411 , n439412 , n439413 , n439414 , n439415 , n439416 , n439417 , n439418 , 
 n439419 , n439420 , n439421 , n439422 , n439423 , n439424 , n439425 , n439426 , n439427 , n439428 , 
 n439429 , n439430 , n439431 , n439432 , n439433 , n439434 , n439435 , n439436 , n439437 , n439438 , 
 n439439 , n439440 , n439441 , n439442 , n439443 , n439444 , n439445 , n439446 , n439447 , n439448 , 
 n439449 , n439450 , n439451 , n439452 , n439453 , n439454 , n439455 , n439456 , n439457 , n439458 , 
 n439459 , n439460 , n439461 , n439462 , n439463 , n439464 , n439465 , n439466 , n439467 , n439468 , 
 n439469 , n439470 , n439471 , n439472 , n439473 , n439474 , n439475 , n439476 , n439477 , n439478 , 
 n439479 , n439480 , n439481 , n439482 , n439483 , n439484 , n439485 , n439486 , n439487 , n439488 , 
 n439489 , n439490 , n439491 , n439492 , n439493 , n439494 , n439495 , n439496 , n439497 , n439498 , 
 n439499 , n439500 , n439501 , n439502 , n439503 , n439504 , n439505 , n439506 , n439507 , n439508 , 
 n439509 , n439510 , n439511 , n439512 , n439513 , n439514 , n439515 , n439516 , n439517 , n439518 , 
 n439519 , n439520 , n439521 , n439522 , n439523 , n439524 , n439525 , n439526 , n439527 , n439528 , 
 n439529 , n439530 , n439531 , n439532 , n439533 , n439534 , n439535 , n439536 , n439537 , n439538 , 
 n439539 , n439540 , n439541 , n439542 , n439543 , n439544 , n439545 , n439546 , n439547 , n439548 , 
 n439549 , n439550 , n439551 , n439552 , n439553 , n439554 , n439555 , n439556 , n439557 , n439558 , 
 n439559 , n439560 , n439561 , n439562 , n439563 , n439564 , n439565 , n439566 , n439567 , n439568 , 
 n439569 , n439570 , n439571 , n439572 , n439573 , n439574 , n439575 , n439576 , n439577 , n439578 , 
 n439579 , n439580 , n439581 , n439582 , n439583 , n439584 , n439585 , n439586 , n439587 , n439588 , 
 n439589 , n439590 , n439591 , n439592 , n439593 , n439594 , n439595 , n439596 , n439597 , n439598 , 
 n439599 , n439600 , n439601 , n439602 , n439603 , n439604 , n439605 , n439606 , n439607 , n439608 , 
 n439609 , n439610 , n439611 , n439612 , n439613 , n439614 , n439615 , n439616 , n439617 , n439618 , 
 n439619 , n439620 , n439621 , n439622 , n439623 , n439624 , n439625 , n439626 , n439627 , n439628 , 
 n439629 , n439630 , n439631 , n439632 , n439633 , n439634 , n439635 , n439636 , n439637 , n439638 , 
 n439639 , n439640 , n439641 , n439642 , n439643 , n439644 , n439645 , n439646 , n439647 , n439648 , 
 n439649 , n439650 , n439651 , n439652 , n439653 , n439654 , n439655 , n439656 , n439657 , n439658 , 
 n439659 , n439660 , n439661 , n439662 , n439663 , n439664 , n439665 , n439666 , n439667 , n439668 , 
 n439669 , n439670 , n439671 , n439672 , n439673 , n439674 , n439675 , n439676 , n439677 , n439678 , 
 n439679 , n439680 , n439681 , n439682 , n439683 , n439684 , n439685 , n439686 , n439687 , n439688 , 
 n439689 , n439690 , n439691 , n439692 , n439693 , n439694 , n439695 , n439696 , n439697 , n439698 , 
 n439699 , n439700 , n439701 , n439702 , n439703 , n439704 , n439705 , n439706 , n439707 , n439708 , 
 n439709 , n439710 , n439711 , n439712 , n439713 , n439714 , n439715 , n439716 , n439717 , n439718 , 
 n439719 , n439720 , n439721 , n439722 , n439723 , n439724 , n439725 , n439726 , n439727 , n439728 , 
 n439729 , n439730 , n439731 , n439732 , n439733 , n439734 , n439735 , n439736 , n439737 , n439738 , 
 n439739 , n439740 , n439741 , n439742 , n439743 , n439744 , n439745 , n439746 , n439747 , n439748 , 
 n439749 , n439750 , n439751 , n439752 , n439753 , n439754 , n439755 , n439756 , n439757 , n439758 , 
 n439759 , n439760 , n439761 , n439762 , n439763 , n439764 , n439765 , n439766 , n439767 , n439768 , 
 n439769 , n439770 , n439771 , n439772 , n439773 , n439774 , n439775 , n439776 , n439777 , n439778 , 
 n439779 , n439780 , n439781 , n439782 , n439783 , n439784 , n439785 , n439786 , n439787 , n439788 , 
 n439789 , n439790 , n439791 , n439792 , n439793 , n439794 , n439795 , n439796 , n439797 , n439798 , 
 n439799 , n439800 , n439801 , n439802 , n439803 , n439804 , n439805 , n439806 , n439807 , n439808 , 
 n439809 , n439810 , n439811 , n439812 , n439813 , n439814 , n439815 , n439816 , n439817 , n439818 , 
 n439819 , n439820 , n439821 , n439822 , n439823 , n439824 , n439825 , n439826 , n439827 , n439828 , 
 n439829 , n439830 , n439831 , n439832 , n439833 , n439834 , n439835 , n439836 , n439837 , n439838 , 
 n439839 , n439840 , n439841 , n439842 , n439843 , n439844 , n439845 , n439846 , n439847 , n439848 , 
 n439849 , n439850 , n439851 , n439852 , n439853 , n439854 , n439855 , n439856 , n439857 , n439858 , 
 n439859 , n439860 , n439861 , n439862 , n439863 , n439864 , n439865 , n439866 , n439867 , n439868 , 
 n439869 , n439870 , n439871 , n439872 , n439873 , n439874 , n439875 , n439876 , n439877 , n439878 , 
 n439879 , n439880 , n439881 , n439882 , n439883 , n439884 , n439885 , n439886 , n439887 , n439888 , 
 n439889 , n439890 , n439891 , n439892 , n439893 , n439894 , n439895 , n439896 , n439897 , n439898 , 
 n439899 , n439900 , n439901 , n439902 , n439903 , n439904 , n439905 , n439906 , n439907 , n439908 , 
 n439909 , n439910 , n439911 , n439912 , n439913 , n439914 , n439915 , n439916 , n439917 , n439918 , 
 n439919 , n439920 , n439921 , n439922 , n439923 , n439924 , n439925 , n439926 , n439927 , n439928 , 
 n439929 , n439930 , n439931 , n439932 , n439933 , n439934 , n439935 , n439936 , n439937 , n439938 , 
 n439939 , n439940 , n439941 , n439942 , n439943 , n439944 , n439945 , n439946 , n439947 , n439948 , 
 n439949 , n439950 , n439951 , n439952 , n439953 , n439954 , n439955 , n439956 , n439957 , n439958 , 
 n439959 , n439960 , n439961 , n439962 , n439963 , n439964 , n439965 , n439966 , n439967 , n439968 , 
 n439969 , n439970 , n439971 , n439972 , n439973 , n439974 , n439975 , n439976 , n439977 , n439978 , 
 n439979 , n439980 , n439981 , n439982 , n439983 , n439984 , n439985 , n439986 , n439987 , n439988 , 
 n439989 , n439990 , n439991 , n439992 , n439993 , n439994 , n439995 , n439996 , n439997 , n439998 , 
 n439999 , n440000 , n440001 , n440002 , n440003 , n440004 , n440005 , n440006 , n440007 , n440008 , 
 n440009 , n440010 , n440011 , n440012 , n440013 , n440014 , n440015 , n440016 , n440017 , n440018 , 
 n440019 , n440020 , n440021 , n440022 , n440023 , n440024 , n440025 , n440026 , n440027 , n440028 , 
 n440029 , n440030 , n440031 , n440032 , n440033 , n440034 , n440035 , n440036 , n440037 , n440038 , 
 n440039 , n440040 , n440041 , n440042 , n440043 , n440044 , n440045 , n440046 , n440047 , n440048 , 
 n440049 , n440050 , n440051 , n440052 , n440053 , n440054 , n440055 , n440056 , n440057 , n440058 , 
 n440059 , n440060 , n440061 , n440062 , n440063 , n440064 , n440065 , n440066 , n440067 , n440068 , 
 n440069 , n440070 , n440071 , n440072 , n440073 , n440074 , n440075 , n440076 , n440077 , n440078 , 
 n440079 , n440080 , n440081 , n440082 , n440083 , n440084 , n440085 , n440086 , n440087 , n440088 , 
 n440089 , n440090 , n440091 , n440092 , n440093 , n440094 , n440095 , n440096 , n440097 , n440098 , 
 n440099 , n440100 , n440101 , n440102 , n440103 , n440104 , n440105 , n440106 , n440107 , n440108 , 
 n440109 , n440110 , n440111 , n440112 , n440113 , n440114 , n440115 , n440116 , n440117 , n440118 , 
 n440119 , n440120 , n440121 , n440122 , n440123 , n440124 , n440125 , n440126 , n440127 , n440128 , 
 n440129 , n440130 , n440131 , n440132 , n440133 , n440134 , n440135 , n440136 , n440137 , n440138 , 
 n440139 , n440140 , n440141 , n440142 , n440143 , n440144 , n440145 , n440146 , n440147 , n440148 , 
 n440149 , n440150 , n440151 , n440152 , n440153 , n440154 , n440155 , n440156 , n440157 , n440158 , 
 n440159 , n440160 , n440161 , n440162 , n440163 , n440164 , n440165 , n440166 , n440167 , n440168 , 
 n440169 , n440170 , n440171 , n440172 , n440173 , n440174 , n440175 , n440176 , n440177 , n440178 , 
 n440179 , n440180 , n440181 , n440182 , n440183 , n440184 , n440185 , n440186 , n440187 , n440188 , 
 n440189 , n440190 , n440191 , n440192 , n440193 , n440194 , n440195 , n440196 , n440197 , n440198 , 
 n440199 , n440200 , n440201 , n440202 , n440203 , n440204 , n440205 , n440206 , n440207 , n440208 , 
 n440209 , n440210 , n440211 , n440212 , n440213 , n440214 , n440215 , n440216 , n440217 , n440218 , 
 n440219 , n440220 , n440221 , n440222 , n440223 , n440224 , n440225 , n440226 , n440227 , n440228 , 
 n440229 , n440230 , n440231 , n440232 , n440233 , n440234 , n440235 , n440236 , n440237 , n440238 , 
 n440239 , n440240 , n440241 , n440242 , n440243 , n440244 , n440245 , n440246 , n440247 , n440248 , 
 n440249 , n440250 , n440251 , n440252 , n440253 , n440254 , n440255 , n440256 , n440257 , n440258 , 
 n440259 , n440260 , n440261 , n440262 , n440263 , n440264 , n440265 , n440266 , n440267 , n440268 , 
 n440269 , n440270 , n440271 , n440272 , n440273 , n440274 , n440275 , n440276 , n440277 , n440278 , 
 n440279 , n440280 , n440281 , n440282 , n440283 , n440284 , n440285 , n440286 , n440287 , n440288 , 
 n440289 , n440290 , n440291 , n440292 , n440293 , n440294 , n440295 , n440296 , n440297 , n440298 , 
 n440299 , n440300 , n440301 , n440302 , n440303 , n440304 , n440305 , n440306 , n440307 , n440308 , 
 n440309 , n440310 , n440311 , n440312 , n440313 , n440314 , n440315 , n440316 , n440317 , n440318 , 
 n440319 , n440320 , n440321 , n440322 , n440323 , n440324 , n440325 , n440326 , n440327 , n440328 , 
 n440329 , n440330 , n440331 , n440332 , n440333 , n440334 , n440335 , n440336 , n440337 , n440338 , 
 n440339 , n440340 , n440341 , n440342 , n440343 , n440344 , n440345 , n440346 , n440347 , n440348 , 
 n440349 , n440350 , n440351 , n440352 , n440353 , n440354 , n440355 , n440356 , n440357 , n440358 , 
 n440359 , n440360 , n440361 , n440362 , n440363 , n440364 , n440365 , n440366 , n440367 , n440368 , 
 n440369 , n440370 , n440371 , n440372 , n440373 , n440374 , n440375 , n440376 , n440377 , n440378 , 
 n440379 , n440380 , n440381 , n440382 , n440383 , n440384 , n440385 , n440386 , n440387 , n440388 , 
 n440389 , n440390 , n440391 , n440392 , n440393 , n440394 , n440395 , n440396 , n440397 , n440398 , 
 n440399 , n440400 , n440401 , n440402 , n440403 , n440404 , n440405 , n440406 , n440407 , n440408 , 
 n440409 , n440410 , n440411 , n440412 , n440413 , n440414 , n440415 , n440416 , n440417 , n440418 , 
 n440419 , n440420 , n440421 , n440422 , n440423 , n440424 , n440425 , n440426 , n440427 , n440428 , 
 n440429 , n440430 , n440431 , n440432 , n440433 , n440434 , n440435 , n440436 , n440437 , n440438 , 
 n440439 , n440440 , n440441 , n440442 , n440443 , n440444 , n440445 , n440446 , n440447 , n440448 , 
 n440449 , n440450 , n440451 , n440452 , n440453 , n440454 , n440455 , n440456 , n440457 , n440458 , 
 n440459 , n440460 , n440461 , n440462 , n440463 , n440464 , n440465 , n440466 , n440467 , n440468 , 
 n440469 , n440470 , n440471 , n440472 , n440473 , n440474 , n440475 , n440476 , n440477 , n440478 , 
 n440479 , n440480 , n440481 , n440482 , n440483 , n440484 , n440485 , n440486 , n440487 , n440488 , 
 n440489 , n440490 , n440491 , n440492 , n440493 , n440494 , n440495 , n440496 , n440497 , n440498 , 
 n440499 , n440500 , n440501 , n440502 , n440503 , n440504 , n440505 , n440506 , n440507 , n440508 , 
 n440509 , n440510 , n440511 , n440512 , n440513 , n440514 , n440515 , n440516 , n440517 , n440518 , 
 n440519 , n440520 , n440521 , n440522 , n440523 , n440524 , n440525 , n440526 , n440527 , n440528 , 
 n440529 , n440530 , n440531 , n440532 , n440533 , n440534 , n440535 , n440536 , n440537 , n440538 , 
 n440539 , n440540 , n440541 , n440542 , n440543 , n440544 , n440545 , n440546 , n440547 , n440548 , 
 n440549 , n440550 , n440551 , n440552 , n440553 , n440554 , n440555 , n440556 , n440557 , n440558 , 
 n440559 , n440560 , n440561 , n440562 , n440563 , n440564 , n440565 , n440566 , n440567 , n440568 , 
 n440569 , n440570 , n440571 , n440572 , n440573 , n440574 , n440575 , n440576 , n440577 , n440578 , 
 n440579 , n440580 , n440581 , n440582 , n440583 , n440584 , n440585 , n440586 , n440587 , n440588 , 
 n440589 , n440590 , n440591 , n440592 , n440593 , n440594 , n440595 , n440596 , n440597 , n440598 , 
 n440599 , n440600 , n440601 , n440602 , n440603 , n440604 , n440605 , n440606 , n440607 , n440608 , 
 n440609 , n440610 , n440611 , n440612 , n440613 , n440614 , n440615 , n440616 , n440617 , n440618 , 
 n440619 , n440620 , n440621 , n440622 , n440623 , n440624 , n440625 , n440626 , n440627 , n440628 , 
 n440629 , n440630 , n440631 , n440632 , n440633 , n440634 , n440635 , n440636 , n440637 , n440638 , 
 n440639 , n440640 , n440641 , n440642 , n440643 , n440644 , n440645 , n440646 , n440647 , n440648 , 
 n440649 , n440650 , n440651 , n440652 , n440653 , n440654 , n440655 , n440656 , n440657 , n440658 , 
 n440659 , n440660 , n440661 , n440662 , n440663 , n440664 , n440665 , n440666 , n440667 , n440668 , 
 n440669 , n440670 , n440671 , n440672 , n440673 , n440674 , n440675 , n440676 , n440677 , n440678 , 
 n440679 , n440680 , n440681 , n440682 , n440683 , n440684 , n440685 , n440686 , n440687 , n440688 , 
 n440689 , n440690 , n440691 , n440692 , n440693 , n440694 , n440695 , n440696 , n440697 , n440698 , 
 n440699 , n440700 , n440701 , n440702 , n440703 , n440704 , n440705 , n440706 , n440707 , n440708 , 
 n440709 , n440710 , n440711 , n440712 , n440713 , n440714 , n440715 , n440716 , n440717 , n440718 , 
 n440719 , n440720 , n440721 , n440722 , n440723 , n440724 , n440725 , n440726 , n440727 , n440728 , 
 n440729 , n440730 , n440731 , n440732 , n440733 , n440734 , n440735 , n440736 , n440737 , n440738 , 
 n440739 , n440740 , n440741 , n440742 , n440743 , n440744 , n440745 , n440746 , n440747 , n440748 , 
 n440749 , n440750 , n440751 , n440752 , n440753 , n440754 , n440755 , n440756 , n440757 , n440758 , 
 n440759 , n440760 , n440761 , n440762 , n440763 , n440764 , n440765 , n440766 , n440767 , n440768 , 
 n440769 , n440770 , n440771 , n440772 , n440773 , n440774 , n440775 , n440776 , n440777 , n440778 , 
 n440779 , n440780 , n440781 , n440782 , n440783 , n440784 , n440785 , n440786 , n440787 , n440788 , 
 n440789 , n440790 , n440791 , n440792 , n440793 , n440794 , n440795 , n440796 , n440797 , n440798 , 
 n440799 , n440800 , n440801 , n440802 , n440803 , n440804 , n440805 , n440806 , n440807 , n440808 , 
 n440809 , n440810 , n440811 , n440812 , n440813 , n440814 , n440815 , n440816 , n440817 , n440818 , 
 n440819 , n440820 , n440821 , n440822 , n440823 , n440824 , n440825 , n440826 , n440827 , n440828 , 
 n440829 , n440830 , n440831 , n440832 , n440833 , n440834 , n440835 , n440836 , n440837 , n440838 , 
 n440839 , n440840 , n440841 , n440842 , n440843 , n440844 , n440845 , n440846 , n440847 , n440848 , 
 n440849 , n440850 , n440851 , n440852 , n440853 , n440854 , n440855 , n440856 , n440857 , n440858 , 
 n440859 , n440860 , n440861 , n440862 , n440863 , n440864 , n440865 , n440866 , n440867 , n440868 , 
 n440869 , n440870 , n440871 , n440872 , n440873 , n440874 , n440875 , n440876 , n440877 , n440878 , 
 n440879 , n440880 , n440881 , n440882 , n440883 , n440884 , n440885 , n440886 , n440887 , n440888 , 
 n440889 , n440890 , n440891 , n440892 , n440893 , n440894 , n440895 , n440896 , n440897 , n440898 , 
 n440899 , n440900 , n440901 , n440902 , n440903 , n440904 , n440905 , n440906 , n440907 , n440908 , 
 n440909 , n440910 , n440911 , n440912 , n440913 , n440914 , n440915 , n440916 , n440917 , n440918 , 
 n440919 , n440920 , n440921 , n440922 , n440923 , n440924 , n440925 , n440926 , n440927 , n440928 , 
 n440929 , n440930 , n440931 , n440932 , n440933 , n440934 , n440935 , n440936 , n440937 , n440938 , 
 n440939 , n440940 , n440941 , n440942 , n440943 , n440944 , n440945 , n440946 , n440947 , n440948 , 
 n440949 , n440950 , n440951 , n440952 , n440953 , n440954 , n440955 , n440956 , n440957 , n440958 , 
 n440959 , n440960 , n440961 , n440962 , n440963 , n440964 , n440965 , n440966 , n440967 , n440968 , 
 n440969 , n440970 , n440971 , n440972 , n440973 , n440974 , n440975 , n440976 , n440977 , n440978 , 
 n440979 , n440980 , n440981 , n440982 , n440983 , n440984 , n440985 , n440986 , n440987 , n440988 , 
 n440989 , n440990 , n440991 , n440992 , n440993 , n440994 , n440995 , n440996 , n440997 , n440998 , 
 n440999 , n441000 , n441001 , n441002 , n441003 , n441004 , n441005 , n441006 , n441007 , n441008 , 
 n441009 , n441010 , n441011 , n441012 , n441013 , n441014 , n441015 , n441016 , n441017 , n441018 , 
 n441019 , n441020 , n441021 , n441022 , n441023 , n441024 , n441025 , n441026 , n441027 , n441028 , 
 n441029 , n441030 , n441031 , n441032 , n441033 , n441034 , n441035 , n441036 , n441037 , n441038 , 
 n441039 , n441040 , n441041 , n441042 , n441043 , n441044 , n441045 , n441046 , n441047 , n441048 , 
 n441049 , n441050 , n441051 , n441052 , n441053 , n441054 , n441055 , n441056 , n441057 , n441058 , 
 n441059 , n441060 , n441061 , n441062 , n441063 , n441064 , n441065 , n441066 , n441067 , n441068 , 
 n441069 , n441070 , n441071 , n441072 , n441073 , n441074 , n441075 , n441076 , n441077 , n441078 , 
 n441079 , n441080 , n441081 , n441082 , n441083 , n441084 , n441085 , n441086 , n441087 , n441088 , 
 n441089 , n441090 , n441091 , n441092 , n441093 , n441094 , n441095 , n441096 , n441097 , n441098 , 
 n441099 , n441100 , n441101 , n441102 , n441103 , n441104 , n441105 , n441106 , n441107 , n441108 , 
 n441109 , n441110 , n441111 , n441112 , n441113 , n441114 , n441115 , n441116 , n441117 , n441118 , 
 n441119 , n441120 , n441121 , n441122 , n441123 , n441124 , n441125 , n441126 , n441127 , n441128 , 
 n441129 , n441130 , n441131 , n441132 , n441133 , n441134 , n441135 , n441136 , n441137 , n441138 , 
 n441139 , n441140 , n441141 , n441142 , n441143 , n441144 , n441145 , n441146 , n441147 , n441148 , 
 n441149 , n441150 , n441151 , n441152 , n441153 , n441154 , n441155 , n441156 , n441157 , n441158 , 
 n441159 , n441160 , n441161 , n441162 , n441163 , n441164 , n441165 , n441166 , n441167 , n441168 , 
 n441169 , n441170 , n441171 , n441172 , n441173 , n441174 , n441175 , n441176 , n441177 , n441178 , 
 n441179 , n441180 , n441181 , n441182 , n441183 , n441184 , n441185 , n441186 , n441187 , n441188 , 
 n441189 , n441190 , n441191 , n441192 , n441193 , n441194 , n441195 , n441196 , n441197 , n441198 , 
 n441199 , n441200 , n441201 , n441202 , n441203 , n441204 , n441205 , n441206 , n441207 , n441208 , 
 n441209 , n441210 , n441211 , n441212 , n441213 , n441214 , n441215 , n441216 , n441217 , n441218 , 
 n441219 , n441220 , n441221 , n441222 , n441223 , n441224 , n441225 , n441226 , n441227 , n441228 , 
 n441229 , n441230 , n441231 , n441232 , n441233 , n441234 , n441235 , n441236 , n441237 , n441238 , 
 n441239 , n441240 , n441241 , n441242 , n441243 , n441244 , n441245 , n441246 , n441247 , n441248 , 
 n441249 , n441250 , n441251 , n441252 , n441253 , n441254 , n441255 , n441256 , n441257 , n441258 , 
 n441259 , n441260 , n441261 , n441262 , n441263 , n441264 , n441265 , n441266 , n441267 , n441268 , 
 n441269 , n441270 , n441271 , n441272 , n441273 , n441274 , n441275 , n441276 , n441277 , n441278 , 
 n441279 , n441280 , n441281 , n441282 , n441283 , n441284 , n441285 , n441286 , n441287 , n441288 , 
 n441289 , n441290 , n441291 , n441292 , n441293 , n441294 , n441295 , n441296 , n441297 , n441298 , 
 n441299 , n441300 , n441301 , n441302 , n441303 , n441304 , n441305 , n441306 , n441307 , n441308 , 
 n441309 , n441310 , n441311 , n441312 , n441313 , n441314 , n441315 , n441316 , n441317 , n441318 , 
 n441319 , n441320 , n441321 , n441322 , n441323 , n441324 , n441325 , n441326 , n441327 , n441328 , 
 n441329 , n441330 , n441331 , n441332 , n441333 , n441334 , n441335 , n441336 , n441337 , n441338 , 
 n441339 , n441340 , n441341 , n441342 , n441343 , n441344 , n441345 , n441346 , n441347 , n441348 , 
 n441349 , n441350 , n441351 , n441352 , n441353 , n441354 , n441355 , n441356 , n441357 , n441358 , 
 n441359 , n441360 , n441361 , n441362 , n441363 , n441364 , n441365 , n441366 , n441367 , n441368 , 
 n441369 , n441370 , n441371 , n441372 , n441373 , n441374 , n441375 , n441376 , n441377 , n441378 , 
 n441379 , n441380 , n441381 , n441382 , n441383 , n441384 , n441385 , n441386 , n441387 , n441388 , 
 n441389 , n441390 , n441391 , n441392 , n441393 , n441394 , n441395 , n441396 , n441397 , n441398 , 
 n441399 , n441400 , n441401 , n441402 , n441403 , n441404 , n441405 , n441406 , n441407 , n441408 , 
 n441409 , n441410 , n441411 , n441412 , n441413 , n441414 , n441415 , n441416 , n441417 , n441418 , 
 n441419 , n441420 , n441421 , n441422 , n441423 , n441424 , n441425 , n441426 , n441427 , n441428 , 
 n441429 , n441430 , n441431 , n441432 , n441433 , n441434 , n441435 , n441436 , n441437 , n441438 , 
 n441439 , n441440 , n441441 , n441442 , n441443 , n441444 , n441445 , n441446 , n441447 , n441448 , 
 n441449 , n441450 , n441451 , n441452 , n441453 , n441454 , n441455 , n441456 , n441457 , n441458 , 
 n441459 , n441460 , n441461 , n441462 , n441463 , n441464 , n441465 , n441466 , n441467 , n441468 , 
 n441469 , n441470 , n441471 , n441472 , n441473 , n441474 , n441475 , n441476 , n441477 , n441478 , 
 n441479 , n441480 , n441481 , n441482 , n441483 , n441484 , n441485 , n441486 , n441487 , n441488 , 
 n441489 , n441490 , n441491 , n441492 , n441493 , n441494 , n441495 , n441496 , n441497 , n441498 , 
 n441499 , n441500 , n441501 , n441502 , n441503 , n441504 , n441505 , n441506 , n441507 , n441508 , 
 n441509 , n441510 , n441511 , n441512 , n441513 , n441514 , n441515 , n441516 , n441517 , n441518 , 
 n441519 , n441520 , n441521 , n441522 , n441523 , n441524 , n441525 , n441526 , n441527 , n441528 , 
 n441529 , n441530 , n441531 , n441532 , n441533 , n441534 , n441535 , n441536 , n441537 , n441538 , 
 n441539 , n441540 , n441541 , n441542 , n441543 , n441544 , n441545 , n441546 , n441547 , n441548 , 
 C0n , C0 , C1n , C1 ;
buf ( n544 , n0 );
buf ( n545 , n1 );
buf ( n546 , n2 );
buf ( n547 , n3 );
buf ( n548 , n4 );
buf ( n549 , n5 );
buf ( n550 , n6 );
buf ( n551 , n7 );
buf ( n552 , n8 );
buf ( n553 , n9 );
buf ( n554 , n10 );
buf ( n555 , n11 );
buf ( n556 , n12 );
buf ( n557 , n13 );
buf ( n558 , n14 );
buf ( n559 , n15 );
buf ( n560 , n16 );
buf ( n561 , n17 );
buf ( n562 , n18 );
buf ( n563 , n19 );
buf ( n564 , n20 );
buf ( n565 , n21 );
buf ( n566 , n22 );
buf ( n567 , n23 );
buf ( n568 , n24 );
buf ( n569 , n25 );
buf ( n570 , n26 );
buf ( n571 , n27 );
buf ( n572 , n28 );
buf ( n573 , n29 );
buf ( n574 , n30 );
buf ( n575 , n31 );
buf ( n576 , n32 );
buf ( n577 , n33 );
buf ( n578 , n34 );
buf ( n579 , n35 );
buf ( n580 , n36 );
buf ( n581 , n37 );
buf ( n582 , n38 );
buf ( n583 , n39 );
buf ( n584 , n40 );
buf ( n585 , n41 );
buf ( n586 , n42 );
buf ( n587 , n43 );
buf ( n588 , n44 );
buf ( n589 , n45 );
buf ( n590 , n46 );
buf ( n591 , n47 );
buf ( n592 , n48 );
buf ( n593 , n49 );
buf ( n594 , n50 );
buf ( n595 , n51 );
buf ( n596 , n52 );
buf ( n597 , n53 );
buf ( n598 , n54 );
buf ( n599 , n55 );
buf ( n600 , n56 );
buf ( n601 , n57 );
buf ( n602 , n58 );
buf ( n603 , n59 );
buf ( n604 , n60 );
buf ( n605 , n61 );
buf ( n606 , n62 );
buf ( n607 , n63 );
buf ( n608 , n64 );
buf ( n609 , n65 );
buf ( n610 , n66 );
buf ( n611 , n67 );
buf ( n612 , n68 );
buf ( n613 , n69 );
buf ( n614 , n70 );
buf ( n615 , n71 );
buf ( n616 , n72 );
buf ( n617 , n73 );
buf ( n618 , n74 );
buf ( n619 , n75 );
buf ( n620 , n76 );
buf ( n621 , n77 );
buf ( n622 , n78 );
buf ( n623 , n79 );
buf ( n80 , n624 );
buf ( n81 , n625 );
buf ( n82 , n626 );
buf ( n83 , n627 );
buf ( n84 , n628 );
buf ( n85 , n629 );
buf ( n86 , n630 );
buf ( n87 , n631 );
buf ( n88 , n632 );
buf ( n89 , n633 );
buf ( n90 , n634 );
buf ( n91 , n635 );
buf ( n92 , n636 );
buf ( n93 , n637 );
buf ( n94 , n638 );
buf ( n95 , n639 );
buf ( n96 , n640 );
buf ( n97 , n641 );
buf ( n98 , n642 );
buf ( n99 , n643 );
buf ( n100 , n644 );
buf ( n101 , n645 );
buf ( n102 , n646 );
buf ( n103 , n647 );
buf ( n104 , n648 );
buf ( n105 , n649 );
buf ( n106 , n650 );
buf ( n107 , n651 );
buf ( n108 , n652 );
buf ( n109 , n653 );
buf ( n110 , n654 );
buf ( n111 , n655 );
buf ( n112 , n656 );
buf ( n113 , n657 );
buf ( n114 , n658 );
buf ( n115 , n659 );
buf ( n116 , n660 );
buf ( n117 , n661 );
buf ( n118 , n662 );
buf ( n119 , n663 );
buf ( n120 , n664 );
buf ( n121 , n665 );
buf ( n122 , n666 );
buf ( n123 , n667 );
buf ( n124 , n668 );
buf ( n125 , n669 );
buf ( n126 , n670 );
buf ( n127 , n671 );
buf ( n128 , n672 );
buf ( n129 , n673 );
buf ( n130 , n674 );
buf ( n131 , n675 );
buf ( n132 , n676 );
buf ( n133 , n677 );
buf ( n134 , n678 );
buf ( n135 , n679 );
buf ( n136 , n680 );
buf ( n137 , n681 );
buf ( n138 , n682 );
buf ( n139 , n683 );
buf ( n140 , n684 );
buf ( n141 , n685 );
buf ( n142 , n686 );
buf ( n143 , n687 );
buf ( n144 , n688 );
buf ( n145 , n689 );
buf ( n146 , n690 );
buf ( n147 , n691 );
buf ( n148 , n692 );
buf ( n149 , n693 );
buf ( n150 , n694 );
buf ( n151 , n695 );
buf ( n152 , n696 );
buf ( n153 , n697 );
buf ( n154 , n698 );
buf ( n155 , n699 );
buf ( n156 , n700 );
buf ( n157 , n701 );
buf ( n158 , n702 );
buf ( n159 , n703 );
buf ( n160 , n704 );
buf ( n161 , n705 );
buf ( n162 , n706 );
buf ( n163 , n707 );
buf ( n164 , n708 );
buf ( n165 , n709 );
buf ( n166 , n710 );
buf ( n167 , n711 );
buf ( n168 , n712 );
buf ( n169 , n713 );
buf ( n170 , n714 );
buf ( n171 , n715 );
buf ( n172 , n716 );
buf ( n173 , n717 );
buf ( n174 , n718 );
buf ( n175 , n719 );
buf ( n176 , n720 );
buf ( n177 , n721 );
buf ( n178 , n722 );
buf ( n179 , n723 );
buf ( n180 , n724 );
buf ( n181 , n725 );
buf ( n182 , n726 );
buf ( n183 , n727 );
buf ( n184 , n728 );
buf ( n185 , n729 );
buf ( n186 , n730 );
buf ( n187 , n731 );
buf ( n188 , n732 );
buf ( n189 , n733 );
buf ( n190 , n734 );
buf ( n191 , n735 );
buf ( n192 , n736 );
buf ( n193 , n737 );
buf ( n194 , n738 );
buf ( n195 , n739 );
buf ( n196 , n740 );
buf ( n197 , n741 );
buf ( n198 , n742 );
buf ( n199 , n743 );
buf ( n200 , n744 );
buf ( n201 , n745 );
buf ( n202 , n746 );
buf ( n203 , n747 );
buf ( n204 , n748 );
buf ( n205 , n749 );
buf ( n206 , n750 );
buf ( n207 , n751 );
buf ( n208 , n752 );
buf ( n209 , n753 );
buf ( n210 , n754 );
buf ( n211 , n755 );
buf ( n212 , n756 );
buf ( n213 , n757 );
buf ( n214 , n758 );
buf ( n215 , n759 );
buf ( n216 , n760 );
buf ( n217 , n761 );
buf ( n218 , n762 );
buf ( n219 , n763 );
buf ( n220 , n764 );
buf ( n221 , n765 );
buf ( n222 , n766 );
buf ( n223 , n767 );
buf ( n224 , n768 );
buf ( n225 , n769 );
buf ( n226 , n770 );
buf ( n227 , n771 );
buf ( n228 , n772 );
buf ( n229 , n773 );
buf ( n230 , n774 );
buf ( n231 , n775 );
buf ( n232 , n776 );
buf ( n233 , n777 );
buf ( n234 , n778 );
buf ( n235 , n779 );
buf ( n236 , n780 );
buf ( n237 , n781 );
buf ( n238 , n782 );
buf ( n239 , n783 );
buf ( n240 , n784 );
buf ( n241 , n785 );
buf ( n242 , n786 );
buf ( n243 , n787 );
buf ( n244 , n788 );
buf ( n245 , n789 );
buf ( n246 , n790 );
buf ( n247 , n791 );
buf ( n248 , n792 );
buf ( n249 , n793 );
buf ( n250 , n794 );
buf ( n251 , n795 );
buf ( n252 , n796 );
buf ( n253 , n797 );
buf ( n254 , n798 );
buf ( n255 , n799 );
buf ( n256 , n800 );
buf ( n257 , n801 );
buf ( n258 , n802 );
buf ( n259 , n803 );
buf ( n260 , n804 );
buf ( n261 , n805 );
buf ( n262 , n806 );
buf ( n263 , n807 );
buf ( n264 , n808 );
buf ( n265 , n809 );
buf ( n266 , n810 );
buf ( n267 , n811 );
buf ( n268 , n812 );
buf ( n269 , n813 );
buf ( n270 , n814 );
buf ( n271 , n815 );
buf ( n624 , n372185 );
buf ( n625 , n372203 );
buf ( n626 , n372206 );
buf ( n627 , n372209 );
buf ( n628 , n372212 );
buf ( n629 , n372215 );
buf ( n630 , n372218 );
buf ( n631 , n372221 );
buf ( n632 , n372224 );
buf ( n633 , n372227 );
buf ( n634 , n372230 );
buf ( n635 , n372233 );
buf ( n636 , n372236 );
buf ( n637 , n372239 );
buf ( n638 , n372253 );
buf ( n639 , n372267 );
buf ( n640 , n372281 );
buf ( n641 , n372289 );
buf ( n642 , n372297 );
buf ( n643 , n441530 );
buf ( n644 , n441545 );
buf ( n645 , n372309 );
buf ( n646 , n372317 );
buf ( n647 , n372320 );
buf ( n648 , n372368 );
buf ( n649 , n441532 );
buf ( n650 , n441548 );
buf ( n651 , n372328 );
buf ( n652 , n372331 );
buf ( n653 , n372350 );
buf ( n654 , n372352 );
buf ( n655 , n348025 );
buf ( n656 , n376735 );
buf ( n657 , n376753 );
buf ( n658 , n376756 );
buf ( n659 , n376759 );
buf ( n660 , n376762 );
buf ( n661 , n376765 );
buf ( n662 , n441526 );
buf ( n663 , n441529 );
buf ( n664 , n376984 );
buf ( n665 , n376980 );
buf ( n666 , n376976 );
buf ( n667 , n376972 );
buf ( n668 , n376964 );
buf ( n669 , n376960 );
buf ( n670 , n376783 );
buf ( n671 , n376795 );
buf ( n672 , n376813 );
buf ( n673 , n376827 );
buf ( n674 , n376841 );
buf ( n675 , n441511 );
buf ( n676 , n376853 );
buf ( n677 , n376856 );
buf ( n678 , n376864 );
buf ( n679 , n376872 );
buf ( n680 , n376880 );
buf ( n681 , n376892 );
buf ( n682 , n376895 );
buf ( n683 , n376898 );
buf ( n684 , n376901 );
buf ( n685 , n376904 );
buf ( n686 , n441514 );
buf ( n687 , n348036 );
buf ( n688 , n441396 );
buf ( n689 , n441396 );
buf ( n690 , n441396 );
buf ( n691 , n441396 );
buf ( n692 , n441396 );
buf ( n693 , n441396 );
buf ( n694 , n441396 );
buf ( n695 , n441396 );
buf ( n696 , n441396 );
buf ( n697 , n441396 );
buf ( n698 , n441396 );
buf ( n699 , n441396 );
buf ( n700 , n441396 );
buf ( n701 , n441396 );
buf ( n702 , n441396 );
buf ( n703 , n441396 );
buf ( n704 , n441396 );
buf ( n705 , n441396 );
buf ( n706 , n441396 );
buf ( n707 , n441396 );
buf ( n708 , n441396 );
buf ( n709 , n441396 );
buf ( n710 , n441396 );
buf ( n711 , n441396 );
buf ( n712 , n441396 );
buf ( n713 , n441396 );
buf ( n714 , n441396 );
buf ( n715 , n441396 );
buf ( n716 , n441332 );
buf ( n717 , n441347 );
buf ( n718 , n441544 );
buf ( n719 , n439667 );
buf ( n720 , n441274 );
buf ( n721 , n439702 );
buf ( n722 , n439778 );
buf ( n723 , n439728 );
buf ( n724 , n439887 );
buf ( n725 , n441467 );
buf ( n726 , n439803 );
buf ( n727 , n439759 );
buf ( n728 , n439902 );
buf ( n729 , n439928 );
buf ( n730 , n439958 );
buf ( n731 , n439875 );
buf ( n732 , n440463 );
buf ( n733 , n439989 );
buf ( n734 , n439853 );
buf ( n735 , n440015 );
buf ( n736 , n440045 );
buf ( n737 , n440071 );
buf ( n738 , n441372 );
buf ( n739 , n441359 );
buf ( n740 , n440480 );
buf ( n741 , n440099 );
buf ( n742 , n440121 );
buf ( n743 , n440148 );
buf ( n744 , n440495 );
buf ( n745 , n441293 );
buf ( n746 , n441491 );
buf ( n747 , n440314 );
buf ( n748 , n441198 );
buf ( n749 , n440216 );
buf ( n750 , n440271 );
buf ( n751 , n440289 );
buf ( n752 , n440534 );
buf ( n753 , n440422 );
buf ( n754 , n440521 );
buf ( n755 , n440446 );
buf ( n756 , n440596 );
buf ( n757 , n441393 );
buf ( n758 , n440382 );
buf ( n759 , n440359 );
buf ( n760 , n440584 );
buf ( n761 , n440650 );
buf ( n762 , n440623 );
buf ( n763 , n441307 );
buf ( n764 , n441435 );
buf ( n765 , n441297 );
buf ( n766 , n440569 );
buf ( n767 , n441402 );
buf ( n768 , n441410 );
buf ( n769 , n441232 );
buf ( n770 , n440704 );
buf ( n771 , n440727 );
buf ( n772 , n441236 );
buf ( n773 , n440768 );
buf ( n774 , n440783 );
buf ( n775 , n440809 );
buf ( n776 , n441443 );
buf ( n777 , n441485 );
buf ( n778 , n440840 );
buf ( n779 , n441454 );
buf ( n780 , n441215 );
buf ( n781 , n440866 );
buf ( n782 , n441203 );
buf ( n783 , n441446 );
buf ( n784 , n441211 );
buf ( n785 , n441430 );
buf ( n786 , n440918 );
buf ( n787 , n440933 );
buf ( n788 , n440955 );
buf ( n789 , n441498 );
buf ( n790 , n441382 );
buf ( n791 , n441494 );
buf ( n792 , n440958 );
buf ( n793 , n440972 );
buf ( n794 , n440986 );
buf ( n795 , n441004 );
buf ( n796 , n441240 );
buf ( n797 , n441415 );
buf ( n798 , n441420 );
buf ( n799 , n441523 );
buf ( n800 , n441032 );
buf ( n801 , n441265 );
buf ( n802 , n441049 );
buf ( n803 , n441052 );
buf ( n804 , n441066 );
buf ( n805 , n441505 );
buf ( n806 , n441084 );
buf ( n807 , n441106 );
buf ( n808 , n441109 );
buf ( n809 , n441111 );
buf ( n810 , n441113 );
buf ( n811 , n441123 );
buf ( n812 , n441126 );
buf ( n813 , n441136 );
buf ( n814 , n441186 );
buf ( n815 , n441190 );
buf ( n347310 , n598 );
not ( n347311 , n347310 );
buf ( n347312 , n347311 );
or ( n347313 , n347312 , n597 );
buf ( n347314 , n597 );
not ( n347315 , n347314 );
buf ( n347316 , n347315 );
or ( n347317 , n347316 , n598 );
nand ( n347318 , n347313 , n347317 );
buf ( n347319 , n347318 );
buf ( n347320 , n347319 );
not ( n347321 , n347320 );
buf ( n347322 , n596 );
not ( n347323 , n347322 );
buf ( n347324 , n559 );
buf ( n347325 , n570 );
xor ( n347326 , n347324 , n347325 );
buf ( n347327 , n347326 );
buf ( n347328 , n347327 );
not ( n347329 , n347328 );
buf ( n347330 , n571 );
buf ( n347331 , n572 );
xor ( n347332 , n347330 , n347331 );
buf ( n347333 , n347332 );
buf ( n347334 , n347333 );
not ( n347335 , n347334 );
buf ( n347336 , n347335 );
buf ( n347337 , n347336 );
xor ( n347338 , n571 , n570 );
buf ( n347339 , n347338 );
nand ( n347340 , n347337 , n347339 );
buf ( n347341 , n347340 );
buf ( n347342 , n347341 );
not ( n347343 , n347342 );
buf ( n347344 , n347343 );
buf ( n347345 , n347344 );
not ( n347346 , n347345 );
or ( n347347 , n347329 , n347346 );
buf ( n347348 , n347336 );
not ( n347349 , n347348 );
buf ( n347350 , n347349 );
buf ( n347351 , n347350 );
buf ( n347352 , n558 );
buf ( n347353 , n570 );
xor ( n347354 , n347352 , n347353 );
buf ( n347355 , n347354 );
buf ( n347356 , n347355 );
nand ( n347357 , n347351 , n347356 );
buf ( n347358 , n347357 );
buf ( n347359 , n347358 );
nand ( n347360 , n347347 , n347359 );
buf ( n347361 , n347360 );
buf ( n347362 , n557 );
buf ( n347363 , n572 );
xor ( n347364 , n347362 , n347363 );
buf ( n347365 , n347364 );
buf ( n347366 , n347365 );
not ( n347367 , n347366 );
not ( n347368 , n572 );
nand ( n347369 , n347368 , n573 );
not ( n347370 , n347369 );
not ( n347371 , n573 );
nand ( n347372 , n347371 , n572 );
not ( n347373 , n347372 );
or ( n347374 , n347370 , n347373 );
xor ( n347375 , n573 , n574 );
not ( n347376 , n347375 );
nand ( n347377 , n347374 , n347376 );
not ( n347378 , n347377 );
buf ( n347379 , n347378 );
not ( n347380 , n347379 );
or ( n347381 , n347367 , n347380 );
buf ( n347382 , n347375 );
buf ( n347383 , n347382 );
buf ( n347384 , n556 );
buf ( n347385 , n572 );
xor ( n347386 , n347384 , n347385 );
buf ( n347387 , n347386 );
buf ( n347388 , n347387 );
nand ( n347389 , n347383 , n347388 );
buf ( n347390 , n347389 );
buf ( n347391 , n347390 );
nand ( n347392 , n347381 , n347391 );
buf ( n347393 , n347392 );
xor ( n347394 , n347361 , n347393 );
buf ( n347395 , n574 );
not ( n347396 , n347395 );
buf ( n347397 , n575 );
nor ( n347398 , n347396 , n347397 );
buf ( n347399 , n347398 );
not ( n347400 , n347399 );
buf ( n347401 , n555 );
buf ( n347402 , n574 );
xor ( n347403 , n347401 , n347402 );
buf ( n347404 , n347403 );
not ( n347405 , n347404 );
or ( n347406 , n347400 , n347405 );
buf ( n347407 , n554 );
buf ( n347408 , n574 );
xor ( n347409 , n347407 , n347408 );
buf ( n347410 , n347409 );
buf ( n347411 , n347410 );
buf ( n347412 , n575 );
nand ( n347413 , n347411 , n347412 );
buf ( n347414 , n347413 );
nand ( n347415 , n347406 , n347414 );
or ( n347416 , n559 , n571 );
nand ( n347417 , n347416 , n572 );
buf ( n347418 , n559 );
buf ( n347419 , n571 );
nand ( n347420 , n347418 , n347419 );
buf ( n347421 , n347420 );
nand ( n347422 , n347417 , n347421 , n570 );
not ( n347423 , n347422 );
and ( n347424 , n347415 , n347423 );
not ( n347425 , n347415 );
and ( n347426 , n347425 , n347422 );
nor ( n347427 , n347424 , n347426 );
xor ( n347428 , n347394 , n347427 );
buf ( n347429 , n347428 );
buf ( n347430 , n347399 );
not ( n347431 , n347430 );
buf ( n347432 , n557 );
buf ( n347433 , n574 );
xor ( n347434 , n347432 , n347433 );
buf ( n347435 , n347434 );
buf ( n347436 , n347435 );
not ( n347437 , n347436 );
or ( n347438 , n347431 , n347437 );
buf ( n347439 , n556 );
buf ( n347440 , n574 );
xor ( n347441 , n347439 , n347440 );
buf ( n347442 , n347441 );
buf ( n347443 , n347442 );
buf ( n347444 , n575 );
nand ( n347445 , n347443 , n347444 );
buf ( n347446 , n347445 );
buf ( n347447 , n347446 );
nand ( n347448 , n347438 , n347447 );
buf ( n347449 , n347448 );
buf ( n347450 , n347449 );
buf ( n347451 , n559 );
buf ( n347452 , n573 );
or ( n347453 , n347451 , n347452 );
buf ( n347454 , n574 );
nand ( n347455 , n347453 , n347454 );
buf ( n347456 , n347455 );
buf ( n347457 , n347456 );
buf ( n347458 , n559 );
buf ( n347459 , n573 );
nand ( n347460 , n347458 , n347459 );
buf ( n347461 , n347460 );
buf ( n347462 , n347461 );
buf ( n347463 , n572 );
nand ( n347464 , n347457 , n347462 , n347463 );
buf ( n347465 , n347464 );
buf ( n347466 , n347465 );
not ( n347467 , n347466 );
buf ( n347468 , n347467 );
buf ( n347469 , n347468 );
and ( n347470 , n347450 , n347469 );
buf ( n347471 , n347470 );
buf ( n347472 , n347471 );
xor ( n347473 , n590 , n557 );
buf ( n347474 , n347473 );
not ( n347475 , n347474 );
not ( n347476 , n591 );
nand ( n347477 , n347476 , n590 );
not ( n347478 , n347477 );
buf ( n347479 , n347478 );
not ( n347480 , n347479 );
or ( n347481 , n347475 , n347480 );
and ( n347482 , n556 , n590 );
not ( n347483 , n556 );
not ( n347484 , n590 );
and ( n347485 , n347483 , n347484 );
nor ( n347486 , n347482 , n347485 );
buf ( n347487 , n347486 );
buf ( n347488 , n591 );
nand ( n347489 , n347487 , n347488 );
buf ( n347490 , n347489 );
buf ( n347491 , n347490 );
nand ( n347492 , n347481 , n347491 );
buf ( n347493 , n347492 );
buf ( n347494 , n347493 );
buf ( n347495 , n559 );
buf ( n347496 , n589 );
or ( n347497 , n347495 , n347496 );
buf ( n347498 , n590 );
nand ( n347499 , n347497 , n347498 );
buf ( n347500 , n347499 );
buf ( n347501 , n347500 );
buf ( n347502 , n559 );
buf ( n347503 , n589 );
nand ( n347504 , n347502 , n347503 );
buf ( n347505 , n347504 );
buf ( n347506 , n347505 );
buf ( n347507 , n588 );
nand ( n347508 , n347501 , n347506 , n347507 );
buf ( n347509 , n347508 );
buf ( n347510 , n347509 );
not ( n347511 , n347510 );
buf ( n347512 , n347511 );
buf ( n347513 , n347512 );
and ( n347514 , n347494 , n347513 );
buf ( n347515 , n347514 );
buf ( n347516 , n347515 );
xor ( n347517 , n347472 , n347516 );
not ( n347518 , n590 );
nor ( n347519 , n347518 , n591 );
not ( n347520 , n347519 );
not ( n347521 , n347486 );
or ( n347522 , n347520 , n347521 );
and ( n347523 , n590 , n555 );
not ( n347524 , n590 );
not ( n347525 , n555 );
and ( n347526 , n347524 , n347525 );
nor ( n347527 , n347523 , n347526 );
nand ( n347528 , n347527 , n591 );
nand ( n347529 , n347522 , n347528 );
xor ( n347530 , n587 , n588 );
buf ( n347531 , n347530 );
buf ( n347532 , n559 );
and ( n347533 , n347531 , n347532 );
buf ( n347534 , n347533 );
xor ( n347535 , n347529 , n347534 );
not ( n347536 , n590 );
nand ( n347537 , n347536 , n589 );
buf ( n347538 , n347537 );
buf ( n347539 , n589 );
not ( n347540 , n347539 );
buf ( n347541 , n590 );
nand ( n347542 , n347540 , n347541 );
buf ( n347543 , n347542 );
buf ( n347544 , n347543 );
buf ( n347545 , n588 );
buf ( n347546 , n589 );
xor ( n347547 , n347545 , n347546 );
buf ( n347548 , n347547 );
buf ( n347549 , n347548 );
and ( n347550 , n347538 , n347544 , n347549 );
buf ( n347551 , n347550 );
buf ( n347552 , n347551 );
buf ( n347553 , n347552 );
buf ( n347554 , n347553 );
buf ( n347555 , n347554 );
not ( n347556 , n347555 );
buf ( n347557 , n347556 );
buf ( n347558 , n347557 );
buf ( n347559 , n558 );
buf ( n347560 , n588 );
xnor ( n347561 , n347559 , n347560 );
buf ( n347562 , n347561 );
buf ( n347563 , n347562 );
or ( n347564 , n347558 , n347563 );
xor ( n347565 , n589 , n590 );
buf ( n347566 , n347565 );
buf ( n347567 , n347566 );
buf ( n347568 , n347567 );
buf ( n347569 , n347568 );
buf ( n347570 , n557 );
buf ( n347571 , n588 );
xor ( n347572 , n347570 , n347571 );
buf ( n347573 , n347572 );
buf ( n347574 , n347573 );
nand ( n347575 , n347569 , n347574 );
buf ( n347576 , n347575 );
buf ( n347577 , n347576 );
nand ( n347578 , n347564 , n347577 );
buf ( n347579 , n347578 );
xor ( n347580 , n347535 , n347579 );
buf ( n347581 , n347580 );
and ( n347582 , n347517 , n347581 );
and ( n347583 , n347472 , n347516 );
or ( n347584 , n347582 , n347583 );
buf ( n347585 , n347584 );
buf ( n347586 , n347585 );
xor ( n347587 , n347429 , n347586 );
xor ( n347588 , n347529 , n347534 );
and ( n347589 , n347588 , n347579 );
and ( n347590 , n347529 , n347534 );
or ( n347591 , n347589 , n347590 );
buf ( n347592 , n347591 );
buf ( n347593 , n347350 );
buf ( n347594 , n559 );
and ( n347595 , n347593 , n347594 );
buf ( n347596 , n347595 );
buf ( n347597 , n347596 );
buf ( n347598 , n347442 );
not ( n347599 , n347598 );
buf ( n347600 , n574 );
not ( n347601 , n347600 );
buf ( n347602 , n575 );
nor ( n347603 , n347601 , n347602 );
buf ( n347604 , n347603 );
buf ( n347605 , n347604 );
not ( n347606 , n347605 );
or ( n347607 , n347599 , n347606 );
buf ( n347608 , n347404 );
buf ( n347609 , n575 );
nand ( n347610 , n347608 , n347609 );
buf ( n347611 , n347610 );
buf ( n347612 , n347611 );
nand ( n347613 , n347607 , n347612 );
buf ( n347614 , n347613 );
buf ( n347615 , n347614 );
xor ( n347616 , n347597 , n347615 );
buf ( n347617 , n558 );
buf ( n347618 , n572 );
xor ( n347619 , n347617 , n347618 );
buf ( n347620 , n347619 );
buf ( n347621 , n347620 );
not ( n347622 , n347621 );
buf ( n347623 , n347378 );
not ( n347624 , n347623 );
or ( n347625 , n347622 , n347624 );
buf ( n347626 , n347382 );
buf ( n347627 , n347365 );
nand ( n347628 , n347626 , n347627 );
buf ( n347629 , n347628 );
buf ( n347630 , n347629 );
nand ( n347631 , n347625 , n347630 );
buf ( n347632 , n347631 );
buf ( n347633 , n347632 );
and ( n347634 , n347616 , n347633 );
and ( n347635 , n347597 , n347615 );
or ( n347636 , n347634 , n347635 );
buf ( n347637 , n347636 );
buf ( n347638 , n347637 );
xor ( n347639 , n347592 , n347638 );
buf ( n347640 , n347573 );
not ( n347641 , n347640 );
buf ( n347642 , n347554 );
not ( n347643 , n347642 );
or ( n347644 , n347641 , n347643 );
buf ( n347645 , n347565 );
buf ( n347646 , n556 );
buf ( n347647 , n588 );
xor ( n347648 , n347646 , n347647 );
buf ( n347649 , n347648 );
buf ( n347650 , n347649 );
nand ( n347651 , n347645 , n347650 );
buf ( n347652 , n347651 );
buf ( n347653 , n347652 );
nand ( n347654 , n347644 , n347653 );
buf ( n347655 , n347654 );
buf ( n347656 , n347655 );
buf ( n347657 , n559 );
buf ( n347658 , n586 );
xor ( n347659 , n347657 , n347658 );
buf ( n347660 , n347659 );
buf ( n347661 , n347660 );
not ( n347662 , n347661 );
xor ( n347663 , n587 , n588 );
not ( n347664 , n347663 );
not ( n347665 , n586 );
not ( n347666 , n587 );
and ( n347667 , n347665 , n347666 );
and ( n347668 , n586 , n587 );
nor ( n347669 , n347667 , n347668 );
nand ( n347670 , n347664 , n347669 );
not ( n347671 , n347670 );
buf ( n347672 , n347671 );
not ( n347673 , n347672 );
or ( n347674 , n347662 , n347673 );
buf ( n347675 , n347530 );
buf ( n347676 , n558 );
buf ( n347677 , n586 );
xor ( n347678 , n347676 , n347677 );
buf ( n347679 , n347678 );
buf ( n347680 , n347679 );
nand ( n347681 , n347675 , n347680 );
buf ( n347682 , n347681 );
buf ( n347683 , n347682 );
nand ( n347684 , n347674 , n347683 );
buf ( n347685 , n347684 );
buf ( n347686 , n347685 );
xor ( n347687 , n347656 , n347686 );
buf ( n347688 , n347527 );
not ( n347689 , n347688 );
buf ( n347690 , n347478 );
not ( n347691 , n347690 );
or ( n347692 , n347689 , n347691 );
and ( n347693 , n554 , n590 );
not ( n347694 , n554 );
buf ( n347695 , n590 );
not ( n347696 , n347695 );
buf ( n347697 , n347696 );
and ( n347698 , n347694 , n347697 );
nor ( n347699 , n347693 , n347698 );
buf ( n347700 , n347699 );
buf ( n347701 , n591 );
nand ( n347702 , n347700 , n347701 );
buf ( n347703 , n347702 );
buf ( n347704 , n347703 );
nand ( n347705 , n347692 , n347704 );
buf ( n347706 , n347705 );
or ( n347707 , n559 , n587 );
nand ( n347708 , n347707 , n588 );
nand ( n347709 , n559 , n587 );
and ( n347710 , n347708 , n347709 , n586 );
and ( n347711 , n347706 , n347710 );
not ( n347712 , n347706 );
not ( n347713 , n347710 );
and ( n347714 , n347712 , n347713 );
nor ( n347715 , n347711 , n347714 );
buf ( n347716 , n347715 );
xor ( n347717 , n347687 , n347716 );
buf ( n347718 , n347717 );
buf ( n347719 , n347718 );
xor ( n347720 , n347639 , n347719 );
buf ( n347721 , n347720 );
buf ( n347722 , n347721 );
xor ( n347723 , n347587 , n347722 );
buf ( n347724 , n347723 );
buf ( n347725 , n347724 );
not ( n347726 , n347725 );
xor ( n347727 , n347597 , n347615 );
xor ( n347728 , n347727 , n347633 );
buf ( n347729 , n347728 );
buf ( n347730 , n347729 );
buf ( n347731 , n559 );
buf ( n347732 , n572 );
xor ( n347733 , n347731 , n347732 );
buf ( n347734 , n347733 );
buf ( n347735 , n347734 );
not ( n347736 , n347735 );
not ( n347737 , n347377 );
buf ( n347738 , n347737 );
not ( n347739 , n347738 );
or ( n347740 , n347736 , n347739 );
buf ( n347741 , n347382 );
buf ( n347742 , n347620 );
nand ( n347743 , n347741 , n347742 );
buf ( n347744 , n347743 );
buf ( n347745 , n347744 );
nand ( n347746 , n347740 , n347745 );
buf ( n347747 , n347746 );
buf ( n347748 , n347747 );
buf ( n347749 , n559 );
buf ( n347750 , n588 );
xor ( n347751 , n347749 , n347750 );
buf ( n347752 , n347751 );
buf ( n347753 , n347752 );
not ( n347754 , n347753 );
buf ( n347755 , n347554 );
buf ( n347756 , n347755 );
buf ( n347757 , n347756 );
buf ( n347758 , n347757 );
not ( n347759 , n347758 );
or ( n347760 , n347754 , n347759 );
buf ( n347761 , n347562 );
not ( n347762 , n347761 );
buf ( n347763 , n347568 );
nand ( n347764 , n347762 , n347763 );
buf ( n347765 , n347764 );
buf ( n347766 , n347765 );
nand ( n347767 , n347760 , n347766 );
buf ( n347768 , n347767 );
buf ( n347769 , n347768 );
xor ( n347770 , n347748 , n347769 );
xnor ( n347771 , n347509 , n347493 );
buf ( n347772 , n347771 );
and ( n347773 , n347770 , n347772 );
and ( n347774 , n347748 , n347769 );
or ( n347775 , n347773 , n347774 );
buf ( n347776 , n347775 );
buf ( n347777 , n347776 );
xor ( n347778 , n347730 , n347777 );
xor ( n347779 , n347472 , n347516 );
xor ( n347780 , n347779 , n347581 );
buf ( n347781 , n347780 );
buf ( n347782 , n347781 );
and ( n347783 , n347778 , n347782 );
and ( n347784 , n347730 , n347777 );
or ( n347785 , n347783 , n347784 );
buf ( n347786 , n347785 );
buf ( n347787 , n347786 );
not ( n347788 , n347787 );
buf ( n347789 , n347788 );
buf ( n347790 , n347789 );
nand ( n347791 , n347726 , n347790 );
buf ( n347792 , n347791 );
buf ( n347793 , n347792 );
buf ( n347794 , n347724 );
buf ( n347795 , n347786 );
nand ( n347796 , n347794 , n347795 );
buf ( n347797 , n347796 );
buf ( n347798 , n347797 );
nand ( n347799 , n347793 , n347798 );
buf ( n347800 , n347799 );
xor ( n347801 , n590 , n558 );
buf ( n347802 , n347801 );
not ( n347803 , n347802 );
buf ( n347804 , n347478 );
not ( n347805 , n347804 );
or ( n347806 , n347803 , n347805 );
buf ( n347807 , n347473 );
buf ( n347808 , n591 );
nand ( n347809 , n347807 , n347808 );
buf ( n347810 , n347809 );
buf ( n347811 , n347810 );
nand ( n347812 , n347806 , n347811 );
buf ( n347813 , n347812 );
buf ( n347814 , n347813 );
buf ( n347815 , n347382 );
buf ( n347816 , n559 );
and ( n347817 , n347815 , n347816 );
buf ( n347818 , n347817 );
buf ( n347819 , n347818 );
nand ( n347820 , n347814 , n347819 );
buf ( n347821 , n347820 );
buf ( n347822 , n347821 );
buf ( n347823 , n347449 );
buf ( n347824 , n347468 );
and ( n347825 , n347823 , n347824 );
not ( n347826 , n347823 );
buf ( n347827 , n347465 );
and ( n347828 , n347826 , n347827 );
nor ( n347829 , n347825 , n347828 );
buf ( n347830 , n347829 );
buf ( n347831 , n347830 );
not ( n347832 , n347831 );
buf ( n347833 , n347832 );
buf ( n347834 , n347833 );
nand ( n347835 , n347822 , n347834 );
buf ( n347836 , n347835 );
buf ( n347837 , n347836 );
not ( n347838 , n347837 );
xor ( n347839 , n347748 , n347769 );
xor ( n347840 , n347839 , n347772 );
buf ( n347841 , n347840 );
buf ( n347842 , n347841 );
not ( n347843 , n347842 );
or ( n347844 , n347838 , n347843 );
buf ( n347845 , n347833 );
not ( n347846 , n347845 );
buf ( n347847 , n347821 );
not ( n347848 , n347847 );
buf ( n347849 , n347848 );
buf ( n347850 , n347849 );
nand ( n347851 , n347846 , n347850 );
buf ( n347852 , n347851 );
buf ( n347853 , n347852 );
nand ( n347854 , n347844 , n347853 );
buf ( n347855 , n347854 );
buf ( n347856 , n347855 );
xor ( n347857 , n347730 , n347777 );
xor ( n347858 , n347857 , n347782 );
buf ( n347859 , n347858 );
buf ( n347860 , n347859 );
nor ( n347861 , n347856 , n347860 );
buf ( n347862 , n347861 );
buf ( n347863 , n347862 );
not ( n347864 , n347863 );
buf ( n347865 , n347864 );
buf ( n347866 , n347865 );
not ( n347867 , n347866 );
not ( n347868 , n347841 );
buf ( n347869 , n347849 );
not ( n347870 , n347869 );
buf ( n347871 , n347833 );
not ( n347872 , n347871 );
and ( n347873 , n347870 , n347872 );
buf ( n347874 , n347849 );
buf ( n347875 , n347833 );
and ( n347876 , n347874 , n347875 );
nor ( n347877 , n347873 , n347876 );
buf ( n347878 , n347877 );
not ( n347879 , n347878 );
nand ( n347880 , n347868 , n347879 );
not ( n347881 , n347880 );
nand ( n347882 , n347841 , n347878 );
not ( n347883 , n347882 );
or ( n347884 , n347881 , n347883 );
buf ( n347885 , n558 );
buf ( n347886 , n574 );
xor ( n347887 , n347885 , n347886 );
buf ( n347888 , n347887 );
buf ( n347889 , n347888 );
not ( n347890 , n347889 );
buf ( n347891 , n347399 );
not ( n347892 , n347891 );
or ( n347893 , n347890 , n347892 );
buf ( n347894 , n575 );
buf ( n347895 , n347435 );
nand ( n347896 , n347894 , n347895 );
buf ( n347897 , n347896 );
buf ( n347898 , n347897 );
nand ( n347899 , n347893 , n347898 );
buf ( n347900 , n347899 );
buf ( n347901 , n347900 );
buf ( n347902 , n347901 );
buf ( n347903 , n347568 );
buf ( n347904 , n559 );
and ( n347905 , n347903 , n347904 );
buf ( n347906 , n347905 );
buf ( n347907 , n347906 );
buf ( n347908 , n347907 );
buf ( n347909 , n347908 );
buf ( n347910 , n347909 );
or ( n347911 , n347902 , n347910 );
buf ( n347912 , n347911 );
buf ( n347913 , n347912 );
not ( n347914 , n347913 );
buf ( n347915 , n347818 );
buf ( n347916 , n347813 );
xnor ( n347917 , n347915 , n347916 );
buf ( n347918 , n347917 );
buf ( n347919 , n347918 );
not ( n347920 , n347919 );
buf ( n347921 , n347920 );
buf ( n347922 , n347921 );
not ( n347923 , n347922 );
or ( n347924 , n347914 , n347923 );
buf ( n347925 , n347909 );
buf ( n347926 , n347901 );
nand ( n347927 , n347925 , n347926 );
buf ( n347928 , n347927 );
buf ( n347929 , n347928 );
nand ( n347930 , n347924 , n347929 );
buf ( n347931 , n347930 );
nand ( n347932 , n347884 , n347931 );
buf ( n347933 , n347932 );
not ( n347934 , n347933 );
buf ( n347935 , n347934 );
not ( n347936 , n347935 );
xor ( n347937 , n347900 , n347906 );
buf ( n347938 , n347937 );
not ( n347939 , n347938 );
buf ( n347940 , n347939 );
buf ( n347941 , n347940 );
not ( n347942 , n347941 );
buf ( n347943 , n347921 );
not ( n347944 , n347943 );
or ( n347945 , n347942 , n347944 );
buf ( n347946 , n347937 );
buf ( n347947 , n347918 );
nand ( n347948 , n347946 , n347947 );
buf ( n347949 , n347948 );
buf ( n347950 , n347949 );
nand ( n347951 , n347945 , n347950 );
buf ( n347952 , n347951 );
buf ( n347953 , n347952 );
buf ( n347954 , n559 );
buf ( n347955 , n591 );
nand ( n347956 , n347954 , n347955 );
buf ( n347957 , n347956 );
buf ( n347958 , n347957 );
buf ( n347959 , n590 );
and ( n347960 , n347958 , n347959 );
buf ( n347961 , n347960 );
buf ( n347962 , n347961 );
buf ( n347963 , n347962 );
buf ( n347964 , n347963 );
buf ( n347965 , n347964 );
buf ( n347966 , n559 );
buf ( n347967 , n575 );
nand ( n347968 , n347966 , n347967 );
buf ( n347969 , n347968 );
buf ( n347970 , n347969 );
buf ( n347971 , n574 );
and ( n347972 , n347970 , n347971 );
buf ( n347973 , n347972 );
buf ( n347974 , n347973 );
buf ( n347975 , n347974 );
buf ( n347976 , n347975 );
buf ( n347977 , n347976 );
or ( n347978 , n347965 , n347977 );
buf ( n347979 , n347978 );
buf ( n347980 , n347979 );
not ( n347981 , n347980 );
buf ( n347982 , n559 );
not ( n347983 , n347982 );
buf ( n347984 , n347983 );
buf ( n347985 , n347984 );
not ( n347986 , n347985 );
buf ( n347987 , n347478 );
not ( n347988 , n347987 );
or ( n347989 , n347986 , n347988 );
buf ( n347990 , n591 );
buf ( n347991 , n347801 );
nand ( n347992 , n347990 , n347991 );
buf ( n347993 , n347992 );
buf ( n347994 , n347993 );
nand ( n347995 , n347989 , n347994 );
buf ( n347996 , n347995 );
buf ( n347997 , n347996 );
not ( n347998 , n347997 );
or ( n347999 , n347981 , n347998 );
buf ( n348000 , n347976 );
buf ( n348001 , n347964 );
nand ( n348002 , n348000 , n348001 );
buf ( n348003 , n348002 );
buf ( n348004 , n348003 );
nand ( n348005 , n347999 , n348004 );
buf ( n348006 , n348005 );
buf ( n348007 , n348006 );
nand ( n348008 , n347953 , n348007 );
buf ( n348009 , n348008 );
not ( n348010 , n348009 );
buf ( n348011 , n347952 );
not ( n348012 , n348011 );
buf ( n348013 , n348012 );
buf ( n348014 , n348013 );
buf ( n348015 , n348006 );
not ( n348016 , n348015 );
buf ( n348017 , n348016 );
buf ( n348018 , n348017 );
nand ( n348019 , n348014 , n348018 );
buf ( n348020 , n348019 );
buf ( n348021 , n348020 );
buf ( n348022 , n559 );
buf ( n348023 , n575 );
and ( n348024 , n348022 , n348023 );
buf ( n348025 , n348024 );
buf ( n348026 , n348025 );
not ( n348027 , n348026 );
buf ( n348028 , n348027 );
buf ( n348029 , n348028 );
buf ( n348030 , n559 );
buf ( n348031 , n591 );
and ( n348032 , n348030 , n348031 );
buf ( n348033 , n348032 );
buf ( n348034 , n348033 );
not ( n348035 , n348034 );
buf ( n348036 , n348035 );
buf ( n348037 , n348036 );
nor ( n348038 , n348029 , n348037 );
buf ( n348039 , n348038 );
buf ( n348040 , n348039 );
buf ( n348041 , n347984 );
not ( n348042 , n348041 );
buf ( n348043 , n347399 );
not ( n348044 , n348043 );
or ( n348045 , n348042 , n348044 );
buf ( n348046 , n347888 );
buf ( n348047 , n575 );
nand ( n348048 , n348046 , n348047 );
buf ( n348049 , n348048 );
buf ( n348050 , n348049 );
nand ( n348051 , n348045 , n348050 );
buf ( n348052 , n348051 );
buf ( n348053 , n348052 );
xor ( n348054 , n348040 , n348053 );
buf ( n348055 , n347961 );
buf ( n348056 , n347973 );
xnor ( n348057 , n348055 , n348056 );
buf ( n348058 , n348057 );
xnor ( n348059 , n347996 , n348058 );
buf ( n348060 , n348059 );
and ( n348061 , n348054 , n348060 );
and ( n348062 , n348040 , n348053 );
or ( n348063 , n348061 , n348062 );
buf ( n348064 , n348063 );
buf ( n348065 , n348064 );
nand ( n348066 , n348021 , n348065 );
buf ( n348067 , n348066 );
not ( n348068 , n348067 );
or ( n348069 , n348010 , n348068 );
not ( n348070 , n347931 );
nand ( n348071 , n347841 , n348070 , n347879 );
not ( n348072 , n348071 );
and ( n348073 , n347868 , n348070 , n347878 );
nor ( n348074 , n348072 , n348073 );
nand ( n348075 , n348069 , n348074 );
nand ( n348076 , n347936 , n348075 );
buf ( n348077 , n348076 );
not ( n348078 , n348077 );
or ( n348079 , n347867 , n348078 );
buf ( n348080 , n347859 );
buf ( n348081 , n347855 );
nand ( n348082 , n348080 , n348081 );
buf ( n348083 , n348082 );
buf ( n348084 , n348083 );
nand ( n348085 , n348079 , n348084 );
buf ( n348086 , n348085 );
xor ( n348087 , n347800 , n348086 );
xor ( n348088 , n557 , n558 );
not ( n348089 , n348088 );
not ( n348090 , n348089 );
not ( n348091 , n348090 );
not ( n348092 , n556 );
not ( n348093 , n573 );
not ( n348094 , n589 );
or ( n348095 , n348093 , n348094 );
nor ( n348096 , n574 , n590 );
nor ( n348097 , n573 , n589 );
nor ( n348098 , n348096 , n348097 );
nand ( n348099 , n574 , n590 );
nand ( n348100 , n575 , n591 );
nand ( n348101 , n348099 , n348100 );
nand ( n348102 , n348098 , n348101 );
nand ( n348103 , n348095 , n348102 );
nand ( n348104 , n572 , n588 );
not ( n348105 , n348104 );
nor ( n348106 , n572 , n588 );
nor ( n348107 , n348105 , n348106 );
and ( n348108 , n348103 , n348107 );
not ( n348109 , n348103 );
not ( n348110 , n588 );
nand ( n348111 , n347368 , n348110 );
nand ( n348112 , n348111 , n348104 );
and ( n348113 , n348109 , n348112 );
nor ( n348114 , n348108 , n348113 );
not ( n348115 , n348114 );
not ( n348116 , n348115 );
or ( n348117 , n348092 , n348116 );
buf ( n348118 , n348114 );
not ( n348119 , n556 );
nand ( n348120 , n348118 , n348119 );
nand ( n348121 , n348117 , n348120 );
not ( n348122 , n348121 );
or ( n348123 , n348091 , n348122 );
not ( n348124 , n556 );
nand ( n348125 , n575 , n591 );
not ( n348126 , n348125 );
not ( n348127 , n348126 );
not ( n348128 , n574 );
not ( n348129 , n590 );
nand ( n348130 , n348128 , n348129 );
not ( n348131 , n348130 );
or ( n348132 , n348127 , n348131 );
nand ( n348133 , n574 , n590 );
nand ( n348134 , n348132 , n348133 );
and ( n348135 , n573 , n589 );
not ( n348136 , n573 );
not ( n348137 , n589 );
and ( n348138 , n348136 , n348137 );
nor ( n348139 , n348135 , n348138 );
not ( n348140 , n348139 );
and ( n348141 , n348134 , n348140 );
not ( n348142 , n348134 );
and ( n348143 , n348142 , n348139 );
nor ( n348144 , n348141 , n348143 );
not ( n348145 , n348144 );
not ( n348146 , n348145 );
not ( n348147 , n348146 );
or ( n348148 , n348124 , n348147 );
nand ( n348149 , n348119 , n348145 );
nand ( n348150 , n348148 , n348149 );
xor ( n348151 , n556 , n557 );
nand ( n348152 , n348089 , n348151 );
not ( n348153 , n348152 );
nand ( n348154 , n348150 , n348153 );
nand ( n348155 , n348123 , n348154 );
or ( n348156 , n555 , n556 );
xor ( n348157 , n591 , n575 );
buf ( n348158 , n348157 );
nand ( n348159 , n348156 , n348158 );
nand ( n348160 , n555 , n556 );
and ( n348161 , n348159 , n348160 , n554 );
xor ( n348162 , n556 , n555 );
not ( n348163 , n348162 );
not ( n348164 , n554 );
xor ( n348165 , n574 , n590 );
nand ( n348166 , n575 , n591 );
and ( n348167 , n348165 , n348166 );
not ( n348168 , n348165 );
and ( n348169 , n575 , n591 );
and ( n348170 , n348168 , n348169 );
nor ( n348171 , n348167 , n348170 );
not ( n348172 , n348171 );
or ( n348173 , n348164 , n348172 );
not ( n348174 , n348171 );
not ( n348175 , n554 );
nand ( n348176 , n348174 , n348175 );
nand ( n348177 , n348173 , n348176 );
not ( n348178 , n348177 );
or ( n348179 , n348163 , n348178 );
not ( n348180 , n554 );
not ( n348181 , n348158 );
not ( n348182 , n348181 );
or ( n348183 , n348180 , n348182 );
nand ( n348184 , n348158 , n348175 );
nand ( n348185 , n348183 , n348184 );
xor ( n348186 , n554 , n555 );
not ( n348187 , n348186 );
nor ( n348188 , n348187 , n348162 );
nand ( n348189 , n348185 , n348188 );
nand ( n348190 , n348179 , n348189 );
xor ( n348191 , n348161 , n348190 );
xor ( n348192 , n348155 , n348191 );
not ( n348193 , n558 );
not ( n348194 , n573 );
not ( n348195 , n589 );
and ( n348196 , n348194 , n348195 );
nor ( n348197 , n348196 , n348106 );
not ( n348198 , n348197 );
not ( n348199 , n574 );
not ( n348200 , n590 );
or ( n348201 , n348199 , n348200 );
nor ( n348202 , n574 , n590 );
nand ( n348203 , n575 , n591 );
or ( n348204 , n348202 , n348203 );
nand ( n348205 , n348201 , n348204 );
not ( n348206 , n348205 );
or ( n348207 , n348198 , n348206 );
nor ( n348208 , n572 , n588 );
nand ( n348209 , n573 , n589 );
or ( n348210 , n348208 , n348209 );
nand ( n348211 , n572 , n588 );
nand ( n348212 , n348210 , n348211 );
not ( n348213 , n348212 );
nand ( n348214 , n348207 , n348213 );
not ( n348215 , n571 );
not ( n348216 , n587 );
and ( n348217 , n348215 , n348216 );
nand ( n348218 , n587 , n571 );
not ( n348219 , n348218 );
nor ( n348220 , n348217 , n348219 );
and ( n348221 , n348214 , n348220 );
not ( n348222 , n348214 );
not ( n348223 , n348220 );
and ( n348224 , n348222 , n348223 );
nor ( n348225 , n348221 , n348224 );
buf ( n348226 , n348225 );
not ( n348227 , n348226 );
not ( n348228 , n348227 );
or ( n348229 , n348193 , n348228 );
not ( n348230 , n558 );
nand ( n348231 , n348226 , n348230 );
nand ( n348232 , n348229 , n348231 );
nor ( n348233 , n348230 , n559 );
buf ( n348234 , n348233 );
nand ( n348235 , n348232 , n348234 );
not ( n348236 , n558 );
nand ( n348237 , n348236 , n559 );
not ( n348238 , n348237 );
or ( n348239 , n587 , n571 );
not ( n348240 , n348239 );
not ( n348241 , n348197 );
nor ( n348242 , n574 , n590 );
nand ( n348243 , n575 , n591 );
or ( n348244 , n348242 , n348243 );
nand ( n348245 , n348244 , n348133 );
not ( n348246 , n348245 );
or ( n348247 , n348241 , n348246 );
nand ( n348248 , n348247 , n348213 );
not ( n348249 , n348248 );
or ( n348250 , n348240 , n348249 );
nand ( n348251 , n348250 , n348218 );
nand ( n348252 , n570 , n586 );
not ( n348253 , n348252 );
nor ( n348254 , n570 , n586 );
nor ( n348255 , n348253 , n348254 );
and ( n348256 , n348251 , n348255 );
not ( n348257 , n348251 );
not ( n348258 , n570 );
not ( n348259 , n348258 );
not ( n348260 , n586 );
not ( n348261 , n348260 );
or ( n348262 , n348259 , n348261 );
nand ( n348263 , n348262 , n348252 );
and ( n348264 , n348257 , n348263 );
nor ( n348265 , n348256 , n348264 );
buf ( n348266 , n348265 );
nand ( n348267 , n348238 , n348266 );
nand ( n348268 , n558 , n559 );
not ( n348269 , n348268 );
not ( n348270 , n348266 );
nand ( n348271 , n348269 , n348270 );
nand ( n348272 , n348235 , n348267 , n348271 );
xor ( n348273 , n348192 , n348272 );
and ( n348274 , n348158 , n348162 );
not ( n348275 , n348088 );
not ( n348276 , n348150 );
or ( n348277 , n348275 , n348276 );
and ( n348278 , n556 , n348171 );
not ( n348279 , n556 );
nand ( n348280 , n575 , n591 );
and ( n348281 , n348165 , n348280 );
not ( n348282 , n348165 );
and ( n348283 , n348282 , n348169 );
nor ( n348284 , n348281 , n348283 );
not ( n348285 , n348284 );
and ( n348286 , n348279 , n348285 );
or ( n348287 , n348278 , n348286 );
nand ( n348288 , n348287 , n348153 );
nand ( n348289 , n348277 , n348288 );
xor ( n348290 , n348274 , n348289 );
or ( n348291 , n557 , n558 );
xor ( n348292 , n591 , n575 );
nand ( n348293 , n348291 , n348292 );
nand ( n348294 , n557 , n558 );
and ( n348295 , n348293 , n348294 , n556 );
not ( n348296 , n348088 );
not ( n348297 , n348287 );
or ( n348298 , n348296 , n348297 );
and ( n348299 , n556 , n348158 );
not ( n348300 , n556 );
not ( n348301 , n348292 );
and ( n348302 , n348300 , n348301 );
nor ( n348303 , n348299 , n348302 );
and ( n348304 , n348089 , n348151 );
nand ( n348305 , n348303 , n348304 );
nand ( n348306 , n348298 , n348305 );
and ( n348307 , n348295 , n348306 );
and ( n348308 , n348290 , n348307 );
and ( n348309 , n348274 , n348289 );
or ( n348310 , n348308 , n348309 );
not ( n348311 , n348310 );
and ( n348312 , n348273 , n348311 );
not ( n348313 , n348273 );
and ( n348314 , n348313 , n348310 );
nor ( n348315 , n348312 , n348314 );
xor ( n348316 , n348274 , n348289 );
xor ( n348317 , n348316 , n348307 );
not ( n348318 , n559 );
not ( n348319 , n348232 );
or ( n348320 , n348318 , n348319 );
and ( n348321 , n558 , n348118 );
not ( n348322 , n558 );
and ( n348323 , n348322 , n348115 );
nor ( n348324 , n348321 , n348323 );
nand ( n348325 , n348324 , n348233 );
nand ( n348326 , n348320 , n348325 );
nor ( n348327 , n348317 , n348326 );
not ( n348328 , n559 );
not ( n348329 , n348324 );
or ( n348330 , n348328 , n348329 );
not ( n348331 , n348144 );
not ( n348332 , n348331 );
nand ( n348333 , n348332 , n558 );
not ( n348334 , n348333 );
not ( n348335 , n558 );
nand ( n348336 , n348335 , n348145 );
not ( n348337 , n348336 );
or ( n348338 , n348334 , n348337 );
nand ( n348339 , n348338 , n348234 );
nand ( n348340 , n348330 , n348339 );
xor ( n348341 , n348295 , n348306 );
xor ( n348342 , n348340 , n348341 );
not ( n348343 , n559 );
nand ( n348344 , n348333 , n348336 );
not ( n348345 , n348344 );
or ( n348346 , n348343 , n348345 );
not ( n348347 , n558 );
not ( n348348 , n348284 );
not ( n348349 , n348348 );
not ( n348350 , n348349 );
or ( n348351 , n348347 , n348350 );
not ( n348352 , n558 );
nand ( n348353 , n348352 , n348174 );
nand ( n348354 , n348351 , n348353 );
nand ( n348355 , n348354 , n348234 );
nand ( n348356 , n348346 , n348355 );
not ( n348357 , n348356 );
and ( n348358 , n348158 , n348088 );
not ( n348359 , n348358 );
or ( n348360 , n348357 , n348359 );
nor ( n348361 , n348356 , n348358 );
not ( n348362 , n559 );
not ( n348363 , n348354 );
or ( n348364 , n348362 , n348363 );
nand ( n348365 , n348181 , n348234 );
nand ( n348366 , n348364 , n348365 );
not ( n348367 , n559 );
not ( n348368 , n348158 );
or ( n348369 , n348367 , n348368 );
nand ( n348370 , n348369 , n558 );
not ( n348371 , n348370 );
nand ( n348372 , n348366 , n348371 );
or ( n348373 , n348361 , n348372 );
nand ( n348374 , n348360 , n348373 );
and ( n348375 , n348342 , n348374 );
and ( n348376 , n348340 , n348341 );
or ( n348377 , n348375 , n348376 );
not ( n348378 , n348377 );
or ( n348379 , n348327 , n348378 );
nand ( n348380 , n348317 , n348326 );
nand ( n348381 , n348379 , n348380 );
buf ( n348382 , n348381 );
not ( n348383 , n348382 );
and ( n348384 , n348315 , n348383 );
not ( n348385 , n348315 );
and ( n348386 , n348385 , n348382 );
nor ( n348387 , n348384 , n348386 );
nand ( n348388 , n348087 , n348387 );
buf ( n348389 , n348074 );
buf ( n348390 , n347932 );
nand ( n348391 , n348389 , n348390 );
buf ( n348392 , n348391 );
buf ( n348393 , n348392 );
buf ( n348394 , n348067 );
buf ( n348395 , n348009 );
nand ( n348396 , n348394 , n348395 );
buf ( n348397 , n348396 );
buf ( n348398 , n348397 );
not ( n348399 , n348398 );
buf ( n348400 , n348399 );
buf ( n348401 , n348400 );
and ( n348402 , n348393 , n348401 );
not ( n348403 , n348393 );
buf ( n348404 , n348397 );
and ( n348405 , n348403 , n348404 );
nor ( n348406 , n348402 , n348405 );
buf ( n348407 , n348406 );
xor ( n348408 , n348340 , n348341 );
xor ( n348409 , n348408 , n348374 );
not ( n348410 , n348409 );
nand ( n348411 , n348410 , n348407 );
buf ( n348412 , n348076 );
not ( n348413 , n348412 );
buf ( n348414 , n348413 );
buf ( n348415 , n348414 );
buf ( n348416 , n347859 );
buf ( n348417 , n347855 );
nor ( n348418 , n348416 , n348417 );
buf ( n348419 , n348418 );
buf ( n348420 , n348419 );
not ( n348421 , n348420 );
buf ( n348422 , n348421 );
buf ( n348423 , n348422 );
buf ( n348424 , n348083 );
nand ( n348425 , n348423 , n348424 );
buf ( n348426 , n348425 );
buf ( n348427 , n348426 );
and ( n348428 , n348415 , n348427 );
not ( n348429 , n348415 );
buf ( n348430 , n348426 );
not ( n348431 , n348430 );
buf ( n348432 , n348431 );
buf ( n348433 , n348432 );
and ( n348434 , n348429 , n348433 );
nor ( n348435 , n348428 , n348434 );
buf ( n348436 , n348435 );
not ( n348437 , n348436 );
not ( n348438 , n348327 );
nand ( n348439 , n348438 , n348380 );
and ( n348440 , n348439 , n348378 );
not ( n348441 , n348439 );
and ( n348442 , n348441 , n348377 );
nor ( n348443 , n348440 , n348442 );
nand ( n348444 , n348437 , n348443 );
and ( n348445 , n348388 , C1 , n348444 );
not ( n348446 , n348443 );
nand ( n348447 , n348446 , n348436 );
not ( n348448 , n348447 );
not ( n348449 , n348448 );
not ( n348450 , n348388 );
or ( n348451 , n348449 , n348450 );
not ( n348452 , n348087 );
not ( n348453 , n348387 );
nand ( n348454 , n348452 , n348453 );
nand ( n348455 , n348451 , n348454 );
nor ( n348456 , n348445 , n348455 );
not ( n348457 , n348456 );
xor ( n348458 , n347592 , n347638 );
and ( n348459 , n348458 , n347719 );
and ( n348460 , n347592 , n347638 );
or ( n348461 , n348459 , n348460 );
buf ( n348462 , n348461 );
buf ( n348463 , n347355 );
not ( n348464 , n348463 );
buf ( n348465 , n347341 );
not ( n348466 , n348465 );
buf ( n348467 , n348466 );
buf ( n348468 , n348467 );
not ( n348469 , n348468 );
or ( n348470 , n348464 , n348469 );
buf ( n348471 , n347336 );
not ( n348472 , n348471 );
buf ( n348473 , n348472 );
buf ( n348474 , n348473 );
buf ( n348475 , n348474 );
buf ( n348476 , n348475 );
buf ( n348477 , n348476 );
buf ( n348478 , n557 );
buf ( n348479 , n570 );
xor ( n348480 , n348478 , n348479 );
buf ( n348481 , n348480 );
buf ( n348482 , n348481 );
nand ( n348483 , n348477 , n348482 );
buf ( n348484 , n348483 );
buf ( n348485 , n348484 );
nand ( n348486 , n348470 , n348485 );
buf ( n348487 , n348486 );
buf ( n348488 , n348487 );
buf ( n348489 , n347415 );
buf ( n348490 , n347423 );
and ( n348491 , n348489 , n348490 );
buf ( n348492 , n348491 );
buf ( n348493 , n348492 );
xor ( n348494 , n348488 , n348493 );
xor ( n348495 , n569 , n570 );
buf ( n348496 , n348495 );
buf ( n348497 , n559 );
and ( n348498 , n348496 , n348497 );
buf ( n348499 , n348498 );
not ( n348500 , n347399 );
not ( n348501 , n347410 );
or ( n348502 , n348500 , n348501 );
buf ( n348503 , n553 );
buf ( n348504 , n574 );
xor ( n348505 , n348503 , n348504 );
buf ( n348506 , n348505 );
buf ( n348507 , n348506 );
buf ( n348508 , n575 );
nand ( n348509 , n348507 , n348508 );
buf ( n348510 , n348509 );
nand ( n348511 , n348502 , n348510 );
xor ( n348512 , n348499 , n348511 );
buf ( n348513 , n347387 );
not ( n348514 , n348513 );
buf ( n348515 , n347378 );
not ( n348516 , n348515 );
or ( n348517 , n348514 , n348516 );
buf ( n348518 , n347382 );
buf ( n348519 , n555 );
buf ( n348520 , n572 );
xor ( n348521 , n348519 , n348520 );
buf ( n348522 , n348521 );
buf ( n348523 , n348522 );
nand ( n348524 , n348518 , n348523 );
buf ( n348525 , n348524 );
buf ( n348526 , n348525 );
nand ( n348527 , n348517 , n348526 );
buf ( n348528 , n348527 );
xor ( n348529 , n348512 , n348528 );
buf ( n348530 , n348529 );
xor ( n348531 , n348494 , n348530 );
buf ( n348532 , n348531 );
not ( n348533 , n348532 );
and ( n348534 , n348462 , n348533 );
not ( n348535 , n348462 );
and ( n348536 , n348535 , n348532 );
nor ( n348537 , n348534 , n348536 );
buf ( n348538 , n347393 );
not ( n348539 , n348538 );
buf ( n348540 , n347427 );
not ( n348541 , n348540 );
or ( n348542 , n348539 , n348541 );
buf ( n348543 , n347393 );
buf ( n348544 , n347427 );
or ( n348545 , n348543 , n348544 );
buf ( n348546 , n347361 );
nand ( n348547 , n348545 , n348546 );
buf ( n348548 , n348547 );
buf ( n348549 , n348548 );
nand ( n348550 , n348542 , n348549 );
buf ( n348551 , n348550 );
xor ( n348552 , n347656 , n347686 );
and ( n348553 , n348552 , n347716 );
and ( n348554 , n347656 , n347686 );
or ( n348555 , n348553 , n348554 );
buf ( n348556 , n348555 );
not ( n348557 , n348556 );
xor ( n348558 , n348551 , n348557 );
buf ( n348559 , n347679 );
not ( n348560 , n348559 );
buf ( n348561 , n347671 );
not ( n348562 , n348561 );
or ( n348563 , n348560 , n348562 );
buf ( n348564 , n347530 );
buf ( n348565 , n557 );
buf ( n348566 , n586 );
xor ( n348567 , n348565 , n348566 );
buf ( n348568 , n348567 );
buf ( n348569 , n348568 );
nand ( n348570 , n348564 , n348569 );
buf ( n348571 , n348570 );
buf ( n348572 , n348571 );
nand ( n348573 , n348563 , n348572 );
buf ( n348574 , n348573 );
buf ( n348575 , n348574 );
not ( n348576 , n348575 );
buf ( n348577 , n348576 );
buf ( n348578 , n347706 );
buf ( n348579 , n347710 );
and ( n348580 , n348578 , n348579 );
buf ( n348581 , n348580 );
not ( n348582 , n348581 );
xor ( n835 , n348577 , n348582 );
buf ( n348584 , n835 );
not ( n837 , n348584 );
buf ( n348586 , n837 );
not ( n839 , n348586 );
buf ( n348588 , n347699 );
not ( n841 , n348588 );
buf ( n348590 , n347478 );
not ( n843 , n348590 );
or ( n348592 , n841 , n843 );
and ( n845 , n553 , n590 );
not ( n348594 , n553 );
buf ( n348595 , n590 );
not ( n848 , n348595 );
buf ( n348597 , n848 );
and ( n850 , n348594 , n348597 );
nor ( n851 , n845 , n850 );
nand ( n852 , n851 , n591 );
buf ( n348601 , n852 );
nand ( n854 , n348592 , n348601 );
buf ( n348603 , n854 );
buf ( n348604 , n348603 );
not ( n857 , n348604 );
buf ( n348606 , n347984 );
not ( n859 , n348606 );
buf ( n348608 , n585 );
buf ( n348609 , n586 );
xor ( n348610 , n348608 , n348609 );
buf ( n348611 , n348610 );
buf ( n348612 , n348611 );
not ( n865 , n348612 );
buf ( n348614 , n865 );
buf ( n348615 , n348614 );
not ( n868 , n348615 );
buf ( n348617 , n868 );
buf ( n348618 , n348617 );
nand ( n871 , n859 , n348618 );
buf ( n348620 , n871 );
buf ( n348621 , n348620 );
not ( n874 , n348621 );
and ( n875 , n857 , n874 );
buf ( n348624 , n348614 );
buf ( n348625 , n348624 );
buf ( n348626 , n348625 );
buf ( n348627 , n348626 );
not ( n880 , n348627 );
buf ( n348629 , n880 );
buf ( n348630 , n348629 );
buf ( n348631 , n559 );
nand ( n348632 , n348630 , n348631 );
buf ( n348633 , n348632 );
buf ( n348634 , n348633 );
buf ( n348635 , n348603 );
and ( n888 , n348634 , n348635 );
nor ( n889 , n875 , n888 );
buf ( n348638 , n889 );
buf ( n348639 , n348638 );
buf ( n348640 , n347649 );
not ( n893 , n348640 );
buf ( n348642 , n347554 );
not ( n895 , n348642 );
or ( n348644 , n893 , n895 );
buf ( n348645 , n347568 );
buf ( n348646 , n555 );
buf ( n348647 , n588 );
xor ( n348648 , n348646 , n348647 );
buf ( n348649 , n348648 );
buf ( n348650 , n348649 );
nand ( n903 , n348645 , n348650 );
buf ( n348652 , n903 );
buf ( n348653 , n348652 );
nand ( n906 , n348644 , n348653 );
buf ( n348655 , n906 );
buf ( n348656 , n348655 );
xor ( n909 , n348639 , n348656 );
buf ( n348658 , n909 );
buf ( n348659 , n348658 );
not ( n912 , n348659 );
buf ( n348661 , n912 );
not ( n914 , n348661 );
or ( n915 , n839 , n914 );
buf ( n348664 , n348658 );
buf ( n348665 , n835 );
nand ( n918 , n348664 , n348665 );
buf ( n348667 , n918 );
nand ( n920 , n915 , n348667 );
xnor ( n921 , n348558 , n920 );
not ( n922 , n921 );
and ( n923 , n348537 , n922 );
not ( n924 , n348537 );
and ( n925 , n924 , n921 );
nor ( n926 , n923 , n925 );
buf ( n348675 , n926 );
xor ( n928 , n347429 , n347586 );
and ( n929 , n928 , n347722 );
and ( n930 , n347429 , n347586 );
or ( n931 , n929 , n930 );
buf ( n348680 , n931 );
buf ( n348681 , n348680 );
nand ( n934 , n348675 , n348681 );
buf ( n348683 , n934 );
buf ( n348684 , n348683 );
buf ( n937 , n348684 );
buf ( n348686 , n937 );
not ( n939 , n926 );
buf ( n348688 , n348680 );
not ( n941 , n348688 );
buf ( n348690 , n941 );
nand ( n943 , n939 , n348690 );
nand ( n944 , n348686 , n943 );
not ( n945 , n944 );
buf ( n348694 , n347724 );
buf ( n348695 , n347786 );
nor ( n948 , n348694 , n348695 );
buf ( n348697 , n948 );
or ( n950 , n348697 , n348083 );
nand ( n951 , n950 , n347797 );
not ( n952 , n951 );
buf ( n348701 , n348419 );
not ( n954 , n348701 );
buf ( n348703 , n347792 );
buf ( n348704 , n348076 );
nand ( n957 , n954 , n348703 , n348704 );
buf ( n348706 , n957 );
nand ( n959 , n952 , n348706 );
not ( n960 , n959 );
or ( n961 , n945 , n960 );
nand ( n962 , n952 , n348706 , n348686 , n943 );
nand ( n963 , n961 , n962 );
not ( n964 , n348090 );
not ( n965 , n556 );
not ( n966 , n348226 );
not ( n967 , n966 );
or ( n968 , n965 , n967 );
nand ( n969 , n348226 , n348119 );
nand ( n970 , n968 , n969 );
not ( n971 , n970 );
or ( n972 , n964 , n971 );
nand ( n973 , n348121 , n348153 );
nand ( n974 , n972 , n973 );
not ( n975 , n558 );
or ( n976 , n571 , n587 );
or ( n977 , n570 , n586 );
nand ( n978 , n976 , n977 );
not ( n979 , n978 );
not ( n980 , n979 );
not ( n981 , n348248 );
or ( n982 , n980 , n981 );
nand ( n348731 , n571 , n587 );
or ( n984 , n348254 , n348731 );
nand ( n985 , n984 , n348252 );
not ( n986 , n985 );
nand ( n987 , n982 , n986 );
nor ( n988 , n569 , n585 );
not ( n989 , n988 );
nand ( n990 , n569 , n585 );
nand ( n991 , n989 , n990 );
not ( n992 , n991 );
and ( n993 , n987 , n992 );
not ( n994 , n987 );
and ( n995 , n994 , n991 );
nor ( n348744 , n993 , n995 );
buf ( n997 , n348744 );
not ( n348746 , n997 );
not ( n999 , n348746 );
or ( n1000 , n975 , n999 );
not ( n1001 , n558 );
nand ( n1002 , n1001 , n997 );
nand ( n1003 , n1000 , n1002 );
not ( n1004 , n1003 );
not ( n1005 , n559 );
or ( n1006 , n1004 , n1005 );
not ( n1007 , n348266 );
nand ( n1008 , n1007 , n348234 );
nand ( n348757 , n1006 , n1008 );
xor ( n1010 , n974 , n348757 );
xor ( n1011 , n553 , n554 );
and ( n1012 , n348158 , n1011 );
not ( n1013 , n348162 );
not ( n1014 , n348145 );
not ( n1015 , n348175 );
or ( n1016 , n1014 , n1015 );
nand ( n1017 , n348332 , n554 );
nand ( n1018 , n1016 , n1017 );
not ( n1019 , n1018 );
or ( n1020 , n1013 , n1019 );
xnor ( n1021 , n555 , n556 );
and ( n1022 , n1021 , n348186 );
nand ( n1023 , n348177 , n1022 );
nand ( n348772 , n1020 , n1023 );
xor ( n1025 , n1012 , n348772 );
and ( n1026 , n348161 , n348190 );
xor ( n1027 , n1025 , n1026 );
xor ( n1028 , n1010 , n1027 );
not ( n1029 , n1028 );
not ( n1030 , n1029 );
xor ( n1031 , n348155 , n348191 );
and ( n1032 , n1031 , n348272 );
and ( n1033 , n348155 , n348191 );
or ( n1034 , n1032 , n1033 );
and ( n1035 , n1030 , n1034 );
not ( n1036 , n1030 );
not ( n1037 , n1034 );
and ( n1038 , n1036 , n1037 );
nor ( n1039 , n1035 , n1038 );
not ( n1040 , n348381 );
not ( n1041 , n348273 );
nand ( n1042 , n1041 , n348311 );
not ( n1043 , n1042 );
or ( n1044 , n1040 , n1043 );
nand ( n1045 , n348273 , n348310 );
nand ( n1046 , n1044 , n1045 );
buf ( n1047 , n1046 );
xor ( n1048 , n1039 , n1047 );
not ( n1049 , n1048 );
nor ( n1050 , n963 , n1049 );
not ( n1051 , n1050 );
not ( n1052 , n1048 );
nand ( n1053 , n1052 , n963 );
nand ( n1054 , n1051 , n1053 );
not ( n1055 , n1054 );
not ( n1056 , n1055 );
or ( n1057 , n348457 , n1056 );
not ( n1058 , n348456 );
nand ( n1059 , n1058 , n1054 );
nand ( n1060 , n1057 , n1059 );
nand ( n1061 , n1060 , n585 );
not ( n1062 , n1060 );
not ( n1063 , n585 );
nand ( n1064 , n1062 , n1063 );
nand ( n1065 , n1061 , n1064 );
nand ( n1086 , C1 , n348411 );
not ( n1091 , n1086 );
and ( n1092 , n1091 , C1 );
nor ( n1093 , C0 , n1092 );
not ( n1094 , n1093 );
not ( n1095 , n588 );
nand ( n1096 , n1094 , n1095 );
nand ( n1110 , n348454 , n348388 );
not ( n1111 , n1110 );
not ( n1112 , n1111 );
not ( n1114 , n348444 );
or ( n1115 , C0 , n1114 );
nand ( n1116 , n1115 , n348447 );
not ( n1117 , n1116 );
not ( n1118 , n1117 );
or ( n1119 , n1112 , n1118 );
nand ( n1120 , n1116 , n1110 );
nand ( n1121 , n1119 , n1120 );
not ( n1122 , n1121 );
nand ( n1123 , n1122 , n348260 );
nand ( n1124 , n348444 , n348447 );
not ( n348835 , n1124 );
and ( n1128 , n348835 , C1 );
nor ( n1129 , C0 , n1128 );
not ( n1130 , n1129 );
nand ( n1131 , n1130 , n348216 );
nor ( n1133 , n1121 , n586 );
buf ( n1134 , n1129 );
nand ( n1135 , n1134 , n587 );
or ( n1136 , n1133 , n1135 );
nand ( n1137 , n1121 , n586 );
nand ( n1138 , n1136 , n1137 );
not ( n1139 , n1138 );
nand ( n1140 , C1 , n1139 );
not ( n1141 , n1140 );
and ( n1142 , n1065 , n1141 );
not ( n1143 , n1065 );
and ( n1144 , n1143 , n1140 );
nor ( n1145 , n1142 , n1144 );
buf ( n348853 , n1145 );
buf ( n1147 , n348853 );
buf ( n348855 , n1147 );
buf ( n348856 , n348855 );
not ( n1150 , n348856 );
buf ( n348858 , n1150 );
buf ( n348859 , n348858 );
not ( n1153 , n348859 );
or ( n1154 , n347323 , n1153 );
buf ( n348862 , n348855 );
buf ( n348863 , n596 );
not ( n1157 , n348863 );
buf ( n348865 , n1157 );
buf ( n348866 , n348865 );
nand ( n1160 , n348862 , n348866 );
buf ( n348868 , n1160 );
buf ( n348869 , n348868 );
nand ( n1163 , n1154 , n348869 );
buf ( n348871 , n1163 );
buf ( n348872 , n348871 );
not ( n1166 , n348872 );
or ( n1167 , n347321 , n1166 );
nand ( n1171 , C1 , n1135 );
not ( n1172 , n1171 );
not ( n1173 , n1172 );
nand ( n1174 , n1123 , n1137 );
not ( n1175 , n1174 );
not ( n1176 , n1175 );
or ( n1177 , n1173 , n1176 );
nand ( n348882 , n1174 , n1171 );
nand ( n1179 , n1177 , n348882 );
buf ( n348884 , n1179 );
and ( n1181 , n348884 , n348865 );
not ( n1182 , n348884 );
and ( n1183 , n1182 , n596 );
or ( n1184 , n1181 , n1183 );
buf ( n348889 , n1184 );
buf ( n348890 , n348865 );
buf ( n348891 , n347316 );
and ( n1188 , n348890 , n348891 );
buf ( n348893 , n596 );
buf ( n348894 , n597 );
and ( n1191 , n348893 , n348894 );
buf ( n348896 , n347318 );
nor ( n1193 , n1188 , n1191 , n348896 );
buf ( n348898 , n1193 );
buf ( n348899 , n348898 );
nand ( n1196 , n348889 , n348899 );
buf ( n348901 , n1196 );
buf ( n348902 , n348901 );
nand ( n1199 , n1167 , n348902 );
buf ( n348904 , n1199 );
buf ( n348905 , n348904 );
xnor ( n1202 , C0 , n591 );
buf ( n348907 , n1202 );
buf ( n348908 , n592 );
not ( n1205 , n348908 );
buf ( n348910 , n1205 );
buf ( n348911 , n348910 );
nor ( n1208 , n348907 , n348911 );
buf ( n348913 , n1208 );
buf ( n348914 , n348913 );
buf ( n348915 , n592 );
not ( n1212 , n348915 );
xor ( n1213 , n590 , C0 );
xnor ( n1214 , n1213 , C0 );
not ( n1215 , n1214 );
buf ( n348920 , n1215 );
buf ( n1217 , n348920 );
buf ( n348922 , n1217 );
buf ( n348923 , n348922 );
not ( n1220 , n348923 );
buf ( n348925 , n1220 );
buf ( n348926 , n348925 );
not ( n348927 , n348926 );
or ( n1224 , n1212 , n348927 );
buf ( n348929 , n1215 );
not ( n1226 , n348929 );
buf ( n348931 , n1226 );
buf ( n348932 , n348931 );
not ( n1229 , n348932 );
buf ( n348934 , n1229 );
buf ( n348935 , n348934 );
buf ( n348936 , n348910 );
nand ( n1233 , n348935 , n348936 );
buf ( n348938 , n1233 );
buf ( n348939 , n348938 );
nand ( n1236 , n1224 , n348939 );
buf ( n348941 , n1236 );
buf ( n348942 , n348941 );
buf ( n348943 , n593 );
buf ( n348944 , n594 );
xor ( n348945 , n348943 , n348944 );
buf ( n348946 , n348945 );
buf ( n348947 , n348946 );
and ( n1244 , n348942 , n348947 );
buf ( n348949 , n593 );
not ( n1246 , n348949 );
buf ( n348951 , n1246 );
and ( n1248 , n348910 , n348951 );
and ( n1249 , n592 , n593 );
nor ( n1250 , n1248 , n1249 , n348946 );
buf ( n348955 , n1250 );
not ( n1252 , n348955 );
buf ( n348957 , n1202 );
buf ( n348958 , n592 );
and ( n1255 , n348957 , n348958 );
not ( n1256 , n1202 );
buf ( n348961 , n1256 );
buf ( n348962 , n348910 );
and ( n1259 , n348961 , n348962 );
nor ( n1260 , n1255 , n1259 );
buf ( n348965 , n1260 );
buf ( n348966 , n348965 );
nor ( n1263 , n1252 , n348966 );
buf ( n348968 , n1263 );
buf ( n348969 , n348968 );
nor ( n1266 , n1244 , n348969 );
buf ( n348971 , n1266 );
buf ( n348972 , n348971 );
buf ( n348973 , n594 );
not ( n1270 , n348973 );
buf ( n348975 , n1270 );
buf ( n348976 , n348975 );
buf ( n348977 , n348951 );
or ( n1274 , n348976 , n348977 );
buf ( n348979 , n593 );
buf ( n348980 , n594 );
or ( n1277 , n348979 , n348980 );
buf ( n348982 , n1256 );
nand ( n1279 , n1277 , n348982 );
buf ( n348984 , n1279 );
buf ( n348985 , n348984 );
buf ( n348986 , n592 );
nand ( n1283 , n1274 , n348985 , n348986 );
buf ( n348988 , n1283 );
buf ( n348989 , n348988 );
nor ( n1286 , n348972 , n348989 );
buf ( n348991 , n1286 );
buf ( n348992 , n348991 );
xor ( n348993 , n348914 , n348992 );
buf ( n348994 , n348910 );
not ( n1291 , n348994 );
buf ( n1292 , C0 );
and ( n1296 , C1 , n589 );
nor ( n1297 , C0 , n1296 );
or ( n1300 , n1292 , n1297 );
nand ( n1301 , C1 , n1300 );
buf ( n349001 , n1301 );
not ( n1303 , n349001 );
and ( n1304 , n1291 , n1303 );
buf ( n1305 , n1301 );
buf ( n349005 , n1305 );
buf ( n349006 , n348910 );
and ( n1308 , n349005 , n349006 );
nor ( n1309 , n1304 , n1308 );
buf ( n349009 , n1309 );
buf ( n349010 , n349009 );
buf ( n349011 , n348946 );
not ( n1313 , n349011 );
buf ( n349013 , n1313 );
buf ( n349014 , n349013 );
or ( n1316 , n349010 , n349014 );
buf ( n349016 , n348941 );
buf ( n349017 , n1250 );
nand ( n1319 , n349016 , n349017 );
buf ( n349019 , n1319 );
buf ( n349020 , n349019 );
nand ( n1322 , n1316 , n349020 );
buf ( n349022 , n1322 );
buf ( n349023 , n349022 );
xor ( n1325 , n348993 , n349023 );
buf ( n349025 , n1325 );
buf ( n349026 , n349025 );
not ( n1328 , n596 );
buf ( n349028 , n595 );
not ( n1330 , n349028 );
buf ( n349030 , n1330 );
not ( n1332 , n349030 );
and ( n1333 , n1328 , n1332 );
nor ( n1334 , n348865 , n595 );
nor ( n1335 , n1333 , n1334 );
not ( n349035 , n1335 );
buf ( n349036 , n349035 );
not ( n1338 , n349036 );
nand ( n1340 , n1129 , n587 );
nand ( n1341 , n1131 , n1340 );
not ( n1342 , n1341 );
not ( n1343 , n1342 );
or ( n1344 , C0 , n1343 );
nand ( n1349 , n1344 , C1 );
buf ( n349044 , n1349 );
buf ( n349045 , n349044 );
buf ( n349046 , n349045 );
buf ( n349047 , n349046 );
not ( n1354 , n349047 );
buf ( n349049 , n1354 );
buf ( n349050 , n349049 );
buf ( n1357 , n349050 );
buf ( n349052 , n1357 );
and ( n1359 , n349052 , n594 );
not ( n1360 , n349052 );
and ( n1361 , n1360 , n348975 );
or ( n1362 , n1359 , n1361 );
buf ( n349057 , n1362 );
not ( n1364 , n349057 );
or ( n1365 , n1338 , n1364 );
buf ( n349060 , n594 );
not ( n1367 , n349060 );
nand ( n1368 , n1096 , C1 );
and ( n1372 , n1368 , C1 );
nor ( n1375 , n1372 , C0 );
buf ( n349065 , n1375 );
buf ( n1377 , n349065 );
buf ( n349067 , n1377 );
buf ( n349068 , n349067 );
not ( n1380 , n349068 );
buf ( n349070 , n1380 );
buf ( n349071 , n349070 );
not ( n1383 , n349071 );
or ( n1384 , n1367 , n1383 );
buf ( n349074 , n349067 );
buf ( n349075 , n348975 );
nand ( n1387 , n349074 , n349075 );
buf ( n349077 , n1387 );
buf ( n349078 , n349077 );
nand ( n1390 , n1384 , n349078 );
buf ( n349080 , n1390 );
buf ( n349081 , n349080 );
and ( n1393 , n349030 , n348975 );
and ( n1394 , n595 , n594 );
nor ( n1395 , n1393 , n1394 );
nand ( n1396 , n1335 , n1395 );
not ( n1397 , n1396 );
buf ( n349087 , n1397 );
nand ( n1399 , n349081 , n349087 );
buf ( n349089 , n1399 );
buf ( n349090 , n349089 );
nand ( n1402 , n1365 , n349090 );
buf ( n349092 , n1402 );
buf ( n349093 , n349092 );
xor ( n1405 , n349026 , n349093 );
xor ( n1406 , n348988 , n348971 );
buf ( n349096 , n1406 );
buf ( n349097 , n349035 );
not ( n1409 , n349097 );
buf ( n349099 , n349080 );
not ( n1411 , n349099 );
or ( n349101 , n1409 , n1411 );
buf ( n349102 , n594 );
not ( n1414 , n349102 );
buf ( n349104 , n1301 );
not ( n1416 , n349104 );
buf ( n349106 , n1416 );
buf ( n349107 , n349106 );
not ( n1419 , n349107 );
or ( n1420 , n1414 , n1419 );
buf ( n349110 , n1305 );
buf ( n349111 , n348975 );
nand ( n1423 , n349110 , n349111 );
buf ( n349113 , n1423 );
buf ( n349114 , n349113 );
nand ( n1426 , n1420 , n349114 );
buf ( n349116 , n1426 );
buf ( n349117 , n349116 );
buf ( n349118 , n1397 );
nand ( n1430 , n349117 , n349118 );
buf ( n349120 , n1430 );
buf ( n349121 , n349120 );
nand ( n1433 , n349101 , n349121 );
buf ( n349123 , n1433 );
buf ( n349124 , n349123 );
xor ( n1436 , n349096 , n349124 );
buf ( n349126 , n1202 );
buf ( n349127 , n349013 );
nor ( n1439 , n349126 , n349127 );
buf ( n349129 , n1439 );
buf ( n349130 , n349129 );
buf ( n349131 , n349035 );
not ( n1443 , n349131 );
buf ( n349133 , n594 );
not ( n1445 , n349133 );
buf ( n349135 , n348931 );
not ( n1447 , n349135 );
or ( n1448 , n1445 , n1447 );
buf ( n349138 , n348922 );
buf ( n349139 , n348975 );
nand ( n1451 , n349138 , n349139 );
buf ( n349141 , n1451 );
buf ( n349142 , n349141 );
nand ( n1454 , n1448 , n349142 );
buf ( n349144 , n1454 );
buf ( n349145 , n349144 );
not ( n1457 , n349145 );
or ( n1458 , n1443 , n1457 );
buf ( n349148 , n1256 );
buf ( n349149 , n1397 );
buf ( n349150 , n594 );
not ( n1462 , n349150 );
and ( n1463 , n349149 , n1462 );
buf ( n349153 , n1463 );
buf ( n349154 , n349153 );
and ( n1466 , n349148 , n349154 );
buf ( n349156 , n1202 );
buf ( n349157 , n1397 );
buf ( n349158 , n594 );
nand ( n1470 , n349157 , n349158 );
buf ( n349160 , n1470 );
buf ( n349161 , n349160 );
not ( n1473 , n349161 );
buf ( n349163 , n1473 );
buf ( n349164 , n349163 );
and ( n1476 , n349156 , n349164 );
nor ( n1477 , n1466 , n1476 );
buf ( n349167 , n1477 );
buf ( n349168 , n349167 );
nand ( n1480 , n1458 , n349168 );
buf ( n349170 , n1480 );
buf ( n349171 , n349170 );
not ( n1483 , n349171 );
buf ( n349173 , n348865 );
buf ( n349174 , n349030 );
or ( n1486 , n349173 , n349174 );
buf ( n349176 , n595 );
buf ( n349177 , n596 );
or ( n1489 , n349176 , n349177 );
buf ( n349179 , n1256 );
nand ( n1491 , n1489 , n349179 );
buf ( n349181 , n1491 );
buf ( n349182 , n349181 );
buf ( n349183 , n594 );
nand ( n1495 , n1486 , n349182 , n349183 );
buf ( n349185 , n1495 );
buf ( n349186 , n349185 );
nor ( n1498 , n1483 , n349186 );
buf ( n349188 , n1498 );
buf ( n349189 , n349188 );
xor ( n1501 , n349130 , n349189 );
buf ( n349191 , n349035 );
not ( n1503 , n349191 );
buf ( n349193 , n349116 );
not ( n1505 , n349193 );
or ( n1506 , n1503 , n1505 );
buf ( n349196 , n349144 );
buf ( n349197 , n1397 );
nand ( n1509 , n349196 , n349197 );
buf ( n349199 , n1509 );
buf ( n349200 , n349199 );
nand ( n1512 , n1506 , n349200 );
buf ( n349202 , n1512 );
buf ( n349203 , n349202 );
and ( n1515 , n1501 , n349203 );
or ( n1517 , n1515 , C0 );
buf ( n349206 , n1517 );
buf ( n349207 , n349206 );
and ( n1520 , n1436 , n349207 );
and ( n1521 , n349096 , n349124 );
or ( n1522 , n1520 , n1521 );
buf ( n349211 , n1522 );
buf ( n349212 , n349211 );
xor ( n1525 , n1405 , n349212 );
buf ( n349214 , n1525 );
buf ( n349215 , n349214 );
xor ( n1528 , n348905 , n349215 );
buf ( n349217 , n347319 );
not ( n1530 , n349217 );
buf ( n349219 , n1184 );
not ( n1532 , n349219 );
or ( n1533 , n1530 , n1532 );
buf ( n349222 , n596 );
not ( n1535 , n349222 );
buf ( n349224 , n349052 );
not ( n1537 , n349224 );
or ( n1538 , n1535 , n1537 );
buf ( n349227 , n1349 );
not ( n1540 , n349227 );
buf ( n349229 , n1540 );
buf ( n349230 , n349229 );
buf ( n1543 , n349230 );
buf ( n349232 , n1543 );
buf ( n349233 , n349232 );
not ( n1546 , n349233 );
buf ( n349235 , n348865 );
nand ( n1548 , n1546 , n349235 );
buf ( n349237 , n1548 );
buf ( n349238 , n349237 );
nand ( n1551 , n1538 , n349238 );
buf ( n349240 , n1551 );
buf ( n349241 , n349240 );
buf ( n349242 , n348898 );
nand ( n1555 , n349241 , n349242 );
buf ( n349244 , n1555 );
buf ( n349245 , n349244 );
nand ( n1558 , n1533 , n349245 );
buf ( n349247 , n1558 );
buf ( n349248 , n349247 );
xor ( n1561 , n349096 , n349124 );
xor ( n1562 , n1561 , n349207 );
buf ( n349251 , n1562 );
buf ( n349252 , n349251 );
xor ( n1565 , n349248 , n349252 );
xor ( n1566 , n349130 , n349189 );
xor ( n1567 , n1566 , n349203 );
buf ( n349256 , n1567 );
buf ( n349257 , n349256 );
buf ( n349258 , n347319 );
not ( n349259 , n349258 );
buf ( n349260 , n349240 );
not ( n1573 , n349260 );
or ( n1574 , n349259 , n1573 );
buf ( n349263 , n596 );
not ( n1576 , n349263 );
buf ( n349265 , n349070 );
not ( n1578 , n349265 );
or ( n1579 , n1576 , n1578 );
buf ( n349268 , n349067 );
buf ( n349269 , n348865 );
nand ( n1582 , n349268 , n349269 );
buf ( n349271 , n1582 );
buf ( n349272 , n349271 );
nand ( n1585 , n1579 , n349272 );
buf ( n349274 , n1585 );
buf ( n349275 , n349274 );
buf ( n349276 , n348898 );
nand ( n1589 , n349275 , n349276 );
buf ( n349278 , n1589 );
buf ( n349279 , n349278 );
nand ( n1592 , n1574 , n349279 );
buf ( n349281 , n1592 );
buf ( n349282 , n349281 );
xor ( n1595 , n349257 , n349282 );
buf ( n349284 , n349185 );
not ( n1597 , n349284 );
buf ( n349286 , n349170 );
not ( n1599 , n349286 );
or ( n1600 , n1597 , n1599 );
buf ( n349289 , n349170 );
buf ( n349290 , n349185 );
or ( n1603 , n349289 , n349290 );
nand ( n1604 , n1600 , n1603 );
buf ( n349293 , n1604 );
buf ( n349294 , n349293 );
buf ( n349295 , n347319 );
not ( n1608 , n349295 );
buf ( n349297 , n349274 );
not ( n1610 , n349297 );
or ( n1611 , n1608 , n1610 );
buf ( n349300 , n596 );
not ( n1613 , n349300 );
buf ( n349302 , n349106 );
not ( n1615 , n349302 );
or ( n1616 , n1613 , n1615 );
buf ( n349305 , n1305 );
buf ( n349306 , n348865 );
nand ( n1619 , n349305 , n349306 );
buf ( n349308 , n1619 );
buf ( n349309 , n349308 );
nand ( n1622 , n1616 , n349309 );
buf ( n349311 , n1622 );
buf ( n349312 , n349311 );
buf ( n349313 , n348898 );
nand ( n1626 , n349312 , n349313 );
buf ( n349315 , n1626 );
buf ( n349316 , n349315 );
nand ( n1629 , n1611 , n349316 );
buf ( n349318 , n1629 );
buf ( n349319 , n349318 );
xor ( n1632 , n349294 , n349319 );
buf ( n349321 , n1335 );
buf ( n349322 , n1202 );
nor ( n1635 , n349321 , n349322 );
buf ( n349324 , n1635 );
buf ( n349325 , n349324 );
not ( n1638 , n347318 );
not ( n1639 , n596 );
not ( n1640 , n348925 );
or ( n1641 , n1639 , n1640 );
buf ( n349330 , n348934 );
buf ( n349331 , n348865 );
nand ( n1644 , n349330 , n349331 );
buf ( n349333 , n1644 );
nand ( n1646 , n1641 , n349333 );
not ( n1647 , n1646 );
or ( n1648 , n1638 , n1647 );
and ( n1649 , n348898 , n596 );
and ( n1650 , n1649 , n1202 );
and ( n1651 , n348898 , n348865 );
and ( n1652 , n1651 , n1256 );
nor ( n1653 , n1650 , n1652 );
nand ( n1654 , n1648 , n1653 );
buf ( n349343 , n1654 );
not ( n1656 , n349343 );
buf ( n349345 , n597 );
buf ( n349346 , n598 );
or ( n1659 , n349345 , n349346 );
buf ( n349348 , n1256 );
nand ( n1661 , n1659 , n349348 );
buf ( n349350 , n1661 );
buf ( n349351 , n349350 );
buf ( n349352 , n597 );
buf ( n349353 , n598 );
nand ( n1666 , n349352 , n349353 );
buf ( n349355 , n1666 );
buf ( n349356 , n349355 );
buf ( n349357 , n596 );
nand ( n1670 , n349351 , n349356 , n349357 );
buf ( n349359 , n1670 );
buf ( n349360 , n349359 );
nor ( n349361 , n1656 , n349360 );
buf ( n349362 , n349361 );
buf ( n349363 , n349362 );
xor ( n1676 , n349325 , n349363 );
buf ( n349365 , n347319 );
not ( n1678 , n349365 );
buf ( n349367 , n349311 );
not ( n1680 , n349367 );
or ( n1681 , n1678 , n1680 );
buf ( n349370 , n1646 );
buf ( n349371 , n348898 );
nand ( n1684 , n349370 , n349371 );
buf ( n349373 , n1684 );
buf ( n349374 , n349373 );
nand ( n1687 , n1681 , n349374 );
buf ( n349376 , n1687 );
buf ( n349377 , n349376 );
and ( n1690 , n1676 , n349377 );
or ( n1692 , n1690 , C0 );
buf ( n349380 , n1692 );
buf ( n349381 , n349380 );
and ( n1695 , n1632 , n349381 );
and ( n1696 , n349294 , n349319 );
or ( n1697 , n1695 , n1696 );
buf ( n349385 , n1697 );
buf ( n349386 , n349385 );
and ( n1700 , n1595 , n349386 );
and ( n349388 , n349257 , n349282 );
or ( n1702 , n1700 , n349388 );
buf ( n349390 , n1702 );
buf ( n349391 , n349390 );
and ( n1705 , n1565 , n349391 );
and ( n1706 , n349248 , n349252 );
or ( n1707 , n1705 , n1706 );
buf ( n349395 , n1707 );
buf ( n349396 , n349395 );
and ( n1710 , n1528 , n349396 );
and ( n1711 , n348905 , n349215 );
or ( n1712 , n1710 , n1711 );
buf ( n349400 , n1712 );
buf ( n349401 , n349400 );
and ( n1715 , n601 , n602 );
not ( n1716 , n601 );
buf ( n349404 , n602 );
not ( n1718 , n349404 );
buf ( n349406 , n1718 );
and ( n1720 , n1716 , n349406 );
nor ( n1721 , n1715 , n1720 );
buf ( n1722 , n1721 );
buf ( n349410 , n1722 );
not ( n1724 , n349410 );
buf ( n349412 , n600 );
not ( n1726 , n349412 );
or ( n1727 , n553 , n554 );
nand ( n1728 , n1727 , n348292 );
nand ( n1729 , n553 , n554 );
and ( n1730 , n1728 , n1729 , n552 );
not ( n1731 , n1011 );
not ( n1732 , n552 );
not ( n1733 , n348349 );
or ( n1734 , n1732 , n1733 );
not ( n1735 , n552 );
nand ( n1736 , n1735 , n348285 );
nand ( n1737 , n1734 , n1736 );
not ( n1738 , n1737 );
or ( n1739 , n1731 , n1738 );
and ( n1740 , n552 , n348181 );
not ( n1741 , n552 );
and ( n1742 , n1741 , n348158 );
or ( n1743 , n1740 , n1742 );
xnor ( n1744 , n552 , n553 );
nor ( n1745 , n1011 , n1744 );
nand ( n1746 , n1743 , n1745 );
nand ( n1747 , n1739 , n1746 );
and ( n1748 , n1730 , n1747 );
not ( n1749 , n348153 );
not ( n1750 , n556 );
not ( n1751 , n348266 );
not ( n1752 , n1751 );
or ( n1753 , n1750 , n1752 );
nand ( n1754 , n348266 , n348119 );
nand ( n1755 , n1753 , n1754 );
not ( n1756 , n1755 );
or ( n1757 , n1749 , n1756 );
not ( n1758 , n348088 );
nor ( n1759 , n1758 , n348119 );
nand ( n1760 , n1759 , n348746 );
not ( n1761 , n1760 );
not ( n1762 , n348088 );
nor ( n1763 , n1762 , n556 );
and ( n1764 , n997 , n1763 );
nor ( n1765 , n1761 , n1764 );
nand ( n349453 , n1757 , n1765 );
xor ( n1767 , n1748 , n349453 );
not ( n1768 , n348233 );
and ( n1769 , n568 , n584 );
not ( n1770 , n568 );
not ( n1771 , n584 );
and ( n1772 , n1770 , n1771 );
nor ( n1773 , n1769 , n1772 );
or ( n1774 , n571 , n587 );
or ( n1775 , n570 , n586 );
nand ( n1776 , n1774 , n1775 );
nor ( n1777 , n1776 , n988 );
not ( n1778 , n1777 );
not ( n1779 , n348214 );
or ( n1780 , n1778 , n1779 );
not ( n349468 , n569 );
nand ( n1782 , n349468 , n1063 );
and ( n1783 , n985 , n1782 );
not ( n1784 , n990 );
nor ( n1785 , n1783 , n1784 );
nand ( n1786 , n1780 , n1785 );
xor ( n1787 , n1773 , n1786 );
buf ( n1788 , n1787 );
not ( n1789 , n1788 );
and ( n1790 , n558 , n1789 );
not ( n1791 , n558 );
and ( n1792 , n1791 , n1788 );
or ( n1793 , n1790 , n1792 );
not ( n1794 , n1793 );
or ( n1795 , n1768 , n1794 );
not ( n1796 , n558 );
nand ( n1797 , n567 , n583 );
not ( n1798 , n1797 );
nor ( n1799 , n567 , n583 );
nor ( n1800 , n1798 , n1799 );
not ( n1801 , n585 );
not ( n1802 , n569 );
nand ( n1803 , n1801 , n1802 );
not ( n1804 , n568 );
nand ( n1805 , n1771 , n1804 );
nand ( n1806 , n348111 , n1803 , n1805 );
nor ( n1807 , n1806 , n978 );
not ( n1808 , n1807 );
not ( n1809 , n348101 );
not ( n1810 , n348098 );
or ( n1811 , n1809 , n1810 );
nand ( n1812 , n573 , n589 );
nand ( n1813 , n572 , n588 );
and ( n1814 , n1812 , n1813 );
nand ( n1815 , n1811 , n1814 );
not ( n1816 , n1815 );
or ( n1817 , n1808 , n1816 );
nand ( n1818 , n568 , n584 );
not ( n1819 , n1818 );
not ( n1820 , n584 );
not ( n1821 , n1820 );
not ( n1822 , n568 );
not ( n1823 , n1822 );
or ( n1824 , n1821 , n1823 );
nand ( n1825 , n1824 , n1782 );
not ( n1826 , n1825 );
or ( n1827 , n1819 , n1826 );
nand ( n1828 , n570 , n586 );
nand ( n1829 , n568 , n584 );
nand ( n1830 , n569 , n585 );
nand ( n1831 , n1828 , n1829 , n1830 );
not ( n349519 , n1831 );
not ( n1833 , n348260 );
not ( n1834 , n348258 );
or ( n1835 , n1833 , n1834 );
and ( n1836 , n571 , n587 );
nand ( n1837 , n1835 , n1836 );
nand ( n349525 , n349519 , n1837 );
nand ( n1839 , n1827 , n349525 );
nand ( n349527 , n1817 , n1839 );
buf ( n1841 , n349527 );
xor ( n1842 , n1800 , n1841 );
buf ( n1843 , n1842 );
not ( n1844 , n1843 );
not ( n1845 , n1844 );
or ( n1846 , n1796 , n1845 );
nand ( n1847 , n1843 , n348230 );
nand ( n1848 , n1846 , n1847 );
nand ( n1849 , n1848 , n559 );
nand ( n1850 , n1795 , n1849 );
and ( n1851 , n1767 , n1850 );
and ( n1852 , n1748 , n349453 );
or ( n1853 , n1851 , n1852 );
not ( n1854 , n1011 );
not ( n1855 , n552 );
not ( n1856 , n348118 );
not ( n1857 , n1856 );
or ( n1858 , n1855 , n1857 );
not ( n1859 , n552 );
nand ( n1860 , n1859 , n348118 );
nand ( n1861 , n1858 , n1860 );
not ( n1862 , n1861 );
or ( n1863 , n1854 , n1862 );
not ( n1864 , n552 );
not ( n1865 , n348146 );
or ( n1866 , n1864 , n1865 );
not ( n1867 , n552 );
nand ( n1868 , n1867 , n348145 );
nand ( n1869 , n1866 , n1868 );
nor ( n1870 , n1744 , n1011 );
buf ( n1871 , n1870 );
nand ( n1872 , n1869 , n1871 );
nand ( n1873 , n1863 , n1872 );
xor ( n1874 , n551 , n552 );
buf ( n1875 , n1874 );
not ( n1876 , n1875 );
not ( n1877 , n550 );
not ( n1878 , n348171 );
or ( n1879 , n1877 , n1878 );
not ( n1880 , n550 );
nand ( n1881 , n348174 , n1880 );
nand ( n1882 , n1879 , n1881 );
not ( n1883 , n1882 );
or ( n1884 , n1876 , n1883 );
not ( n1885 , n550 );
not ( n1886 , n348181 );
or ( n1887 , n1885 , n1886 );
nand ( n1888 , n348158 , n1880 );
nand ( n1889 , n1887 , n1888 );
xnor ( n1890 , n550 , n551 );
nor ( n1891 , n1874 , n1890 );
nand ( n1892 , n1889 , n1891 );
nand ( n1893 , n1884 , n1892 );
or ( n1894 , n551 , n552 );
not ( n1895 , n1894 );
not ( n1896 , n348158 );
or ( n1897 , n1895 , n1896 );
nand ( n1898 , n551 , n552 );
and ( n1899 , n1898 , n550 );
nand ( n1900 , n1897 , n1899 );
and ( n1901 , n1893 , n1900 );
not ( n1902 , n1893 );
not ( n1903 , n1900 );
and ( n1904 , n1902 , n1903 );
or ( n1905 , n1901 , n1904 );
xor ( n1906 , n1873 , n1905 );
not ( n1907 , n348090 );
not ( n1908 , n556 );
not ( n1909 , n1789 );
or ( n1910 , n1908 , n1909 );
not ( n1911 , n1789 );
nand ( n1912 , n1911 , n348119 );
nand ( n1913 , n1910 , n1912 );
not ( n349601 , n1913 );
or ( n1915 , n1907 , n349601 );
and ( n1916 , n348304 , n556 );
and ( n1917 , n348746 , n1916 );
not ( n1918 , n348746 );
and ( n1919 , n348153 , n348119 );
and ( n349607 , n1918 , n1919 );
nor ( n1921 , n1917 , n349607 );
nand ( n349609 , n1915 , n1921 );
xor ( n1923 , n1906 , n349609 );
xor ( n1924 , n1853 , n1923 );
buf ( n1925 , n348162 );
not ( n1926 , n1925 );
not ( n1927 , n554 );
not ( n1928 , n1751 );
or ( n1929 , n1927 , n1928 );
nand ( n1930 , n348266 , n348175 );
nand ( n1931 , n1929 , n1930 );
not ( n1932 , n1931 );
or ( n1933 , n1926 , n1932 );
not ( n1934 , n554 );
not ( n1935 , n348227 );
or ( n1936 , n1934 , n1935 );
nand ( n1937 , n348226 , n348175 );
nand ( n1938 , n1936 , n1937 );
nand ( n1939 , n1938 , n1022 );
nand ( n1940 , n1933 , n1939 );
and ( n1941 , n348158 , n1874 );
not ( n1942 , n1011 );
not ( n1943 , n1869 );
or ( n1944 , n1942 , n1943 );
nand ( n1945 , n1737 , n1870 );
nand ( n1946 , n1944 , n1945 );
xor ( n1947 , n1941 , n1946 );
not ( n1948 , n348162 );
not ( n1949 , n1938 );
or ( n1950 , n1948 , n1949 );
and ( n1951 , n348115 , n554 );
not ( n1952 , n348115 );
and ( n1953 , n1952 , n348175 );
or ( n1954 , n1951 , n1953 );
nand ( n1955 , n1954 , n1022 );
nand ( n1956 , n1950 , n1955 );
and ( n1957 , n1947 , n1956 );
and ( n1958 , n1941 , n1946 );
or ( n1959 , n1957 , n1958 );
xor ( n1960 , n1940 , n1959 );
not ( n1961 , n559 );
not ( n1962 , n558 );
not ( n1963 , n1799 );
not ( n1964 , n1963 );
not ( n1965 , n349527 );
or ( n1966 , n1964 , n1965 );
nand ( n1967 , n1966 , n1797 );
xnor ( n1968 , n566 , n582 );
not ( n1969 , n1968 );
and ( n1970 , n1967 , n1969 );
not ( n1971 , n1967 );
and ( n1972 , n1971 , n1968 );
nor ( n1973 , n1970 , n1972 );
buf ( n1974 , n1973 );
not ( n1975 , n1974 );
not ( n1976 , n1975 );
or ( n1977 , n1962 , n1976 );
not ( n1978 , n558 );
nand ( n1979 , n1978 , n1974 );
nand ( n1980 , n1977 , n1979 );
not ( n1981 , n1980 );
or ( n1982 , n1961 , n1981 );
nand ( n1983 , n1848 , n348233 );
nand ( n1984 , n1982 , n1983 );
xor ( n1985 , n1960 , n1984 );
and ( n1986 , n1924 , n1985 );
and ( n1987 , n1853 , n1923 );
or ( n1988 , n1986 , n1987 );
and ( n1989 , n1893 , n1903 );
not ( n1990 , n348153 );
not ( n1991 , n1913 );
or ( n1992 , n1990 , n1991 );
and ( n1993 , n1843 , n348119 );
not ( n1994 , n1843 );
and ( n1995 , n1994 , n556 );
or ( n1996 , n1993 , n1995 );
nand ( n1997 , n1996 , n348088 );
nand ( n1998 , n1992 , n1997 );
xor ( n1999 , n1989 , n1998 );
not ( n2000 , n1925 );
not ( n2001 , n554 );
not ( n2002 , n997 );
not ( n2003 , n2002 );
or ( n2004 , n2001 , n2003 );
not ( n2005 , n2002 );
nand ( n2006 , n2005 , n348175 );
nand ( n2007 , n2004 , n2006 );
not ( n2008 , n2007 );
or ( n2009 , n2000 , n2008 );
nand ( n2010 , n1931 , n1022 );
nand ( n2011 , n2009 , n2010 );
xor ( n2012 , n1999 , n2011 );
xor ( n2013 , n1940 , n1959 );
and ( n349701 , n2013 , n1984 );
and ( n2015 , n1940 , n1959 );
or ( n2016 , n349701 , n2015 );
xor ( n2017 , n2012 , n2016 );
not ( n2018 , n348158 );
xor ( n2019 , n549 , n550 );
not ( n2020 , n2019 );
nor ( n2021 , n2018 , n2020 );
not ( n2022 , n1875 );
not ( n2023 , n550 );
not ( n2024 , n348146 );
or ( n2025 , n2023 , n2024 );
nand ( n2026 , n348145 , n1880 );
nand ( n2027 , n2025 , n2026 );
not ( n2028 , n2027 );
or ( n2029 , n2022 , n2028 );
nand ( n2030 , n1882 , n1891 );
nand ( n2031 , n2029 , n2030 );
xor ( n2032 , n2021 , n2031 );
not ( n2033 , n1011 );
not ( n2034 , n552 );
not ( n2035 , n348227 );
or ( n2036 , n2034 , n2035 );
not ( n2037 , n552 );
nand ( n2038 , n2037 , n348226 );
nand ( n2039 , n2036 , n2038 );
not ( n2040 , n2039 );
or ( n2041 , n2033 , n2040 );
nand ( n2042 , n1861 , n1871 );
nand ( n2043 , n2041 , n2042 );
xor ( n2044 , n2032 , n2043 );
not ( n2045 , n559 );
not ( n2046 , n566 );
not ( n2047 , n582 );
and ( n2048 , n2046 , n2047 );
nor ( n2049 , n2048 , n1799 );
not ( n2050 , n2049 );
not ( n2051 , n349527 );
or ( n2052 , n2050 , n2051 );
not ( n2053 , n566 );
not ( n2054 , n582 );
or ( n2055 , n2053 , n2054 );
nor ( n2056 , n566 , n582 );
nand ( n2057 , n567 , n583 );
or ( n2058 , n2056 , n2057 );
nand ( n2059 , n2055 , n2058 );
buf ( n2060 , n2059 );
not ( n2061 , n2060 );
nand ( n2062 , n2052 , n2061 );
or ( n2063 , n565 , n581 );
nand ( n2064 , n565 , n581 );
nand ( n2065 , n2063 , n2064 );
not ( n2066 , n2065 );
and ( n349754 , n2062 , n2066 );
not ( n2068 , n2062 );
and ( n2069 , n2068 , n2065 );
nor ( n2070 , n349754 , n2069 );
buf ( n2071 , n2070 );
not ( n2072 , n2071 );
and ( n2073 , n2072 , n558 );
not ( n2074 , n2072 );
and ( n2075 , n2074 , n348230 );
or ( n2076 , n2073 , n2075 );
not ( n2077 , n2076 );
or ( n2078 , n2045 , n2077 );
nand ( n2079 , n1980 , n348233 );
nand ( n2080 , n2078 , n2079 );
xor ( n2081 , n2044 , n2080 );
xor ( n2082 , n1873 , n1905 );
and ( n2083 , n2082 , n349609 );
and ( n2084 , n1873 , n1905 );
or ( n2085 , n2083 , n2084 );
xor ( n2086 , n2081 , n2085 );
xor ( n2087 , n2017 , n2086 );
buf ( n2088 , n2087 );
not ( n2089 , n2088 );
xor ( n2090 , n1988 , n2089 );
xor ( n2091 , n1941 , n1946 );
xor ( n2092 , n2091 , n1956 );
not ( n2093 , n348162 );
not ( n2094 , n1954 );
or ( n2095 , n2093 , n2094 );
nand ( n2096 , n1018 , n1022 );
nand ( n2097 , n2095 , n2096 );
xor ( n2098 , n1730 , n1747 );
xor ( n2099 , n2097 , n2098 );
not ( n2100 , n348090 );
not ( n2101 , n1755 );
or ( n2102 , n2100 , n2101 );
nand ( n2103 , n970 , n348153 );
nand ( n2104 , n2102 , n2103 );
and ( n2105 , n2099 , n2104 );
and ( n2106 , n2097 , n2098 );
or ( n2107 , n2105 , n2106 );
xor ( n2108 , n2092 , n2107 );
xor ( n2109 , n1748 , n349453 );
xor ( n2110 , n2109 , n1850 );
and ( n2111 , n2108 , n2110 );
and ( n2112 , n2092 , n2107 );
or ( n2113 , n2111 , n2112 );
not ( n2114 , n2113 );
xor ( n2115 , n1853 , n1923 );
xor ( n2116 , n2115 , n1985 );
not ( n2117 , n2116 );
or ( n2118 , n2114 , n2117 );
xor ( n2119 , n2092 , n2107 );
xor ( n2120 , n2119 , n2110 );
not ( n2121 , n559 );
not ( n2122 , n1793 );
or ( n2123 , n2121 , n2122 );
nand ( n2124 , n1003 , n348233 );
nand ( n2125 , n2123 , n2124 );
xor ( n2126 , n1012 , n348772 );
and ( n2127 , n2126 , n1026 );
and ( n2128 , n1012 , n348772 );
or ( n2129 , n2127 , n2128 );
xor ( n2130 , n2125 , n2129 );
xor ( n2131 , n2097 , n2098 );
xor ( n2132 , n2131 , n2104 );
and ( n2133 , n2130 , n2132 );
and ( n2134 , n2125 , n2129 );
or ( n2135 , n2133 , n2134 );
nand ( n2136 , n2120 , n2135 );
nand ( n2137 , n2118 , n2136 );
not ( n2138 , n2137 );
not ( n2139 , n2116 );
not ( n2140 , n2113 );
nand ( n2141 , n2139 , n2140 );
not ( n2142 , n2141 );
or ( n2143 , n2138 , n2142 );
not ( n2144 , n2116 );
nand ( n2145 , n2144 , n2140 );
xor ( n2146 , n2125 , n2129 );
xor ( n2147 , n2146 , n2132 );
not ( n2148 , n2147 );
xor ( n2149 , n974 , n348757 );
and ( n2150 , n2149 , n1027 );
and ( n2151 , n974 , n348757 );
or ( n2152 , n2150 , n2151 );
not ( n2153 , n2152 );
nand ( n2154 , n2148 , n2153 );
not ( n2155 , n2154 );
not ( n2156 , n1030 );
not ( n349844 , n1034 );
or ( n2158 , n2156 , n349844 );
not ( n2159 , n1029 );
not ( n2160 , n1037 );
or ( n2161 , n2159 , n2160 );
nand ( n2162 , n2161 , n1046 );
nand ( n2163 , n2158 , n2162 );
not ( n2164 , n2163 );
or ( n2165 , n2155 , n2164 );
buf ( n2166 , n2147 );
nand ( n2167 , n2166 , n2152 );
nand ( n2168 , n2165 , n2167 );
not ( n2169 , n2120 );
not ( n2170 , n2135 );
nand ( n2171 , n2169 , n2170 );
nand ( n2172 , n2145 , n2168 , n2171 );
nand ( n2173 , n2143 , n2172 );
buf ( n2174 , n2173 );
xnor ( n2175 , n2090 , n2174 );
not ( n2176 , n2175 );
xor ( n2177 , n348499 , n348511 );
and ( n2178 , n2177 , n348528 );
and ( n2179 , n348499 , n348511 );
or ( n2180 , n2178 , n2179 );
buf ( n349868 , n348506 );
not ( n2182 , n349868 );
buf ( n349870 , n347604 );
not ( n2184 , n349870 );
or ( n349872 , n2182 , n2184 );
buf ( n349873 , n552 );
buf ( n349874 , n574 );
xor ( n2188 , n349873 , n349874 );
buf ( n349876 , n2188 );
buf ( n349877 , n349876 );
buf ( n349878 , n575 );
nand ( n2192 , n349877 , n349878 );
buf ( n349880 , n2192 );
buf ( n349881 , n349880 );
nand ( n2195 , n349872 , n349881 );
buf ( n349883 , n2195 );
buf ( n349884 , n349883 );
buf ( n349885 , n559 );
buf ( n349886 , n569 );
or ( n2200 , n349885 , n349886 );
buf ( n349888 , n570 );
nand ( n2202 , n2200 , n349888 );
buf ( n349890 , n2202 );
buf ( n349891 , n349890 );
buf ( n349892 , n559 );
buf ( n349893 , n569 );
nand ( n2207 , n349892 , n349893 );
buf ( n349895 , n2207 );
buf ( n349896 , n349895 );
buf ( n349897 , n568 );
nand ( n2211 , n349891 , n349896 , n349897 );
buf ( n349899 , n2211 );
buf ( n349900 , n349899 );
and ( n2214 , n349884 , n349900 );
not ( n2215 , n349884 );
buf ( n349903 , n349899 );
not ( n2217 , n349903 );
buf ( n349905 , n2217 );
buf ( n349906 , n349905 );
and ( n2220 , n2215 , n349906 );
nor ( n2221 , n2214 , n2220 );
buf ( n349909 , n2221 );
xor ( n2223 , n2180 , n349909 );
buf ( n349911 , n559 );
buf ( n349912 , n568 );
xor ( n2226 , n349911 , n349912 );
buf ( n349914 , n2226 );
buf ( n349915 , n349914 );
not ( n2229 , n349915 );
not ( n2230 , n348495 );
not ( n2231 , n568 );
nand ( n2232 , n2231 , n569 );
not ( n2233 , n569 );
nand ( n2234 , n2233 , n568 );
nand ( n2235 , n2232 , n2234 );
and ( n2236 , n2230 , n2235 );
buf ( n349924 , n2236 );
not ( n2238 , n349924 );
or ( n2239 , n2229 , n2238 );
and ( n2240 , n569 , n570 );
not ( n2241 , n569 );
and ( n2242 , n2241 , n348258 );
nor ( n2243 , n2240 , n2242 );
buf ( n349931 , n2243 );
buf ( n2245 , n349931 );
buf ( n349933 , n2245 );
buf ( n349934 , n349933 );
buf ( n349935 , n558 );
buf ( n349936 , n568 );
xor ( n2250 , n349935 , n349936 );
buf ( n349938 , n2250 );
buf ( n349939 , n349938 );
nand ( n2253 , n349934 , n349939 );
buf ( n349941 , n2253 );
buf ( n349942 , n349941 );
nand ( n2256 , n2239 , n349942 );
buf ( n349944 , n2256 );
buf ( n349945 , n349944 );
not ( n2259 , n349945 );
buf ( n349947 , n348522 );
not ( n2261 , n349947 );
buf ( n349949 , n347378 );
not ( n2263 , n349949 );
or ( n2264 , n2261 , n2263 );
buf ( n349952 , n347382 );
buf ( n349953 , n554 );
buf ( n349954 , n572 );
xor ( n2268 , n349953 , n349954 );
buf ( n349956 , n2268 );
buf ( n349957 , n349956 );
nand ( n2271 , n349952 , n349957 );
buf ( n349959 , n2271 );
buf ( n349960 , n349959 );
nand ( n2274 , n2264 , n349960 );
buf ( n349962 , n2274 );
buf ( n349963 , n349962 );
not ( n2277 , n349963 );
buf ( n349965 , n2277 );
buf ( n349966 , n349965 );
not ( n2280 , n349966 );
or ( n2281 , n2259 , n2280 );
buf ( n349969 , n349962 );
buf ( n349970 , n349944 );
not ( n2284 , n349970 );
buf ( n349972 , n2284 );
buf ( n349973 , n349972 );
nand ( n2287 , n349969 , n349973 );
buf ( n349975 , n2287 );
buf ( n349976 , n349975 );
nand ( n2290 , n2281 , n349976 );
buf ( n349978 , n2290 );
buf ( n349979 , n349978 );
buf ( n349980 , n348481 );
not ( n2294 , n349980 );
buf ( n349982 , n347344 );
not ( n2296 , n349982 );
or ( n2297 , n2294 , n2296 );
buf ( n349985 , n347350 );
buf ( n349986 , n556 );
buf ( n349987 , n570 );
xor ( n2301 , n349986 , n349987 );
buf ( n349989 , n2301 );
buf ( n349990 , n349989 );
nand ( n2304 , n349985 , n349990 );
buf ( n349992 , n2304 );
buf ( n349993 , n349992 );
nand ( n2307 , n2297 , n349993 );
buf ( n349995 , n2307 );
buf ( n349996 , n349995 );
and ( n2310 , n349979 , n349996 );
not ( n2311 , n349979 );
buf ( n349999 , n349995 );
not ( n2313 , n349999 );
buf ( n350001 , n2313 );
buf ( n350002 , n350001 );
and ( n2316 , n2311 , n350002 );
nor ( n2317 , n2310 , n2316 );
buf ( n350005 , n2317 );
and ( n2319 , n2223 , n350005 );
not ( n2320 , n2223 );
not ( n2321 , n350005 );
and ( n2322 , n2320 , n2321 );
or ( n2323 , n2319 , n2322 );
buf ( n350011 , n2323 );
buf ( n2325 , n348551 );
not ( n2326 , n2325 );
not ( n2327 , n348556 );
or ( n2328 , n2326 , n2327 );
not ( n2329 , n2325 );
not ( n2330 , n2329 );
not ( n2331 , n348557 );
or ( n350019 , n2330 , n2331 );
nand ( n2333 , n350019 , n920 );
nand ( n2334 , n2328 , n2333 );
buf ( n350022 , n2334 );
xor ( n2336 , n350011 , n350022 );
xor ( n2337 , n348488 , n348493 );
and ( n2338 , n2337 , n348530 );
and ( n2339 , n348488 , n348493 );
or ( n2340 , n2338 , n2339 );
buf ( n350028 , n2340 );
buf ( n350029 , n350028 );
not ( n2343 , n348581 );
and ( n2344 , n348577 , n2343 );
not ( n350032 , n2344 );
buf ( n350033 , n350032 );
not ( n2347 , n350033 );
buf ( n350035 , n348661 );
not ( n2349 , n350035 );
or ( n2350 , n2347 , n2349 );
buf ( n350038 , n348581 );
buf ( n350039 , n348574 );
nand ( n2353 , n350038 , n350039 );
buf ( n350041 , n2353 );
buf ( n350042 , n350041 );
nand ( n2356 , n2350 , n350042 );
buf ( n350044 , n2356 );
buf ( n350045 , n350044 );
xor ( n2359 , n350029 , n350045 );
buf ( n350047 , n559 );
buf ( n350048 , n585 );
or ( n2362 , n350047 , n350048 );
buf ( n350050 , n586 );
nand ( n2364 , n2362 , n350050 );
buf ( n350052 , n2364 );
buf ( n350053 , n350052 );
buf ( n350054 , n559 );
buf ( n350055 , n585 );
nand ( n2369 , n350054 , n350055 );
buf ( n350057 , n2369 );
buf ( n350058 , n350057 );
buf ( n350059 , n584 );
nand ( n2373 , n350053 , n350058 , n350059 );
buf ( n350061 , n2373 );
buf ( n350062 , n350061 );
not ( n2376 , n350062 );
buf ( n350064 , n851 );
not ( n2378 , n350064 );
buf ( n350066 , n347478 );
not ( n2380 , n350066 );
or ( n2381 , n2378 , n2380 );
buf ( n350069 , n552 );
buf ( n350070 , n590 );
xor ( n2384 , n350069 , n350070 );
buf ( n350072 , n2384 );
buf ( n350073 , n350072 );
buf ( n350074 , n591 );
nand ( n2388 , n350073 , n350074 );
buf ( n350076 , n2388 );
buf ( n350077 , n350076 );
nand ( n2391 , n2381 , n350077 );
buf ( n350079 , n2391 );
buf ( n350080 , n350079 );
not ( n2394 , n350080 );
or ( n2395 , n2376 , n2394 );
buf ( n350083 , n350079 );
buf ( n350084 , n350061 );
or ( n2398 , n350083 , n350084 );
nand ( n2399 , n2395 , n2398 );
buf ( n350087 , n2399 );
buf ( n350088 , n350087 );
buf ( n350089 , n348603 );
not ( n2403 , n350089 );
buf ( n350091 , n2403 );
nand ( n2405 , n350091 , n348633 );
not ( n2406 , n2405 );
not ( n2407 , n348655 );
or ( n2408 , n2406 , n2407 );
not ( n2409 , n348633 );
nand ( n2410 , n2409 , n348603 );
nand ( n2411 , n2408 , n2410 );
buf ( n350099 , n2411 );
xor ( n2413 , n350088 , n350099 );
buf ( n350101 , n348568 );
not ( n2415 , n350101 );
buf ( n350103 , n586 );
buf ( n350104 , n587 );
xnor ( n2418 , n350103 , n350104 );
buf ( n350106 , n2418 );
buf ( n350107 , n350106 );
buf ( n350108 , n347663 );
nor ( n2422 , n350107 , n350108 );
buf ( n350110 , n2422 );
buf ( n350111 , n350110 );
not ( n2425 , n350111 );
or ( n2426 , n2415 , n2425 );
buf ( n350114 , n347530 );
buf ( n350115 , n556 );
buf ( n350116 , n586 );
xor ( n2430 , n350115 , n350116 );
buf ( n350118 , n2430 );
buf ( n350119 , n350118 );
nand ( n2433 , n350114 , n350119 );
buf ( n350121 , n2433 );
buf ( n350122 , n350121 );
nand ( n2436 , n2426 , n350122 );
buf ( n350124 , n2436 );
buf ( n350125 , n350124 );
buf ( n350126 , n348649 );
not ( n2440 , n350126 );
buf ( n350128 , n347551 );
not ( n2442 , n350128 );
buf ( n350130 , n2442 );
buf ( n350131 , n350130 );
not ( n2445 , n350131 );
buf ( n350133 , n2445 );
buf ( n350134 , n350133 );
not ( n2448 , n350134 );
or ( n2449 , n2440 , n2448 );
buf ( n350137 , n347565 );
buf ( n350138 , n554 );
buf ( n350139 , n588 );
xor ( n2453 , n350138 , n350139 );
buf ( n350141 , n2453 );
buf ( n350142 , n350141 );
nand ( n2456 , n350137 , n350142 );
buf ( n350144 , n2456 );
buf ( n350145 , n350144 );
nand ( n2459 , n2449 , n350145 );
buf ( n350147 , n2459 );
buf ( n350148 , n350147 );
xor ( n2462 , n350125 , n350148 );
buf ( n350150 , n559 );
buf ( n350151 , n584 );
xor ( n2465 , n350150 , n350151 );
buf ( n350153 , n2465 );
buf ( n350154 , n350153 );
not ( n2468 , n350154 );
xor ( n2469 , n585 , n584 );
nand ( n2470 , n2469 , n348614 );
not ( n2471 , n2470 );
buf ( n350159 , n2471 );
not ( n2473 , n350159 );
or ( n2474 , n2468 , n2473 );
buf ( n350162 , n348617 );
buf ( n350163 , n558 );
buf ( n350164 , n584 );
xor ( n2478 , n350163 , n350164 );
buf ( n350166 , n2478 );
buf ( n350167 , n350166 );
nand ( n2481 , n350162 , n350167 );
buf ( n350169 , n2481 );
buf ( n350170 , n350169 );
nand ( n2484 , n2474 , n350170 );
buf ( n350172 , n2484 );
buf ( n350173 , n350172 );
xor ( n2487 , n2462 , n350173 );
buf ( n350175 , n2487 );
buf ( n350176 , n350175 );
xor ( n2490 , n2413 , n350176 );
buf ( n350178 , n2490 );
buf ( n350179 , n350178 );
xor ( n2493 , n2359 , n350179 );
buf ( n350181 , n2493 );
buf ( n350182 , n350181 );
xor ( n2496 , n2336 , n350182 );
buf ( n350184 , n2496 );
buf ( n350185 , n350184 );
not ( n2499 , n350185 );
not ( n2500 , n921 );
not ( n2501 , n348462 );
nand ( n2502 , n2501 , n348533 );
not ( n2503 , n2502 );
or ( n2504 , n2500 , n2503 );
nand ( n2505 , n348462 , n348532 );
nand ( n2506 , n2504 , n2505 );
buf ( n350194 , n2506 );
not ( n2508 , n350194 );
buf ( n350196 , n2508 );
buf ( n350197 , n350196 );
nand ( n2511 , n2499 , n350197 );
buf ( n350199 , n2511 );
buf ( n350200 , n350199 );
buf ( n350201 , n347792 );
buf ( n350202 , n348076 );
buf ( n350203 , n348422 );
and ( n2517 , n350201 , n350202 , n350203 );
buf ( n350205 , n2517 );
buf ( n350206 , n350205 );
buf ( n350207 , n943 );
nand ( n2521 , n350200 , n350206 , n350207 );
buf ( n350209 , n2521 );
buf ( n350210 , n350184 );
not ( n2524 , n350210 );
buf ( n350212 , n2524 );
buf ( n350213 , n350212 );
buf ( n350214 , n350196 );
nand ( n2528 , n350213 , n350214 );
buf ( n350216 , n2528 );
nand ( n2530 , n350216 , n943 , n951 );
buf ( n350218 , n350216 );
buf ( n350219 , n348683 );
not ( n2533 , n350219 );
buf ( n350221 , n2533 );
buf ( n350222 , n350221 );
and ( n2536 , n350218 , n350222 );
buf ( n350224 , n350184 );
buf ( n350225 , n2506 );
nand ( n2539 , n350224 , n350225 );
buf ( n350227 , n2539 );
buf ( n350228 , n350227 );
not ( n2542 , n350228 );
buf ( n350230 , n2542 );
buf ( n350231 , n350230 );
nor ( n2545 , n2536 , n350231 );
buf ( n350233 , n2545 );
nand ( n2547 , n350209 , n2530 , n350233 );
buf ( n2548 , n2547 );
not ( n2549 , n2548 );
xor ( n2550 , n567 , n568 );
buf ( n350238 , n2550 );
buf ( n350239 , n559 );
and ( n2553 , n350238 , n350239 );
buf ( n350241 , n2553 );
buf ( n350242 , n350241 );
buf ( n350243 , n349876 );
not ( n2557 , n350243 );
buf ( n350245 , n347604 );
not ( n2559 , n350245 );
or ( n2560 , n2557 , n2559 );
buf ( n350248 , n551 );
buf ( n350249 , n574 );
xor ( n2563 , n350248 , n350249 );
buf ( n350251 , n2563 );
buf ( n350252 , n350251 );
buf ( n350253 , n575 );
nand ( n2567 , n350252 , n350253 );
buf ( n350255 , n2567 );
buf ( n350256 , n350255 );
nand ( n2570 , n2560 , n350256 );
buf ( n350258 , n2570 );
buf ( n350259 , n350258 );
xor ( n2573 , n350242 , n350259 );
buf ( n350261 , n349938 );
not ( n2575 , n350261 );
buf ( n350263 , n2236 );
not ( n2577 , n350263 );
or ( n2578 , n2575 , n2577 );
xor ( n2579 , n570 , n569 );
buf ( n350267 , n2579 );
buf ( n350268 , n557 );
buf ( n350269 , n568 );
xor ( n2583 , n350268 , n350269 );
buf ( n350271 , n2583 );
buf ( n350272 , n350271 );
nand ( n2586 , n350267 , n350272 );
buf ( n350274 , n2586 );
buf ( n350275 , n350274 );
nand ( n2589 , n2578 , n350275 );
buf ( n350277 , n2589 );
buf ( n350278 , n350277 );
xor ( n2592 , n2573 , n350278 );
buf ( n350280 , n2592 );
buf ( n350281 , n350280 );
not ( n2595 , n349962 );
not ( n2596 , n349944 );
or ( n2597 , n2595 , n2596 );
not ( n2598 , n349972 );
not ( n2599 , n349965 );
or ( n2600 , n2598 , n2599 );
nand ( n2601 , n2600 , n349995 );
nand ( n2602 , n2597 , n2601 );
buf ( n350290 , n2602 );
xor ( n2604 , n350281 , n350290 );
buf ( n350292 , n349956 );
not ( n2606 , n350292 );
buf ( n350294 , n347737 );
not ( n2608 , n350294 );
or ( n2609 , n2606 , n2608 );
buf ( n350297 , n347382 );
buf ( n350298 , n553 );
buf ( n350299 , n572 );
xor ( n2613 , n350298 , n350299 );
buf ( n350301 , n2613 );
buf ( n350302 , n350301 );
nand ( n2616 , n350297 , n350302 );
buf ( n350304 , n2616 );
buf ( n350305 , n350304 );
nand ( n2619 , n2609 , n350305 );
buf ( n350307 , n2619 );
buf ( n350308 , n350307 );
buf ( n350309 , n349989 );
not ( n2623 , n350309 );
buf ( n350311 , n348467 );
not ( n2625 , n350311 );
or ( n2626 , n2623 , n2625 );
buf ( n350314 , n347350 );
buf ( n350315 , n555 );
buf ( n350316 , n570 );
xor ( n2630 , n350315 , n350316 );
buf ( n350318 , n2630 );
buf ( n350319 , n350318 );
nand ( n2633 , n350314 , n350319 );
buf ( n350321 , n2633 );
buf ( n350322 , n350321 );
nand ( n2636 , n2626 , n350322 );
buf ( n350324 , n2636 );
buf ( n350325 , n350324 );
xor ( n2639 , n350308 , n350325 );
buf ( n350327 , n349883 );
buf ( n350328 , n349905 );
and ( n2642 , n350327 , n350328 );
buf ( n350330 , n2642 );
buf ( n350331 , n350330 );
xor ( n2645 , n2639 , n350331 );
buf ( n350333 , n2645 );
buf ( n350334 , n350333 );
xor ( n2648 , n2604 , n350334 );
buf ( n350336 , n2648 );
not ( n2650 , n350336 );
xor ( n2651 , n350029 , n350045 );
and ( n2652 , n2651 , n350179 );
and ( n2653 , n350029 , n350045 );
or ( n2654 , n2652 , n2653 );
buf ( n350342 , n2654 );
not ( n2656 , n350342 );
not ( n2657 , n2656 );
or ( n2658 , n2650 , n2657 );
not ( n2659 , n350336 );
nand ( n2660 , n350342 , n2659 );
nand ( n2661 , n2658 , n2660 );
not ( n2662 , n2180 );
nand ( n2663 , n2662 , n349909 );
not ( n2664 , n2663 );
not ( n2665 , n350005 );
or ( n2666 , n2664 , n2665 );
buf ( n350354 , n349909 );
not ( n2668 , n350354 );
buf ( n350356 , n2180 );
nand ( n2670 , n2668 , n350356 );
buf ( n350358 , n2670 );
nand ( n2672 , n2666 , n350358 );
buf ( n350360 , n2672 );
xor ( n2674 , n350088 , n350099 );
and ( n2675 , n2674 , n350176 );
and ( n2676 , n350088 , n350099 );
or ( n2677 , n2675 , n2676 );
buf ( n350365 , n2677 );
buf ( n350366 , n350365 );
xor ( n2680 , n350360 , n350366 );
buf ( n350368 , n583 );
buf ( n350369 , n584 );
xor ( n2683 , n350368 , n350369 );
buf ( n350371 , n2683 );
buf ( n350372 , n350371 );
not ( n2686 , n350372 );
buf ( n350374 , n2686 );
buf ( n350375 , n350374 );
not ( n2689 , n350375 );
buf ( n350377 , n2689 );
buf ( n350378 , n350377 );
buf ( n350379 , n559 );
and ( n2693 , n350378 , n350379 );
buf ( n350381 , n2693 );
buf ( n350382 , n350381 );
buf ( n350383 , n350072 );
not ( n2697 , n350383 );
buf ( n350385 , n347478 );
not ( n2699 , n350385 );
or ( n2700 , n2697 , n2699 );
buf ( n350388 , n551 );
buf ( n350389 , n590 );
xor ( n2703 , n350388 , n350389 );
buf ( n350391 , n2703 );
buf ( n350392 , n350391 );
buf ( n350393 , n591 );
nand ( n2707 , n350392 , n350393 );
buf ( n350395 , n2707 );
buf ( n350396 , n350395 );
nand ( n2710 , n2700 , n350396 );
buf ( n350398 , n2710 );
buf ( n350399 , n350398 );
xor ( n2713 , n350382 , n350399 );
buf ( n350401 , n350166 );
not ( n2715 , n350401 );
buf ( n350403 , n2471 );
not ( n2717 , n350403 );
or ( n2718 , n2715 , n2717 );
buf ( n350406 , n348617 );
buf ( n350407 , n557 );
buf ( n350408 , n584 );
xor ( n2722 , n350407 , n350408 );
buf ( n350410 , n2722 );
buf ( n350411 , n350410 );
nand ( n2725 , n350406 , n350411 );
buf ( n350413 , n2725 );
buf ( n350414 , n350413 );
nand ( n2728 , n2718 , n350414 );
buf ( n350416 , n2728 );
buf ( n350417 , n350416 );
xor ( n2731 , n2713 , n350417 );
buf ( n350419 , n2731 );
buf ( n350420 , n350419 );
xor ( n2734 , n350125 , n350148 );
and ( n2735 , n2734 , n350173 );
and ( n2736 , n350125 , n350148 );
or ( n2737 , n2735 , n2736 );
buf ( n350425 , n2737 );
buf ( n350426 , n350425 );
xor ( n2740 , n350420 , n350426 );
buf ( n350428 , n350118 );
not ( n2742 , n350428 );
buf ( n350430 , n347671 );
not ( n2744 , n350430 );
or ( n2745 , n2742 , n2744 );
buf ( n350433 , n347530 );
buf ( n350434 , n555 );
buf ( n350435 , n586 );
xor ( n2749 , n350434 , n350435 );
buf ( n350437 , n2749 );
buf ( n350438 , n350437 );
nand ( n2752 , n350433 , n350438 );
buf ( n350440 , n2752 );
buf ( n350441 , n350440 );
nand ( n2755 , n2745 , n350441 );
buf ( n350443 , n2755 );
buf ( n350444 , n350443 );
not ( n2758 , n350444 );
buf ( n350446 , n2758 );
buf ( n350447 , n350446 );
not ( n2761 , n350447 );
buf ( n350449 , n350141 );
not ( n2763 , n350449 );
buf ( n350451 , n347757 );
not ( n2765 , n350451 );
or ( n2766 , n2763 , n2765 );
buf ( n350454 , n347568 );
buf ( n350455 , n553 );
buf ( n350456 , n588 );
xor ( n2770 , n350455 , n350456 );
buf ( n350458 , n2770 );
buf ( n350459 , n350458 );
nand ( n2773 , n350454 , n350459 );
buf ( n350461 , n2773 );
buf ( n350462 , n350461 );
nand ( n2776 , n2766 , n350462 );
buf ( n350464 , n2776 );
buf ( n350465 , n350464 );
not ( n2779 , n350465 );
or ( n2780 , n2761 , n2779 );
buf ( n350468 , n350141 );
not ( n2782 , n350468 );
buf ( n350470 , n347757 );
not ( n2784 , n350470 );
or ( n2785 , n2782 , n2784 );
buf ( n350473 , n350461 );
nand ( n2787 , n2785 , n350473 );
buf ( n350475 , n2787 );
buf ( n350476 , n350475 );
buf ( n350477 , n350446 );
or ( n2791 , n350476 , n350477 );
nand ( n2792 , n2780 , n2791 );
buf ( n350480 , n2792 );
buf ( n350481 , n350480 );
buf ( n350482 , n350061 );
not ( n2796 , n350482 );
buf ( n350484 , n350079 );
nand ( n2798 , n2796 , n350484 );
buf ( n350486 , n2798 );
buf ( n350487 , n350486 );
not ( n2801 , n350487 );
buf ( n350489 , n2801 );
buf ( n350490 , n350489 );
xor ( n2804 , n350481 , n350490 );
buf ( n350492 , n2804 );
buf ( n350493 , n350492 );
xor ( n2807 , n2740 , n350493 );
buf ( n350495 , n2807 );
buf ( n350496 , n350495 );
xor ( n2810 , n2680 , n350496 );
buf ( n350498 , n2810 );
and ( n2812 , n2661 , n350498 );
not ( n2813 , n2661 );
not ( n2814 , n350498 );
and ( n2815 , n2813 , n2814 );
nor ( n2816 , n2812 , n2815 );
not ( n2817 , n2816 );
xor ( n2818 , n350011 , n350022 );
and ( n2819 , n2818 , n350182 );
and ( n2820 , n350011 , n350022 );
or ( n2821 , n2819 , n2820 );
buf ( n350509 , n2821 );
not ( n2823 , n350509 );
and ( n2824 , n2817 , n2823 );
buf ( n350512 , n350271 );
not ( n2826 , n350512 );
nand ( n2827 , n2230 , n2235 );
not ( n2828 , n2827 );
buf ( n350516 , n2828 );
not ( n2830 , n350516 );
or ( n2831 , n2826 , n2830 );
buf ( n350519 , n2579 );
and ( n2833 , n556 , n568 );
not ( n2834 , n556 );
and ( n2835 , n2834 , n1822 );
nor ( n2836 , n2833 , n2835 );
buf ( n350524 , n2836 );
nand ( n2838 , n350519 , n350524 );
buf ( n350526 , n2838 );
buf ( n350527 , n350526 );
nand ( n2841 , n2831 , n350527 );
buf ( n350529 , n2841 );
buf ( n350530 , n559 );
buf ( n350531 , n566 );
xor ( n2845 , n350530 , n350531 );
buf ( n350533 , n2845 );
buf ( n350534 , n350533 );
not ( n2848 , n350534 );
xor ( n2849 , n567 , n566 );
xnor ( n2850 , n567 , n568 );
and ( n2851 , n2849 , n2850 );
buf ( n350539 , n2851 );
not ( n2853 , n350539 );
or ( n2854 , n2848 , n2853 );
buf ( n350542 , n2550 );
buf ( n350543 , n558 );
buf ( n350544 , n566 );
xor ( n2858 , n350543 , n350544 );
buf ( n350546 , n2858 );
buf ( n350547 , n350546 );
nand ( n2861 , n350542 , n350547 );
buf ( n350549 , n2861 );
buf ( n350550 , n350549 );
nand ( n2864 , n2854 , n350550 );
buf ( n350552 , n2864 );
xor ( n2866 , n350529 , n350552 );
buf ( n350554 , n350251 );
not ( n2868 , n350554 );
buf ( n350556 , n347604 );
not ( n2870 , n350556 );
or ( n2871 , n2868 , n2870 );
buf ( n350559 , n550 );
buf ( n350560 , n574 );
xor ( n2874 , n350559 , n350560 );
buf ( n350562 , n2874 );
buf ( n350563 , n350562 );
buf ( n350564 , n575 );
nand ( n2878 , n350563 , n350564 );
buf ( n350566 , n2878 );
buf ( n350567 , n350566 );
nand ( n2881 , n2871 , n350567 );
buf ( n350569 , n2881 );
xor ( n2883 , n2866 , n350569 );
buf ( n350571 , n2883 );
xor ( n2885 , n350308 , n350325 );
and ( n2886 , n2885 , n350331 );
and ( n2887 , n350308 , n350325 );
or ( n2888 , n2886 , n2887 );
buf ( n350576 , n2888 );
buf ( n350577 , n350576 );
xor ( n2891 , n350571 , n350577 );
buf ( n350579 , n350318 );
not ( n2893 , n350579 );
buf ( n350581 , n348467 );
not ( n2895 , n350581 );
or ( n2896 , n2893 , n2895 );
buf ( n350584 , n348476 );
buf ( n350585 , n554 );
buf ( n350586 , n570 );
xor ( n2900 , n350585 , n350586 );
buf ( n350588 , n2900 );
buf ( n350589 , n350588 );
nand ( n2903 , n350584 , n350589 );
buf ( n350591 , n2903 );
buf ( n350592 , n350591 );
nand ( n2906 , n2896 , n350592 );
buf ( n350594 , n2906 );
buf ( n350595 , n350594 );
not ( n2909 , n350301 );
not ( n2910 , n347737 );
or ( n2911 , n2909 , n2910 );
buf ( n350599 , n347382 );
buf ( n350600 , n552 );
buf ( n350601 , n572 );
xor ( n2915 , n350600 , n350601 );
buf ( n350603 , n2915 );
buf ( n350604 , n350603 );
nand ( n2918 , n350599 , n350604 );
buf ( n350606 , n2918 );
nand ( n2920 , n2911 , n350606 );
buf ( n350608 , n559 );
buf ( n350609 , n567 );
nand ( n2923 , n350608 , n350609 );
buf ( n350611 , n2923 );
or ( n2925 , n559 , n567 );
nand ( n2926 , n2925 , n568 );
nand ( n2927 , n350611 , n2926 , n566 );
and ( n2928 , n2920 , n2927 );
not ( n2929 , n2920 );
not ( n2930 , n2927 );
and ( n2931 , n2929 , n2930 );
or ( n2932 , n2928 , n2931 );
buf ( n350620 , n2932 );
xor ( n2934 , n350595 , n350620 );
xor ( n2935 , n350242 , n350259 );
and ( n2936 , n2935 , n350278 );
and ( n2937 , n350242 , n350259 );
or ( n2938 , n2936 , n2937 );
buf ( n350626 , n2938 );
buf ( n350627 , n350626 );
xor ( n2941 , n2934 , n350627 );
buf ( n350629 , n2941 );
buf ( n350630 , n350629 );
xor ( n2944 , n2891 , n350630 );
buf ( n350632 , n2944 );
buf ( n350633 , n350632 );
xor ( n2947 , n350360 , n350366 );
and ( n2948 , n2947 , n350496 );
and ( n2949 , n350360 , n350366 );
or ( n2950 , n2948 , n2949 );
buf ( n350638 , n2950 );
buf ( n350639 , n350638 );
xor ( n2953 , n350633 , n350639 );
xor ( n2954 , n350281 , n350290 );
and ( n2955 , n2954 , n350334 );
and ( n2956 , n350281 , n350290 );
or ( n2957 , n2955 , n2956 );
buf ( n350645 , n2957 );
buf ( n350646 , n350645 );
xor ( n2960 , n350420 , n350426 );
and ( n2961 , n2960 , n350493 );
and ( n2962 , n350420 , n350426 );
or ( n2963 , n2961 , n2962 );
buf ( n350651 , n2963 );
buf ( n350652 , n350651 );
xor ( n2966 , n350646 , n350652 );
buf ( n350654 , n350446 );
not ( n2968 , n350654 );
buf ( n350656 , n350486 );
not ( n2970 , n350656 );
or ( n2971 , n2968 , n2970 );
buf ( n350659 , n350475 );
nand ( n2973 , n2971 , n350659 );
buf ( n350661 , n2973 );
buf ( n350662 , n350661 );
buf ( n350663 , n350489 );
buf ( n350664 , n350443 );
nand ( n2978 , n350663 , n350664 );
buf ( n350666 , n2978 );
buf ( n350667 , n350666 );
nand ( n2981 , n350662 , n350667 );
buf ( n350669 , n2981 );
buf ( n350670 , n350669 );
buf ( n350671 , n350391 );
not ( n2985 , n350671 );
buf ( n350673 , n347478 );
not ( n2987 , n350673 );
or ( n2988 , n2985 , n2987 );
buf ( n350676 , n550 );
buf ( n350677 , n590 );
xor ( n2991 , n350676 , n350677 );
buf ( n350679 , n2991 );
buf ( n350680 , n350679 );
buf ( n350681 , n591 );
nand ( n2995 , n350680 , n350681 );
buf ( n350683 , n2995 );
buf ( n350684 , n350683 );
nand ( n2998 , n2988 , n350684 );
buf ( n350686 , n2998 );
buf ( n350687 , n350686 );
buf ( n350688 , n559 );
buf ( n350689 , n582 );
xor ( n3003 , n350688 , n350689 );
buf ( n350691 , n3003 );
buf ( n350692 , n350691 );
not ( n3006 , n350692 );
xnor ( n3007 , n583 , n584 );
xor ( n3008 , n583 , n582 );
nand ( n3009 , n3007 , n3008 );
buf ( n350697 , n3009 );
not ( n3011 , n350697 );
buf ( n350699 , n3011 );
buf ( n350700 , n350699 );
not ( n3014 , n350700 );
or ( n3015 , n3006 , n3014 );
buf ( n350703 , n350371 );
buf ( n3017 , n350703 );
buf ( n350705 , n3017 );
buf ( n350706 , n350705 );
buf ( n350707 , n558 );
buf ( n350708 , n582 );
xor ( n3022 , n350707 , n350708 );
buf ( n350710 , n3022 );
buf ( n350711 , n350710 );
nand ( n3025 , n350706 , n350711 );
buf ( n350713 , n3025 );
buf ( n350714 , n350713 );
nand ( n3028 , n3015 , n350714 );
buf ( n350716 , n3028 );
buf ( n350717 , n350716 );
xor ( n3031 , n350687 , n350717 );
buf ( n350719 , n350410 );
not ( n3033 , n350719 );
buf ( n350721 , n2471 );
not ( n3035 , n350721 );
or ( n3036 , n3033 , n3035 );
buf ( n350724 , n348626 );
not ( n3038 , n350724 );
buf ( n350726 , n3038 );
buf ( n350727 , n350726 );
buf ( n350728 , n556 );
buf ( n350729 , n584 );
xor ( n3043 , n350728 , n350729 );
buf ( n350731 , n3043 );
buf ( n350732 , n350731 );
nand ( n3046 , n350727 , n350732 );
buf ( n350734 , n3046 );
buf ( n350735 , n350734 );
nand ( n3049 , n3036 , n350735 );
buf ( n350737 , n3049 );
buf ( n350738 , n350737 );
xor ( n3052 , n3031 , n350738 );
buf ( n350740 , n3052 );
buf ( n350741 , n350740 );
xor ( n3055 , n350670 , n350741 );
buf ( n350743 , n350437 );
not ( n3057 , n350743 );
buf ( n350745 , n347671 );
not ( n3059 , n350745 );
or ( n3060 , n3057 , n3059 );
buf ( n350748 , n347530 );
and ( n3062 , n586 , n554 );
not ( n3063 , n586 );
not ( n3064 , n554 );
and ( n3065 , n3063 , n3064 );
nor ( n3066 , n3062 , n3065 );
buf ( n350754 , n3066 );
nand ( n3068 , n350748 , n350754 );
buf ( n350756 , n3068 );
buf ( n350757 , n350756 );
nand ( n3071 , n3060 , n350757 );
buf ( n350759 , n3071 );
buf ( n350760 , n350759 );
buf ( n350761 , n559 );
buf ( n350762 , n583 );
or ( n3076 , n350761 , n350762 );
buf ( n350764 , n584 );
nand ( n3078 , n3076 , n350764 );
buf ( n350766 , n3078 );
buf ( n350767 , n350766 );
buf ( n350768 , n559 );
buf ( n350769 , n583 );
nand ( n3083 , n350768 , n350769 );
buf ( n350771 , n3083 );
buf ( n350772 , n350771 );
buf ( n350773 , n582 );
and ( n3087 , n350767 , n350772 , n350773 );
buf ( n350775 , n3087 );
buf ( n350776 , n350458 );
not ( n3090 , n350776 );
not ( n3091 , n590 );
nand ( n3092 , n3091 , n589 );
and ( n3093 , n347543 , n347548 , n3092 );
buf ( n350781 , n3093 );
not ( n3095 , n350781 );
or ( n3096 , n3090 , n3095 );
buf ( n350784 , n347565 );
buf ( n350785 , n552 );
buf ( n350786 , n588 );
xor ( n3100 , n350785 , n350786 );
buf ( n350788 , n3100 );
buf ( n350789 , n350788 );
nand ( n3103 , n350784 , n350789 );
buf ( n350791 , n3103 );
buf ( n350792 , n350791 );
nand ( n3106 , n3096 , n350792 );
buf ( n350794 , n3106 );
xor ( n3108 , n350775 , n350794 );
buf ( n350796 , n3108 );
xor ( n3110 , n350760 , n350796 );
xor ( n3111 , n350382 , n350399 );
and ( n3112 , n3111 , n350417 );
and ( n3113 , n350382 , n350399 );
or ( n3114 , n3112 , n3113 );
buf ( n350802 , n3114 );
buf ( n350803 , n350802 );
xor ( n3117 , n3110 , n350803 );
buf ( n350805 , n3117 );
buf ( n350806 , n350805 );
xor ( n3120 , n3055 , n350806 );
buf ( n350808 , n3120 );
buf ( n350809 , n350808 );
xor ( n3123 , n2966 , n350809 );
buf ( n350811 , n3123 );
buf ( n350812 , n350811 );
xor ( n3126 , n2953 , n350812 );
buf ( n350814 , n3126 );
buf ( n350815 , n350814 );
nand ( n3129 , n2659 , n2656 );
not ( n3130 , n3129 );
not ( n3131 , n350498 );
or ( n3132 , n3130 , n3131 );
nand ( n3133 , n350336 , n350342 );
nand ( n3134 , n3132 , n3133 );
buf ( n350822 , n3134 );
nor ( n3136 , n350815 , n350822 );
buf ( n350824 , n3136 );
nor ( n3138 , n2824 , n350824 );
not ( n3139 , n3138 );
or ( n3140 , n2549 , n3139 );
buf ( n350828 , n2816 );
buf ( n350829 , n350509 );
nand ( n3143 , n350828 , n350829 );
buf ( n350831 , n3143 );
buf ( n350832 , n350831 );
buf ( n350833 , n350824 );
or ( n3147 , n350832 , n350833 );
buf ( n350835 , n350814 );
buf ( n350836 , n3134 );
nand ( n3150 , n350835 , n350836 );
buf ( n350838 , n3150 );
buf ( n350839 , n350838 );
nand ( n3153 , n3147 , n350839 );
buf ( n350841 , n3153 );
buf ( n350842 , n350841 );
not ( n3156 , n350842 );
buf ( n350844 , n3156 );
nand ( n3158 , n3140 , n350844 );
xor ( n3159 , n350633 , n350639 );
and ( n3160 , n3159 , n350812 );
and ( n3161 , n350633 , n350639 );
or ( n3162 , n3160 , n3161 );
buf ( n350850 , n3162 );
not ( n3164 , n350850 );
buf ( n350852 , n350562 );
not ( n3166 , n350852 );
buf ( n350854 , n347604 );
not ( n3168 , n350854 );
or ( n3169 , n3166 , n3168 );
and ( n3170 , n574 , n549 );
not ( n3171 , n574 );
not ( n3172 , n549 );
and ( n3173 , n3171 , n3172 );
nor ( n3174 , n3170 , n3173 );
buf ( n350862 , n3174 );
buf ( n350863 , n575 );
nand ( n3177 , n350862 , n350863 );
buf ( n350865 , n3177 );
buf ( n350866 , n350865 );
nand ( n3180 , n3169 , n350866 );
buf ( n350868 , n3180 );
buf ( n350869 , n350546 );
not ( n3183 , n350869 );
nand ( n3184 , n2850 , n2849 );
buf ( n350872 , n3184 );
not ( n3186 , n350872 );
buf ( n350874 , n3186 );
buf ( n350875 , n350874 );
not ( n3189 , n350875 );
or ( n3190 , n3183 , n3189 );
not ( n3191 , n2850 );
xor ( n3192 , n566 , n557 );
nand ( n3193 , n3191 , n3192 );
buf ( n350881 , n3193 );
nand ( n3195 , n3190 , n350881 );
buf ( n350883 , n3195 );
xor ( n3197 , n350868 , n350883 );
buf ( n350885 , n350588 );
not ( n3199 , n350885 );
buf ( n350887 , n347344 );
not ( n3201 , n350887 );
or ( n3202 , n3199 , n3201 );
buf ( n350890 , n347350 );
buf ( n350891 , n553 );
buf ( n350892 , n570 );
xor ( n3206 , n350891 , n350892 );
buf ( n350894 , n3206 );
buf ( n350895 , n350894 );
nand ( n3209 , n350890 , n350895 );
buf ( n350897 , n3209 );
buf ( n350898 , n350897 );
nand ( n3212 , n3202 , n350898 );
buf ( n350900 , n3212 );
xor ( n3214 , n3197 , n350900 );
buf ( n350902 , n3214 );
xor ( n3216 , n350595 , n350620 );
and ( n3217 , n3216 , n350627 );
and ( n3218 , n350595 , n350620 );
or ( n3219 , n3217 , n3218 );
buf ( n350907 , n3219 );
buf ( n350908 , n350907 );
xor ( n3222 , n350902 , n350908 );
nand ( n3223 , n2920 , n2930 );
not ( n3224 , n350569 );
not ( n3225 , n350529 );
or ( n3226 , n3224 , n3225 );
buf ( n350914 , n350569 );
buf ( n350915 , n350529 );
or ( n3229 , n350914 , n350915 );
buf ( n350917 , n350552 );
nand ( n3231 , n3229 , n350917 );
buf ( n350919 , n3231 );
nand ( n3233 , n3226 , n350919 );
xor ( n3234 , n3223 , n3233 );
xor ( n3235 , n565 , n566 );
buf ( n350923 , n3235 );
buf ( n350924 , n559 );
and ( n3238 , n350923 , n350924 );
buf ( n350926 , n3238 );
not ( n3240 , n350603 );
nand ( n3241 , n347369 , n347372 );
and ( n3242 , n347376 , n3241 );
not ( n3243 , n3242 );
or ( n3244 , n3240 , n3243 );
buf ( n350932 , n551 );
buf ( n350933 , n572 );
xor ( n3247 , n350932 , n350933 );
buf ( n350935 , n3247 );
nand ( n3249 , n347382 , n350935 );
nand ( n3250 , n3244 , n3249 );
xor ( n3251 , n350926 , n3250 );
not ( n3252 , n2836 );
not ( n3253 , n2236 );
or ( n3254 , n3252 , n3253 );
buf ( n350942 , n2579 );
buf ( n350943 , n555 );
buf ( n350944 , n568 );
xor ( n3258 , n350943 , n350944 );
buf ( n350946 , n3258 );
buf ( n350947 , n350946 );
nand ( n3261 , n350942 , n350947 );
buf ( n350949 , n3261 );
nand ( n3263 , n3254 , n350949 );
xnor ( n3264 , n3251 , n3263 );
buf ( n350952 , n3264 );
not ( n3266 , n350952 );
buf ( n350954 , n3266 );
xnor ( n3268 , n3234 , n350954 );
buf ( n350956 , n3268 );
xor ( n3270 , n3222 , n350956 );
buf ( n350958 , n3270 );
buf ( n350959 , n350958 );
xor ( n3273 , n350646 , n350652 );
and ( n3274 , n3273 , n350809 );
and ( n3275 , n350646 , n350652 );
or ( n3276 , n3274 , n3275 );
buf ( n350964 , n3276 );
buf ( n350965 , n350964 );
xor ( n3279 , n350959 , n350965 );
xor ( n3280 , n350571 , n350577 );
and ( n3281 , n3280 , n350630 );
and ( n3282 , n350571 , n350577 );
or ( n3283 , n3281 , n3282 );
buf ( n350971 , n3283 );
buf ( n350972 , n350971 );
xor ( n3286 , n350670 , n350741 );
and ( n3287 , n3286 , n350806 );
and ( n3288 , n350670 , n350741 );
or ( n3289 , n3287 , n3288 );
buf ( n350977 , n3289 );
buf ( n350978 , n350977 );
xor ( n3292 , n350972 , n350978 );
xor ( n3293 , n586 , n553 );
not ( n3294 , n3293 );
not ( n3295 , n347530 );
or ( n3296 , n3294 , n3295 );
nand ( n3297 , n347664 , n347669 , n3066 );
nand ( n3298 , n3296 , n3297 );
not ( n3299 , n347478 );
not ( n3300 , n350679 );
or ( n3301 , n3299 , n3300 );
and ( n3302 , n590 , n549 );
not ( n3303 , n590 );
and ( n3304 , n3303 , n3172 );
nor ( n3305 , n3302 , n3304 );
buf ( n350993 , n3305 );
buf ( n350994 , n591 );
nand ( n3308 , n350993 , n350994 );
buf ( n350996 , n3308 );
nand ( n3310 , n3301 , n350996 );
nor ( n3311 , n3298 , n3310 );
nand ( n3312 , n3008 , n350374 );
not ( n3313 , n3312 );
nand ( n3314 , n350710 , n3313 );
buf ( n351002 , n350705 );
buf ( n351003 , n557 );
buf ( n351004 , n582 );
xor ( n3318 , n351003 , n351004 );
buf ( n351006 , n3318 );
buf ( n351007 , n351006 );
nand ( n3321 , n351002 , n351007 );
buf ( n351009 , n3321 );
and ( n3323 , n3314 , n351009 );
not ( n3324 , n3323 );
nand ( n3325 , n3311 , n3324 );
nand ( n3326 , n3324 , n3298 , n3310 );
not ( n3327 , n3310 );
nand ( n3328 , n3323 , n3298 , n3327 );
not ( n3329 , n3298 );
nand ( n3330 , n3323 , n3329 , n3310 );
nand ( n3331 , n3325 , n3326 , n3328 , n3330 );
buf ( n351019 , n3331 );
xor ( n3333 , n350760 , n350796 );
and ( n3334 , n3333 , n350803 );
and ( n3335 , n350760 , n350796 );
or ( n3336 , n3334 , n3335 );
buf ( n351024 , n3336 );
buf ( n351025 , n351024 );
xor ( n3339 , n351019 , n351025 );
buf ( n351027 , n350794 );
buf ( n351028 , n350775 );
and ( n3342 , n351027 , n351028 );
buf ( n351030 , n3342 );
buf ( n351031 , n351030 );
xor ( n3345 , n581 , n582 );
buf ( n351033 , n3345 );
not ( n3347 , n351033 );
buf ( n351035 , n3347 );
buf ( n351036 , n351035 );
not ( n3350 , n351036 );
buf ( n351038 , n3350 );
buf ( n351039 , n351038 );
buf ( n351040 , n559 );
and ( n3354 , n351039 , n351040 );
buf ( n351042 , n3354 );
buf ( n351043 , n350788 );
not ( n3357 , n351043 );
buf ( n351045 , n3093 );
not ( n3359 , n351045 );
or ( n3360 , n3357 , n3359 );
nand ( n3361 , n348137 , n590 );
nand ( n3362 , n3091 , n589 );
nand ( n3363 , n3361 , n3362 );
buf ( n351051 , n551 );
buf ( n351052 , n588 );
xor ( n3366 , n351051 , n351052 );
buf ( n351054 , n3366 );
nand ( n3368 , n3363 , n351054 );
buf ( n351056 , n3368 );
nand ( n3370 , n3360 , n351056 );
buf ( n351058 , n3370 );
xor ( n3372 , n351042 , n351058 );
buf ( n351060 , n350731 );
not ( n3374 , n351060 );
buf ( n351062 , n2471 );
not ( n3376 , n351062 );
or ( n3377 , n3374 , n3376 );
buf ( n351065 , n350726 );
buf ( n351066 , n555 );
buf ( n351067 , n584 );
xor ( n3381 , n351066 , n351067 );
buf ( n351069 , n3381 );
buf ( n351070 , n351069 );
nand ( n3384 , n351065 , n351070 );
buf ( n351072 , n3384 );
buf ( n351073 , n351072 );
nand ( n3387 , n3377 , n351073 );
buf ( n351075 , n3387 );
xor ( n3389 , n3372 , n351075 );
buf ( n351077 , n3389 );
xor ( n3391 , n351031 , n351077 );
xor ( n3392 , n350687 , n350717 );
and ( n3393 , n3392 , n350738 );
and ( n3394 , n350687 , n350717 );
or ( n3395 , n3393 , n3394 );
buf ( n351083 , n3395 );
buf ( n351084 , n351083 );
xor ( n3398 , n3391 , n351084 );
buf ( n351086 , n3398 );
buf ( n351087 , n351086 );
xor ( n3401 , n3339 , n351087 );
buf ( n351089 , n3401 );
buf ( n351090 , n351089 );
xor ( n3404 , n3292 , n351090 );
buf ( n351092 , n3404 );
buf ( n351093 , n351092 );
xor ( n3407 , n3279 , n351093 );
buf ( n351095 , n3407 );
not ( n3409 , n351095 );
or ( n3410 , n3164 , n3409 );
buf ( n351098 , n351095 );
not ( n3412 , n351098 );
buf ( n351100 , n3412 );
buf ( n351101 , n350850 );
not ( n3415 , n351101 );
buf ( n351103 , n3415 );
nand ( n3417 , n351100 , n351103 );
nand ( n3418 , n3410 , n3417 );
and ( n3419 , n3158 , n3418 );
not ( n3420 , n3158 );
not ( n3421 , n3418 );
and ( n3422 , n3420 , n3421 );
nor ( n3423 , n3419 , n3422 );
not ( n3424 , n3423 );
nand ( n3425 , n2176 , n3424 );
nand ( n3426 , n2175 , n3423 );
nand ( n3427 , n3425 , n3426 );
or ( n3428 , n348445 , n348455 );
buf ( n351116 , n926 );
not ( n3430 , n351116 );
buf ( n351118 , n348690 );
nand ( n3432 , n3430 , n351118 );
buf ( n351120 , n3432 );
nand ( n3434 , n351120 , n951 );
buf ( n351122 , n926 );
not ( n3436 , n351122 );
buf ( n351124 , n348690 );
nand ( n3438 , n3436 , n351124 );
buf ( n351126 , n3438 );
buf ( n351127 , n348697 );
buf ( n351128 , n347862 );
nor ( n3442 , n351127 , n351128 );
buf ( n351130 , n3442 );
nand ( n3444 , n351126 , n351130 , n348076 );
nand ( n3445 , n3434 , n3444 , n348686 );
not ( n3446 , n350230 );
nand ( n3447 , n3446 , n350199 );
not ( n3448 , n3447 );
and ( n3449 , n3445 , n3448 );
not ( n3450 , n3445 );
and ( n3451 , n3450 , n3447 );
nor ( n3452 , n3449 , n3451 );
not ( n3453 , n3452 );
not ( n3454 , n2166 );
nand ( n3455 , n3454 , n2153 );
nand ( n3456 , n3455 , n2167 );
buf ( n3457 , n2163 );
and ( n3458 , n3456 , n3457 );
not ( n3459 , n3456 );
not ( n3460 , n3457 );
and ( n3461 , n3459 , n3460 );
nor ( n3462 , n3458 , n3461 );
not ( n3463 , n3462 );
nand ( n3464 , n3453 , n3463 );
nand ( n3465 , n3428 , n3464 , n1051 );
nand ( n3466 , n3452 , n3462 );
not ( n3467 , n3466 );
not ( n3468 , n3452 );
and ( n3469 , n3468 , n3463 );
nor ( n3470 , n3469 , n1053 );
nor ( n3471 , n3467 , n3470 );
nand ( n3472 , n3465 , n3471 );
buf ( n3473 , n3472 );
not ( n3474 , n3473 );
and ( n3475 , n2139 , n2140 );
not ( n3476 , n2139 );
and ( n3477 , n3476 , n2113 );
or ( n3478 , n3475 , n3477 );
not ( n3479 , n3478 );
not ( n3480 , n2120 );
nand ( n3481 , n3480 , n2170 );
not ( n3482 , n3481 );
buf ( n3483 , n2168 );
not ( n3484 , n3483 );
or ( n3485 , n3482 , n3484 );
nand ( n3486 , n2120 , n2135 );
nand ( n3487 , n3485 , n3486 );
not ( n3488 , n3487 );
or ( n3489 , n3479 , n3488 );
or ( n3490 , n3478 , n3487 );
nand ( n3491 , n3489 , n3490 );
buf ( n351179 , n350814 );
not ( n3493 , n351179 );
buf ( n351181 , n3134 );
not ( n3495 , n351181 );
buf ( n351183 , n3495 );
buf ( n351184 , n351183 );
nand ( n3498 , n3493 , n351184 );
buf ( n351186 , n3498 );
nand ( n3500 , n350838 , n351186 );
not ( n3501 , n3500 );
not ( n3502 , n350509 );
not ( n3503 , n2816 );
nand ( n3504 , n3502 , n3503 );
not ( n3505 , n3504 );
not ( n3506 , n2547 );
or ( n3507 , n3505 , n3506 );
nand ( n3508 , n3507 , n350831 );
not ( n3509 , n3508 );
and ( n3510 , n3501 , n3509 );
and ( n3511 , n3500 , n3508 );
nor ( n3512 , n3510 , n3511 );
nand ( n3513 , n3491 , n3512 );
buf ( n351201 , n2548 );
buf ( n351202 , n3504 );
buf ( n351203 , n350831 );
and ( n3517 , n351202 , n351203 );
buf ( n351205 , n3517 );
buf ( n351206 , n351205 );
xor ( n3520 , n351201 , n351206 );
buf ( n351208 , n3520 );
not ( n3522 , n351208 );
nand ( n3523 , n3481 , n3486 );
not ( n3524 , n3523 );
not ( n3525 , n3483 );
or ( n3526 , n3524 , n3525 );
or ( n3527 , n3483 , n3523 );
nand ( n3528 , n3526 , n3527 );
nand ( n3529 , n3522 , n3528 );
and ( n3530 , n3513 , n3529 );
not ( n3531 , n3530 );
or ( n3532 , n3474 , n3531 );
not ( n3533 , n3528 );
nand ( n3534 , n3533 , n351208 );
not ( n3535 , n3534 );
not ( n3536 , n3535 );
not ( n3537 , n3513 );
or ( n3538 , n3536 , n3537 );
not ( n3539 , n3491 );
not ( n3540 , n3512 );
nand ( n3541 , n3539 , n3540 );
nand ( n3542 , n3538 , n3541 );
not ( n3543 , n3542 );
nand ( n3544 , n3532 , n3543 );
xor ( n3545 , n3427 , n3544 );
not ( n3546 , n581 );
nand ( n3547 , n3545 , n3546 );
nand ( n3551 , C1 , n1139 );
nand ( n3552 , n1051 , n348455 );
nand ( n3553 , n1051 , n348445 );
nand ( n3554 , n3552 , n3553 , n1053 );
and ( n3555 , n3464 , n3466 );
and ( n3556 , n3554 , n3555 );
not ( n3557 , n3554 );
not ( n3558 , n3555 );
and ( n3559 , n3557 , n3558 );
nor ( n3560 , n3556 , n3559 );
not ( n3561 , n3560 );
nand ( n3562 , n3561 , n1820 );
nand ( n3563 , n3551 , n3562 , n1064 );
not ( n3564 , n3561 );
nand ( n3565 , n3564 , n584 );
not ( n3566 , n1061 );
nand ( n3567 , n3566 , n3562 );
nand ( n3568 , n3563 , n3565 , n3567 );
and ( n3569 , n3529 , n3534 );
and ( n3570 , n3569 , n3473 );
not ( n3571 , n3569 );
not ( n3572 , n3473 );
and ( n3573 , n3571 , n3572 );
nor ( n3574 , n3570 , n3573 );
not ( n3575 , n3574 );
not ( n3576 , n583 );
and ( n3577 , n3575 , n3576 );
not ( n3578 , n3529 );
not ( n3579 , n3472 );
or ( n3580 , n3578 , n3579 );
nand ( n3581 , n3580 , n3534 );
not ( n3582 , n3581 );
nand ( n3583 , n3513 , n3541 );
not ( n3584 , n3583 );
nand ( n3585 , n3582 , n3584 );
nand ( n3586 , n3581 , n3583 );
not ( n3587 , n582 );
and ( n3588 , n3585 , n3586 , n3587 );
nor ( n3589 , n3577 , n3588 );
nand ( n3590 , n3547 , n3568 , n3589 );
buf ( n351275 , n583 );
not ( n3592 , n351275 );
buf ( n351277 , n3592 );
not ( n3594 , n351277 );
nand ( n3595 , n3594 , n3574 );
or ( n3596 , n3588 , n3595 );
not ( n3597 , n3586 );
not ( n3598 , n3585 );
or ( n3599 , n3597 , n3598 );
nand ( n3600 , n3599 , n582 );
nand ( n3601 , n3596 , n3600 );
nand ( n3602 , n3601 , n3547 );
not ( n3603 , n3545 );
nand ( n3604 , n3603 , n581 );
nand ( n3605 , n3590 , n3602 , n3604 );
nand ( n3606 , n3542 , n3426 );
nand ( n3607 , n3423 , n2175 );
nand ( n3608 , n3530 , n3607 , n3473 );
nand ( n3609 , n3606 , n3608 , n3425 );
not ( n3610 , n3609 );
buf ( n351295 , n351186 );
buf ( n351296 , n3504 );
nand ( n3613 , n351295 , n351296 );
buf ( n351298 , n3613 );
buf ( n351299 , n351298 );
buf ( n351300 , n351095 );
buf ( n351301 , n350850 );
nor ( n3618 , n351300 , n351301 );
buf ( n351303 , n3618 );
buf ( n351304 , n351303 );
nor ( n3621 , n351299 , n351304 );
buf ( n351306 , n3621 );
not ( n3623 , n351306 );
not ( n3624 , n2548 );
or ( n3625 , n3623 , n3624 );
and ( n3626 , n350841 , n3417 );
and ( n3627 , n351095 , n350850 );
nor ( n3628 , n3626 , n3627 );
nand ( n3629 , n3625 , n3628 );
buf ( n351314 , n559 );
buf ( n351315 , n564 );
xor ( n3632 , n351314 , n351315 );
buf ( n351317 , n3632 );
buf ( n351318 , n351317 );
not ( n3635 , n351318 );
buf ( n351320 , n3235 );
not ( n3637 , n351320 );
buf ( n351322 , n3637 );
buf ( n351323 , n351322 );
xor ( n3640 , n564 , n565 );
buf ( n351325 , n3640 );
nand ( n3642 , n351323 , n351325 );
buf ( n351327 , n3642 );
buf ( n351328 , n351327 );
not ( n3645 , n351328 );
buf ( n351330 , n3645 );
buf ( n351331 , n351330 );
not ( n3648 , n351331 );
or ( n3649 , n3635 , n3648 );
buf ( n3650 , n3235 );
buf ( n351335 , n3650 );
buf ( n351336 , n558 );
buf ( n351337 , n564 );
xor ( n3654 , n351336 , n351337 );
buf ( n351339 , n3654 );
buf ( n351340 , n351339 );
nand ( n3657 , n351335 , n351340 );
buf ( n351342 , n3657 );
buf ( n351343 , n351342 );
nand ( n3660 , n3649 , n351343 );
buf ( n351345 , n3660 );
buf ( n351346 , n351345 );
buf ( n351347 , n350894 );
not ( n3664 , n351347 );
buf ( n351349 , n348467 );
not ( n3666 , n351349 );
or ( n3667 , n3664 , n3666 );
buf ( n351352 , n348476 );
buf ( n351353 , n552 );
buf ( n351354 , n570 );
xor ( n3671 , n351353 , n351354 );
buf ( n351356 , n3671 );
buf ( n351357 , n351356 );
nand ( n3674 , n351352 , n351357 );
buf ( n351359 , n3674 );
buf ( n351360 , n351359 );
nand ( n3677 , n3667 , n351360 );
buf ( n351362 , n3677 );
buf ( n351363 , n351362 );
xor ( n3680 , n351346 , n351363 );
buf ( n351365 , n559 );
buf ( n351366 , n565 );
or ( n3683 , n351365 , n351366 );
buf ( n351368 , n566 );
nand ( n3685 , n3683 , n351368 );
buf ( n351370 , n3685 );
buf ( n351371 , n351370 );
buf ( n351372 , n559 );
buf ( n351373 , n565 );
nand ( n3690 , n351372 , n351373 );
buf ( n351375 , n3690 );
buf ( n351376 , n351375 );
buf ( n351377 , n564 );
and ( n3694 , n351371 , n351376 , n351377 );
buf ( n351379 , n3694 );
buf ( n351380 , n351379 );
buf ( n351381 , n350935 );
not ( n3698 , n351381 );
buf ( n351383 , n347378 );
not ( n3700 , n351383 );
or ( n3701 , n3698 , n3700 );
buf ( n351386 , n347382 );
xor ( n3703 , n572 , n550 );
buf ( n351388 , n3703 );
nand ( n3705 , n351386 , n351388 );
buf ( n351390 , n3705 );
buf ( n351391 , n351390 );
nand ( n3708 , n3701 , n351391 );
buf ( n351393 , n3708 );
buf ( n351394 , n351393 );
xor ( n3711 , n351380 , n351394 );
buf ( n351396 , n3711 );
buf ( n351397 , n351396 );
xor ( n3714 , n3680 , n351397 );
buf ( n351399 , n3714 );
buf ( n351400 , n351399 );
not ( n3717 , n3223 );
not ( n3718 , n3717 );
not ( n3719 , n350954 );
or ( n3720 , n3718 , n3719 );
not ( n3721 , n3223 );
not ( n3722 , n3264 );
or ( n3723 , n3721 , n3722 );
nand ( n3724 , n3723 , n3233 );
nand ( n3725 , n3720 , n3724 );
buf ( n351410 , n3725 );
xor ( n3727 , n351400 , n351410 );
buf ( n351412 , n350868 );
not ( n3729 , n351412 );
buf ( n351414 , n350883 );
not ( n3731 , n351414 );
or ( n3732 , n3729 , n3731 );
buf ( n351417 , n350883 );
buf ( n351418 , n350868 );
or ( n3735 , n351417 , n351418 );
buf ( n351420 , n350900 );
nand ( n3737 , n3735 , n351420 );
buf ( n351422 , n3737 );
buf ( n351423 , n351422 );
nand ( n3740 , n3732 , n351423 );
buf ( n351425 , n3740 );
buf ( n351426 , n351425 );
buf ( n351427 , n350926 );
not ( n3744 , n351427 );
buf ( n351429 , n3250 );
not ( n3746 , n351429 );
or ( n3747 , n3744 , n3746 );
or ( n3748 , n3250 , n350926 );
nand ( n3749 , n3748 , n3263 );
buf ( n351434 , n3749 );
nand ( n3751 , n3747 , n351434 );
buf ( n351436 , n3751 );
buf ( n351437 , n351436 );
xor ( n3754 , n351426 , n351437 );
not ( n3755 , n575 );
buf ( n351440 , n548 );
buf ( n351441 , n574 );
xor ( n3758 , n351440 , n351441 );
buf ( n351443 , n3758 );
not ( n3760 , n351443 );
or ( n3761 , n3755 , n3760 );
not ( n3762 , n574 );
nor ( n3763 , n3762 , n575 );
nand ( n3764 , n3763 , n3174 );
nand ( n3765 , n3761 , n3764 );
buf ( n351450 , n3765 );
not ( n3767 , n350946 );
not ( n3768 , n2827 );
not ( n3769 , n3768 );
or ( n3770 , n3767 , n3769 );
buf ( n351455 , n348495 );
buf ( n351456 , n554 );
buf ( n351457 , n568 );
xor ( n3774 , n351456 , n351457 );
buf ( n351459 , n3774 );
buf ( n351460 , n351459 );
nand ( n3777 , n351455 , n351460 );
buf ( n351462 , n3777 );
nand ( n3779 , n3770 , n351462 );
buf ( n351464 , n3779 );
xor ( n3781 , n351450 , n351464 );
buf ( n351466 , n3192 );
not ( n3783 , n351466 );
buf ( n351468 , n350874 );
not ( n3785 , n351468 );
or ( n3786 , n3783 , n3785 );
buf ( n351471 , n2550 );
xor ( n3788 , n566 , n556 );
buf ( n351473 , n3788 );
nand ( n3790 , n351471 , n351473 );
buf ( n351475 , n3790 );
buf ( n351476 , n351475 );
nand ( n3793 , n3786 , n351476 );
buf ( n351478 , n3793 );
buf ( n351479 , n351478 );
xor ( n3796 , n3781 , n351479 );
buf ( n351481 , n3796 );
buf ( n351482 , n351481 );
xor ( n3799 , n3754 , n351482 );
buf ( n351484 , n3799 );
buf ( n351485 , n351484 );
xor ( n3802 , n3727 , n351485 );
buf ( n351487 , n3802 );
buf ( n351488 , n351487 );
xor ( n3805 , n350972 , n350978 );
and ( n3806 , n3805 , n351090 );
and ( n3807 , n350972 , n350978 );
or ( n3808 , n3806 , n3807 );
buf ( n351493 , n3808 );
buf ( n351494 , n351493 );
xor ( n3811 , n351488 , n351494 );
xor ( n3812 , n350902 , n350908 );
and ( n3813 , n3812 , n350956 );
and ( n3814 , n350902 , n350908 );
or ( n3815 , n3813 , n3814 );
buf ( n351500 , n3815 );
buf ( n351501 , n351500 );
xor ( n3818 , n351019 , n351025 );
and ( n3819 , n3818 , n351087 );
and ( n3820 , n351019 , n351025 );
or ( n3821 , n3819 , n3820 );
buf ( n351506 , n3821 );
buf ( n351507 , n351506 );
xor ( n3824 , n351501 , n351507 );
buf ( n351509 , n559 );
buf ( n351510 , n581 );
or ( n3827 , n351509 , n351510 );
buf ( n351512 , n582 );
nand ( n3829 , n3827 , n351512 );
buf ( n351514 , n3829 );
buf ( n351515 , n351514 );
buf ( n351516 , n559 );
buf ( n351517 , n581 );
nand ( n3834 , n351516 , n351517 );
buf ( n351519 , n3834 );
buf ( n351520 , n351519 );
buf ( n351521 , n580 );
and ( n3838 , n351515 , n351520 , n351521 );
buf ( n351523 , n3838 );
buf ( n351524 , n351054 );
not ( n3841 , n351524 );
buf ( n351526 , n347554 );
not ( n3843 , n351526 );
or ( n3844 , n3841 , n3843 );
buf ( n351529 , n347565 );
buf ( n351530 , n550 );
buf ( n351531 , n588 );
xor ( n3848 , n351530 , n351531 );
buf ( n351533 , n3848 );
buf ( n351534 , n351533 );
nand ( n3851 , n351529 , n351534 );
buf ( n351536 , n3851 );
buf ( n351537 , n351536 );
nand ( n3854 , n3844 , n351537 );
buf ( n351539 , n3854 );
xor ( n3856 , n351523 , n351539 );
not ( n3857 , n3856 );
buf ( n351542 , n559 );
buf ( n351543 , n580 );
xor ( n3860 , n351542 , n351543 );
buf ( n351545 , n3860 );
not ( n3862 , n351545 );
not ( n3863 , n580 );
not ( n3864 , n3546 );
or ( n3865 , n3863 , n3864 );
not ( n3866 , n580 );
nand ( n3867 , n3866 , n581 );
nand ( n3868 , n3865 , n3867 );
nand ( n3869 , n3868 , n351035 );
not ( n3870 , n3869 );
not ( n3871 , n3870 );
or ( n3872 , n3862 , n3871 );
buf ( n351557 , n351038 );
buf ( n3874 , n351557 );
buf ( n351559 , n3874 );
buf ( n351560 , n351559 );
buf ( n351561 , n558 );
buf ( n351562 , n580 );
xor ( n3879 , n351561 , n351562 );
buf ( n351564 , n3879 );
buf ( n351565 , n351564 );
nand ( n3882 , n351560 , n351565 );
buf ( n351567 , n3882 );
nand ( n3884 , n3872 , n351567 );
not ( n3885 , n3293 );
not ( n3886 , n347671 );
or ( n3887 , n3885 , n3886 );
buf ( n351572 , n347530 );
buf ( n351573 , n552 );
buf ( n351574 , n586 );
xor ( n3891 , n351573 , n351574 );
buf ( n351576 , n3891 );
buf ( n351577 , n351576 );
nand ( n3894 , n351572 , n351577 );
buf ( n351579 , n3894 );
nand ( n3896 , n3887 , n351579 );
not ( n3897 , n3896 );
and ( n3898 , n3884 , n3897 );
not ( n3899 , n3884 );
and ( n3900 , n3899 , n3896 );
nor ( n3901 , n3898 , n3900 );
not ( n3902 , n3901 );
or ( n3903 , n3857 , n3902 );
or ( n3904 , n3856 , n3901 );
nand ( n3905 , n3903 , n3904 );
buf ( n351590 , n3905 );
xor ( n3907 , n351031 , n351077 );
and ( n3908 , n3907 , n351084 );
and ( n3909 , n351031 , n351077 );
or ( n3910 , n3908 , n3909 );
buf ( n351595 , n3910 );
buf ( n351596 , n351595 );
xor ( n3913 , n351590 , n351596 );
not ( n3914 , n3327 );
not ( n3915 , n3329 );
or ( n3916 , n3914 , n3915 );
nand ( n3917 , n3916 , n3324 );
nand ( n3918 , n3298 , n3310 );
nand ( n3919 , n3917 , n3918 );
xor ( n3920 , n351042 , n351058 );
and ( n3921 , n3920 , n351075 );
and ( n3922 , n351042 , n351058 );
or ( n3923 , n3921 , n3922 );
xor ( n3924 , n3919 , n3923 );
not ( n3925 , n3305 );
not ( n3926 , n347478 );
or ( n3927 , n3925 , n3926 );
xor ( n3928 , n590 , n548 );
nand ( n3929 , n3928 , n591 );
nand ( n3930 , n3927 , n3929 );
not ( n3931 , n351069 );
not ( n3932 , n2471 );
or ( n3933 , n3931 , n3932 );
buf ( n351618 , n348617 );
buf ( n351619 , n554 );
buf ( n351620 , n584 );
xor ( n3937 , n351619 , n351620 );
buf ( n351622 , n3937 );
buf ( n351623 , n351622 );
nand ( n3940 , n351618 , n351623 );
buf ( n351625 , n3940 );
nand ( n3942 , n3933 , n351625 );
xor ( n3943 , n3930 , n3942 );
buf ( n351628 , n556 );
buf ( n351629 , n582 );
xor ( n3946 , n351628 , n351629 );
buf ( n351631 , n3946 );
and ( n3948 , n350705 , n351631 );
and ( n3949 , n350699 , n351006 );
nor ( n3950 , n3948 , n3949 );
not ( n3951 , n3950 );
xor ( n3952 , n3943 , n3951 );
xor ( n3953 , n3924 , n3952 );
buf ( n351638 , n3953 );
xor ( n3955 , n3913 , n351638 );
buf ( n351640 , n3955 );
buf ( n351641 , n351640 );
xor ( n3958 , n3824 , n351641 );
buf ( n351643 , n3958 );
buf ( n351644 , n351643 );
xor ( n3961 , n3811 , n351644 );
buf ( n351646 , n3961 );
buf ( n351647 , n351646 );
not ( n3964 , n351647 );
buf ( n351649 , n3964 );
xor ( n3966 , n350959 , n350965 );
and ( n3967 , n3966 , n351093 );
and ( n3968 , n350959 , n350965 );
or ( n3969 , n3967 , n3968 );
buf ( n351654 , n3969 );
buf ( n351655 , n351654 );
not ( n3972 , n351655 );
buf ( n351657 , n3972 );
nand ( n3974 , n351649 , n351657 );
not ( n3975 , n3974 );
nand ( n3976 , n351646 , n351654 );
not ( n3977 , n3976 );
nor ( n3978 , n3975 , n3977 );
buf ( n3979 , n3978 );
and ( n3980 , n3629 , n3979 );
not ( n3981 , n3629 );
buf ( n351666 , n3978 );
not ( n3983 , n351666 );
buf ( n351668 , n3983 );
and ( n3985 , n3981 , n351668 );
or ( n3986 , n3980 , n3985 );
xor ( n3987 , n2012 , n2016 );
and ( n3988 , n3987 , n2086 );
and ( n3989 , n2012 , n2016 );
or ( n3990 , n3988 , n3989 );
not ( n3991 , n3990 );
not ( n3992 , n1022 );
not ( n3993 , n2007 );
or ( n3994 , n3992 , n3993 );
not ( n3995 , n554 );
not ( n3996 , n1788 );
not ( n3997 , n3996 );
or ( n3998 , n3995 , n3997 );
not ( n3999 , n554 );
nand ( n4000 , n3999 , n1788 );
nand ( n4001 , n3998 , n4000 );
nand ( n4002 , n4001 , n1925 );
nand ( n4003 , n3994 , n4002 );
xor ( n4004 , n2021 , n2031 );
and ( n4005 , n4004 , n2043 );
and ( n4006 , n2021 , n2031 );
or ( n4007 , n4005 , n4006 );
xor ( n4008 , n4003 , n4007 );
not ( n4009 , n348090 );
not ( n4010 , n556 );
not ( n4011 , n1974 );
not ( n4012 , n4011 );
or ( n4013 , n4010 , n4012 );
nand ( n4014 , n1974 , n348119 );
nand ( n4015 , n4013 , n4014 );
not ( n4016 , n4015 );
or ( n4017 , n4009 , n4016 );
nand ( n4018 , n1996 , n348153 );
nand ( n4019 , n4017 , n4018 );
xor ( n4020 , n4008 , n4019 );
xor ( n4021 , n2044 , n2080 );
and ( n4022 , n4021 , n2085 );
and ( n4023 , n2044 , n2080 );
or ( n4024 , n4022 , n4023 );
xor ( n4025 , n4020 , n4024 );
not ( n4026 , n559 );
not ( n4027 , n558 );
nand ( n4028 , n564 , n580 );
not ( n4029 , n4028 );
nor ( n4030 , n564 , n580 );
nor ( n4031 , n4029 , n4030 );
not ( n4032 , n4031 );
and ( n4033 , n2049 , n2063 );
not ( n4034 , n4033 );
not ( n4035 , n1815 );
not ( n4036 , n1807 );
or ( n4037 , n4035 , n4036 );
not ( n4038 , n349519 );
not ( n4039 , n1837 );
or ( n4040 , n4038 , n4039 );
nand ( n351725 , n1825 , n1818 );
nand ( n351726 , n4040 , n351725 );
nand ( n351727 , n4037 , n351726 );
not ( n351728 , n351727 );
or ( n4045 , n4034 , n351728 );
and ( n351730 , n2063 , n2059 );
not ( n351731 , n2064 );
nor ( n4048 , n351730 , n351731 );
nand ( n351733 , n4045 , n4048 );
not ( n351734 , n351733 );
not ( n4051 , n351734 );
or ( n351736 , n4032 , n4051 );
not ( n351737 , n4028 );
or ( n4054 , n351737 , n4030 );
nand ( n351739 , n4054 , n351733 );
nand ( n351740 , n351736 , n351739 );
not ( n4057 , n351740 );
not ( n351742 , n4057 );
or ( n351743 , n4027 , n351742 );
not ( n4060 , n4057 );
nand ( n351745 , n4060 , n348230 );
nand ( n351746 , n351743 , n351745 );
not ( n4063 , n351746 );
or ( n351748 , n4026 , n4063 );
nand ( n351749 , n2076 , n348233 );
nand ( n4066 , n351748 , n351749 );
not ( n351751 , n1875 );
not ( n351752 , n550 );
not ( n4069 , n1856 );
or ( n351754 , n351752 , n4069 );
not ( n351755 , n348115 );
nand ( n4072 , n351755 , n1880 );
nand ( n351757 , n351754 , n4072 );
not ( n351758 , n351757 );
or ( n4075 , n351751 , n351758 );
not ( n351760 , n1890 );
not ( n351761 , n1874 );
and ( n4078 , n351760 , n351761 );
nand ( n351763 , n2027 , n4078 );
nand ( n351764 , n4075 , n351763 );
or ( n4081 , n549 , n550 );
nand ( n351766 , n4081 , n348158 );
nand ( n351767 , n549 , n550 );
and ( n4084 , n351766 , n351767 , n548 );
not ( n351769 , n2019 );
not ( n351770 , n548 );
not ( n4087 , n348171 );
or ( n351772 , n351770 , n4087 );
not ( n351773 , n548 );
nand ( n4090 , n348174 , n351773 );
nand ( n4091 , n351772 , n4090 );
not ( n4092 , n4091 );
or ( n4093 , n351769 , n4092 );
not ( n4094 , n548 );
not ( n4095 , n348181 );
or ( n4096 , n4094 , n4095 );
nand ( n4097 , n348158 , n351773 );
nand ( n4098 , n4096 , n4097 );
xnor ( n4099 , n548 , n549 );
and ( n4100 , n549 , n1880 );
not ( n4101 , n549 );
and ( n4102 , n4101 , n550 );
or ( n4103 , n4100 , n4102 );
nor ( n4104 , n4099 , n4103 );
nand ( n4105 , n4098 , n4104 );
nand ( n4106 , n4093 , n4105 );
xor ( n4107 , n4084 , n4106 );
xor ( n4108 , n351764 , n4107 );
buf ( n4109 , n1011 );
not ( n4110 , n4109 );
not ( n4111 , n552 );
not ( n4112 , n348270 );
or ( n4113 , n4111 , n4112 );
not ( n4114 , n348266 );
or ( n4115 , n4114 , n552 );
nand ( n4116 , n4113 , n4115 );
not ( n4117 , n4116 );
or ( n4118 , n4110 , n4117 );
nand ( n4119 , n1871 , n2039 );
nand ( n4120 , n4118 , n4119 );
xor ( n4121 , n4108 , n4120 );
xor ( n4122 , n4066 , n4121 );
xor ( n4123 , n1989 , n1998 );
and ( n4124 , n4123 , n2011 );
and ( n4125 , n1989 , n1998 );
or ( n4126 , n4124 , n4125 );
xor ( n4127 , n4122 , n4126 );
xor ( n4128 , n4025 , n4127 );
not ( n4129 , n4128 );
or ( n4130 , n3991 , n4129 );
nor ( n4131 , n4128 , n3990 );
not ( n4132 , n4131 );
nand ( n4133 , n4130 , n4132 );
not ( n4134 , n4133 );
not ( n4135 , n2087 );
not ( n351820 , n1988 );
nand ( n351821 , n4135 , n351820 );
nand ( n4138 , n2173 , n351821 );
not ( n351823 , n4138 );
not ( n4140 , n351823 );
nand ( n351825 , n2088 , n1988 );
nand ( n4142 , n4140 , n351825 );
not ( n4143 , n4142 );
or ( n351828 , n4134 , n4143 );
not ( n4145 , n351823 );
nand ( n4146 , n4145 , n351825 );
or ( n4147 , n4146 , n4133 );
nand ( n4148 , n351828 , n4147 );
nor ( n4149 , n3986 , n4148 );
not ( n4150 , n4149 );
and ( n4151 , n3629 , n3979 );
not ( n4152 , n3629 );
and ( n4153 , n4152 , n351668 );
nor ( n4154 , n4151 , n4153 );
not ( n4155 , n4154 );
not ( n4156 , n4133 );
not ( n4157 , n4142 );
or ( n4158 , n4156 , n4157 );
or ( n4159 , n4133 , n4146 );
nand ( n351844 , n4158 , n4159 );
nand ( n351845 , n4155 , n351844 );
nand ( n4162 , n4150 , n351845 );
and ( n351847 , n3610 , n4162 );
not ( n4164 , n3610 );
not ( n351849 , n4162 );
and ( n4166 , n4164 , n351849 );
nor ( n4167 , n351847 , n4166 );
nor ( n4168 , n580 , n4167 );
not ( n4169 , n4168 );
and ( n4170 , n3610 , n4162 );
not ( n4171 , n3610 );
and ( n4172 , n4171 , n351849 );
nor ( n4173 , n4170 , n4172 );
nand ( n4174 , n4173 , n580 );
nand ( n4175 , n4169 , n4174 );
or ( n4176 , n3605 , n4175 );
nand ( n4177 , n3605 , n4175 );
nand ( n4178 , n4176 , n4177 );
not ( n4179 , n4178 );
buf ( n351864 , n4179 );
not ( n4181 , n351864 );
or ( n4182 , n1726 , n4181 );
buf ( n4183 , n4178 );
buf ( n351868 , n4183 );
not ( n4185 , n351868 );
buf ( n351870 , n4185 );
buf ( n351871 , n351870 );
not ( n4188 , n351871 );
buf ( n351873 , n4188 );
buf ( n351874 , n351873 );
not ( n351875 , n600 );
buf ( n4192 , n351875 );
buf ( n4193 , n4192 );
buf ( n351878 , n4193 );
nand ( n4195 , n351874 , n351878 );
buf ( n351880 , n4195 );
buf ( n351881 , n351880 );
nand ( n4198 , n4182 , n351881 );
buf ( n351883 , n4198 );
buf ( n351884 , n351883 );
not ( n351885 , n351884 );
or ( n4202 , n1724 , n351885 );
buf ( n351887 , n600 );
not ( n4204 , n351887 );
nand ( n4205 , n3545 , n3546 );
nand ( n4206 , n4205 , n3604 );
not ( n4207 , n4206 );
not ( n4208 , n3589 );
not ( n4209 , n3568 );
or ( n4210 , n4208 , n4209 );
not ( n4211 , n3601 );
nand ( n4212 , n4210 , n4211 );
not ( n4213 , n4212 );
or ( n4214 , n4207 , n4213 );
or ( n4215 , n4212 , n4206 );
nand ( n4216 , n4214 , n4215 );
not ( n351901 , n4216 );
buf ( n351902 , n351901 );
not ( n351903 , n351902 );
or ( n4220 , n4204 , n351903 );
buf ( n4221 , n4216 );
buf ( n351906 , n4221 );
buf ( n351907 , n4193 );
nand ( n4224 , n351906 , n351907 );
buf ( n351909 , n4224 );
buf ( n351910 , n351909 );
nand ( n4227 , n4220 , n351910 );
buf ( n351912 , n4227 );
buf ( n351913 , n351912 );
buf ( n351914 , n600 );
buf ( n351915 , n601 );
and ( n351916 , n351914 , n351915 );
buf ( n351917 , n1721 );
buf ( n351918 , n600 );
buf ( n351919 , n601 );
nor ( n4236 , n351918 , n351919 );
buf ( n351921 , n4236 );
buf ( n351922 , n351921 );
nor ( n4239 , n351916 , n351917 , n351922 );
buf ( n351924 , n4239 );
buf ( n351925 , n351924 );
nand ( n4242 , n351913 , n351925 );
buf ( n351927 , n4242 );
buf ( n351928 , n351927 );
nand ( n4245 , n4202 , n351928 );
buf ( n351930 , n4245 );
buf ( n351931 , n351930 );
xor ( n4248 , n349401 , n351931 );
buf ( n351933 , n347319 );
not ( n4250 , n351933 );
buf ( n351935 , n596 );
not ( n4252 , n351935 );
not ( n4253 , n1139 );
or ( n351938 , n4253 , C0 );
or ( n4256 , n1060 , n585 );
nand ( n4257 , n351938 , n4256 );
nand ( n4258 , n4257 , n1061 );
not ( n4259 , n4258 );
not ( n4260 , n4259 );
nand ( n4261 , n3565 , n3562 );
not ( n4262 , n4261 );
not ( n4263 , n4262 );
or ( n4264 , n4260 , n4263 );
nand ( n4265 , n4261 , n4258 );
nand ( n4266 , n4264 , n4265 );
buf ( n351950 , n4266 );
not ( n4268 , n351950 );
buf ( n351952 , n4268 );
buf ( n351953 , n351952 );
not ( n4271 , n351953 );
or ( n4272 , n4252 , n4271 );
buf ( n351956 , n4266 );
buf ( n4274 , n351956 );
buf ( n351958 , n4274 );
buf ( n351959 , n351958 );
buf ( n351960 , n348865 );
nand ( n4278 , n351959 , n351960 );
buf ( n351962 , n4278 );
buf ( n351963 , n351962 );
nand ( n351964 , n4272 , n351963 );
buf ( n351965 , n351964 );
buf ( n351966 , n351965 );
not ( n4284 , n351966 );
or ( n4285 , n4250 , n4284 );
buf ( n351969 , n348871 );
buf ( n351970 , n348898 );
nand ( n4288 , n351969 , n351970 );
buf ( n351972 , n4288 );
buf ( n351973 , n351972 );
nand ( n4291 , n4285 , n351973 );
buf ( n351975 , n4291 );
buf ( n351976 , n351975 );
buf ( n351977 , n349035 );
not ( n4295 , n351977 );
buf ( n351979 , n594 );
not ( n4297 , n351979 );
not ( n4298 , n1179 );
buf ( n351982 , n4298 );
not ( n4300 , n351982 );
or ( n4301 , n4297 , n4300 );
buf ( n351985 , n348884 );
buf ( n351986 , n348975 );
nand ( n4304 , n351985 , n351986 );
buf ( n351988 , n4304 );
buf ( n351989 , n351988 );
nand ( n4307 , n4301 , n351989 );
buf ( n351991 , n4307 );
buf ( n351992 , n351991 );
not ( n4310 , n351992 );
or ( n4311 , n4295 , n4310 );
buf ( n351995 , n1362 );
buf ( n351996 , n1397 );
nand ( n351997 , n351995 , n351996 );
buf ( n351998 , n351997 );
buf ( n351999 , n351998 );
nand ( n4317 , n4311 , n351999 );
buf ( n352001 , n4317 );
buf ( n352002 , n352001 );
buf ( n352003 , n348934 );
buf ( n352004 , n592 );
and ( n4322 , n352003 , n352004 );
buf ( n352006 , n4322 );
buf ( n352007 , n352006 );
xor ( n4325 , n348914 , n348992 );
and ( n4326 , n4325 , n349023 );
or ( n4328 , n4326 , C0 );
buf ( n352011 , n4328 );
buf ( n352012 , n352011 );
xor ( n4331 , n352007 , n352012 );
and ( n4332 , n349067 , n348910 );
not ( n4333 , n349067 );
and ( n4334 , n4333 , n592 );
nor ( n4335 , n4332 , n4334 );
or ( n4336 , n4335 , n349013 );
buf ( n352019 , n349009 );
not ( n4338 , n352019 );
buf ( n352021 , n1250 );
nand ( n4340 , n4338 , n352021 );
buf ( n352023 , n4340 );
nand ( n4342 , n4336 , n352023 );
buf ( n352025 , n4342 );
xor ( n4344 , n4331 , n352025 );
buf ( n352027 , n4344 );
buf ( n352028 , n352027 );
xor ( n4347 , n352002 , n352028 );
xor ( n4348 , n349026 , n349093 );
and ( n4349 , n4348 , n349212 );
and ( n4350 , n349026 , n349093 );
or ( n4351 , n4349 , n4350 );
buf ( n352034 , n4351 );
buf ( n352035 , n352034 );
xor ( n4354 , n4347 , n352035 );
buf ( n352037 , n4354 );
buf ( n352038 , n352037 );
xor ( n4357 , n351976 , n352038 );
and ( n4358 , n599 , n600 );
not ( n4359 , n599 );
and ( n4360 , n4359 , n351875 );
nor ( n4361 , n4358 , n4360 );
buf ( n4362 , n4361 );
buf ( n352045 , n4362 );
not ( n4364 , n352045 );
buf ( n352047 , n598 );
not ( n4366 , n352047 );
and ( n4367 , n3569 , n3572 );
not ( n4368 , n3569 );
and ( n4369 , n4368 , n3473 );
nor ( n4370 , n4367 , n4369 );
nand ( n4371 , n351277 , n4370 );
not ( n4372 , n4371 );
not ( n4373 , n3568 );
or ( n4374 , n4372 , n4373 );
buf ( n4375 , n3595 );
nand ( n4376 , n4374 , n4375 );
not ( n4377 , n3588 );
nand ( n4378 , n4377 , n3600 );
not ( n4379 , n4378 );
and ( n4380 , n4376 , n4379 );
not ( n4381 , n4376 );
and ( n4382 , n4381 , n4378 );
nor ( n352065 , n4380 , n4382 );
not ( n352066 , n352065 );
buf ( n352067 , n352066 );
not ( n4386 , n352067 );
or ( n4387 , n4366 , n4386 );
buf ( n4388 , n352065 );
buf ( n352071 , n4388 );
buf ( n352072 , n347312 );
nand ( n4391 , n352071 , n352072 );
buf ( n352074 , n4391 );
buf ( n352075 , n352074 );
nand ( n4394 , n4387 , n352075 );
buf ( n352077 , n4394 );
buf ( n352078 , n352077 );
not ( n4397 , n352078 );
or ( n4398 , n4364 , n4397 );
buf ( n352081 , n598 );
not ( n4400 , n352081 );
not ( n4401 , n583 );
not ( n352084 , n3574 );
or ( n4403 , n4401 , n352084 );
nand ( n352086 , n4403 , n4371 );
nand ( n4405 , n3563 , n3565 , n3567 );
and ( n4406 , n352086 , n4405 );
not ( n4407 , n352086 );
not ( n4408 , n4405 );
and ( n4409 , n4407 , n4408 );
nor ( n4410 , n4406 , n4409 );
buf ( n352093 , n4410 );
buf ( n4412 , n352093 );
buf ( n352095 , n4412 );
buf ( n352096 , n352095 );
not ( n4415 , n352096 );
or ( n4416 , n4400 , n4415 );
buf ( n352099 , n352095 );
not ( n352100 , n352099 );
buf ( n352101 , n352100 );
buf ( n352102 , n352101 );
buf ( n352103 , n347312 );
nand ( n4422 , n352102 , n352103 );
buf ( n352105 , n4422 );
buf ( n352106 , n352105 );
nand ( n4425 , n4416 , n352106 );
buf ( n352108 , n4425 );
buf ( n352109 , n352108 );
buf ( n352110 , n4361 );
not ( n4429 , n352110 );
buf ( n352112 , n4429 );
buf ( n352113 , n352112 );
buf ( n352114 , n599 );
buf ( n352115 , n598 );
and ( n4434 , n352114 , n352115 );
not ( n352117 , n352114 );
buf ( n352118 , n347312 );
and ( n4437 , n352117 , n352118 );
nor ( n4438 , n4434 , n4437 );
buf ( n352121 , n4438 );
buf ( n352122 , n352121 );
and ( n4441 , n352113 , n352122 );
buf ( n352124 , n4441 );
buf ( n4443 , n352124 );
buf ( n352126 , n4443 );
nand ( n4445 , n352109 , n352126 );
buf ( n352128 , n4445 );
buf ( n352129 , n352128 );
nand ( n4448 , n4398 , n352129 );
buf ( n352131 , n4448 );
buf ( n352132 , n352131 );
xor ( n4451 , n4357 , n352132 );
buf ( n352134 , n4451 );
buf ( n352135 , n352134 );
and ( n4454 , n4248 , n352135 );
and ( n4455 , n349401 , n351931 );
or ( n4456 , n4454 , n4455 );
buf ( n352139 , n4456 );
buf ( n352140 , n352139 );
or ( n4459 , n603 , n604 );
buf ( n352142 , n603 );
buf ( n352143 , n604 );
nand ( n4462 , n352142 , n352143 );
buf ( n352145 , n4462 );
nand ( n4464 , n4459 , n352145 );
buf ( n352147 , n4464 );
not ( n4466 , n352147 );
buf ( n352149 , n4466 );
buf ( n352150 , n352149 );
not ( n4469 , n352150 );
buf ( n352152 , n602 );
not ( n4471 , n352152 );
xor ( n4472 , n351346 , n351363 );
and ( n4473 , n4472 , n351397 );
and ( n4474 , n351346 , n351363 );
or ( n4475 , n4473 , n4474 );
buf ( n352158 , n4475 );
not ( n4477 , n352158 );
buf ( n352160 , n547 );
buf ( n352161 , n574 );
xor ( n4480 , n352160 , n352161 );
buf ( n352163 , n4480 );
not ( n4482 , n352163 );
not ( n4483 , n575 );
or ( n4484 , n4482 , n4483 );
nand ( n4485 , n351443 , n3763 );
nand ( n4486 , n4484 , n4485 );
not ( n4487 , n351339 );
not ( n4488 , n3640 );
xor ( n4489 , n565 , n566 );
nor ( n4490 , n4488 , n4489 );
not ( n4491 , n4490 );
or ( n4492 , n4487 , n4491 );
buf ( n352175 , n3650 );
buf ( n352176 , n557 );
buf ( n352177 , n564 );
xor ( n4496 , n352176 , n352177 );
buf ( n352179 , n4496 );
buf ( n352180 , n352179 );
nand ( n4499 , n352175 , n352180 );
buf ( n352182 , n4499 );
nand ( n4501 , n4492 , n352182 );
xor ( n4502 , n4486 , n4501 );
not ( n4503 , n3788 );
not ( n4504 , n350874 );
or ( n4505 , n4503 , n4504 );
buf ( n352188 , n2550 );
buf ( n352189 , n555 );
buf ( n352190 , n566 );
xor ( n4509 , n352189 , n352190 );
buf ( n352192 , n4509 );
buf ( n352193 , n352192 );
nand ( n352194 , n352188 , n352193 );
buf ( n352195 , n352194 );
nand ( n4514 , n4505 , n352195 );
xor ( n4515 , n4502 , n4514 );
not ( n4516 , n4515 );
buf ( n352199 , n563 );
buf ( n352200 , n564 );
xor ( n4519 , n352199 , n352200 );
buf ( n352202 , n4519 );
buf ( n352203 , n352202 );
not ( n352204 , n352203 );
buf ( n352205 , n347984 );
nor ( n4524 , n352204 , n352205 );
buf ( n352207 , n4524 );
buf ( n352208 , n352207 );
buf ( n352209 , n3703 );
not ( n4528 , n352209 );
buf ( n352211 , n3242 );
not ( n4530 , n352211 );
or ( n4531 , n4528 , n4530 );
buf ( n352214 , n347382 );
xor ( n4533 , n572 , n549 );
buf ( n352216 , n4533 );
nand ( n4535 , n352214 , n352216 );
buf ( n352218 , n4535 );
buf ( n352219 , n352218 );
nand ( n4538 , n4531 , n352219 );
buf ( n352221 , n4538 );
buf ( n352222 , n352221 );
xor ( n4541 , n352208 , n352222 );
buf ( n352224 , n351459 );
not ( n4543 , n352224 );
buf ( n352226 , n2828 );
not ( n4545 , n352226 );
or ( n352228 , n4543 , n4545 );
buf ( n352229 , n2243 );
xor ( n352230 , n568 , n553 );
buf ( n352231 , n352230 );
nand ( n4550 , n352229 , n352231 );
buf ( n352233 , n4550 );
buf ( n352234 , n352233 );
nand ( n4553 , n352228 , n352234 );
buf ( n352236 , n4553 );
buf ( n352237 , n352236 );
xor ( n4556 , n4541 , n352237 );
buf ( n352239 , n4556 );
not ( n4558 , n352239 );
nand ( n4559 , n4516 , n4558 );
not ( n4560 , n4559 );
or ( n4561 , n4477 , n4560 );
nand ( n4562 , n4515 , n352239 );
nand ( n4563 , n4561 , n4562 );
buf ( n4564 , n4563 );
xor ( n4565 , n352208 , n352222 );
and ( n4566 , n4565 , n352237 );
and ( n4567 , n352208 , n352222 );
or ( n4568 , n4566 , n4567 );
buf ( n352251 , n4568 );
buf ( n352252 , n352163 );
not ( n4571 , n352252 );
buf ( n352254 , n347604 );
not ( n4573 , n352254 );
or ( n4574 , n4571 , n4573 );
xor ( n4575 , n546 , n574 );
nand ( n4576 , n4575 , n575 );
buf ( n352259 , n4576 );
nand ( n4578 , n4574 , n352259 );
buf ( n352261 , n4578 );
buf ( n352262 , n352261 );
buf ( n352263 , n559 );
buf ( n352264 , n563 );
nand ( n4583 , n352263 , n352264 );
buf ( n352266 , n4583 );
or ( n4585 , n559 , n563 );
nand ( n4586 , n4585 , n564 );
nand ( n4587 , n352266 , n4586 , n562 );
not ( n4588 , n4587 );
buf ( n352271 , n4588 );
and ( n4590 , n352262 , n352271 );
not ( n4591 , n352262 );
buf ( n352274 , n4587 );
and ( n4593 , n4591 , n352274 );
nor ( n4594 , n4590 , n4593 );
buf ( n352277 , n4594 );
not ( n4596 , n352277 );
and ( n4597 , n352251 , n4596 );
not ( n4598 , n352251 );
and ( n4599 , n4598 , n352277 );
nor ( n4600 , n4597 , n4599 );
xor ( n4601 , n4486 , n4501 );
and ( n4602 , n4601 , n4514 );
and ( n4603 , n4486 , n4501 );
or ( n4604 , n4602 , n4603 );
xor ( n4605 , n4600 , n4604 );
not ( n4606 , n4605 );
and ( n4607 , n4564 , n4606 );
not ( n4608 , n4564 );
and ( n4609 , n4608 , n4605 );
nor ( n4610 , n4607 , n4609 );
buf ( n352293 , n352202 );
buf ( n4612 , n352293 );
buf ( n352295 , n4612 );
not ( n4614 , n352295 );
buf ( n352297 , n558 );
buf ( n352298 , n562 );
xor ( n4617 , n352297 , n352298 );
buf ( n352300 , n4617 );
not ( n4619 , n352300 );
or ( n4620 , n4614 , n4619 );
not ( n4621 , n563 );
or ( n4622 , n4621 , n564 );
not ( n4623 , n564 );
or ( n4624 , n4623 , n563 );
nand ( n4625 , n4622 , n4624 );
not ( n4626 , n4625 );
buf ( n352309 , n562 );
buf ( n352310 , n563 );
xnor ( n4629 , n352309 , n352310 );
buf ( n352312 , n4629 );
not ( n4631 , n352312 );
xor ( n4632 , n559 , n562 );
nand ( n4633 , n4626 , n4631 , n4632 );
nand ( n4634 , n4620 , n4633 );
buf ( n352317 , n4634 );
buf ( n352318 , n551 );
buf ( n352319 , n570 );
xor ( n4638 , n352318 , n352319 );
buf ( n352321 , n4638 );
buf ( n352322 , n352321 );
not ( n4641 , n352322 );
buf ( n352324 , n347344 );
not ( n4643 , n352324 );
or ( n4644 , n4641 , n4643 );
buf ( n352327 , n348473 );
buf ( n352328 , n550 );
buf ( n352329 , n570 );
xor ( n4648 , n352328 , n352329 );
buf ( n352331 , n4648 );
buf ( n352332 , n352331 );
nand ( n4651 , n352327 , n352332 );
buf ( n352334 , n4651 );
buf ( n352335 , n352334 );
nand ( n4654 , n4644 , n352335 );
buf ( n352337 , n4654 );
buf ( n352338 , n352337 );
xor ( n4657 , n352317 , n352338 );
buf ( n352340 , n352179 );
not ( n4659 , n352340 );
buf ( n352342 , n351330 );
not ( n352343 , n352342 );
or ( n4662 , n4659 , n352343 );
buf ( n352345 , n3650 );
buf ( n352346 , n556 );
buf ( n352347 , n564 );
xor ( n4666 , n352346 , n352347 );
buf ( n352349 , n4666 );
buf ( n352350 , n352349 );
nand ( n4669 , n352345 , n352350 );
buf ( n352352 , n4669 );
buf ( n352353 , n352352 );
nand ( n4672 , n4662 , n352353 );
buf ( n352355 , n4672 );
buf ( n352356 , n352355 );
xor ( n4675 , n4657 , n352356 );
buf ( n352358 , n4675 );
buf ( n352359 , n352358 );
not ( n4678 , n2579 );
xor ( n4679 , n552 , n568 );
not ( n4680 , n4679 );
or ( n4681 , n4678 , n4680 );
nand ( n4682 , n3768 , n352230 );
nand ( n4683 , n4681 , n4682 );
buf ( n352366 , n4683 );
not ( n4685 , n4533 );
not ( n4686 , n347378 );
or ( n4687 , n4685 , n4686 );
buf ( n352370 , n548 );
buf ( n352371 , n572 );
xor ( n4690 , n352370 , n352371 );
buf ( n352373 , n4690 );
nand ( n4692 , n352373 , n347382 );
nand ( n4693 , n4687 , n4692 );
buf ( n352376 , n4693 );
xor ( n4695 , n352366 , n352376 );
buf ( n352378 , n352192 );
not ( n4697 , n352378 );
buf ( n352380 , n350874 );
not ( n4699 , n352380 );
or ( n4700 , n4697 , n4699 );
buf ( n352383 , n2550 );
buf ( n352384 , n554 );
buf ( n352385 , n566 );
xor ( n4704 , n352384 , n352385 );
buf ( n352387 , n4704 );
buf ( n352388 , n352387 );
nand ( n4707 , n352383 , n352388 );
buf ( n352390 , n4707 );
buf ( n352391 , n352390 );
nand ( n4710 , n4700 , n352391 );
buf ( n352393 , n4710 );
buf ( n352394 , n352393 );
xor ( n4713 , n4695 , n352394 );
buf ( n352396 , n4713 );
buf ( n352397 , n352396 );
xor ( n4716 , n352359 , n352397 );
buf ( n352399 , n351356 );
not ( n4718 , n352399 );
buf ( n352401 , n347344 );
not ( n4720 , n352401 );
or ( n4721 , n4718 , n4720 );
buf ( n352404 , n348476 );
buf ( n352405 , n352321 );
nand ( n4724 , n352404 , n352405 );
buf ( n352407 , n4724 );
buf ( n352408 , n352407 );
nand ( n4727 , n4721 , n352408 );
buf ( n352410 , n4727 );
buf ( n352411 , n352410 );
xor ( n4730 , n351450 , n351464 );
and ( n4731 , n4730 , n351479 );
and ( n4732 , n351450 , n351464 );
or ( n4733 , n4731 , n4732 );
buf ( n352416 , n4733 );
buf ( n352417 , n352416 );
xor ( n4736 , n352411 , n352417 );
and ( n4737 , n351380 , n351394 );
buf ( n352420 , n4737 );
buf ( n352421 , n352420 );
and ( n4740 , n4736 , n352421 );
and ( n4741 , n352411 , n352417 );
or ( n4742 , n4740 , n4741 );
buf ( n352425 , n4742 );
buf ( n352426 , n352425 );
xor ( n4745 , n4716 , n352426 );
buf ( n352428 , n4745 );
and ( n4747 , n4610 , n352428 );
not ( n4748 , n4610 );
not ( n4749 , n352428 );
and ( n4750 , n4748 , n4749 );
nor ( n4751 , n4747 , n4750 );
buf ( n352434 , n4751 );
xor ( n4753 , n351400 , n351410 );
and ( n4754 , n4753 , n351485 );
and ( n4755 , n351400 , n351410 );
or ( n4756 , n4754 , n4755 );
buf ( n352439 , n4756 );
buf ( n352440 , n352439 );
xor ( n4759 , n351590 , n351596 );
and ( n4760 , n4759 , n351638 );
and ( n4761 , n351590 , n351596 );
or ( n4762 , n4760 , n4761 );
buf ( n352445 , n4762 );
buf ( n352446 , n352445 );
xor ( n4765 , n352440 , n352446 );
buf ( n352448 , n351576 );
not ( n4767 , n352448 );
buf ( n352450 , n347671 );
not ( n4769 , n352450 );
or ( n4770 , n4767 , n4769 );
buf ( n352453 , n347530 );
buf ( n352454 , n551 );
buf ( n352455 , n586 );
xor ( n4774 , n352454 , n352455 );
buf ( n352457 , n4774 );
buf ( n352458 , n352457 );
nand ( n4777 , n352453 , n352458 );
buf ( n352460 , n4777 );
buf ( n352461 , n352460 );
nand ( n4780 , n4770 , n352461 );
buf ( n352463 , n4780 );
buf ( n352464 , n352463 );
buf ( n352465 , n351539 );
buf ( n352466 , n351523 );
nand ( n352467 , n352465 , n352466 );
buf ( n352468 , n352467 );
buf ( n352469 , n352468 );
xor ( n4788 , n352464 , n352469 );
not ( n4789 , n3930 );
not ( n4790 , n4789 );
not ( n4791 , n3950 );
or ( n4792 , n4790 , n4791 );
nand ( n4793 , n4792 , n3942 );
nand ( n4794 , n3951 , n3930 );
nand ( n4795 , n4793 , n4794 );
buf ( n352478 , n4795 );
xnor ( n4797 , n4788 , n352478 );
buf ( n352480 , n4797 );
buf ( n352481 , n352480 );
xor ( n4800 , n3919 , n3923 );
and ( n4801 , n4800 , n3952 );
and ( n4802 , n3919 , n3923 );
or ( n4803 , n4801 , n4802 );
buf ( n352486 , n4803 );
xor ( n4805 , n352481 , n352486 );
buf ( n352488 , n579 );
buf ( n352489 , n580 );
xor ( n4808 , n352488 , n352489 );
buf ( n352491 , n4808 );
buf ( n352492 , n352491 );
buf ( n352493 , n559 );
and ( n4812 , n352492 , n352493 );
buf ( n352495 , n4812 );
buf ( n352496 , n352495 );
not ( n4815 , n352496 );
buf ( n352498 , n351533 );
not ( n4817 , n352498 );
buf ( n352500 , n3093 );
not ( n4819 , n352500 );
or ( n4820 , n4817 , n4819 );
buf ( n352503 , n549 );
buf ( n352504 , n588 );
xor ( n4823 , n352503 , n352504 );
buf ( n352506 , n4823 );
nand ( n4825 , n352506 , n3363 );
buf ( n352508 , n4825 );
nand ( n4827 , n4820 , n352508 );
buf ( n352510 , n4827 );
buf ( n352511 , n352510 );
not ( n4830 , n352511 );
buf ( n352513 , n4830 );
buf ( n352514 , n352513 );
not ( n4833 , n352514 );
or ( n4834 , n4815 , n4833 );
buf ( n352517 , n352510 );
buf ( n352518 , n352491 );
buf ( n352519 , n559 );
nand ( n4838 , n352518 , n352519 );
buf ( n352521 , n4838 );
buf ( n352522 , n352521 );
nand ( n4841 , n352517 , n352522 );
buf ( n352524 , n4841 );
buf ( n352525 , n352524 );
nand ( n4844 , n4834 , n352525 );
buf ( n352527 , n4844 );
buf ( n352528 , n352527 );
buf ( n352529 , n351622 );
not ( n4848 , n352529 );
buf ( n352531 , n2471 );
not ( n4850 , n352531 );
or ( n4851 , n4848 , n4850 );
buf ( n352534 , n348629 );
and ( n4853 , n553 , n584 );
not ( n4854 , n553 );
and ( n4855 , n4854 , n1771 );
nor ( n4856 , n4853 , n4855 );
buf ( n352539 , n4856 );
nand ( n4858 , n352534 , n352539 );
buf ( n352541 , n4858 );
buf ( n352542 , n352541 );
nand ( n4861 , n4851 , n352542 );
buf ( n352544 , n4861 );
buf ( n352545 , n352544 );
not ( n4864 , n352545 );
buf ( n352547 , n4864 );
buf ( n352548 , n352547 );
and ( n4867 , n352528 , n352548 );
not ( n4868 , n352528 );
buf ( n352551 , n352544 );
and ( n4870 , n4868 , n352551 );
nor ( n4871 , n4867 , n4870 );
buf ( n352554 , n4871 );
not ( n4873 , n352554 );
not ( n4874 , n4873 );
buf ( n352557 , n3928 );
not ( n4876 , n352557 );
buf ( n352559 , n347478 );
not ( n4878 , n352559 );
or ( n4879 , n4876 , n4878 );
buf ( n352562 , n547 );
buf ( n352563 , n590 );
xor ( n4882 , n352562 , n352563 );
buf ( n352565 , n4882 );
buf ( n352566 , n352565 );
buf ( n352567 , n591 );
nand ( n4886 , n352566 , n352567 );
buf ( n352569 , n4886 );
buf ( n352570 , n352569 );
nand ( n4889 , n4879 , n352570 );
buf ( n352572 , n4889 );
buf ( n352573 , n352572 );
buf ( n352574 , n351631 );
not ( n4893 , n352574 );
buf ( n352576 , n3313 );
not ( n4895 , n352576 );
or ( n4896 , n4893 , n4895 );
buf ( n352579 , n350377 );
buf ( n352580 , n555 );
buf ( n352581 , n582 );
xor ( n4900 , n352580 , n352581 );
buf ( n352583 , n4900 );
buf ( n352584 , n352583 );
nand ( n4903 , n352579 , n352584 );
buf ( n352586 , n4903 );
buf ( n352587 , n352586 );
nand ( n4906 , n4896 , n352587 );
buf ( n352589 , n4906 );
buf ( n352590 , n352589 );
xor ( n4909 , n352573 , n352590 );
buf ( n352592 , n351564 );
not ( n4911 , n352592 );
buf ( n352594 , n3870 );
not ( n4913 , n352594 );
or ( n352596 , n4911 , n4913 );
buf ( n352597 , n351038 );
buf ( n352598 , n557 );
buf ( n352599 , n580 );
xor ( n4918 , n352598 , n352599 );
buf ( n352601 , n4918 );
buf ( n352602 , n352601 );
nand ( n4921 , n352597 , n352602 );
buf ( n352604 , n4921 );
buf ( n352605 , n352604 );
nand ( n352606 , n352596 , n352605 );
buf ( n352607 , n352606 );
buf ( n352608 , n352607 );
xor ( n4927 , n4909 , n352608 );
buf ( n352610 , n4927 );
not ( n4929 , n352610 );
or ( n4930 , n4874 , n4929 );
not ( n4931 , n352610 );
nand ( n4932 , n4931 , n352554 );
nand ( n4933 , n4930 , n4932 );
buf ( n352616 , n3884 );
not ( n4935 , n352616 );
buf ( n352618 , n3897 );
nand ( n4937 , n4935 , n352618 );
buf ( n352620 , n4937 );
buf ( n352621 , n352620 );
not ( n4940 , n352621 );
buf ( n352623 , n3856 );
not ( n4942 , n352623 );
or ( n4943 , n4940 , n4942 );
buf ( n352626 , n3896 );
buf ( n352627 , n3884 );
nand ( n4946 , n352626 , n352627 );
buf ( n352629 , n4946 );
buf ( n352630 , n352629 );
nand ( n352631 , n4943 , n352630 );
buf ( n352632 , n352631 );
not ( n4951 , n352632 );
and ( n4952 , n4933 , n4951 );
not ( n4953 , n4933 );
and ( n4954 , n4953 , n352632 );
nor ( n4955 , n4952 , n4954 );
buf ( n352638 , n4955 );
xor ( n4957 , n4805 , n352638 );
buf ( n352640 , n4957 );
buf ( n352641 , n352640 );
and ( n4960 , n4765 , n352641 );
and ( n4961 , n352440 , n352446 );
or ( n4962 , n4960 , n4961 );
buf ( n352645 , n4962 );
buf ( n352646 , n352645 );
xor ( n4965 , n352434 , n352646 );
xor ( n4966 , n351426 , n351437 );
and ( n4967 , n4966 , n351482 );
and ( n4968 , n351426 , n351437 );
or ( n4969 , n4967 , n4968 );
buf ( n352652 , n4969 );
not ( n4971 , n352652 );
xor ( n4972 , n352411 , n352417 );
xor ( n4973 , n4972 , n352421 );
buf ( n352656 , n4973 );
not ( n4975 , n352656 );
nand ( n4976 , n4971 , n4975 );
not ( n4977 , n4976 );
buf ( n4978 , n352158 );
not ( n4979 , n4978 );
not ( n4980 , n4516 );
not ( n4981 , n352239 );
and ( n4982 , n4980 , n4981 );
and ( n4983 , n4516 , n352239 );
nor ( n4984 , n4982 , n4983 );
not ( n4985 , n4984 );
or ( n4986 , n4979 , n4985 );
or ( n4987 , n4984 , n4978 );
nand ( n4988 , n4986 , n4987 );
not ( n4989 , n4988 );
or ( n4990 , n4977 , n4989 );
nand ( n4991 , n352656 , n352652 );
nand ( n4992 , n4990 , n4991 );
buf ( n352675 , n4992 );
xor ( n4994 , n352481 , n352486 );
and ( n4995 , n4994 , n352638 );
and ( n4996 , n352481 , n352486 );
or ( n4997 , n4995 , n4996 );
buf ( n352680 , n4997 );
buf ( n352681 , n352680 );
xor ( n5000 , n352675 , n352681 );
buf ( n352683 , n352554 );
not ( n5002 , n352683 );
buf ( n352685 , n4931 );
not ( n5004 , n352685 );
or ( n5005 , n5002 , n5004 );
buf ( n352688 , n352632 );
nand ( n5007 , n5005 , n352688 );
buf ( n352690 , n5007 );
buf ( n352691 , n352690 );
buf ( n352692 , n352554 );
not ( n5011 , n352692 );
buf ( n352694 , n352610 );
nand ( n5013 , n5011 , n352694 );
buf ( n352696 , n5013 );
buf ( n352697 , n352696 );
nand ( n5016 , n352691 , n352697 );
buf ( n352699 , n5016 );
buf ( n352700 , n352699 );
buf ( n352701 , n352521 );
not ( n5020 , n352701 );
buf ( n352703 , n352513 );
not ( n5022 , n352703 );
or ( n5023 , n5020 , n5022 );
buf ( n352706 , n352544 );
nand ( n5025 , n5023 , n352706 );
buf ( n352708 , n5025 );
buf ( n352709 , n352708 );
buf ( n352710 , n352513 );
not ( n5029 , n352710 );
buf ( n352712 , n352495 );
nand ( n5031 , n5029 , n352712 );
buf ( n352714 , n5031 );
buf ( n352715 , n352714 );
nand ( n5034 , n352709 , n352715 );
buf ( n352717 , n5034 );
buf ( n352718 , n559 );
buf ( n352719 , n579 );
or ( n5038 , n352718 , n352719 );
buf ( n352721 , n580 );
nand ( n5040 , n5038 , n352721 );
buf ( n352723 , n5040 );
buf ( n352724 , n559 );
buf ( n352725 , n579 );
nand ( n5044 , n352724 , n352725 );
buf ( n352727 , n5044 );
and ( n5046 , n352723 , n352727 , n578 );
buf ( n352729 , n352565 );
not ( n5048 , n352729 );
buf ( n352731 , n347478 );
not ( n5050 , n352731 );
or ( n5051 , n5048 , n5050 );
buf ( n352734 , n546 );
buf ( n352735 , n590 );
xor ( n5054 , n352734 , n352735 );
buf ( n352737 , n5054 );
buf ( n352738 , n352737 );
buf ( n352739 , n591 );
nand ( n5058 , n352738 , n352739 );
buf ( n352741 , n5058 );
buf ( n352742 , n352741 );
nand ( n5061 , n5051 , n352742 );
buf ( n352744 , n5061 );
xor ( n5063 , n5046 , n352744 );
buf ( n5064 , n5063 );
xor ( n5065 , n352573 , n352590 );
and ( n5066 , n5065 , n352608 );
and ( n5067 , n352573 , n352590 );
or ( n5068 , n5066 , n5067 );
buf ( n352751 , n5068 );
nand ( n5070 , n352717 , n5064 , n352751 );
buf ( n352753 , n352708 );
buf ( n352754 , n352714 );
nand ( n5073 , n352753 , n352754 );
buf ( n352756 , n5073 );
nor ( n5075 , n352756 , n5064 );
nand ( n5076 , n5075 , n352751 );
not ( n5077 , n352717 );
not ( n5078 , n352751 );
nand ( n5079 , n5077 , n5078 , n5064 );
not ( n5080 , n5064 );
nand ( n5081 , n5080 , n5078 , n352717 );
nand ( n5082 , n5070 , n5076 , n5079 , n5081 );
buf ( n352765 , n5082 );
xor ( n5084 , n352700 , n352765 );
not ( n5085 , n352506 );
not ( n5086 , n3093 );
or ( n5087 , n5085 , n5086 );
buf ( n352770 , n548 );
buf ( n352771 , n588 );
xor ( n5090 , n352770 , n352771 );
buf ( n352773 , n5090 );
nand ( n5092 , n3363 , n352773 );
nand ( n5093 , n5087 , n5092 );
not ( n5094 , n348611 );
buf ( n352777 , n552 );
buf ( n352778 , n584 );
xor ( n5097 , n352777 , n352778 );
buf ( n352780 , n5097 );
not ( n5099 , n352780 );
or ( n5100 , n5094 , n5099 );
nand ( n5101 , n2469 , n348614 , n4856 );
nand ( n5102 , n5100 , n5101 );
not ( n5103 , n5102 );
xor ( n5104 , n5093 , n5103 );
not ( n5105 , n352583 );
not ( n5106 , n3313 );
or ( n5107 , n5105 , n5106 );
buf ( n352790 , n350705 );
buf ( n352791 , n554 );
buf ( n352792 , n582 );
xor ( n5111 , n352791 , n352792 );
buf ( n352794 , n5111 );
buf ( n352795 , n352794 );
nand ( n5114 , n352790 , n352795 );
buf ( n352797 , n5114 );
nand ( n5116 , n5107 , n352797 );
xor ( n5117 , n5104 , n5116 );
not ( n5118 , n350110 );
not ( n5119 , n352457 );
or ( n5120 , n5118 , n5119 );
and ( n5121 , n586 , n550 );
not ( n5122 , n586 );
not ( n5123 , n550 );
and ( n5124 , n5122 , n5123 );
nor ( n5125 , n5121 , n5124 );
nand ( n5126 , n5125 , n347530 );
nand ( n5127 , n5120 , n5126 );
buf ( n352810 , n5127 );
buf ( n352811 , n352601 );
not ( n5130 , n352811 );
buf ( n352813 , n3870 );
not ( n5132 , n352813 );
or ( n5133 , n5130 , n5132 );
buf ( n352816 , n351038 );
buf ( n352817 , n556 );
buf ( n352818 , n580 );
xor ( n5137 , n352817 , n352818 );
buf ( n352820 , n5137 );
buf ( n352821 , n352820 );
nand ( n5140 , n352816 , n352821 );
buf ( n352823 , n5140 );
buf ( n352824 , n352823 );
nand ( n5143 , n5133 , n352824 );
buf ( n352826 , n5143 );
buf ( n352827 , n352826 );
xor ( n5146 , n352810 , n352827 );
buf ( n352829 , n559 );
buf ( n352830 , n578 );
xor ( n5149 , n352829 , n352830 );
buf ( n352832 , n5149 );
buf ( n352833 , n352832 );
not ( n5152 , n352833 );
and ( n5153 , n579 , n580 );
not ( n5154 , n579 );
and ( n5155 , n5154 , n3866 );
nor ( n5156 , n5153 , n5155 );
not ( n5157 , n578 );
and ( n5158 , n579 , n5157 );
not ( n5159 , n579 );
and ( n5160 , n5159 , n578 );
nor ( n5161 , n5158 , n5160 );
nor ( n5162 , n5156 , n5161 );
buf ( n352845 , n5162 );
not ( n5164 , n352845 );
or ( n5165 , n5152 , n5164 );
buf ( n352848 , n352491 );
buf ( n352849 , n558 );
buf ( n352850 , n578 );
xor ( n5169 , n352849 , n352850 );
buf ( n352852 , n5169 );
buf ( n352853 , n352852 );
nand ( n5172 , n352848 , n352853 );
buf ( n352855 , n5172 );
buf ( n352856 , n352855 );
nand ( n5175 , n5165 , n352856 );
buf ( n352858 , n5175 );
buf ( n352859 , n352858 );
xor ( n5178 , n5146 , n352859 );
buf ( n352861 , n5178 );
xnor ( n5180 , n5117 , n352861 );
buf ( n352863 , n352463 );
not ( n5182 , n352863 );
buf ( n352865 , n352468 );
not ( n5184 , n352865 );
buf ( n352867 , n5184 );
buf ( n352868 , n352867 );
not ( n5187 , n352868 );
or ( n5188 , n5182 , n5187 );
buf ( n352871 , n352463 );
not ( n5190 , n352871 );
buf ( n352873 , n5190 );
buf ( n352874 , n352873 );
not ( n5193 , n352874 );
buf ( n352876 , n352468 );
not ( n5195 , n352876 );
or ( n5196 , n5193 , n5195 );
buf ( n352879 , n4795 );
nand ( n5198 , n5196 , n352879 );
buf ( n352881 , n5198 );
buf ( n352882 , n352881 );
nand ( n5201 , n5188 , n352882 );
buf ( n352884 , n5201 );
xor ( n5203 , n5180 , n352884 );
buf ( n352886 , n5203 );
xor ( n5205 , n5084 , n352886 );
buf ( n352888 , n5205 );
buf ( n352889 , n352888 );
xor ( n5208 , n5000 , n352889 );
buf ( n352891 , n5208 );
buf ( n352892 , n352891 );
xor ( n5211 , n4965 , n352892 );
buf ( n352894 , n5211 );
not ( n5213 , n4988 );
nand ( n5214 , n4991 , n4976 );
not ( n5215 , n5214 );
or ( n5216 , n5213 , n5215 );
not ( n5217 , n4988 );
xor ( n5218 , n352652 , n352656 );
nand ( n5219 , n5217 , n5218 );
nand ( n5220 , n5216 , n5219 );
buf ( n352903 , n5220 );
xor ( n5222 , n351501 , n351507 );
and ( n5223 , n5222 , n351641 );
and ( n5224 , n351501 , n351507 );
or ( n5225 , n5223 , n5224 );
buf ( n352908 , n5225 );
buf ( n352909 , n352908 );
xor ( n5228 , n352903 , n352909 );
xor ( n5229 , n352440 , n352446 );
xor ( n5230 , n5229 , n352641 );
buf ( n352913 , n5230 );
buf ( n352914 , n352913 );
and ( n5233 , n5228 , n352914 );
and ( n5234 , n352903 , n352909 );
or ( n5235 , n5233 , n5234 );
buf ( n352918 , n5235 );
nor ( n5237 , n352894 , n352918 );
xor ( n5238 , n352903 , n352909 );
xor ( n5239 , n5238 , n352914 );
buf ( n352922 , n5239 );
xor ( n5241 , n351488 , n351494 );
and ( n5242 , n5241 , n351644 );
and ( n5243 , n351488 , n351494 );
or ( n5244 , n5242 , n5243 );
buf ( n352927 , n5244 );
nand ( n5246 , n352922 , n352927 );
or ( n5247 , n5237 , n5246 );
nand ( n5248 , n352894 , n352918 );
nand ( n5249 , n5247 , n5248 );
buf ( n352932 , n5249 );
not ( n5251 , n352932 );
nand ( n5252 , n3417 , n3974 , n3138 );
not ( n5253 , n5252 );
buf ( n352936 , n5253 );
not ( n5255 , n352894 );
not ( n5256 , n352918 );
and ( n5257 , n5255 , n5256 );
not ( n5258 , n352922 );
not ( n5259 , n352927 );
and ( n5260 , n5258 , n5259 );
nor ( n5261 , n5257 , n5260 );
buf ( n352944 , n5261 );
buf ( n5263 , n352944 );
buf ( n352946 , n5263 );
buf ( n352947 , n352946 );
buf ( n5266 , n2548 );
buf ( n352949 , n5266 );
nand ( n5268 , n352936 , n352947 , n352949 );
buf ( n352951 , n5268 );
buf ( n352952 , n352951 );
not ( n5271 , n350841 );
not ( n5272 , n351646 );
not ( n5273 , n351654 );
and ( n5274 , n5272 , n5273 );
nor ( n5275 , n5274 , n351303 );
not ( n5276 , n5275 );
or ( n5277 , n5271 , n5276 );
nor ( n5278 , n351100 , n351103 );
and ( n5279 , n5278 , n3974 );
nor ( n5280 , n5279 , n3977 );
nand ( n5281 , n5277 , n5280 );
not ( n5282 , n5281 );
not ( n5283 , n5282 );
nand ( n5284 , n352946 , n5283 );
buf ( n352967 , n5284 );
nand ( n5286 , n5251 , n352952 , n352967 );
buf ( n352969 , n5286 );
buf ( n352970 , n352969 );
buf ( n352971 , n352300 );
not ( n5290 , n352971 );
nor ( n5291 , n352312 , n4625 );
buf ( n352974 , n5291 );
not ( n5293 , n352974 );
or ( n5294 , n5290 , n5293 );
buf ( n352977 , n352295 );
buf ( n352978 , n557 );
buf ( n352979 , n562 );
xor ( n5298 , n352978 , n352979 );
buf ( n352981 , n5298 );
buf ( n352982 , n352981 );
nand ( n5301 , n352977 , n352982 );
buf ( n352984 , n5301 );
buf ( n352985 , n352984 );
nand ( n5304 , n5294 , n352985 );
buf ( n352987 , n5304 );
buf ( n352988 , n352987 );
buf ( n352989 , n352349 );
not ( n5308 , n352989 );
buf ( n352991 , n351330 );
not ( n5310 , n352991 );
or ( n5311 , n5308 , n5310 );
buf ( n352994 , n3650 );
buf ( n352995 , n555 );
buf ( n352996 , n564 );
xor ( n5315 , n352995 , n352996 );
buf ( n352998 , n5315 );
buf ( n352999 , n352998 );
nand ( n5318 , n352994 , n352999 );
buf ( n353001 , n5318 );
buf ( n353002 , n353001 );
nand ( n5321 , n5311 , n353002 );
buf ( n353004 , n5321 );
buf ( n353005 , n353004 );
xor ( n5324 , n352988 , n353005 );
buf ( n353007 , n352261 );
buf ( n353008 , n4588 );
and ( n5327 , n353007 , n353008 );
buf ( n353010 , n5327 );
buf ( n353011 , n353010 );
xor ( n5330 , n5324 , n353011 );
buf ( n353013 , n5330 );
not ( n5332 , n353013 );
xor ( n5333 , n568 , n551 );
not ( n5334 , n5333 );
not ( n5335 , n2579 );
or ( n5336 , n5334 , n5335 );
nand ( n5337 , n2232 , n2234 );
nand ( n5338 , n2230 , n4679 , n5337 );
nand ( n5339 , n5336 , n5338 );
not ( n5340 , n352331 );
not ( n5341 , n347344 );
or ( n5342 , n5340 , n5341 );
buf ( n353025 , n347350 );
buf ( n353026 , n549 );
buf ( n353027 , n570 );
xor ( n5346 , n353026 , n353027 );
buf ( n353029 , n5346 );
buf ( n353030 , n353029 );
nand ( n5349 , n353025 , n353030 );
buf ( n353032 , n5349 );
nand ( n5351 , n5342 , n353032 );
xor ( n5352 , n5339 , n5351 );
not ( n5353 , n352387 );
not ( n5354 , n2851 );
or ( n5355 , n5353 , n5354 );
buf ( n353038 , n2550 );
buf ( n353039 , n553 );
buf ( n353040 , n566 );
xor ( n5359 , n353039 , n353040 );
buf ( n353042 , n5359 );
buf ( n353043 , n353042 );
nand ( n5362 , n353038 , n353043 );
buf ( n353045 , n5362 );
nand ( n5364 , n5355 , n353045 );
xnor ( n5365 , n5352 , n5364 );
not ( n5366 , n5365 );
or ( n5367 , n5332 , n5366 );
not ( n5368 , n353013 );
not ( n5369 , n5365 );
nand ( n5370 , n5368 , n5369 );
nand ( n5371 , n5367 , n5370 );
not ( n5372 , n352251 );
not ( n5373 , n352277 );
or ( n5374 , n5372 , n5373 );
buf ( n353057 , n352251 );
buf ( n353058 , n352277 );
or ( n5377 , n353057 , n353058 );
buf ( n353060 , n4604 );
nand ( n5379 , n5377 , n353060 );
buf ( n353062 , n5379 );
nand ( n5381 , n5374 , n353062 );
and ( n5382 , n5371 , n5381 );
not ( n5383 , n5371 );
not ( n5384 , n5381 );
and ( n5385 , n5383 , n5384 );
nor ( n5386 , n5382 , n5385 );
buf ( n353069 , n5386 );
xor ( n5388 , n352366 , n352376 );
and ( n5389 , n5388 , n352394 );
and ( n5390 , n352366 , n352376 );
or ( n5391 , n5389 , n5390 );
buf ( n353074 , n5391 );
buf ( n353075 , n353074 );
not ( n5394 , n353075 );
buf ( n353077 , n5394 );
buf ( n353078 , n353077 );
not ( n5397 , n347399 );
not ( n5398 , n4575 );
or ( n5399 , n5397 , n5398 );
and ( n5400 , n574 , n545 );
not ( n5401 , n574 );
not ( n5402 , n545 );
and ( n5403 , n5401 , n5402 );
nor ( n5404 , n5400 , n5403 );
nand ( n5405 , n5404 , n575 );
nand ( n5406 , n5399 , n5405 );
xor ( n5407 , n561 , n562 );
buf ( n353090 , n5407 );
buf ( n353091 , n559 );
nand ( n5410 , n353090 , n353091 );
buf ( n353093 , n5410 );
xor ( n5412 , n5406 , n353093 );
buf ( n353095 , n352373 );
not ( n5414 , n353095 );
buf ( n353097 , n347378 );
not ( n5416 , n353097 );
or ( n5417 , n5414 , n5416 );
buf ( n353100 , n347382 );
buf ( n353101 , n547 );
buf ( n353102 , n572 );
xor ( n5421 , n353101 , n353102 );
buf ( n353104 , n5421 );
buf ( n353105 , n353104 );
nand ( n5424 , n353100 , n353105 );
buf ( n353107 , n5424 );
buf ( n353108 , n353107 );
nand ( n5427 , n5417 , n353108 );
buf ( n353110 , n5427 );
xor ( n5429 , n5412 , n353110 );
buf ( n353112 , n5429 );
and ( n5431 , n353078 , n353112 );
not ( n5432 , n353078 );
buf ( n353115 , n5429 );
not ( n5434 , n353115 );
buf ( n353117 , n5434 );
buf ( n353118 , n353117 );
and ( n5437 , n5432 , n353118 );
nor ( n5438 , n5431 , n5437 );
buf ( n353121 , n5438 );
buf ( n353122 , n353121 );
xor ( n5441 , n352317 , n352338 );
and ( n5442 , n5441 , n352356 );
and ( n5443 , n352317 , n352338 );
or ( n5444 , n5442 , n5443 );
buf ( n353127 , n5444 );
buf ( n353128 , n353127 );
and ( n5447 , n353122 , n353128 );
not ( n5448 , n353122 );
buf ( n353131 , n353127 );
not ( n5450 , n353131 );
buf ( n353133 , n5450 );
buf ( n353134 , n353133 );
and ( n5453 , n5448 , n353134 );
nor ( n5454 , n5447 , n5453 );
buf ( n353137 , n5454 );
buf ( n353138 , n353137 );
and ( n5457 , n353069 , n353138 );
not ( n5458 , n353069 );
buf ( n353141 , n353137 );
not ( n5460 , n353141 );
buf ( n353143 , n5460 );
buf ( n353144 , n353143 );
and ( n5463 , n5458 , n353144 );
nor ( n5464 , n5457 , n5463 );
buf ( n353147 , n5464 );
xor ( n5466 , n352359 , n352397 );
and ( n5467 , n5466 , n352426 );
and ( n5468 , n352359 , n352397 );
or ( n5469 , n5467 , n5468 );
buf ( n353152 , n5469 );
xor ( n5471 , n353147 , n353152 );
buf ( n353154 , n5471 );
xor ( n5473 , n352675 , n352681 );
and ( n5474 , n5473 , n352889 );
and ( n5475 , n352675 , n352681 );
or ( n5476 , n5474 , n5475 );
buf ( n353159 , n5476 );
buf ( n353160 , n353159 );
xor ( n5479 , n353154 , n353160 );
not ( n5480 , n4563 );
nand ( n5481 , n5480 , n4605 );
not ( n5482 , n5481 );
not ( n5483 , n352428 );
or ( n5484 , n5482 , n5483 );
nand ( n5485 , n4564 , n4606 );
nand ( n5486 , n5484 , n5485 );
xor ( n5487 , n352700 , n352765 );
and ( n5488 , n5487 , n352886 );
and ( n5489 , n352700 , n352765 );
or ( n5490 , n5488 , n5489 );
buf ( n353173 , n5490 );
xor ( n5492 , n5486 , n353173 );
buf ( n353175 , n352861 );
not ( n5494 , n353175 );
buf ( n353177 , n5494 );
nand ( n5496 , n353177 , n5117 );
nand ( n5497 , n5496 , n352884 );
buf ( n353180 , n5497 );
buf ( n353181 , n5117 );
not ( n5500 , n353181 );
buf ( n353183 , n352861 );
nand ( n5502 , n5500 , n353183 );
buf ( n353185 , n5502 );
buf ( n353186 , n353185 );
nand ( n5505 , n353180 , n353186 );
buf ( n353188 , n5505 );
buf ( n353189 , n353188 );
buf ( n353190 , n577 );
buf ( n353191 , n578 );
xor ( n5510 , n353190 , n353191 );
buf ( n353193 , n5510 );
buf ( n353194 , n353193 );
buf ( n353195 , n559 );
and ( n5514 , n353194 , n353195 );
buf ( n353197 , n5514 );
buf ( n353198 , n353197 );
not ( n5517 , n591 );
buf ( n353200 , n545 );
buf ( n353201 , n590 );
xor ( n5520 , n353200 , n353201 );
buf ( n353203 , n5520 );
not ( n5522 , n353203 );
or ( n5523 , n5517 , n5522 );
nand ( n5524 , n352737 , n347478 );
nand ( n5525 , n5523 , n5524 );
buf ( n353208 , n5525 );
xor ( n5527 , n353198 , n353208 );
buf ( n353210 , n352773 );
not ( n5529 , n353210 );
buf ( n353212 , n3093 );
not ( n5531 , n353212 );
or ( n5532 , n5529 , n5531 );
buf ( n353215 , n547 );
buf ( n353216 , n588 );
xor ( n5535 , n353215 , n353216 );
buf ( n353218 , n5535 );
nand ( n5537 , n353218 , n3363 );
buf ( n353220 , n5537 );
nand ( n5539 , n5532 , n353220 );
buf ( n353222 , n5539 );
buf ( n353223 , n353222 );
xor ( n5542 , n5527 , n353223 );
buf ( n353225 , n5542 );
buf ( n353226 , n353225 );
nor ( n5545 , n5116 , n5093 );
or ( n5546 , n5545 , n5103 );
nand ( n5547 , n5116 , n5093 );
nand ( n5548 , n5546 , n5547 );
buf ( n353231 , n5548 );
xor ( n5550 , n353226 , n353231 );
xor ( n5551 , n352810 , n352827 );
and ( n5552 , n5551 , n352859 );
and ( n5553 , n352810 , n352827 );
or ( n5554 , n5552 , n5553 );
buf ( n353237 , n5554 );
buf ( n353238 , n353237 );
xor ( n5557 , n5550 , n353238 );
buf ( n353240 , n5557 );
buf ( n353241 , n353240 );
xor ( n5560 , n353189 , n353241 );
not ( n5561 , n352751 );
not ( n5562 , n5075 );
not ( n5563 , n5562 );
or ( n5564 , n5561 , n5563 );
nand ( n5565 , n352756 , n5064 );
nand ( n5566 , n5564 , n5565 );
not ( n5567 , n5566 );
buf ( n353250 , n352780 );
not ( n5569 , n353250 );
and ( n5570 , n2469 , n348614 );
buf ( n353253 , n5570 );
not ( n5572 , n353253 );
or ( n5573 , n5569 , n5572 );
buf ( n353256 , n348617 );
buf ( n353257 , n551 );
buf ( n353258 , n584 );
xor ( n5577 , n353257 , n353258 );
buf ( n353260 , n5577 );
buf ( n353261 , n353260 );
nand ( n5580 , n353256 , n353261 );
buf ( n353263 , n5580 );
buf ( n353264 , n353263 );
nand ( n5583 , n5573 , n353264 );
buf ( n353266 , n5583 );
buf ( n353267 , n352794 );
not ( n5586 , n353267 );
buf ( n353269 , n3313 );
not ( n5588 , n353269 );
or ( n5589 , n5586 , n5588 );
buf ( n353272 , n350705 );
buf ( n353273 , n553 );
buf ( n353274 , n582 );
xor ( n5593 , n353273 , n353274 );
buf ( n353276 , n5593 );
buf ( n353277 , n353276 );
nand ( n5596 , n353272 , n353277 );
buf ( n353279 , n5596 );
buf ( n353280 , n353279 );
nand ( n5599 , n5589 , n353280 );
buf ( n353282 , n5599 );
buf ( n353283 , n353282 );
not ( n5602 , n353283 );
buf ( n353285 , n5602 );
and ( n5604 , n353266 , n353285 );
not ( n5605 , n353266 );
and ( n5606 , n5605 , n353282 );
or ( n5607 , n5604 , n5606 );
not ( n5608 , n347530 );
buf ( n353291 , n549 );
buf ( n353292 , n586 );
xor ( n5611 , n353291 , n353292 );
buf ( n353294 , n5611 );
not ( n5613 , n353294 );
or ( n5614 , n5608 , n5613 );
nand ( n5615 , n347669 , n347664 , n5125 );
nand ( n5616 , n5614 , n5615 );
not ( n5617 , n5616 );
and ( n5618 , n5607 , n5617 );
not ( n5619 , n5607 );
and ( n5620 , n5619 , n5616 );
or ( n5621 , n5618 , n5620 );
buf ( n353304 , n352852 );
not ( n5623 , n353304 );
buf ( n353306 , n5162 );
not ( n5625 , n353306 );
or ( n5626 , n5623 , n5625 );
buf ( n353309 , n352491 );
buf ( n353310 , n557 );
buf ( n353311 , n578 );
xor ( n5630 , n353310 , n353311 );
buf ( n353313 , n5630 );
buf ( n353314 , n353313 );
nand ( n5633 , n353309 , n353314 );
buf ( n353316 , n5633 );
buf ( n353317 , n353316 );
nand ( n5636 , n5626 , n353317 );
buf ( n353319 , n5636 );
buf ( n353320 , n352744 );
buf ( n353321 , n5046 );
and ( n5640 , n353320 , n353321 );
buf ( n353323 , n5640 );
and ( n5642 , n353319 , n353323 );
not ( n5643 , n353319 );
not ( n5644 , n353323 );
and ( n5645 , n5643 , n5644 );
or ( n5646 , n5642 , n5645 );
buf ( n353329 , n352820 );
not ( n5648 , n353329 );
buf ( n353331 , n3870 );
not ( n5650 , n353331 );
or ( n5651 , n5648 , n5650 );
not ( n5652 , n580 );
not ( n5653 , n347525 );
or ( n5654 , n5652 , n5653 );
not ( n5655 , n580 );
nand ( n5656 , n5655 , n555 );
nand ( n5657 , n5654 , n5656 );
nand ( n5658 , n5657 , n351559 );
buf ( n353341 , n5658 );
nand ( n5660 , n5651 , n353341 );
buf ( n353343 , n5660 );
not ( n5662 , n353343 );
and ( n5663 , n5646 , n5662 );
not ( n5664 , n5646 );
and ( n5665 , n5664 , n353343 );
nor ( n5666 , n5663 , n5665 );
not ( n5667 , n5666 );
and ( n5668 , n5621 , n5667 );
not ( n5669 , n5621 );
and ( n5670 , n5669 , n5666 );
nor ( n5671 , n5668 , n5670 );
not ( n5672 , n5671 );
or ( n5673 , n5567 , n5672 );
or ( n5674 , n5566 , n5671 );
nand ( n5675 , n5673 , n5674 );
buf ( n353358 , n5675 );
xor ( n5677 , n5560 , n353358 );
buf ( n353360 , n5677 );
xor ( n5679 , n5492 , n353360 );
buf ( n353362 , n5679 );
xor ( n5681 , n5479 , n353362 );
buf ( n353364 , n5681 );
buf ( n353365 , n353364 );
xor ( n5684 , n352434 , n352646 );
and ( n5685 , n5684 , n352892 );
and ( n5686 , n352434 , n352646 );
or ( n5687 , n5685 , n5686 );
buf ( n353370 , n5687 );
buf ( n353371 , n353370 );
nor ( n5690 , n353365 , n353371 );
buf ( n353373 , n5690 );
buf ( n353374 , n353373 );
not ( n5693 , n353374 );
buf ( n353376 , n5693 );
buf ( n353377 , n353376 );
buf ( n353378 , n353364 );
buf ( n353379 , n353370 );
nand ( n5698 , n353378 , n353379 );
buf ( n353381 , n5698 );
buf ( n353382 , n353381 );
buf ( n5701 , n353382 );
buf ( n353384 , n5701 );
buf ( n353385 , n353384 );
nand ( n5704 , n353377 , n353385 );
buf ( n353387 , n5704 );
buf ( n353388 , n353387 );
not ( n5707 , n353388 );
buf ( n353390 , n5707 );
buf ( n353391 , n353390 );
and ( n5710 , n352970 , n353391 );
not ( n5711 , n352970 );
buf ( n353394 , n353387 );
and ( n5713 , n5711 , n353394 );
nor ( n5714 , n5710 , n5713 );
buf ( n353397 , n5714 );
not ( n5716 , n353397 );
not ( n5717 , n1022 );
not ( n5718 , n5717 );
not ( n5719 , n5718 );
buf ( n5720 , n1974 );
and ( n5721 , n5720 , n348175 );
not ( n5722 , n5720 );
and ( n5723 , n5722 , n554 );
or ( n5724 , n5721 , n5723 );
not ( n5725 , n5724 );
or ( n5726 , n5719 , n5725 );
not ( n5727 , n554 );
not ( n5728 , n2072 );
or ( n5729 , n5727 , n5728 );
not ( n5730 , n2072 );
nand ( n5731 , n5730 , n348175 );
nand ( n5732 , n5729 , n5731 );
nand ( n5733 , n5732 , n1925 );
nand ( n5734 , n5726 , n5733 );
not ( n5735 , n2020 );
not ( n5736 , n5735 );
not ( n5737 , n548 );
not ( n5738 , n348115 );
or ( n5739 , n5737 , n5738 );
nand ( n5740 , n348118 , n351773 );
nand ( n5741 , n5739 , n5740 );
not ( n5742 , n5741 );
or ( n5743 , n5736 , n5742 );
not ( n5744 , n348332 );
not ( n5745 , n5744 );
not ( n5746 , n351773 );
or ( n5747 , n5745 , n5746 );
nand ( n5748 , n548 , n348146 );
nand ( n5749 , n5747 , n5748 );
nor ( n5750 , n4099 , n4103 );
buf ( n5751 , n5750 );
nand ( n5752 , n5749 , n5751 );
nand ( n5753 , n5743 , n5752 );
buf ( n5754 , n348348 );
not ( n5755 , n5754 );
not ( n5756 , n5755 );
xor ( n5757 , n547 , n548 );
and ( n5758 , n5757 , n546 );
not ( n5759 , n5758 );
or ( n5760 , n5756 , n5759 );
not ( n5761 , n546 );
nand ( n5762 , n348285 , n5757 , n5761 );
not ( n5763 , n546 );
nand ( n5764 , n5763 , n548 , n547 );
not ( n5765 , n5764 );
and ( n5766 , n348158 , n5765 );
not ( n5767 , n348158 );
not ( n5768 , n546 );
nor ( n5769 , n5768 , n548 , n547 );
and ( n5770 , n5767 , n5769 );
nor ( n5771 , n5766 , n5770 );
and ( n5772 , n5762 , n5771 );
nand ( n5773 , n5760 , n5772 );
or ( n5774 , n547 , n548 );
not ( n5775 , n5774 );
not ( n5776 , n348158 );
or ( n5777 , n5775 , n5776 );
nand ( n5778 , n547 , n548 );
and ( n5779 , n5778 , n546 );
nand ( n5780 , n5777 , n5779 );
not ( n5781 , n5780 );
and ( n5782 , n5773 , n5781 );
not ( n353465 , n5773 );
and ( n353466 , n353465 , n5780 );
nor ( n5785 , n5782 , n353466 );
xor ( n5786 , n5753 , n5785 );
not ( n5787 , n1875 );
not ( n353470 , n550 );
not ( n353471 , n1751 );
or ( n5790 , n353470 , n353471 );
nand ( n353473 , n348266 , n1880 );
nand ( n353474 , n5790 , n353473 );
not ( n5793 , n353474 );
or ( n5794 , n5787 , n5793 );
not ( n5795 , n550 );
not ( n353478 , n966 );
or ( n353479 , n5795 , n353478 );
nand ( n5798 , n348226 , n1880 );
nand ( n353481 , n353479 , n5798 );
nand ( n353482 , n353481 , n4078 );
nand ( n5801 , n5794 , n353482 );
and ( n5802 , n5786 , n5801 );
and ( n5803 , n5753 , n5785 );
or ( n353486 , n5802 , n5803 );
xor ( n353487 , n5734 , n353486 );
not ( n5806 , n5735 );
and ( n353489 , n348226 , n351773 );
not ( n353490 , n348226 );
and ( n5809 , n353490 , n548 );
or ( n5810 , n353489 , n5809 );
not ( n5811 , n5810 );
or ( n353494 , n5806 , n5811 );
nand ( n353495 , n5741 , n5751 );
nand ( n5814 , n353494 , n353495 );
not ( n353497 , n4078 );
not ( n353498 , n353474 );
or ( n5817 , n353497 , n353498 );
and ( n5818 , n997 , n550 );
not ( n5819 , n997 );
and ( n353502 , n5819 , n1880 );
nor ( n353503 , n5818 , n353502 );
nand ( n5822 , n353503 , n1875 );
nand ( n353505 , n5817 , n5822 );
xor ( n353506 , n5814 , n353505 );
not ( n5825 , n1011 );
not ( n5826 , n552 );
not ( n5827 , n1843 );
not ( n353510 , n5827 );
or ( n353511 , n5826 , n353510 );
not ( n5830 , n552 );
nand ( n353513 , n5830 , n1843 );
nand ( n353514 , n353511 , n353513 );
not ( n5833 , n353514 );
or ( n5834 , n5825 , n5833 );
and ( n5835 , n552 , n1789 );
not ( n353518 , n552 );
and ( n353519 , n353518 , n1788 );
or ( n5838 , n5835 , n353519 );
not ( n353521 , n5838 );
not ( n353522 , n1871 );
or ( n5841 , n353521 , n353522 );
nand ( n5842 , n5834 , n5841 );
xor ( n5843 , n353506 , n5842 );
xor ( n353526 , n353487 , n5843 );
not ( n353527 , n1875 );
not ( n5846 , n353481 );
or ( n353529 , n353527 , n5846 );
nand ( n353530 , n351757 , n4078 );
nand ( n5849 , n353529 , n353530 );
not ( n5850 , n1022 );
not ( n5851 , n4001 );
or ( n353534 , n5850 , n5851 );
not ( n353535 , n554 );
not ( n5854 , n5827 );
or ( n353537 , n353535 , n5854 );
nand ( n353538 , n1843 , n348175 );
nand ( n5857 , n353537 , n353538 );
nand ( n5858 , n5857 , n1925 );
nand ( n5859 , n353534 , n5858 );
xor ( n353542 , n5849 , n5859 );
not ( n353543 , n1871 );
not ( n5862 , n4116 );
or ( n353545 , n353543 , n5862 );
not ( n353546 , n552 );
not ( n5865 , n348746 );
or ( n5866 , n353546 , n5865 );
not ( n5867 , n552 );
nand ( n353550 , n5867 , n2005 );
nand ( n353551 , n5866 , n353550 );
nand ( n5870 , n353551 , n1011 );
nand ( n353553 , n353545 , n5870 );
and ( n353554 , n353542 , n353553 );
and ( n5873 , n5849 , n5859 );
or ( n5874 , n353554 , n5873 );
not ( n5875 , n348153 );
not ( n353558 , n4015 );
or ( n353559 , n5875 , n353558 );
or ( n5878 , n348119 , n2071 );
nand ( n353561 , n2071 , n348119 );
nand ( n353562 , n5878 , n353561 );
buf ( n5881 , n348088 );
nand ( n5882 , n353562 , n5881 );
nand ( n5883 , n353559 , n5882 );
not ( n353566 , n5757 );
nor ( n353567 , n353566 , n348181 );
not ( n5886 , n4103 );
not ( n353569 , n5749 );
or ( n353570 , n5886 , n353569 );
nand ( n5889 , n4091 , n5750 );
nand ( n5890 , n353570 , n5889 );
xor ( n5891 , n353567 , n5890 );
and ( n353574 , n4106 , n4084 );
xor ( n353575 , n5891 , n353574 );
xor ( n5894 , n5883 , n353575 );
not ( n353577 , n348233 );
not ( n353578 , n351746 );
or ( n5897 , n353577 , n353578 );
not ( n5898 , n558 );
or ( n5899 , n566 , n582 );
or ( n353582 , n567 , n583 );
nand ( n353583 , n5899 , n353582 );
not ( n5902 , n353583 );
not ( n353585 , n565 );
not ( n353586 , n581 );
and ( n5905 , n353585 , n353586 );
nor ( n5906 , n5905 , n4030 );
nand ( n5907 , n5902 , n5906 );
not ( n353590 , n5907 );
not ( n353591 , n353590 );
not ( n5910 , n351727 );
or ( n353593 , n353591 , n5910 );
not ( n353594 , n565 );
not ( n5913 , n581 );
and ( n5914 , n353594 , n5913 );
nor ( n5915 , n564 , n580 );
nor ( n353598 , n5914 , n5915 );
not ( n353599 , n353598 );
not ( n5918 , n2059 );
or ( n353601 , n353599 , n5918 );
not ( n353602 , n5915 );
not ( n5921 , n2064 );
and ( n5922 , n353602 , n5921 );
nor ( n5923 , n5922 , n351737 );
nand ( n353606 , n353601 , n5923 );
not ( n353607 , n353606 );
nand ( n5926 , n353593 , n353607 );
not ( n353609 , n5926 );
and ( n353610 , n563 , n579 );
nor ( n5929 , n563 , n579 );
nor ( n5930 , n353610 , n5929 );
buf ( n5931 , n5930 );
nand ( n353614 , n353609 , n5931 );
not ( n353615 , n5931 );
nand ( n5934 , n5926 , n353615 );
nand ( n353617 , n353614 , n5934 );
buf ( n353618 , n353617 );
not ( n5937 , n353618 );
not ( n5938 , n5937 );
or ( n5939 , n5898 , n5938 );
not ( n353622 , n5934 );
not ( n353623 , n353614 );
or ( n5942 , n353622 , n353623 );
nand ( n353625 , n5942 , n348230 );
nand ( n353626 , n5939 , n353625 );
nand ( n5945 , n353626 , n559 );
nand ( n5946 , n5897 , n5945 );
and ( n5947 , n5894 , n5946 );
and ( n353630 , n5883 , n353575 );
or ( n353631 , n5947 , n353630 );
xor ( n5950 , n5874 , n353631 );
not ( n353633 , n4109 );
not ( n353634 , n5838 );
or ( n5953 , n353633 , n353634 );
nand ( n5954 , n353551 , n1871 );
nand ( n5955 , n5953 , n5954 );
not ( n353638 , n348153 );
not ( n353639 , n353562 );
or ( n5958 , n353638 , n353639 );
buf ( n353641 , n351740 );
nand ( n353642 , n353641 , n348119 );
not ( n5961 , n353642 );
not ( n5962 , n353641 );
nand ( n5963 , n5962 , n556 );
not ( n353646 , n5963 );
or ( n353647 , n5961 , n353646 );
nand ( n5966 , n353647 , n5881 );
nand ( n353649 , n5958 , n5966 );
xor ( n353650 , n5955 , n353649 );
xor ( n5969 , n353567 , n5890 );
and ( n5970 , n5969 , n353574 );
and ( n5971 , n353567 , n5890 );
or ( n353654 , n5970 , n5971 );
xor ( n353655 , n353650 , n353654 );
and ( n5974 , n5950 , n353655 );
and ( n353657 , n5874 , n353631 );
or ( n353658 , n5974 , n353657 );
xor ( n5977 , n353526 , n353658 );
xor ( n5978 , n5955 , n353649 );
and ( n5979 , n5978 , n353654 );
and ( n353662 , n5955 , n353649 );
or ( n353663 , n5979 , n353662 );
xor ( n5982 , n545 , n546 );
and ( n353665 , n348158 , n5982 );
not ( n353666 , n546 );
not ( n5985 , n348332 );
or ( n5986 , n353666 , n5985 );
nand ( n5987 , n348331 , n5761 );
nand ( n353670 , n5986 , n5987 );
not ( n353671 , n353670 );
not ( n5990 , n5757 );
not ( n353673 , n5990 );
not ( n353674 , n353673 );
or ( n5993 , n353671 , n353674 );
and ( n5994 , n348285 , n5765 );
not ( n5995 , n348285 );
not ( n353678 , n546 );
nor ( n353679 , n353678 , n547 , n548 );
and ( n5998 , n5995 , n353679 );
nor ( n353681 , n5994 , n5998 );
nand ( n353682 , n5993 , n353681 );
xor ( n6001 , n353665 , n353682 );
and ( n6002 , n5755 , n5758 );
not ( n6003 , n5762 );
not ( n353686 , n5771 );
nor ( n353687 , n6002 , n6003 , n353686 );
nor ( n6006 , n353687 , n5780 );
xor ( n353689 , n6001 , n6006 );
not ( n353690 , n353641 );
nand ( n6009 , n353690 , n1916 );
not ( n6010 , n348119 );
nand ( n6011 , n6010 , n348090 );
not ( n353694 , n6011 );
not ( n353695 , n353618 );
nand ( n6014 , n353694 , n353695 );
nand ( n353697 , n353641 , n1919 );
nand ( n353698 , n353618 , n1763 );
nand ( n6017 , n6009 , n6014 , n353697 , n353698 );
xor ( n6018 , n353689 , n6017 );
not ( n6019 , n348233 );
not ( n353702 , n558 );
xor ( n353703 , n562 , n578 );
nor ( n6022 , n5907 , n5929 );
not ( n353705 , n6022 );
not ( n353706 , n1841 );
or ( n6025 , n353705 , n353706 );
not ( n6026 , n5929 );
not ( n6027 , n6026 );
not ( n6028 , n353606 );
or ( n6029 , n6027 , n6028 );
nand ( n6030 , n563 , n579 );
nand ( n6031 , n6029 , n6030 );
not ( n6032 , n6031 );
nand ( n6033 , n6025 , n6032 );
xor ( n6034 , n353703 , n6033 );
not ( n6035 , n6034 );
not ( n6036 , n6035 );
or ( n6037 , n353702 , n6036 );
nand ( n6038 , n6034 , n348230 );
nand ( n6039 , n6037 , n6038 );
not ( n6040 , n6039 );
or ( n6041 , n6019 , n6040 );
not ( n6042 , n558 );
or ( n6043 , n577 , n561 );
nand ( n6044 , n577 , n561 );
nand ( n6045 , n6043 , n6044 );
not ( n6046 , n6045 );
not ( n6047 , n6046 );
not ( n6048 , n562 );
not ( n6049 , n578 );
and ( n6050 , n6048 , n6049 );
nor ( n6051 , n6050 , n5929 );
not ( n6052 , n580 );
nand ( n6053 , n4623 , n6052 );
and ( n6054 , n6051 , n2049 , n2063 , n6053 );
not ( n6055 , n6054 );
not ( n6056 , n351727 );
or ( n6057 , n6055 , n6056 );
not ( n6058 , n2059 );
not ( n6059 , n353598 );
or ( n6060 , n6058 , n6059 );
nand ( n6061 , n6060 , n5923 );
not ( n6062 , n562 );
not ( n6063 , n578 );
and ( n6064 , n6062 , n6063 );
nor ( n6065 , n6064 , n5929 );
and ( n6066 , n6061 , n6065 );
nor ( n6067 , n562 , n578 );
or ( n6068 , n6067 , n6030 );
nand ( n6069 , n562 , n578 );
nand ( n6070 , n6068 , n6069 );
nor ( n6071 , n6066 , n6070 );
nand ( n6072 , n6057 , n6071 );
not ( n6073 , n6072 );
not ( n6074 , n6073 );
or ( n6075 , n6047 , n6074 );
not ( n6076 , n6044 );
nor ( n6077 , n561 , n577 );
nor ( n6078 , n6076 , n6077 );
not ( n6079 , n6078 );
nand ( n6080 , n6079 , n6072 );
nand ( n6081 , n6075 , n6080 );
not ( n6082 , n6081 );
not ( n6083 , n6082 );
or ( n6084 , n6042 , n6083 );
and ( n6085 , n6072 , n6078 );
not ( n6086 , n6072 );
and ( n6087 , n6086 , n6045 );
nor ( n6088 , n6085 , n6087 );
nand ( n6089 , n6088 , n348230 );
nand ( n6090 , n6084 , n6089 );
nand ( n6091 , n6090 , n559 );
nand ( n6092 , n6041 , n6091 );
xor ( n6093 , n6018 , n6092 );
xor ( n6094 , n353663 , n6093 );
not ( n6095 , n559 );
not ( n6096 , n6039 );
or ( n6097 , n6095 , n6096 );
nand ( n6098 , n353626 , n348233 );
nand ( n6099 , n6097 , n6098 );
not ( n6100 , n1925 );
not ( n6101 , n5724 );
or ( n6102 , n6100 , n6101 );
nand ( n6103 , n5857 , n5718 );
nand ( n6104 , n6102 , n6103 );
xor ( n6105 , n6099 , n6104 );
xor ( n6106 , n5753 , n5785 );
xor ( n6107 , n6106 , n5801 );
and ( n6108 , n6105 , n6107 );
and ( n6109 , n6099 , n6104 );
or ( n6110 , n6108 , n6109 );
xor ( n6111 , n6094 , n6110 );
xor ( n6112 , n5977 , n6111 );
buf ( n6113 , n6112 );
xor ( n6114 , n6099 , n6104 );
xor ( n6115 , n6114 , n6107 );
xor ( n6116 , n351764 , n4107 );
and ( n6117 , n6116 , n4120 );
and ( n6118 , n351764 , n4107 );
or ( n6119 , n6117 , n6118 );
xor ( n6120 , n5849 , n5859 );
xor ( n353803 , n6120 , n353553 );
xor ( n353804 , n6119 , n353803 );
xor ( n353805 , n4003 , n4007 );
and ( n353806 , n353805 , n4019 );
and ( n353807 , n4003 , n4007 );
or ( n353808 , n353806 , n353807 );
and ( n353809 , n353804 , n353808 );
and ( n353810 , n6119 , n353803 );
or ( n353811 , n353809 , n353810 );
xor ( n353812 , n6115 , n353811 );
xor ( n353813 , n5874 , n353631 );
xor ( n353814 , n353813 , n353655 );
and ( n353815 , n353812 , n353814 );
and ( n353816 , n6115 , n353811 );
or ( n353817 , n353815 , n353816 );
nand ( n353818 , n6113 , n353817 );
not ( n353819 , n353818 );
nor ( n353820 , n6113 , n353817 );
nor ( n353821 , n353819 , n353820 );
not ( n353822 , n3990 );
not ( n353823 , n4128 );
or ( n353824 , n353822 , n353823 );
nand ( n353825 , n1988 , n2087 );
nand ( n353826 , n353824 , n353825 );
or ( n353827 , n351823 , n353826 );
xor ( n353828 , n5883 , n353575 );
xor ( n353829 , n353828 , n5946 );
xor ( n353830 , n4066 , n4121 );
and ( n353831 , n353830 , n4126 );
and ( n353832 , n4066 , n4121 );
or ( n353833 , n353831 , n353832 );
xor ( n353834 , n353829 , n353833 );
xor ( n353835 , n6119 , n353803 );
xor ( n353836 , n353835 , n353808 );
xor ( n353837 , n353834 , n353836 );
xor ( n353838 , n4020 , n4024 );
and ( n353839 , n353838 , n4127 );
and ( n353840 , n4020 , n4024 );
or ( n353841 , n353839 , n353840 );
nor ( n353842 , n353837 , n353841 );
nor ( n353843 , n353842 , n4131 );
nand ( n353844 , n353827 , n353843 );
xor ( n353845 , n6115 , n353811 );
xor ( n353846 , n353845 , n353814 );
xor ( n353847 , n353829 , n353833 );
and ( n353848 , n353847 , n353836 );
and ( n353849 , n353829 , n353833 );
or ( n353850 , n353848 , n353849 );
nand ( n353851 , n353846 , n353850 );
buf ( n353852 , n353837 );
nand ( n353853 , n353852 , n353841 );
nand ( n353854 , n353844 , n353851 , n353853 );
or ( n353855 , n353846 , n353850 );
nand ( n353856 , n353854 , n353855 );
and ( n353857 , n353821 , n353856 );
not ( n353858 , n353821 );
not ( n353859 , n353856 );
and ( n353860 , n353858 , n353859 );
nor ( n353861 , n353857 , n353860 );
not ( n353862 , n353861 );
nand ( n353863 , n5716 , n353862 );
not ( n353864 , n353863 );
nand ( n353865 , n353397 , n353861 );
not ( n353866 , n353865 );
nor ( n353867 , n353864 , n353866 );
not ( n353868 , n353867 );
not ( n353869 , n353868 );
not ( n353870 , n353869 );
not ( n353871 , n351844 );
not ( n353872 , n4155 );
or ( n353873 , n353871 , n353872 );
nand ( n353874 , n353873 , n3607 );
not ( n353875 , n353874 );
and ( n353876 , n353875 , n3530 );
not ( n353877 , n353876 );
not ( n353878 , n353877 );
not ( n353879 , n4132 );
not ( n353880 , n353826 );
or ( n353881 , n353879 , n353880 );
nand ( n353882 , n2089 , n351820 );
nand ( n353883 , n2174 , n353882 , n4132 );
nand ( n353884 , n353881 , n353883 );
not ( n353885 , n353842 );
nand ( n353886 , n353885 , n353853 );
xnor ( n353887 , n353884 , n353886 );
not ( n353888 , n353887 );
not ( n353889 , n5266 );
not ( n353890 , n5253 );
or ( n353891 , n353889 , n353890 );
nand ( n353892 , n353891 , n5282 );
or ( n353893 , n352927 , n352922 );
not ( n353894 , n353893 );
not ( n353895 , n5246 );
nor ( n353896 , n353894 , n353895 );
and ( n353897 , n353892 , n353896 );
not ( n353898 , n353892 );
not ( n353899 , n353895 );
nand ( n353900 , n353893 , n353899 );
and ( n353901 , n353898 , n353900 );
nor ( n353902 , n353897 , n353901 );
nor ( n353903 , n353888 , n353902 );
not ( n353904 , n353903 );
nor ( n353905 , n352894 , n352918 );
buf ( n353906 , n353905 );
not ( n353907 , n353906 );
buf ( n353908 , n5248 );
nand ( n353909 , n353907 , n353908 );
buf ( n353910 , n353909 );
not ( n353911 , n353910 );
not ( n353912 , n353911 );
nand ( n353913 , n5283 , n353893 );
nand ( n353914 , n5266 , n353893 );
not ( n353915 , n353914 );
nand ( n353916 , n353915 , n5253 );
nand ( n353917 , n353913 , n353916 , n353899 );
not ( n353918 , n353917 );
or ( n353919 , n353912 , n353918 );
nand ( n353920 , n353913 , n353910 , n353916 , n353899 );
nand ( n353921 , n353919 , n353920 );
not ( n353922 , n353885 );
not ( n353923 , n353884 );
or ( n353924 , n353922 , n353923 );
buf ( n353925 , n353853 );
nand ( n353926 , n353924 , n353925 );
nand ( n353927 , n353855 , n353851 );
not ( n353928 , n353927 );
and ( n353929 , n353926 , n353928 );
not ( n353930 , n353926 );
and ( n353931 , n353930 , n353927 );
nor ( n353932 , n353929 , n353931 );
nand ( n353933 , n353921 , n353932 );
and ( n353934 , n353904 , n353933 );
buf ( n353935 , n3473 );
nand ( n353936 , n353878 , n353934 , n353935 );
not ( n353937 , n353933 );
nand ( n353938 , n353902 , n353888 );
not ( n353939 , n353938 );
not ( n353940 , n353939 );
or ( n353941 , n353937 , n353940 );
not ( n353942 , n353932 );
not ( n353943 , n353921 );
nand ( n353944 , n353942 , n353943 );
nand ( n353945 , n353941 , n353944 );
not ( n353946 , n353945 );
not ( n353947 , n3542 );
not ( n353948 , n353875 );
or ( n353949 , n353947 , n353948 );
nor ( n353950 , n2175 , n3423 );
nand ( n353951 , n4155 , n351844 );
and ( n353952 , n353950 , n353951 );
nor ( n353953 , n353952 , n4149 );
nand ( n353954 , n353949 , n353953 );
buf ( n353955 , n353954 );
not ( n353956 , n353933 );
nor ( n353957 , n353888 , n353902 );
nor ( n353958 , n353956 , n353957 );
nand ( n353959 , n353955 , n353958 );
nand ( n353960 , n353936 , n353946 , n353959 );
not ( n353961 , n353960 );
not ( n353962 , n353961 );
or ( n353963 , n353870 , n353962 );
not ( n353964 , n353867 );
nand ( n353965 , n353964 , n353960 );
nand ( n353966 , n353963 , n353965 );
not ( n353967 , n353966 );
not ( n353968 , n577 );
and ( n353969 , n353967 , n353968 );
and ( n353970 , n353966 , n577 );
nor ( n353971 , n353969 , n353970 );
not ( n353972 , n353957 );
not ( n353973 , n353939 );
nand ( n353974 , n353972 , n353973 );
and ( n353975 , n3513 , n3581 );
not ( n353976 , n353975 );
not ( n353977 , n353875 );
or ( n353978 , n353976 , n353977 );
not ( n353979 , n3541 );
and ( n353980 , n353875 , n353979 );
not ( n353981 , n353950 );
not ( n353982 , n351845 );
or ( n353983 , n353981 , n353982 );
not ( n353984 , n4149 );
nand ( n353985 , n353983 , n353984 );
nor ( n353986 , n353980 , n353985 );
nand ( n353987 , n353978 , n353986 );
and ( n353988 , n353974 , n353987 );
not ( n353989 , n353974 );
not ( n353990 , n353987 );
and ( n353991 , n353989 , n353990 );
nor ( n353992 , n353988 , n353991 );
not ( n353993 , n353992 );
nor ( n353994 , n353993 , n579 );
not ( n6311 , n353956 );
nand ( n6312 , n6311 , n353944 );
and ( n353997 , n6312 , n5157 );
not ( n353998 , n353997 );
nand ( n6315 , n353876 , n353904 , n353935 );
nand ( n6316 , n353972 , n353954 );
nand ( n354001 , n6315 , n6316 , n353973 );
not ( n354002 , n354001 );
not ( n6319 , n354002 );
or ( n6320 , n353998 , n6319 );
nor ( n354005 , n6312 , n578 );
nand ( n354006 , n354001 , n354005 );
nand ( n6323 , n6320 , n354006 );
nor ( n6324 , n353994 , n6323 );
not ( n354009 , n6324 );
not ( n354010 , n4168 );
buf ( n6327 , n3589 );
buf ( n6328 , n3568 );
nand ( n354013 , n354010 , n6327 , n3547 , n6328 );
not ( n354014 , n354013 );
not ( n6331 , n354014 );
or ( n6332 , n354009 , n6331 );
not ( n354017 , n3601 );
not ( n354018 , n4167 );
not ( n6335 , n580 );
and ( n6336 , n354018 , n6335 );
not ( n354021 , n4205 );
nor ( n354022 , n6336 , n354021 );
not ( n6339 , n354022 );
or ( n6340 , n354017 , n6339 );
not ( n354025 , n4174 );
not ( n354026 , n4167 );
not ( n6343 , n580 );
and ( n6344 , n354026 , n6343 );
nor ( n354029 , n6344 , n3604 );
nor ( n354030 , n354025 , n354029 );
nand ( n6347 , n6340 , n354030 );
and ( n6348 , n6324 , n6347 );
not ( n354033 , n6323 );
not ( n354034 , n354033 );
not ( n6351 , n353992 );
nand ( n6352 , n6351 , n579 );
not ( n354037 , n6352 );
not ( n354038 , n354037 );
or ( n6355 , n354034 , n354038 );
nand ( n6356 , n354001 , n6312 );
not ( n354041 , n6356 );
not ( n354042 , n6312 );
nand ( n6359 , n354002 , n354042 );
not ( n6360 , n6359 );
or ( n354045 , n354041 , n6360 );
nand ( n354046 , n354045 , n578 );
nand ( n6363 , n6355 , n354046 );
nor ( n6364 , n6348 , n6363 );
nand ( n354049 , n6332 , n6364 );
xor ( n354050 , n353971 , n354049 );
buf ( n354051 , n354050 );
buf ( n6368 , n354051 );
buf ( n354053 , n6368 );
buf ( n354054 , n354053 );
not ( n6371 , n354054 );
buf ( n354056 , n6371 );
buf ( n354057 , n354056 );
not ( n354058 , n354057 );
or ( n6375 , n4471 , n354058 );
buf ( n354060 , n354053 );
buf ( n354061 , n349406 );
nand ( n354062 , n354060 , n354061 );
buf ( n354063 , n354062 );
buf ( n354064 , n354063 );
nand ( n6381 , n6375 , n354064 );
buf ( n354066 , n6381 );
buf ( n354067 , n354066 );
not ( n354068 , n354067 );
or ( n354069 , n4469 , n354068 );
buf ( n354070 , n602 );
not ( n6387 , n354070 );
not ( n6388 , n579 );
not ( n354073 , n353993 );
nand ( n354074 , n6388 , n354073 );
nand ( n354075 , n6347 , n354074 );
not ( n6392 , n353994 );
nand ( n6393 , n6392 , n354022 , n6327 , n6328 );
nand ( n6394 , n353993 , n579 );
nand ( n354079 , n354075 , n6393 , n6394 );
not ( n354080 , n354079 );
not ( n354081 , n354080 );
nand ( n6398 , n354046 , n354033 );
not ( n6399 , n6398 );
not ( n6400 , n6399 );
and ( n354085 , n354081 , n6400 );
and ( n354086 , n354080 , n6399 );
nor ( n354087 , n354085 , n354086 );
buf ( n354088 , n354087 );
not ( n6405 , n354088 );
or ( n6406 , n6387 , n6405 );
buf ( n354091 , n354087 );
not ( n354092 , n354091 );
buf ( n354093 , n354092 );
buf ( n354094 , n354093 );
buf ( n354095 , n349406 );
nand ( n6412 , n354094 , n354095 );
buf ( n354097 , n6412 );
buf ( n354098 , n354097 );
nand ( n354099 , n6406 , n354098 );
buf ( n354100 , n354099 );
buf ( n354101 , n354100 );
buf ( n354102 , n4464 );
buf ( n354103 , n603 );
buf ( n354104 , n602 );
and ( n354105 , n354103 , n354104 );
not ( n6422 , n354103 );
buf ( n354107 , n349406 );
and ( n6424 , n6422 , n354107 );
nor ( n354109 , n354105 , n6424 );
buf ( n354110 , n354109 );
buf ( n354111 , n354110 );
and ( n6428 , n354102 , n354111 );
buf ( n354113 , n6428 );
buf ( n354114 , n354113 );
nand ( n354115 , n354101 , n354114 );
buf ( n354116 , n354115 );
buf ( n354117 , n354116 );
nand ( n6434 , n354069 , n354117 );
buf ( n354119 , n6434 );
buf ( n354120 , n354119 );
xor ( n354121 , n352140 , n354120 );
xor ( n354122 , n351976 , n352038 );
and ( n354123 , n354122 , n352132 );
and ( n6440 , n351976 , n352038 );
or ( n6441 , n354123 , n6440 );
buf ( n354126 , n6441 );
buf ( n354127 , n354126 );
not ( n354128 , n351924 );
not ( n354129 , n351883 );
or ( n6446 , n354128 , n354129 );
not ( n6447 , n6347 );
nand ( n6448 , n6447 , n354013 );
not ( n354133 , n6388 );
not ( n354134 , n354073 );
or ( n354135 , n354133 , n354134 );
nand ( n6452 , n354135 , n6394 );
not ( n6453 , n6452 );
and ( n6454 , n6448 , n6453 );
not ( n354139 , n6448 );
and ( n354140 , n354139 , n6452 );
nor ( n354141 , n6454 , n354140 );
buf ( n6458 , n354141 );
or ( n6459 , n6458 , n351875 );
not ( n6460 , n600 );
nand ( n354145 , n354141 , n6460 );
nand ( n354146 , n6459 , n354145 );
nand ( n354147 , n354146 , n1722 );
nand ( n6464 , n6446 , n354147 );
buf ( n354149 , n6464 );
xor ( n6466 , n354127 , n354149 );
xor ( n6467 , n352002 , n352028 );
and ( n6468 , n6467 , n352035 );
and ( n6469 , n352002 , n352028 );
or ( n6470 , n6468 , n6469 );
buf ( n354155 , n6470 );
buf ( n354156 , n354155 );
buf ( n354157 , n4362 );
not ( n6474 , n354157 );
buf ( n354159 , n598 );
not ( n6476 , n354159 );
buf ( n354161 , n351901 );
not ( n6478 , n354161 );
or ( n6479 , n6476 , n6478 );
buf ( n354164 , n4221 );
buf ( n354165 , n347312 );
nand ( n6482 , n354164 , n354165 );
buf ( n354167 , n6482 );
buf ( n354168 , n354167 );
nand ( n6485 , n6479 , n354168 );
buf ( n354170 , n6485 );
buf ( n354171 , n354170 );
not ( n6488 , n354171 );
or ( n6489 , n6474 , n6488 );
buf ( n354174 , n4443 );
buf ( n354175 , n352077 );
nand ( n6492 , n354174 , n354175 );
buf ( n354177 , n6492 );
buf ( n354178 , n354177 );
nand ( n6495 , n6489 , n354178 );
buf ( n354180 , n6495 );
buf ( n354181 , n354180 );
xor ( n6498 , n354156 , n354181 );
buf ( n354183 , n349035 );
not ( n6500 , n354183 );
and ( n6501 , n348855 , n348975 );
not ( n6502 , n348855 );
and ( n6503 , n6502 , n594 );
or ( n6504 , n6501 , n6503 );
buf ( n354189 , n6504 );
not ( n6506 , n354189 );
or ( n6507 , n6500 , n6506 );
buf ( n354192 , n351991 );
buf ( n354193 , n1397 );
nand ( n6510 , n354192 , n354193 );
buf ( n354195 , n6510 );
buf ( n354196 , n354195 );
nand ( n6513 , n6507 , n354196 );
buf ( n354198 , n6513 );
buf ( n354199 , n354198 );
buf ( n354200 , n1305 );
buf ( n354201 , n592 );
and ( n6518 , n354200 , n354201 );
buf ( n354203 , n6518 );
buf ( n354204 , n354203 );
not ( n6521 , n348946 );
buf ( n354206 , n592 );
not ( n6523 , n354206 );
buf ( n354208 , n349229 );
not ( n6525 , n354208 );
or ( n6526 , n6523 , n6525 );
buf ( n354211 , n349229 );
not ( n6528 , n354211 );
buf ( n354213 , n6528 );
buf ( n354214 , n354213 );
buf ( n354215 , n348910 );
nand ( n6532 , n354214 , n354215 );
buf ( n354217 , n6532 );
buf ( n354218 , n354217 );
nand ( n6535 , n6526 , n354218 );
buf ( n354220 , n6535 );
not ( n6537 , n354220 );
or ( n6538 , n6521 , n6537 );
not ( n6539 , n4335 );
nand ( n6540 , n6539 , n1250 );
nand ( n6541 , n6538 , n6540 );
buf ( n354226 , n6541 );
xor ( n6543 , n354204 , n354226 );
xor ( n6544 , n352007 , n352012 );
and ( n6545 , n6544 , n352025 );
and ( n6546 , n352007 , n352012 );
or ( n6547 , n6545 , n6546 );
buf ( n354232 , n6547 );
buf ( n354233 , n354232 );
xor ( n6550 , n6543 , n354233 );
buf ( n354235 , n6550 );
buf ( n354236 , n354235 );
xor ( n6553 , n354199 , n354236 );
buf ( n354238 , n347319 );
not ( n6555 , n354238 );
buf ( n354240 , n596 );
not ( n6557 , n354240 );
buf ( n354242 , n352095 );
not ( n6559 , n354242 );
or ( n6560 , n6557 , n6559 );
not ( n6561 , n4410 );
buf ( n354246 , n6561 );
not ( n6563 , n354246 );
buf ( n354248 , n6563 );
buf ( n354249 , n354248 );
not ( n6566 , n354249 );
buf ( n354251 , n6566 );
buf ( n354252 , n354251 );
buf ( n354253 , n348865 );
nand ( n6570 , n354252 , n354253 );
buf ( n354255 , n6570 );
buf ( n354256 , n354255 );
nand ( n6573 , n6560 , n354256 );
buf ( n354258 , n6573 );
buf ( n354259 , n354258 );
not ( n6576 , n354259 );
or ( n6577 , n6555 , n6576 );
buf ( n354262 , n351965 );
buf ( n354263 , n348898 );
nand ( n6580 , n354262 , n354263 );
buf ( n354265 , n6580 );
buf ( n354266 , n354265 );
nand ( n6583 , n6577 , n354266 );
buf ( n354268 , n6583 );
buf ( n354269 , n354268 );
xor ( n6586 , n6553 , n354269 );
buf ( n354271 , n6586 );
buf ( n354272 , n354271 );
xor ( n6589 , n6498 , n354272 );
buf ( n354274 , n6589 );
buf ( n354275 , n354274 );
xor ( n6592 , n6466 , n354275 );
buf ( n354277 , n6592 );
buf ( n354278 , n354277 );
xor ( n6595 , n354121 , n354278 );
buf ( n354280 , n6595 );
buf ( n354281 , n354280 );
xor ( n6598 , n605 , n606 );
buf ( n6599 , n6598 );
buf ( n6600 , n6599 );
buf ( n354285 , n6600 );
not ( n6602 , n354285 );
nand ( n6603 , n353867 , n353961 );
not ( n6604 , n577 );
nand ( n6605 , n6603 , n353965 , n6604 );
not ( n6606 , n6605 );
not ( n6607 , n6363 );
or ( n6608 , n6606 , n6607 );
not ( n6609 , n6604 );
nand ( n6610 , n6609 , n353966 );
nand ( n6611 , n6608 , n6610 );
not ( n6612 , n6611 );
or ( n6613 , n354014 , n6347 );
and ( n6614 , n6605 , n6324 );
nand ( n6615 , n6613 , n6614 );
nand ( n6616 , n6612 , n6615 );
buf ( n354301 , n576 );
not ( n354302 , n354301 );
buf ( n354303 , n354302 );
not ( n354304 , n354303 );
buf ( n354305 , n353376 );
not ( n6618 , n354305 );
buf ( n354307 , n5249 );
not ( n354308 , n354307 );
or ( n6621 , n6618 , n354308 );
buf ( n354310 , n353384 );
nand ( n354311 , n6621 , n354310 );
buf ( n354312 , n354311 );
not ( n354313 , n354312 );
buf ( n354314 , n5253 );
buf ( n354315 , n352946 );
buf ( n354316 , n353376 );
buf ( n354317 , n5266 );
nand ( n6630 , n354314 , n354315 , n354316 , n354317 );
buf ( n354319 , n6630 );
nand ( n354320 , n5283 , n352946 , n353376 );
nand ( n6633 , n354313 , n354319 , n354320 );
not ( n354322 , n5381 );
not ( n354323 , n5369 );
nand ( n6636 , n354323 , n5368 );
not ( n354325 , n6636 );
or ( n354326 , n354322 , n354325 );
not ( n6639 , n5368 );
nand ( n354328 , n6639 , n5369 );
nand ( n354329 , n354326 , n354328 );
not ( n6642 , n5351 );
not ( n354331 , n5364 );
or ( n354332 , n6642 , n354331 );
or ( n6645 , n5364 , n5351 );
nand ( n354334 , n6645 , n5339 );
nand ( n354335 , n354332 , n354334 );
buf ( n354336 , n354335 );
not ( n354337 , n354336 );
buf ( n354338 , n354337 );
not ( n6651 , n354338 );
buf ( n354340 , n353042 );
not ( n354341 , n354340 );
buf ( n354342 , n2851 );
not ( n354343 , n354342 );
or ( n354344 , n354341 , n354343 );
buf ( n354345 , n2550 );
buf ( n354346 , n552 );
buf ( n354347 , n566 );
xor ( n6660 , n354346 , n354347 );
buf ( n354349 , n6660 );
buf ( n354350 , n354349 );
nand ( n6663 , n354345 , n354350 );
buf ( n354352 , n6663 );
buf ( n354353 , n354352 );
nand ( n6666 , n354344 , n354353 );
buf ( n354355 , n6666 );
buf ( n354356 , n354355 );
not ( n6669 , n354356 );
buf ( n354358 , n6669 );
buf ( n354359 , n354358 );
not ( n6672 , n354359 );
buf ( n354361 , n353029 );
not ( n354362 , n354361 );
buf ( n354363 , n347336 );
buf ( n354364 , n347338 );
and ( n354365 , n354363 , n354364 );
buf ( n354366 , n354365 );
buf ( n354367 , n354366 );
not ( n354368 , n354367 );
or ( n6681 , n354362 , n354368 );
buf ( n354370 , n348473 );
buf ( n354371 , n548 );
buf ( n354372 , n570 );
xor ( n354373 , n354371 , n354372 );
buf ( n354374 , n354373 );
buf ( n354375 , n354374 );
nand ( n354376 , n354370 , n354375 );
buf ( n354377 , n354376 );
buf ( n354378 , n354377 );
nand ( n354379 , n6681 , n354378 );
buf ( n354380 , n354379 );
buf ( n354381 , n354380 );
not ( n354382 , n354381 );
and ( n354383 , n6672 , n354382 );
buf ( n354384 , n354380 );
buf ( n354385 , n354358 );
and ( n354386 , n354384 , n354385 );
nor ( n6699 , n354383 , n354386 );
buf ( n354388 , n6699 );
buf ( n354389 , n352998 );
not ( n6702 , n354389 );
buf ( n354391 , n351330 );
not ( n354392 , n354391 );
or ( n6705 , n6702 , n354392 );
buf ( n354394 , n3650 );
xor ( n354395 , n564 , n554 );
buf ( n354396 , n354395 );
nand ( n354397 , n354394 , n354396 );
buf ( n354398 , n354397 );
buf ( n354399 , n354398 );
nand ( n354400 , n6705 , n354399 );
buf ( n354401 , n354400 );
and ( n6714 , n354388 , n354401 );
not ( n354403 , n354388 );
buf ( n354404 , n354401 );
not ( n6717 , n354404 );
buf ( n354406 , n6717 );
and ( n354407 , n354403 , n354406 );
nor ( n6720 , n6714 , n354407 );
not ( n354409 , n6720 );
not ( n354410 , n354409 );
or ( n6723 , n6651 , n354410 );
nand ( n354412 , n354335 , n6720 );
nand ( n354413 , n6723 , n354412 );
buf ( n354414 , n353104 );
not ( n354415 , n354414 );
buf ( n354416 , n3242 );
not ( n6729 , n354416 );
or ( n354418 , n354415 , n6729 );
buf ( n354419 , n347382 );
xor ( n6732 , n572 , n546 );
buf ( n354421 , n6732 );
nand ( n354422 , n354419 , n354421 );
buf ( n354423 , n354422 );
buf ( n354424 , n354423 );
nand ( n354425 , n354418 , n354424 );
buf ( n354426 , n354425 );
buf ( n354427 , n5333 );
not ( n354428 , n354427 );
buf ( n354429 , n2828 );
not ( n354430 , n354429 );
or ( n354431 , n354428 , n354430 );
buf ( n354432 , n2243 );
buf ( n354433 , n550 );
buf ( n354434 , n568 );
xor ( n6747 , n354433 , n354434 );
buf ( n354436 , n6747 );
buf ( n354437 , n354436 );
nand ( n6750 , n354432 , n354437 );
buf ( n354439 , n6750 );
buf ( n354440 , n354439 );
nand ( n6753 , n354431 , n354440 );
buf ( n354442 , n6753 );
xor ( n354443 , n354426 , n354442 );
buf ( n354444 , n354443 );
not ( n354445 , n5407 );
buf ( n354446 , n558 );
buf ( n354447 , n560 );
xor ( n354448 , n354446 , n354447 );
buf ( n354449 , n354448 );
not ( n6762 , n354449 );
or ( n354451 , n354445 , n6762 );
not ( n354452 , n560 );
nor ( n6765 , n561 , n562 );
not ( n354454 , n6765 );
or ( n354455 , n354452 , n354454 );
not ( n6768 , n560 );
nand ( n354457 , n6768 , n561 , n562 );
nand ( n354458 , n354455 , n354457 );
xor ( n6771 , n560 , n559 );
nand ( n354460 , n354458 , n6771 );
nand ( n354461 , n354451 , n354460 );
buf ( n354462 , n354461 );
xor ( n354463 , n354444 , n354462 );
buf ( n354464 , n354463 );
xnor ( n6777 , n354413 , n354464 );
xor ( n354466 , n354329 , n6777 );
xor ( n354467 , n352988 , n353005 );
and ( n6780 , n354467 , n353011 );
and ( n354469 , n352988 , n353005 );
or ( n354470 , n6780 , n354469 );
buf ( n354471 , n354470 );
buf ( n354472 , n354471 );
buf ( n354473 , n352981 );
not ( n6786 , n354473 );
buf ( n354475 , n352312 );
buf ( n354476 , n4625 );
nor ( n6789 , n354475 , n354476 );
buf ( n354478 , n6789 );
buf ( n354479 , n354478 );
not ( n6792 , n354479 );
or ( n354481 , n6786 , n6792 );
buf ( n354482 , n352295 );
buf ( n354483 , n556 );
buf ( n354484 , n562 );
xor ( n354485 , n354483 , n354484 );
buf ( n354486 , n354485 );
buf ( n354487 , n354486 );
nand ( n354488 , n354482 , n354487 );
buf ( n354489 , n354488 );
buf ( n354490 , n354489 );
nand ( n354491 , n354481 , n354490 );
buf ( n354492 , n354491 );
buf ( n354493 , n354492 );
buf ( n354494 , n559 );
buf ( n354495 , n561 );
or ( n354496 , n354494 , n354495 );
buf ( n354497 , n562 );
nand ( n6810 , n354496 , n354497 );
buf ( n354499 , n6810 );
buf ( n354500 , n354499 );
buf ( n354501 , n559 );
buf ( n354502 , n561 );
nand ( n354503 , n354501 , n354502 );
buf ( n354504 , n354503 );
buf ( n354505 , n354504 );
buf ( n354506 , n560 );
nand ( n6819 , n354500 , n354505 , n354506 );
buf ( n354508 , n6819 );
buf ( n354509 , n354508 );
not ( n6822 , n354509 );
buf ( n354511 , n5404 );
not ( n354512 , n354511 );
buf ( n354513 , n3763 );
not ( n354514 , n354513 );
or ( n354515 , n354512 , n354514 );
buf ( n354516 , n544 );
buf ( n354517 , n574 );
xor ( n354518 , n354516 , n354517 );
buf ( n354519 , n354518 );
buf ( n354520 , n354519 );
buf ( n354521 , n575 );
nand ( n6834 , n354520 , n354521 );
buf ( n354523 , n6834 );
buf ( n354524 , n354523 );
nand ( n6837 , n354515 , n354524 );
buf ( n354526 , n6837 );
buf ( n354527 , n354526 );
not ( n6840 , n354527 );
or ( n354529 , n6822 , n6840 );
buf ( n354530 , n354526 );
buf ( n354531 , n354508 );
or ( n354532 , n354530 , n354531 );
nand ( n354533 , n354529 , n354532 );
buf ( n354534 , n354533 );
buf ( n354535 , n354534 );
xor ( n354536 , n354493 , n354535 );
buf ( n354537 , n353093 );
not ( n354538 , n354537 );
buf ( n354539 , n5406 );
not ( n6852 , n354539 );
buf ( n354541 , n6852 );
buf ( n354542 , n354541 );
not ( n6855 , n354542 );
or ( n354544 , n354538 , n6855 );
buf ( n354545 , n353110 );
nand ( n6858 , n354544 , n354545 );
buf ( n354547 , n6858 );
buf ( n354548 , n354547 );
buf ( n354549 , n353093 );
not ( n354550 , n354549 );
buf ( n354551 , n5406 );
nand ( n6864 , n354550 , n354551 );
buf ( n354553 , n6864 );
buf ( n354554 , n354553 );
nand ( n6867 , n354548 , n354554 );
buf ( n354556 , n6867 );
buf ( n354557 , n354556 );
xor ( n6870 , n354536 , n354557 );
buf ( n354559 , n6870 );
buf ( n354560 , n354559 );
xor ( n6873 , n354472 , n354560 );
buf ( n354562 , n5429 );
not ( n354563 , n354562 );
buf ( n354564 , n353077 );
not ( n354565 , n354564 );
or ( n354566 , n354563 , n354565 );
buf ( n354567 , n353127 );
nand ( n354568 , n354566 , n354567 );
buf ( n354569 , n354568 );
buf ( n354570 , n354569 );
buf ( n354571 , n353074 );
buf ( n354572 , n353117 );
nand ( n6885 , n354571 , n354572 );
buf ( n354574 , n6885 );
buf ( n354575 , n354574 );
nand ( n6888 , n354570 , n354575 );
buf ( n354577 , n6888 );
buf ( n354578 , n354577 );
xor ( n6891 , n6873 , n354578 );
buf ( n354580 , n6891 );
xnor ( n354581 , n354466 , n354580 );
buf ( n354582 , n354581 );
xor ( n354583 , n5486 , n353173 );
and ( n354584 , n354583 , n353360 );
and ( n6897 , n5486 , n353173 );
or ( n354586 , n354584 , n6897 );
buf ( n354587 , n354586 );
xor ( n6900 , n354582 , n354587 );
buf ( n354589 , n353152 );
not ( n354590 , n354589 );
buf ( n354591 , n5386 );
not ( n354592 , n354591 );
or ( n354593 , n354590 , n354592 );
buf ( n354594 , n353152 );
buf ( n354595 , n5386 );
or ( n354596 , n354594 , n354595 );
buf ( n354597 , n353137 );
nand ( n354598 , n354596 , n354597 );
buf ( n354599 , n354598 );
buf ( n354600 , n354599 );
nand ( n354601 , n354593 , n354600 );
buf ( n354602 , n354601 );
buf ( n354603 , n354602 );
xor ( n354604 , n353189 , n353241 );
and ( n354605 , n354604 , n353358 );
and ( n6918 , n353189 , n353241 );
or ( n354607 , n354605 , n6918 );
buf ( n354608 , n354607 );
buf ( n354609 , n354608 );
xor ( n354610 , n354603 , n354609 );
not ( n354611 , n3345 );
and ( n6924 , n580 , n3064 );
not ( n354613 , n580 );
and ( n354614 , n354613 , n554 );
or ( n6927 , n6924 , n354614 );
not ( n354616 , n6927 );
or ( n354617 , n354611 , n354616 );
nand ( n6930 , n3868 , n5657 , n351035 );
nand ( n354619 , n354617 , n6930 );
buf ( n354620 , n353294 );
not ( n6933 , n354620 );
buf ( n354622 , n350110 );
not ( n354623 , n354622 );
or ( n6936 , n6933 , n354623 );
and ( n354625 , n548 , n586 );
not ( n354626 , n548 );
and ( n6939 , n354626 , n348260 );
nor ( n354628 , n354625 , n6939 );
nand ( n354629 , n347663 , n354628 );
buf ( n354630 , n354629 );
nand ( n354631 , n6936 , n354630 );
buf ( n354632 , n354631 );
xor ( n6945 , n354619 , n354632 );
buf ( n354634 , n353276 );
not ( n354635 , n354634 );
buf ( n354636 , n350699 );
not ( n354637 , n354636 );
or ( n354638 , n354635 , n354637 );
buf ( n354639 , n350705 );
buf ( n354640 , n552 );
buf ( n354641 , n582 );
xor ( n354642 , n354640 , n354641 );
buf ( n354643 , n354642 );
buf ( n354644 , n354643 );
nand ( n354645 , n354639 , n354644 );
buf ( n354646 , n354645 );
buf ( n354647 , n354646 );
nand ( n6960 , n354638 , n354647 );
buf ( n354649 , n6960 );
xor ( n354650 , n6945 , n354649 );
not ( n6963 , n354650 );
not ( n6964 , n5616 );
not ( n354653 , n353282 );
or ( n354654 , n6964 , n354653 );
not ( n6967 , n5617 );
not ( n6968 , n353285 );
or ( n354657 , n6967 , n6968 );
nand ( n354658 , n354657 , n353266 );
nand ( n6971 , n354654 , n354658 );
not ( n6972 , n6971 );
not ( n354661 , n6972 );
or ( n354662 , n6963 , n354661 );
or ( n6975 , n6972 , n354650 );
nand ( n6976 , n354662 , n6975 );
buf ( n354665 , n6976 );
not ( n354666 , n353218 );
not ( n6979 , n3093 );
or ( n6980 , n354666 , n6979 );
not ( n354669 , n3362 );
not ( n354670 , n3361 );
or ( n6983 , n354669 , n354670 );
buf ( n354672 , n546 );
buf ( n354673 , n588 );
xor ( n354674 , n354672 , n354673 );
buf ( n354675 , n354674 );
nand ( n6988 , n6983 , n354675 );
nand ( n354677 , n6980 , n6988 );
buf ( n354678 , n559 );
buf ( n354679 , n576 );
xor ( n6992 , n354678 , n354679 );
buf ( n354681 , n6992 );
not ( n354682 , n354681 );
buf ( n354683 , n353193 );
buf ( n354684 , n576 );
buf ( n354685 , n577 );
xnor ( n354686 , n354684 , n354685 );
buf ( n354687 , n354686 );
buf ( n354688 , n354687 );
nor ( n354689 , n354683 , n354688 );
buf ( n354690 , n354689 );
not ( n7003 , n354690 );
or ( n7004 , n354682 , n7003 );
buf ( n354693 , n353193 );
buf ( n354694 , n558 );
buf ( n354695 , n576 );
xor ( n7008 , n354694 , n354695 );
buf ( n354697 , n7008 );
buf ( n354698 , n354697 );
nand ( n354699 , n354693 , n354698 );
buf ( n354700 , n354699 );
nand ( n354701 , n7004 , n354700 );
xor ( n354702 , n354677 , n354701 );
not ( n7015 , n353260 );
not ( n7016 , n2471 );
or ( n7017 , n7015 , n7016 );
buf ( n354706 , n348629 );
buf ( n354707 , n550 );
buf ( n354708 , n584 );
xor ( n7021 , n354707 , n354708 );
buf ( n354710 , n7021 );
buf ( n354711 , n354710 );
nand ( n7024 , n354706 , n354711 );
buf ( n354713 , n7024 );
nand ( n7026 , n7017 , n354713 );
xnor ( n7027 , n354702 , n7026 );
buf ( n354716 , n7027 );
buf ( n7029 , n354716 );
buf ( n354718 , n7029 );
buf ( n354719 , n354718 );
xnor ( n7032 , n354665 , n354719 );
buf ( n354721 , n7032 );
buf ( n354722 , n354721 );
not ( n7035 , n352751 );
not ( n7036 , n5562 );
or ( n7037 , n7035 , n7036 );
nand ( n7038 , n7037 , n5565 );
not ( n7039 , n7038 );
not ( n7040 , n5621 );
nand ( n7041 , n7040 , n5667 );
not ( n7042 , n7041 );
or ( n7043 , n7039 , n7042 );
nand ( n7044 , n5621 , n5666 );
nand ( n7045 , n7043 , n7044 );
buf ( n354734 , n7045 );
xor ( n7047 , n354722 , n354734 );
not ( n7048 , n353319 );
nand ( n7049 , n7048 , n5644 );
not ( n7050 , n7049 );
not ( n7051 , n353343 );
or ( n7052 , n7050 , n7051 );
not ( n7053 , n5644 );
nand ( n7054 , n7053 , n353319 );
nand ( n7055 , n7052 , n7054 );
buf ( n354744 , n7055 );
buf ( n354745 , n559 );
buf ( n354746 , n577 );
or ( n7059 , n354745 , n354746 );
buf ( n354748 , n578 );
nand ( n7061 , n7059 , n354748 );
buf ( n354750 , n7061 );
buf ( n354751 , n354750 );
buf ( n354752 , n559 );
buf ( n354753 , n577 );
nand ( n7066 , n354752 , n354753 );
buf ( n354755 , n7066 );
buf ( n354756 , n354755 );
buf ( n354757 , n576 );
and ( n7070 , n354751 , n354756 , n354757 );
buf ( n354759 , n7070 );
buf ( n354760 , n354759 );
buf ( n354761 , n353203 );
not ( n7074 , n354761 );
buf ( n354763 , n347478 );
not ( n7076 , n354763 );
or ( n7077 , n7074 , n7076 );
buf ( n354766 , n544 );
buf ( n354767 , n590 );
xor ( n7080 , n354766 , n354767 );
buf ( n354769 , n7080 );
buf ( n354770 , n354769 );
buf ( n354771 , n591 );
nand ( n7084 , n354770 , n354771 );
buf ( n354773 , n7084 );
buf ( n354774 , n354773 );
nand ( n7087 , n7077 , n354774 );
buf ( n354776 , n7087 );
buf ( n354777 , n354776 );
xor ( n7090 , n354760 , n354777 );
buf ( n354779 , n7090 );
buf ( n354780 , n354779 );
buf ( n354781 , n353313 );
not ( n7094 , n354781 );
buf ( n354783 , n5162 );
not ( n7096 , n354783 );
or ( n7097 , n7094 , n7096 );
buf ( n354786 , n352491 );
buf ( n7099 , n354786 );
buf ( n354788 , n7099 );
buf ( n354789 , n354788 );
xor ( n7102 , n578 , n556 );
buf ( n354791 , n7102 );
nand ( n7104 , n354789 , n354791 );
buf ( n354793 , n7104 );
buf ( n354794 , n354793 );
nand ( n7107 , n7097 , n354794 );
buf ( n354796 , n7107 );
buf ( n354797 , n354796 );
xor ( n7110 , n354780 , n354797 );
xor ( n7111 , n353198 , n353208 );
and ( n7112 , n7111 , n353223 );
and ( n7113 , n353198 , n353208 );
or ( n7114 , n7112 , n7113 );
buf ( n354803 , n7114 );
buf ( n354804 , n354803 );
xor ( n7117 , n7110 , n354804 );
buf ( n354806 , n7117 );
buf ( n354807 , n354806 );
xor ( n7120 , n354744 , n354807 );
xor ( n7121 , n353226 , n353231 );
and ( n7122 , n7121 , n353238 );
and ( n7123 , n353226 , n353231 );
or ( n7124 , n7122 , n7123 );
buf ( n354813 , n7124 );
buf ( n354814 , n354813 );
xor ( n7127 , n7120 , n354814 );
buf ( n354816 , n7127 );
buf ( n354817 , n354816 );
xor ( n7130 , n7047 , n354817 );
buf ( n354819 , n7130 );
buf ( n354820 , n354819 );
xor ( n7133 , n354610 , n354820 );
buf ( n354822 , n7133 );
buf ( n354823 , n354822 );
xor ( n7136 , n6900 , n354823 );
buf ( n354825 , n7136 );
buf ( n354826 , n354825 );
xor ( n7139 , n353154 , n353160 );
and ( n7140 , n7139 , n353362 );
and ( n7141 , n353154 , n353160 );
or ( n7142 , n7140 , n7141 );
buf ( n354831 , n7142 );
buf ( n354832 , n354831 );
and ( n7145 , n354826 , n354832 );
buf ( n354834 , n7145 );
not ( n7147 , n354834 );
buf ( n354836 , n354825 );
not ( n7149 , n354836 );
buf ( n354838 , n7149 );
buf ( n354839 , n354838 );
buf ( n354840 , n354831 );
not ( n7153 , n354840 );
buf ( n354842 , n7153 );
buf ( n354843 , n354842 );
nand ( n7156 , n354839 , n354843 );
buf ( n354845 , n7156 );
nand ( n7158 , n7147 , n354845 );
not ( n7159 , n7158 );
and ( n7160 , n6633 , n7159 );
not ( n7161 , n6633 );
and ( n7162 , n7161 , n7158 );
nor ( n7163 , n7160 , n7162 );
not ( n7164 , n7163 );
xor ( n7165 , n5734 , n353486 );
and ( n7166 , n7165 , n5843 );
and ( n7167 , n5734 , n353486 );
or ( n7168 , n7166 , n7167 );
xor ( n7169 , n353663 , n6093 );
and ( n7170 , n7169 , n6110 );
and ( n7171 , n353663 , n6093 );
or ( n7172 , n7170 , n7171 );
xor ( n7173 , n7168 , n7172 );
not ( n7174 , n348090 );
not ( n7175 , n556 );
not ( n7176 , n6035 );
or ( n7177 , n7175 , n7176 );
not ( n7178 , n556 );
nand ( n7179 , n7178 , n6034 );
nand ( n7180 , n7177 , n7179 );
not ( n7181 , n7180 );
or ( n7182 , n7174 , n7181 );
and ( n7183 , n353618 , n1919 );
and ( n7184 , n5937 , n1916 );
nor ( n7185 , n7183 , n7184 );
nand ( n7186 , n7182 , n7185 );
xor ( n7187 , n353665 , n353682 );
and ( n7188 , n7187 , n6006 );
and ( n7189 , n353665 , n353682 );
or ( n7190 , n7188 , n7189 );
xor ( n7191 , n7186 , n7190 );
not ( n7192 , n1925 );
not ( n7193 , n554 );
not ( n7194 , n4057 );
or ( n7195 , n7193 , n7194 );
nand ( n7196 , n353641 , n348175 );
nand ( n7197 , n7195 , n7196 );
not ( n7198 , n7197 );
or ( n7199 , n7192 , n7198 );
nand ( n7200 , n5732 , n5718 );
nand ( n7201 , n7199 , n7200 );
xor ( n7202 , n7191 , n7201 );
not ( n7203 , n1875 );
and ( n7204 , n1788 , n1880 );
not ( n7205 , n1788 );
and ( n7206 , n7205 , n550 );
or ( n7207 , n7204 , n7206 );
not ( n7208 , n7207 );
or ( n7209 , n7203 , n7208 );
nand ( n7210 , n353503 , n4078 );
nand ( n7211 , n7209 , n7210 );
nand ( n7212 , n353514 , n1871 );
not ( n7213 , n1974 );
and ( n7214 , n1011 , n552 );
nand ( n7215 , n7213 , n7214 );
not ( n7216 , n552 );
nand ( n7217 , n7216 , n1011 , n1974 );
nand ( n7218 , n7212 , n7215 , n7217 );
xor ( n7219 , n7211 , n7218 );
not ( n7220 , n559 );
not ( n7221 , n558 );
nand ( n7222 , n6051 , n6043 );
nor ( n7223 , n5907 , n7222 );
not ( n7224 , n7223 );
not ( n7225 , n349527 );
or ( n7226 , n7224 , n7225 );
not ( n7227 , n7222 );
and ( n7228 , n6061 , n7227 );
nor ( n7229 , n577 , n561 );
not ( n7230 , n7229 );
or ( n7231 , n578 , n562 );
nand ( n7232 , n7230 , n7231 , n353610 );
or ( n7233 , n7229 , n6069 );
nand ( n7234 , n7232 , n7233 , n6044 );
nor ( n7235 , n7228 , n7234 );
nand ( n7236 , n7226 , n7235 );
nor ( n7237 , n560 , n576 );
not ( n7238 , n7237 );
nand ( n7239 , n560 , n576 );
nand ( n7240 , n7238 , n7239 );
and ( n7241 , n7236 , n7240 );
not ( n7242 , n7236 );
not ( n7243 , n7240 );
and ( n7244 , n7242 , n7243 );
nor ( n7245 , n7241 , n7244 );
not ( n7246 , n7245 );
not ( n7247 , n7246 );
not ( n7248 , n7247 );
or ( n7249 , n7221 , n7248 );
nand ( n7250 , n7246 , n348230 );
nand ( n7251 , n7249 , n7250 );
not ( n7252 , n7251 );
or ( n7253 , n7220 , n7252 );
nand ( n7254 , n6090 , n348233 );
nand ( n7255 , n7253 , n7254 );
xor ( n7256 , n7219 , n7255 );
xor ( n7257 , n7202 , n7256 );
xor ( n7258 , n5814 , n353505 );
and ( n7259 , n7258 , n5842 );
and ( n7260 , n5814 , n353505 );
or ( n7261 , n7259 , n7260 );
not ( n7262 , n5757 );
not ( n7263 , n546 );
not ( n7264 , n1856 );
or ( n7265 , n7263 , n7264 );
nand ( n7266 , n351755 , n5761 );
nand ( n7267 , n7265 , n7266 );
not ( n7268 , n7267 );
or ( n7269 , n7262 , n7268 );
xor ( n7270 , n546 , n547 );
not ( n7271 , n7270 );
nor ( n7272 , n7271 , n5757 );
nand ( n7273 , n353670 , n7272 );
nand ( n7274 , n7269 , n7273 );
or ( n7275 , n545 , n546 );
nand ( n7276 , n7275 , n348158 );
nand ( n7277 , n545 , n546 );
and ( n7278 , n7276 , n7277 , n544 );
not ( n7279 , n5982 );
not ( n7280 , n544 );
not ( n7281 , n348171 );
or ( n7282 , n7280 , n7281 );
not ( n7283 , n544 );
nand ( n7284 , n348174 , n7283 );
nand ( n7285 , n7282 , n7284 );
not ( n7286 , n7285 );
or ( n7287 , n7279 , n7286 );
not ( n7288 , n544 );
not ( n7289 , n348181 );
or ( n7290 , n7288 , n7289 );
nand ( n7291 , n348292 , n7283 );
nand ( n7292 , n7290 , n7291 );
xnor ( n7293 , n544 , n545 );
nor ( n7294 , n5982 , n7293 );
nand ( n7295 , n7292 , n7294 );
nand ( n7296 , n7287 , n7295 );
xor ( n7297 , n7278 , n7296 );
xor ( n7298 , n7274 , n7297 );
not ( n7299 , n5735 );
not ( n7300 , n548 );
not ( n7301 , n4114 );
or ( n7302 , n7300 , n7301 );
nand ( n7303 , n348266 , n351773 );
nand ( n7304 , n7302 , n7303 );
not ( n7305 , n7304 );
or ( n7306 , n7299 , n7305 );
nand ( n7307 , n5810 , n5751 );
nand ( n7308 , n7306 , n7307 );
xor ( n7309 , n7298 , n7308 );
xor ( n7310 , n7261 , n7309 );
xor ( n7311 , n353689 , n6017 );
and ( n7312 , n7311 , n6092 );
and ( n7313 , n353689 , n6017 );
or ( n7314 , n7312 , n7313 );
xor ( n7315 , n7310 , n7314 );
xor ( n7316 , n7257 , n7315 );
xor ( n7317 , n7173 , n7316 );
not ( n7318 , n7317 );
xor ( n7319 , n353526 , n353658 );
and ( n7320 , n7319 , n6111 );
and ( n7321 , n353526 , n353658 );
or ( n7322 , n7320 , n7321 );
not ( n7323 , n7322 );
nand ( n7324 , n7318 , n7323 );
buf ( n7325 , n7324 );
buf ( n7326 , n7317 );
nand ( n7327 , n7326 , n7322 );
nand ( n7328 , n7325 , n7327 );
not ( n7329 , n7328 );
or ( n7330 , n353856 , n353820 );
nand ( n7331 , n7330 , n353818 );
not ( n7332 , n7331 );
or ( n7333 , n7329 , n7332 );
or ( n7334 , n7328 , n7331 );
nand ( n7335 , n7333 , n7334 );
nor ( n7336 , n7164 , n7335 );
not ( n7337 , n7336 );
nand ( n7338 , n7164 , n7335 );
nand ( n7339 , n7337 , n7338 );
and ( n7340 , n353945 , n353863 );
nor ( n7341 , n7340 , n353866 );
nand ( n7342 , n353955 , n353863 , n353958 );
not ( n7343 , n353935 );
nor ( n7344 , n7343 , n353877 );
nand ( n7345 , n7344 , n353863 , n353958 );
nand ( n7346 , n7341 , n7342 , n7345 );
xor ( n7347 , n7339 , n7346 );
not ( n7348 , n7347 );
not ( n7349 , n7348 );
not ( n7350 , n7349 );
or ( n7351 , n354304 , n7350 );
nand ( n7352 , n7348 , n576 );
nand ( n7353 , n7351 , n7352 );
not ( n7354 , n7353 );
and ( n7355 , n6616 , n7354 );
not ( n7356 , n6616 );
and ( n7357 , n7356 , n7353 );
nor ( n7358 , n7355 , n7357 );
buf ( n7359 , n7358 );
not ( n7360 , n7359 );
and ( n7361 , n604 , n7360 );
not ( n7362 , n604 );
not ( n7363 , n7360 );
and ( n7364 , n7362 , n7363 );
or ( n7365 , n7361 , n7364 );
buf ( n355054 , n7365 );
not ( n7367 , n355054 );
or ( n7368 , n6602 , n7367 );
and ( n7369 , n604 , n354056 );
not ( n7370 , n604 );
and ( n7371 , n7370 , n354053 );
or ( n7372 , n7369 , n7371 );
buf ( n355061 , n7372 );
buf ( n355062 , n604 );
buf ( n355063 , n605 );
and ( n7376 , n355062 , n355063 );
buf ( n355065 , n6598 );
buf ( n355066 , n604 );
buf ( n355067 , n605 );
nor ( n7380 , n355066 , n355067 );
buf ( n355069 , n7380 );
buf ( n355070 , n355069 );
nor ( n7383 , n7376 , n355065 , n355070 );
buf ( n355072 , n7383 );
buf ( n355073 , n355072 );
buf ( n7386 , n355073 );
buf ( n355075 , n7386 );
buf ( n355076 , n355075 );
nand ( n7389 , n355061 , n355076 );
buf ( n355078 , n7389 );
buf ( n355079 , n355078 );
nand ( n7392 , n7368 , n355079 );
buf ( n355081 , n7392 );
buf ( n355082 , n355081 );
buf ( n355083 , n4362 );
not ( n7396 , n355083 );
buf ( n355085 , n598 );
not ( n7398 , n355085 );
buf ( n355087 , n351958 );
not ( n7400 , n355087 );
buf ( n355089 , n7400 );
buf ( n355090 , n355089 );
not ( n7403 , n355090 );
or ( n7404 , n7398 , n7403 );
buf ( n355093 , n351952 );
not ( n7406 , n355093 );
buf ( n355095 , n347312 );
nand ( n7408 , n7406 , n355095 );
buf ( n355097 , n7408 );
buf ( n355098 , n355097 );
nand ( n7411 , n7404 , n355098 );
buf ( n355100 , n7411 );
buf ( n355101 , n355100 );
not ( n7414 , n355101 );
or ( n7415 , n7396 , n7414 );
buf ( n355104 , n598 );
not ( n7417 , n355104 );
buf ( n355106 , n348858 );
not ( n7419 , n355106 );
or ( n7420 , n7417 , n7419 );
buf ( n355109 , n348855 );
buf ( n355110 , n347312 );
nand ( n7423 , n355109 , n355110 );
buf ( n355112 , n7423 );
buf ( n355113 , n355112 );
nand ( n7426 , n7420 , n355113 );
buf ( n355115 , n7426 );
buf ( n355116 , n355115 );
buf ( n355117 , n4443 );
nand ( n7430 , n355116 , n355117 );
buf ( n355119 , n7430 );
buf ( n355120 , n355119 );
nand ( n7433 , n7415 , n355120 );
buf ( n355122 , n7433 );
buf ( n355123 , n355122 );
xor ( n7436 , n349248 , n349252 );
xor ( n7437 , n7436 , n349391 );
buf ( n355126 , n7437 );
buf ( n355127 , n355126 );
xor ( n7440 , n355123 , n355127 );
buf ( n355129 , n1722 );
not ( n7442 , n355129 );
buf ( n355131 , n600 );
not ( n7444 , n355131 );
not ( n7445 , n4388 );
buf ( n355134 , n7445 );
not ( n7447 , n355134 );
or ( n7448 , n7444 , n7447 );
buf ( n355137 , n4388 );
buf ( n355138 , n4193 );
nand ( n7451 , n355137 , n355138 );
buf ( n355140 , n7451 );
buf ( n355141 , n355140 );
nand ( n7454 , n7448 , n355141 );
buf ( n355143 , n7454 );
buf ( n355144 , n355143 );
not ( n7457 , n355144 );
or ( n7458 , n7442 , n7457 );
buf ( n355147 , n600 );
not ( n7460 , n355147 );
buf ( n355149 , n352095 );
not ( n7462 , n355149 );
or ( n7463 , n7460 , n7462 );
buf ( n355152 , n354251 );
buf ( n355153 , n4192 );
nand ( n7466 , n355152 , n355153 );
buf ( n355155 , n7466 );
buf ( n355156 , n355155 );
nand ( n7469 , n7463 , n355156 );
buf ( n355158 , n7469 );
buf ( n355159 , n355158 );
buf ( n355160 , n351924 );
nand ( n7473 , n355159 , n355160 );
buf ( n355162 , n7473 );
buf ( n355163 , n355162 );
nand ( n7476 , n7458 , n355163 );
buf ( n355165 , n7476 );
buf ( n355166 , n355165 );
and ( n7479 , n7440 , n355166 );
and ( n7480 , n355123 , n355127 );
or ( n7481 , n7479 , n7480 );
buf ( n355170 , n7481 );
buf ( n355171 , n355170 );
buf ( n355172 , n352149 );
not ( n7485 , n355172 );
buf ( n355174 , n602 );
not ( n7487 , n355174 );
buf ( n355176 , n6458 );
not ( n7489 , n355176 );
buf ( n355178 , n7489 );
buf ( n355179 , n355178 );
not ( n7492 , n355179 );
or ( n7493 , n7487 , n7492 );
buf ( n355182 , n6458 );
buf ( n355183 , n349406 );
nand ( n7496 , n355182 , n355183 );
buf ( n355185 , n7496 );
buf ( n355186 , n355185 );
nand ( n7499 , n7493 , n355186 );
buf ( n355188 , n7499 );
buf ( n355189 , n355188 );
not ( n7502 , n355189 );
or ( n7503 , n7485 , n7502 );
buf ( n355192 , n602 );
not ( n7505 , n355192 );
buf ( n355194 , n351870 );
not ( n7507 , n355194 );
or ( n7508 , n7505 , n7507 );
buf ( n355197 , n351873 );
buf ( n355198 , n349406 );
nand ( n7511 , n355197 , n355198 );
buf ( n355200 , n7511 );
buf ( n355201 , n355200 );
nand ( n7514 , n7508 , n355201 );
buf ( n355203 , n7514 );
buf ( n355204 , n355203 );
buf ( n355205 , n354113 );
nand ( n7518 , n355204 , n355205 );
buf ( n355207 , n7518 );
buf ( n355208 , n355207 );
nand ( n7521 , n7503 , n355208 );
buf ( n355210 , n7521 );
buf ( n355211 , n355210 );
xor ( n7524 , n355171 , n355211 );
buf ( n355213 , n4362 );
not ( n7526 , n355213 );
buf ( n355215 , n352108 );
not ( n7528 , n355215 );
or ( n7529 , n7526 , n7528 );
buf ( n355218 , n355100 );
buf ( n355219 , n4443 );
nand ( n7532 , n355218 , n355219 );
buf ( n355221 , n7532 );
buf ( n355222 , n355221 );
nand ( n7535 , n7529 , n355222 );
buf ( n355224 , n7535 );
buf ( n355225 , n355224 );
buf ( n355226 , n1722 );
not ( n7539 , n355226 );
buf ( n355228 , n351912 );
not ( n7541 , n355228 );
or ( n7542 , n7539 , n7541 );
buf ( n355231 , n355143 );
buf ( n355232 , n351924 );
nand ( n7545 , n355231 , n355232 );
buf ( n355234 , n7545 );
buf ( n355235 , n355234 );
nand ( n7548 , n7542 , n355235 );
buf ( n355237 , n7548 );
buf ( n355238 , n355237 );
xor ( n7551 , n355225 , n355238 );
xor ( n7552 , n348905 , n349215 );
xor ( n7553 , n7552 , n349396 );
buf ( n355242 , n7553 );
buf ( n355243 , n355242 );
xor ( n7556 , n7551 , n355243 );
buf ( n355245 , n7556 );
buf ( n355246 , n355245 );
and ( n7559 , n7524 , n355246 );
and ( n7560 , n355171 , n355211 );
or ( n7561 , n7559 , n7560 );
buf ( n355250 , n7561 );
buf ( n355251 , n355250 );
xor ( n7564 , n355082 , n355251 );
xor ( n7565 , n355225 , n355238 );
and ( n7566 , n7565 , n355243 );
and ( n7567 , n355225 , n355238 );
or ( n7568 , n7566 , n7567 );
buf ( n355257 , n7568 );
buf ( n355258 , n355257 );
xor ( n7571 , n349401 , n351931 );
xor ( n7572 , n7571 , n352135 );
buf ( n355261 , n7572 );
buf ( n355262 , n355261 );
xor ( n7575 , n355258 , n355262 );
buf ( n355264 , n352149 );
not ( n7577 , n355264 );
buf ( n355266 , n354100 );
not ( n7579 , n355266 );
or ( n7580 , n7577 , n7579 );
buf ( n355269 , n355188 );
buf ( n355270 , n354113 );
nand ( n7583 , n355269 , n355270 );
buf ( n355272 , n7583 );
buf ( n355273 , n355272 );
nand ( n7586 , n7580 , n355273 );
buf ( n355275 , n7586 );
buf ( n355276 , n355275 );
xor ( n7589 , n7575 , n355276 );
buf ( n355278 , n7589 );
buf ( n355279 , n355278 );
and ( n7592 , n7564 , n355279 );
and ( n7593 , n355082 , n355251 );
or ( n7594 , n7592 , n7593 );
buf ( n355283 , n7594 );
buf ( n355284 , n355283 );
xor ( n7597 , n354281 , n355284 );
xor ( n7598 , n355258 , n355262 );
and ( n7599 , n7598 , n355276 );
and ( n7600 , n355258 , n355262 );
or ( n7601 , n7599 , n7600 );
buf ( n355290 , n7601 );
buf ( n355291 , n355290 );
buf ( n355292 , n6600 );
not ( n7605 , n355292 );
xor ( n7606 , n354493 , n354535 );
and ( n7607 , n7606 , n354557 );
and ( n7608 , n354493 , n354535 );
or ( n7609 , n7607 , n7608 );
buf ( n355298 , n7609 );
buf ( n355299 , n355298 );
buf ( n355300 , n354526 );
not ( n7613 , n355300 );
buf ( n355302 , n354508 );
nor ( n7615 , n7613 , n355302 );
buf ( n355304 , n7615 );
buf ( n355305 , n354461 );
not ( n7618 , n355305 );
buf ( n355307 , n354426 );
not ( n7620 , n355307 );
or ( n7621 , n7618 , n7620 );
buf ( n355310 , n354426 );
buf ( n355311 , n354461 );
or ( n7624 , n355310 , n355311 );
buf ( n355313 , n354442 );
nand ( n7626 , n7624 , n355313 );
buf ( n355315 , n7626 );
buf ( n355316 , n355315 );
nand ( n7629 , n7621 , n355316 );
buf ( n355318 , n7629 );
xor ( n7631 , n355304 , n355318 );
not ( n7632 , n354380 );
buf ( n355321 , n352998 );
not ( n7634 , n355321 );
buf ( n355323 , n351330 );
not ( n7636 , n355323 );
or ( n7637 , n7634 , n7636 );
buf ( n355326 , n354398 );
nand ( n7639 , n7637 , n355326 );
buf ( n355328 , n7639 );
not ( n7641 , n355328 );
or ( n7642 , n7632 , n7641 );
buf ( n355331 , n354380 );
buf ( n355332 , n355328 );
nor ( n7645 , n355331 , n355332 );
buf ( n355334 , n7645 );
or ( n7647 , n355334 , n354358 );
nand ( n7648 , n7642 , n7647 );
xor ( n7649 , n7631 , n7648 );
buf ( n355338 , n7649 );
xor ( n7651 , n355299 , n355338 );
not ( n7652 , n354409 );
not ( n7653 , n354335 );
or ( n7654 , n7652 , n7653 );
not ( n7655 , n354338 );
not ( n7656 , n6720 );
or ( n7657 , n7655 , n7656 );
nand ( n7658 , n7657 , n354464 );
nand ( n7659 , n7654 , n7658 );
buf ( n355348 , n7659 );
xor ( n7661 , n7651 , n355348 );
buf ( n355350 , n7661 );
xor ( n7663 , n354472 , n354560 );
and ( n7664 , n7663 , n354578 );
and ( n7665 , n354472 , n354560 );
or ( n7666 , n7664 , n7665 );
buf ( n355355 , n7666 );
xor ( n7668 , n355350 , n355355 );
buf ( n355357 , n574 );
buf ( n355358 , n575 );
and ( n7671 , n355357 , n355358 );
buf ( n355360 , n3763 );
buf ( n355361 , n354519 );
and ( n7674 , n355360 , n355361 );
nor ( n7675 , n7671 , n7674 );
buf ( n355364 , n7675 );
buf ( n355365 , n355364 );
not ( n7678 , n355365 );
buf ( n355367 , n7678 );
buf ( n355368 , n559 );
buf ( n355369 , n560 );
nand ( n7682 , n355368 , n355369 );
buf ( n355371 , n7682 );
and ( n7684 , n355367 , n355371 );
not ( n7685 , n355367 );
buf ( n355374 , n355371 );
not ( n7687 , n355374 );
buf ( n355376 , n7687 );
and ( n7689 , n7685 , n355376 );
or ( n7690 , n7684 , n7689 );
buf ( n355379 , n6732 );
not ( n7692 , n355379 );
buf ( n355381 , n347737 );
not ( n7694 , n355381 );
or ( n7695 , n7692 , n7694 );
buf ( n355384 , n347382 );
buf ( n355385 , n545 );
buf ( n355386 , n572 );
xor ( n7699 , n355385 , n355386 );
buf ( n355388 , n7699 );
buf ( n355389 , n355388 );
nand ( n7702 , n355384 , n355389 );
buf ( n355391 , n7702 );
buf ( n355392 , n355391 );
nand ( n7705 , n7695 , n355392 );
buf ( n355394 , n7705 );
and ( n7707 , n7690 , n355394 );
not ( n7708 , n7690 );
not ( n7709 , n355394 );
and ( n7710 , n7708 , n7709 );
nor ( n7711 , n7707 , n7710 );
not ( n7712 , n7711 );
not ( n7713 , n7712 );
not ( n7714 , n354486 );
not ( n7715 , n5291 );
or ( n7716 , n7714 , n7715 );
buf ( n355405 , n352295 );
buf ( n355406 , n555 );
buf ( n355407 , n562 );
xor ( n7720 , n355406 , n355407 );
buf ( n355409 , n7720 );
buf ( n355410 , n355409 );
nand ( n7723 , n355405 , n355410 );
buf ( n355412 , n7723 );
nand ( n7725 , n7716 , n355412 );
buf ( n355414 , n354374 );
not ( n7727 , n355414 );
buf ( n355416 , n354366 );
not ( n7729 , n355416 );
or ( n7730 , n7727 , n7729 );
buf ( n355419 , n348473 );
buf ( n355420 , n547 );
buf ( n355421 , n570 );
xor ( n7734 , n355420 , n355421 );
buf ( n355423 , n7734 );
buf ( n355424 , n355423 );
nand ( n7737 , n355419 , n355424 );
buf ( n355426 , n7737 );
buf ( n355427 , n355426 );
nand ( n7740 , n7730 , n355427 );
buf ( n355429 , n7740 );
xor ( n7742 , n7725 , n355429 );
buf ( n355431 , n354395 );
not ( n7744 , n355431 );
buf ( n355433 , n4490 );
not ( n7746 , n355433 );
or ( n7747 , n7744 , n7746 );
buf ( n355436 , n3650 );
buf ( n355437 , n553 );
buf ( n355438 , n564 );
xor ( n7751 , n355437 , n355438 );
buf ( n355440 , n7751 );
buf ( n355441 , n355440 );
nand ( n7754 , n355436 , n355441 );
buf ( n355443 , n7754 );
buf ( n355444 , n355443 );
nand ( n7757 , n7747 , n355444 );
buf ( n355446 , n7757 );
xnor ( n7759 , n7742 , n355446 );
buf ( n355448 , n7759 );
not ( n7761 , n355448 );
buf ( n355450 , n7761 );
not ( n7763 , n355450 );
or ( n7764 , n7713 , n7763 );
buf ( n355453 , n7759 );
buf ( n355454 , n7711 );
nand ( n7767 , n355453 , n355454 );
buf ( n355456 , n7767 );
nand ( n7769 , n7764 , n355456 );
buf ( n355458 , n7769 );
not ( n7771 , n5407 );
and ( n7772 , n557 , n560 );
not ( n7773 , n557 );
and ( n7774 , n7773 , n6768 );
nor ( n7775 , n7772 , n7774 );
not ( n7776 , n7775 );
or ( n7777 , n7771 , n7776 );
nand ( n7778 , n354449 , n354458 );
nand ( n7779 , n7777 , n7778 );
buf ( n355468 , n7779 );
not ( n7781 , n354436 );
not ( n7782 , n3768 );
or ( n7783 , n7781 , n7782 );
and ( n7784 , n549 , n568 );
not ( n7785 , n549 );
and ( n7786 , n7785 , n1822 );
nor ( n7787 , n7784 , n7786 );
nand ( n7788 , n2243 , n7787 );
nand ( n7789 , n7783 , n7788 );
buf ( n355478 , n7789 );
xor ( n7791 , n355468 , n355478 );
buf ( n355480 , n354349 );
not ( n7793 , n355480 );
buf ( n355482 , n350874 );
not ( n7795 , n355482 );
or ( n7796 , n7793 , n7795 );
buf ( n355485 , n2550 );
buf ( n355486 , n551 );
buf ( n355487 , n566 );
xor ( n7800 , n355486 , n355487 );
buf ( n355489 , n7800 );
buf ( n355490 , n355489 );
nand ( n7803 , n355485 , n355490 );
buf ( n355492 , n7803 );
buf ( n355493 , n355492 );
nand ( n7806 , n7796 , n355493 );
buf ( n355495 , n7806 );
buf ( n355496 , n355495 );
xor ( n7809 , n7791 , n355496 );
buf ( n355498 , n7809 );
buf ( n355499 , n355498 );
xor ( n7812 , n355458 , n355499 );
buf ( n355501 , n7812 );
xor ( n7814 , n7668 , n355501 );
not ( n7815 , n7814 );
not ( n7816 , n7815 );
xor ( n7817 , n354603 , n354609 );
and ( n7818 , n7817 , n354820 );
and ( n7819 , n354603 , n354609 );
or ( n7820 , n7818 , n7819 );
buf ( n355509 , n7820 );
not ( n7822 , n355509 );
or ( n7823 , n7816 , n7822 );
not ( n7824 , n355509 );
nand ( n7825 , n7824 , n7814 );
nand ( n7826 , n7823 , n7825 );
xor ( n7827 , n354722 , n354734 );
and ( n7828 , n7827 , n354817 );
and ( n7829 , n354722 , n354734 );
or ( n7830 , n7828 , n7829 );
buf ( n355519 , n7830 );
buf ( n355520 , n6777 );
not ( n7833 , n355520 );
buf ( n355522 , n7833 );
buf ( n355523 , n355522 );
not ( n7836 , n355523 );
buf ( n355525 , n354580 );
not ( n7838 , n355525 );
or ( n7839 , n7836 , n7838 );
buf ( n355528 , n354580 );
buf ( n355529 , n355522 );
or ( n7842 , n355528 , n355529 );
buf ( n355531 , n354329 );
nand ( n7844 , n7842 , n355531 );
buf ( n355533 , n7844 );
buf ( n355534 , n355533 );
nand ( n7847 , n7839 , n355534 );
buf ( n355536 , n7847 );
xor ( n7849 , n355519 , n355536 );
buf ( n355538 , n7102 );
not ( n7851 , n355538 );
buf ( n355540 , n5161 );
buf ( n355541 , n5156 );
nor ( n7854 , n355540 , n355541 );
buf ( n355543 , n7854 );
buf ( n355544 , n355543 );
not ( n7857 , n355544 );
or ( n7858 , n7851 , n7857 );
buf ( n355547 , n352491 );
xor ( n7860 , n578 , n555 );
buf ( n355549 , n7860 );
nand ( n7862 , n355547 , n355549 );
buf ( n355551 , n7862 );
buf ( n355552 , n355551 );
nand ( n7865 , n7858 , n355552 );
buf ( n355554 , n7865 );
not ( n7867 , n354628 );
not ( n7868 , n347671 );
or ( n7869 , n7867 , n7868 );
buf ( n355558 , n347530 );
buf ( n355559 , n547 );
buf ( n355560 , n586 );
xor ( n7873 , n355559 , n355560 );
buf ( n355562 , n7873 );
buf ( n355563 , n355562 );
nand ( n7876 , n355558 , n355563 );
buf ( n355565 , n7876 );
nand ( n7878 , n7869 , n355565 );
xor ( n7879 , n355554 , n7878 );
not ( n7880 , n6927 );
not ( n7881 , n3870 );
or ( n7882 , n7880 , n7881 );
buf ( n355571 , n351038 );
xor ( n7884 , n580 , n553 );
buf ( n355573 , n7884 );
nand ( n7886 , n355571 , n355573 );
buf ( n355575 , n7886 );
nand ( n7888 , n7882 , n355575 );
xor ( n7889 , n7879 , n7888 );
buf ( n355578 , n354769 );
not ( n7891 , n355578 );
buf ( n355580 , n347478 );
not ( n7893 , n355580 );
or ( n7894 , n7891 , n7893 );
buf ( n355583 , n590 );
buf ( n355584 , n591 );
nand ( n7897 , n355583 , n355584 );
buf ( n355586 , n7897 );
buf ( n355587 , n355586 );
nand ( n7900 , n7894 , n355587 );
buf ( n355589 , n7900 );
buf ( n355590 , n559 );
buf ( n355591 , n576 );
nand ( n7904 , n355590 , n355591 );
buf ( n355593 , n7904 );
xor ( n7906 , n355589 , n355593 );
buf ( n355595 , n354675 );
not ( n7908 , n355595 );
buf ( n355597 , n350133 );
not ( n7910 , n355597 );
or ( n7911 , n7908 , n7910 );
buf ( n355600 , n545 );
buf ( n355601 , n588 );
xor ( n7914 , n355600 , n355601 );
buf ( n355603 , n7914 );
buf ( n355604 , n355603 );
buf ( n355605 , n347565 );
nand ( n7918 , n355604 , n355605 );
buf ( n355607 , n7918 );
buf ( n355608 , n355607 );
nand ( n7921 , n7911 , n355608 );
buf ( n355610 , n7921 );
xor ( n7923 , n7906 , n355610 );
not ( n7924 , n7923 );
xor ( n7925 , n7889 , n7924 );
buf ( n355614 , n354697 );
not ( n7927 , n355614 );
buf ( n355616 , n354690 );
not ( n7929 , n355616 );
or ( n7930 , n7927 , n7929 );
buf ( n355619 , n353193 );
buf ( n355620 , n557 );
buf ( n355621 , n576 );
xor ( n7934 , n355620 , n355621 );
buf ( n355623 , n7934 );
buf ( n355624 , n355623 );
nand ( n7937 , n355619 , n355624 );
buf ( n355626 , n7937 );
buf ( n355627 , n355626 );
nand ( n7940 , n7930 , n355627 );
buf ( n355629 , n7940 );
buf ( n355630 , n355629 );
buf ( n355631 , n354643 );
not ( n7944 , n355631 );
buf ( n355633 , n3313 );
not ( n7946 , n355633 );
or ( n7947 , n7944 , n7946 );
buf ( n355636 , n350377 );
buf ( n355637 , n551 );
buf ( n355638 , n582 );
xor ( n7951 , n355637 , n355638 );
buf ( n355640 , n7951 );
buf ( n355641 , n355640 );
nand ( n7954 , n355636 , n355641 );
buf ( n355643 , n7954 );
buf ( n355644 , n355643 );
nand ( n7957 , n7947 , n355644 );
buf ( n355646 , n7957 );
buf ( n355647 , n355646 );
xor ( n7960 , n355630 , n355647 );
buf ( n355649 , n354710 );
not ( n7962 , n355649 );
buf ( n355651 , n2471 );
not ( n7964 , n355651 );
or ( n7965 , n7962 , n7964 );
buf ( n355654 , n350726 );
buf ( n355655 , n549 );
buf ( n355656 , n584 );
xor ( n7969 , n355655 , n355656 );
buf ( n355658 , n7969 );
buf ( n355659 , n355658 );
nand ( n7972 , n355654 , n355659 );
buf ( n355661 , n7972 );
buf ( n355662 , n355661 );
nand ( n7975 , n7965 , n355662 );
buf ( n355664 , n7975 );
buf ( n355665 , n355664 );
xnor ( n7978 , n7960 , n355665 );
buf ( n355667 , n7978 );
buf ( n355668 , n355667 );
not ( n7981 , n355668 );
buf ( n355670 , n7981 );
xor ( n7983 , n7925 , n355670 );
buf ( n355672 , n7983 );
xor ( n7985 , n354744 , n354807 );
and ( n7986 , n7985 , n354814 );
and ( n7987 , n354744 , n354807 );
or ( n7988 , n7986 , n7987 );
buf ( n355677 , n7988 );
buf ( n355678 , n355677 );
xor ( n7991 , n355672 , n355678 );
xor ( n7992 , n354780 , n354797 );
and ( n7993 , n7992 , n354804 );
and ( n7994 , n354780 , n354797 );
or ( n7995 , n7993 , n7994 );
buf ( n355684 , n7995 );
buf ( n355685 , n355684 );
buf ( n355686 , n6972 );
not ( n7999 , n355686 );
buf ( n355688 , n7027 );
not ( n8001 , n355688 );
or ( n8002 , n7999 , n8001 );
buf ( n355691 , n354650 );
nand ( n8004 , n8002 , n355691 );
buf ( n355693 , n8004 );
buf ( n355694 , n355693 );
buf ( n355695 , n7027 );
not ( n8008 , n355695 );
buf ( n355697 , n6971 );
nand ( n8010 , n8008 , n355697 );
buf ( n355699 , n8010 );
buf ( n355700 , n355699 );
nand ( n8013 , n355694 , n355700 );
buf ( n355702 , n8013 );
buf ( n355703 , n355702 );
xor ( n8016 , n355685 , n355703 );
and ( n8017 , n354760 , n354777 );
buf ( n355706 , n8017 );
buf ( n355707 , n355706 );
xor ( n8020 , n354619 , n354632 );
and ( n8021 , n8020 , n354649 );
and ( n8022 , n354619 , n354632 );
or ( n8023 , n8021 , n8022 );
buf ( n355712 , n8023 );
xor ( n8025 , n355707 , n355712 );
not ( n8026 , n354677 );
not ( n8027 , n354701 );
or ( n8028 , n8026 , n8027 );
or ( n8029 , n354677 , n354701 );
nand ( n8030 , n8029 , n7026 );
nand ( n8031 , n8028 , n8030 );
buf ( n355720 , n8031 );
xor ( n8033 , n8025 , n355720 );
buf ( n355722 , n8033 );
buf ( n355723 , n355722 );
xor ( n8036 , n8016 , n355723 );
buf ( n355725 , n8036 );
buf ( n355726 , n355725 );
xor ( n8039 , n7991 , n355726 );
buf ( n355728 , n8039 );
xor ( n8041 , n7849 , n355728 );
and ( n8042 , n7826 , n8041 );
not ( n8043 , n7826 );
not ( n8044 , n8041 );
and ( n8045 , n8043 , n8044 );
nor ( n8046 , n8042 , n8045 );
xor ( n8047 , n354582 , n354587 );
and ( n8048 , n8047 , n354823 );
and ( n8049 , n354582 , n354587 );
or ( n8050 , n8048 , n8049 );
buf ( n355739 , n8050 );
nor ( n8052 , n8046 , n355739 );
not ( n8053 , n8052 );
nand ( n8054 , n355739 , n8046 );
and ( n8055 , n8053 , n8054 );
not ( n8056 , n8055 );
not ( n8057 , n8056 );
buf ( n355746 , n5249 );
not ( n8059 , n355746 );
buf ( n355748 , n354825 );
buf ( n355749 , n354831 );
nor ( n8062 , n355748 , n355749 );
buf ( n355751 , n8062 );
buf ( n355752 , n355751 );
buf ( n355753 , n353373 );
nor ( n8066 , n355752 , n355753 );
buf ( n355755 , n8066 );
buf ( n355756 , n355755 );
not ( n8069 , n355756 );
or ( n8070 , n8059 , n8069 );
buf ( n355759 , n354845 );
buf ( n355760 , n353381 );
not ( n8073 , n355760 );
buf ( n355762 , n8073 );
buf ( n355763 , n355762 );
and ( n8076 , n355759 , n355763 );
buf ( n355765 , n354834 );
nor ( n8078 , n8076 , n355765 );
buf ( n355767 , n8078 );
buf ( n355768 , n355767 );
nand ( n8081 , n8070 , n355768 );
buf ( n355770 , n8081 );
buf ( n355771 , n355770 );
not ( n8084 , n355771 );
buf ( n355773 , n8084 );
buf ( n355774 , n355773 );
buf ( n355775 , n355751 );
buf ( n355776 , n353373 );
nor ( n8089 , n355775 , n355776 );
buf ( n355778 , n8089 );
nand ( n8091 , n5281 , n355778 , n5261 );
buf ( n355780 , n8091 );
buf ( n355781 , n5253 );
buf ( n355782 , n355778 );
buf ( n355783 , n5261 );
buf ( n355784 , n5266 );
nand ( n8097 , n355781 , n355782 , n355783 , n355784 );
buf ( n355786 , n8097 );
buf ( n355787 , n355786 );
and ( n8100 , n355774 , n355780 , n355787 );
buf ( n355789 , n8100 );
buf ( n355790 , n355789 );
buf ( n8103 , n355790 );
buf ( n355792 , n8103 );
buf ( n355793 , n355792 );
not ( n8106 , n355793 );
buf ( n355795 , n8106 );
not ( n8108 , n355795 );
or ( n8109 , n8057 , n8108 );
nand ( n8110 , n8055 , n355792 );
nand ( n8111 , n8109 , n8110 );
xor ( n8112 , n7211 , n7218 );
and ( n8113 , n8112 , n7255 );
and ( n8114 , n7211 , n7218 );
or ( n8115 , n8113 , n8114 );
and ( n8116 , n7278 , n7296 );
not ( n8117 , n1875 );
not ( n8118 , n1880 );
not ( n8119 , n1843 );
or ( n8120 , n8118 , n8119 );
nand ( n8121 , n1844 , n550 );
nand ( n8122 , n8120 , n8121 );
not ( n8123 , n8122 );
or ( n8124 , n8117 , n8123 );
not ( n8125 , n1788 );
not ( n8126 , n1880 );
or ( n8127 , n8125 , n8126 );
or ( n8128 , n1880 , n1788 );
nand ( n8129 , n8127 , n8128 );
nand ( n8130 , n8129 , n4078 );
nand ( n8131 , n8124 , n8130 );
xor ( n8132 , n8116 , n8131 );
buf ( n8133 , n2019 );
not ( n8134 , n8133 );
not ( n8135 , n548 );
not ( n8136 , n348746 );
or ( n8137 , n8135 , n8136 );
nand ( n8138 , n997 , n351773 );
nand ( n8139 , n8137 , n8138 );
not ( n8140 , n8139 );
or ( n8141 , n8134 , n8140 );
nand ( n8142 , n7304 , n5751 );
nand ( n8143 , n8141 , n8142 );
xor ( n8144 , n8132 , n8143 );
xor ( n8145 , n8115 , n8144 );
xor ( n8146 , n7186 , n7190 );
and ( n8147 , n8146 , n7201 );
and ( n8148 , n7186 , n7190 );
or ( n8149 , n8147 , n8148 );
xor ( n8150 , n8145 , n8149 );
not ( n8151 , n1871 );
not ( n8152 , n552 );
not ( n8153 , n4011 );
or ( n8154 , n8152 , n8153 );
not ( n8155 , n552 );
nand ( n8156 , n8155 , n1974 );
nand ( n8157 , n8154 , n8156 );
not ( n8158 , n8157 );
or ( n8159 , n8151 , n8158 );
xor ( n8160 , n2071 , n552 );
nand ( n8161 , n8160 , n4109 );
nand ( n8162 , n8159 , n8161 );
not ( n8163 , n348233 );
not ( n8164 , n7251 );
or ( n8165 , n8163 , n8164 );
not ( n8166 , n348230 );
nor ( n8167 , n7237 , n6077 );
nand ( n8168 , n6065 , n8167 );
nor ( n8169 , n8168 , n5907 );
not ( n8170 , n8169 );
not ( n8171 , n1841 );
or ( n8172 , n8170 , n8171 );
and ( n8173 , n6065 , n8167 );
and ( n8174 , n353606 , n8173 );
not ( n8175 , n8167 );
not ( n8176 , n6070 );
or ( n8177 , n8175 , n8176 );
or ( n8178 , n7237 , n6044 );
nand ( n8179 , n8178 , n7239 );
not ( n8180 , n8179 );
nand ( n8181 , n8177 , n8180 );
nor ( n8182 , n8174 , n8181 );
nand ( n8183 , n8172 , n8182 );
not ( n8184 , n8183 );
not ( n8185 , n8184 );
not ( n8186 , n8185 );
or ( n8187 , n8166 , n8186 );
not ( n8188 , n8185 );
nand ( n8189 , n8188 , n558 );
nand ( n8190 , n8187 , n8189 );
nand ( n8191 , n559 , n8190 );
nand ( n8192 , n8165 , n8191 );
xor ( n8193 , n8162 , n8192 );
not ( n8194 , n7180 );
or ( n8195 , n8194 , n348152 );
and ( n8196 , n6088 , n348119 );
not ( n8197 , n6088 );
and ( n8198 , n8197 , n556 );
or ( n8199 , n8196 , n8198 );
not ( n8200 , n8199 );
or ( n8201 , n8200 , n348089 );
nand ( n8202 , n8195 , n8201 );
xor ( n8203 , n8193 , n8202 );
not ( n8204 , n5718 );
not ( n8205 , n7197 );
or ( n8206 , n8204 , n8205 );
not ( n8207 , n554 );
not ( n8208 , n5937 );
or ( n8209 , n8207 , n8208 );
nand ( n8210 , n353618 , n348175 );
nand ( n8211 , n8209 , n8210 );
nand ( n8212 , n8211 , n1925 );
nand ( n8213 , n8206 , n8212 );
nor ( n8214 , n348181 , n7283 );
buf ( n8215 , n5982 );
not ( n8216 , n8215 );
and ( n8217 , n348146 , n544 );
not ( n8218 , n348146 );
and ( n8219 , n8218 , n7283 );
or ( n8220 , n8217 , n8219 );
not ( n8221 , n8220 );
or ( n8222 , n8216 , n8221 );
nor ( n8223 , n7293 , n5982 );
nand ( n8224 , n7285 , n8223 );
nand ( n8225 , n8222 , n8224 );
xor ( n8226 , n8214 , n8225 );
not ( n8227 , n5757 );
and ( n8228 , n966 , n546 );
not ( n8229 , n966 );
and ( n8230 , n8229 , n5761 );
or ( n8231 , n8228 , n8230 );
not ( n8232 , n8231 );
or ( n8233 , n8227 , n8232 );
nand ( n8234 , n7267 , n7272 );
nand ( n8235 , n8233 , n8234 );
xor ( n8236 , n8226 , n8235 );
xor ( n8237 , n8213 , n8236 );
xor ( n8238 , n7274 , n7297 );
and ( n8239 , n8238 , n7308 );
and ( n8240 , n7274 , n7297 );
or ( n8241 , n8239 , n8240 );
xor ( n8242 , n8237 , n8241 );
xor ( n8243 , n8203 , n8242 );
xor ( n8244 , n7261 , n7309 );
and ( n8245 , n8244 , n7314 );
and ( n8246 , n7261 , n7309 );
or ( n8247 , n8245 , n8246 );
xor ( n8248 , n8243 , n8247 );
xor ( n8249 , n8150 , n8248 );
xor ( n8250 , n7202 , n7256 );
and ( n8251 , n8250 , n7315 );
and ( n8252 , n7202 , n7256 );
or ( n8253 , n8251 , n8252 );
xor ( n8254 , n8249 , n8253 );
xor ( n8255 , n7168 , n7172 );
and ( n8256 , n8255 , n7316 );
and ( n8257 , n7168 , n7172 );
or ( n8258 , n8256 , n8257 );
or ( n8259 , n8254 , n8258 );
nand ( n8260 , n8254 , n8258 );
nand ( n8261 , n8259 , n8260 );
not ( n8262 , n8261 );
not ( n8263 , n6112 );
not ( n8264 , n353817 );
and ( n8265 , n8263 , n8264 );
nor ( n8266 , n353846 , n353850 );
nor ( n8267 , n8265 , n8266 );
nand ( n8268 , n7324 , n353854 , n8267 );
or ( n8269 , n7326 , n7322 );
and ( n8270 , n6112 , n353817 );
nand ( n8271 , n8269 , n8270 );
nand ( n8272 , n8268 , n7327 , n8271 );
buf ( n8273 , n8272 );
not ( n8274 , n8273 );
not ( n8275 , n8274 );
or ( n8276 , n8262 , n8275 );
or ( n8277 , n8261 , n8274 );
nand ( n8278 , n8276 , n8277 );
nand ( n8279 , n8111 , n8278 );
buf ( n8280 , n8279 );
not ( n8281 , n8111 );
not ( n8282 , n8278 );
nand ( n8283 , n8281 , n8282 );
buf ( n8284 , n8283 );
nand ( n8285 , n8280 , n8284 );
not ( n8286 , n8285 );
not ( n8287 , n353397 );
not ( n8288 , n353861 );
and ( n8289 , n8287 , n8288 );
not ( n8290 , n7163 );
and ( n8291 , n7335 , n8290 );
nor ( n8292 , n8289 , n8291 );
nand ( n8293 , n8292 , n353934 , n353987 );
nand ( n8294 , n8292 , n353945 );
and ( n8295 , n7338 , n353866 );
nor ( n8296 , n8295 , n7336 );
nand ( n8297 , n8293 , n8294 , n8296 );
buf ( n8298 , n8297 );
not ( n8299 , n8298 );
or ( n8300 , n8286 , n8299 );
or ( n8301 , n8285 , n8298 );
nand ( n8302 , n8300 , n8301 );
buf ( n8303 , n8302 );
not ( n8304 , n8303 );
not ( n8305 , n8304 );
nand ( n8306 , n7347 , n354303 );
nand ( n8307 , n8306 , n354014 );
not ( n8308 , n8307 );
buf ( n8309 , n6605 );
buf ( n8310 , n6324 );
nand ( n8311 , n8308 , n8309 , n8310 );
not ( n8312 , n6364 );
not ( n8313 , n6605 );
not ( n8314 , n7347 );
nor ( n8315 , n8314 , n576 );
nor ( n8316 , n8313 , n8315 );
and ( n8317 , n8312 , n8316 );
nor ( n8318 , n7348 , n576 );
or ( n8319 , n8318 , n6610 );
nand ( n8320 , n8319 , n7352 );
nor ( n8321 , n8317 , n8320 );
nand ( n8322 , n8311 , n8321 );
buf ( n8323 , n8322 );
not ( n8324 , n8323 );
or ( n8325 , n8305 , n8324 );
not ( n8326 , n8322 );
not ( n8327 , n8326 );
or ( n8328 , n8327 , n8304 );
nand ( n8329 , n8325 , n8328 );
not ( n8330 , n8329 );
and ( n8331 , n604 , n8330 );
not ( n8332 , n604 );
buf ( n8333 , n8329 );
and ( n8334 , n8332 , n8333 );
or ( n8335 , n8331 , n8334 );
buf ( n356024 , n8335 );
not ( n8337 , n356024 );
or ( n8338 , n7605 , n8337 );
buf ( n356027 , n7365 );
buf ( n356028 , n355075 );
nand ( n8341 , n356027 , n356028 );
buf ( n356030 , n8341 );
buf ( n356031 , n356030 );
nand ( n8344 , n8338 , n356031 );
buf ( n356033 , n8344 );
buf ( n356034 , n356033 );
xor ( n8347 , n355291 , n356034 );
buf ( n356036 , n607 );
not ( n8349 , n356036 );
buf ( n356038 , n606 );
not ( n8351 , n356038 );
not ( n8352 , n8326 );
not ( n8353 , n8284 );
buf ( n8354 , n8297 );
not ( n8355 , n8354 );
or ( n8356 , n8353 , n8355 );
nand ( n8357 , n8356 , n8280 );
not ( n8358 , n8259 );
not ( n8359 , n8273 );
or ( n8360 , n8358 , n8359 );
nand ( n8361 , n8360 , n8260 );
xor ( n8362 , n8150 , n8248 );
and ( n8363 , n8362 , n8253 );
and ( n8364 , n8150 , n8248 );
or ( n8365 , n8363 , n8364 );
xor ( n8366 , n8162 , n8192 );
and ( n8367 , n8366 , n8202 );
and ( n8368 , n8162 , n8192 );
or ( n8369 , n8367 , n8368 );
not ( n8370 , n5751 );
not ( n8371 , n8139 );
or ( n8372 , n8370 , n8371 );
not ( n8373 , n548 );
not ( n8374 , n3996 );
or ( n8375 , n8373 , n8374 );
nand ( n8376 , n1788 , n351773 );
nand ( n8377 , n8375 , n8376 );
nand ( n8378 , n8377 , n2019 );
nand ( n8379 , n8372 , n8378 );
not ( n8380 , n8231 );
and ( n8381 , n5990 , n7270 );
not ( n8382 , n8381 );
or ( n8383 , n8380 , n8382 );
not ( n8384 , n4114 );
not ( n8385 , n5761 );
and ( n8386 , n8384 , n8385 );
and ( n8387 , n4114 , n5761 );
nor ( n8388 , n8386 , n8387 );
nand ( n8389 , n8388 , n5757 );
nand ( n8390 , n8383 , n8389 );
xor ( n8391 , n8379 , n8390 );
xnor ( n8392 , n4060 , n552 );
not ( n8393 , n4109 );
or ( n8394 , n8392 , n8393 );
nand ( n8395 , n8160 , n1871 );
nand ( n8396 , n8394 , n8395 );
xor ( n8397 , n8391 , n8396 );
xor ( n8398 , n8369 , n8397 );
nand ( n8399 , n7246 , n348119 , n5881 );
nand ( n8400 , n348153 , n8199 );
nand ( n8401 , n7247 , n5881 , n556 );
nand ( n8402 , n8399 , n8400 , n8401 );
not ( n8403 , n8122 );
not ( n8404 , n4078 );
or ( n8405 , n8403 , n8404 );
and ( n8406 , n1974 , n550 );
not ( n8407 , n1974 );
and ( n8408 , n8407 , n1880 );
nor ( n8409 , n8406 , n8408 );
not ( n8410 , n8409 );
not ( n8411 , n1875 );
or ( n8412 , n8410 , n8411 );
nand ( n8413 , n8405 , n8412 );
xor ( n8414 , n8402 , n8413 );
xor ( n8415 , n8214 , n8225 );
and ( n8416 , n8415 , n8235 );
and ( n8417 , n8214 , n8225 );
or ( n8418 , n8416 , n8417 );
xor ( n8419 , n8414 , n8418 );
xor ( n8420 , n8398 , n8419 );
not ( n8421 , n1022 );
not ( n8422 , n8211 );
or ( n8423 , n8421 , n8422 );
not ( n8424 , n1925 );
not ( n8425 , n8424 );
not ( n8426 , n554 );
not ( n8427 , n6035 );
or ( n8428 , n8426 , n8427 );
nand ( n8429 , n6034 , n348175 );
nand ( n8430 , n8428 , n8429 );
nand ( n8431 , n8425 , n8430 );
nand ( n8432 , n8423 , n8431 );
not ( n8433 , n8215 );
not ( n8434 , n544 );
not ( n8435 , n348115 );
or ( n8436 , n8434 , n8435 );
nand ( n8437 , n351755 , n7283 );
nand ( n8438 , n8436 , n8437 );
not ( n8439 , n8438 );
or ( n8440 , n8433 , n8439 );
nand ( n8441 , n8223 , n8220 );
nand ( n8442 , n8440 , n8441 );
not ( n8443 , n544 );
nor ( n8444 , n8443 , n348171 );
xor ( n8445 , n8442 , n8444 );
not ( n8446 , n348233 );
not ( n8447 , n8190 );
or ( n8448 , n8446 , n8447 );
nand ( n8449 , n8448 , n348268 );
xor ( n8450 , n8445 , n8449 );
xor ( n8451 , n8432 , n8450 );
xor ( n8452 , n8116 , n8131 );
and ( n8453 , n8452 , n8143 );
and ( n8454 , n8116 , n8131 );
or ( n8455 , n8453 , n8454 );
xor ( n8456 , n8451 , n8455 );
xor ( n8457 , n8213 , n8236 );
and ( n8458 , n8457 , n8241 );
and ( n8459 , n8213 , n8236 );
or ( n8460 , n8458 , n8459 );
xor ( n8461 , n8456 , n8460 );
xor ( n8462 , n8115 , n8144 );
and ( n8463 , n8462 , n8149 );
and ( n8464 , n8115 , n8144 );
or ( n8465 , n8463 , n8464 );
xor ( n8466 , n8461 , n8465 );
xor ( n8467 , n8420 , n8466 );
xor ( n8468 , n8203 , n8242 );
and ( n8469 , n8468 , n8247 );
and ( n8470 , n8203 , n8242 );
or ( n8471 , n8469 , n8470 );
xor ( n8472 , n8467 , n8471 );
nor ( n8473 , n8365 , n8472 );
not ( n8474 , n8473 );
not ( n8475 , n8472 );
not ( n8476 , n8365 );
nor ( n8477 , n8475 , n8476 );
not ( n8478 , n8477 );
and ( n8479 , n8474 , n8478 );
and ( n8480 , n8361 , n8479 );
not ( n8481 , n8361 );
not ( n8482 , n8479 );
and ( n8483 , n8481 , n8482 );
nor ( n8484 , n8480 , n8483 );
not ( n8485 , n8484 );
not ( n8486 , n8053 );
nand ( n8487 , n355773 , n8091 , n355786 );
not ( n8488 , n8487 );
or ( n8489 , n8486 , n8488 );
nand ( n8490 , n8489 , n8054 );
xor ( n8491 , n355299 , n355338 );
and ( n8492 , n8491 , n355348 );
and ( n8493 , n355299 , n355338 );
or ( n8494 , n8492 , n8493 );
buf ( n356183 , n8494 );
buf ( n356184 , n574 );
buf ( n356185 , n558 );
buf ( n356186 , n560 );
nand ( n8499 , n356185 , n356186 );
buf ( n356188 , n8499 );
buf ( n356189 , n356188 );
xor ( n8502 , n356184 , n356189 );
not ( n8503 , n5407 );
buf ( n356192 , n556 );
buf ( n356193 , n560 );
xor ( n8506 , n356192 , n356193 );
buf ( n356195 , n8506 );
not ( n8508 , n356195 );
or ( n8509 , n8503 , n8508 );
nand ( n8510 , n354458 , n7775 );
nand ( n8511 , n8509 , n8510 );
buf ( n356200 , n8511 );
xnor ( n8513 , n8502 , n356200 );
buf ( n356202 , n8513 );
buf ( n356203 , n356202 );
not ( n8516 , n356203 );
buf ( n356205 , n8516 );
buf ( n356206 , n356205 );
not ( n8519 , n356206 );
buf ( n356208 , n355388 );
not ( n8521 , n356208 );
buf ( n356210 , n347737 );
not ( n8523 , n356210 );
or ( n8524 , n8521 , n8523 );
buf ( n356213 , n347382 );
buf ( n356214 , n544 );
buf ( n356215 , n572 );
xor ( n8528 , n356214 , n356215 );
buf ( n356217 , n8528 );
buf ( n356218 , n356217 );
nand ( n8531 , n356213 , n356218 );
buf ( n356220 , n8531 );
buf ( n356221 , n356220 );
nand ( n8534 , n8524 , n356221 );
buf ( n356223 , n8534 );
buf ( n356224 , n355423 );
not ( n8537 , n356224 );
buf ( n356226 , n348467 );
not ( n8539 , n356226 );
or ( n8540 , n8537 , n8539 );
buf ( n356229 , n348473 );
buf ( n356230 , n546 );
buf ( n356231 , n570 );
xor ( n8544 , n356230 , n356231 );
buf ( n356233 , n8544 );
buf ( n356234 , n356233 );
nand ( n8547 , n356229 , n356234 );
buf ( n356236 , n8547 );
buf ( n356237 , n356236 );
nand ( n8550 , n8540 , n356237 );
buf ( n356239 , n8550 );
xor ( n8552 , n356223 , n356239 );
buf ( n356241 , n355489 );
not ( n8554 , n356241 );
buf ( n356243 , n350874 );
not ( n8556 , n356243 );
or ( n8557 , n8554 , n8556 );
buf ( n356246 , n2550 );
xor ( n8559 , n566 , n550 );
buf ( n356248 , n8559 );
nand ( n8561 , n356246 , n356248 );
buf ( n356250 , n8561 );
buf ( n356251 , n356250 );
nand ( n8564 , n8557 , n356251 );
buf ( n356253 , n8564 );
not ( n8566 , n356253 );
and ( n8567 , n8552 , n8566 );
not ( n8568 , n8552 );
and ( n8569 , n8568 , n356253 );
nor ( n8570 , n8567 , n8569 );
buf ( n356259 , n8570 );
not ( n8572 , n356259 );
or ( n8573 , n8519 , n8572 );
not ( n8574 , n8570 );
nand ( n8575 , n8574 , n356202 );
buf ( n356264 , n8575 );
nand ( n8577 , n8573 , n356264 );
buf ( n356266 , n8577 );
buf ( n356267 , n356266 );
xor ( n8580 , n355304 , n355318 );
and ( n8581 , n8580 , n7648 );
and ( n8582 , n355304 , n355318 );
or ( n8583 , n8581 , n8582 );
buf ( n356272 , n8583 );
not ( n8585 , n356272 );
buf ( n356274 , n8585 );
buf ( n356275 , n356274 );
and ( n8588 , n356267 , n356275 );
not ( n8589 , n356267 );
buf ( n356278 , n8583 );
and ( n8591 , n8589 , n356278 );
nor ( n8592 , n8588 , n8591 );
buf ( n356281 , n8592 );
and ( n8594 , n356183 , n356281 );
not ( n8595 , n356183 );
buf ( n356284 , n356281 );
not ( n8597 , n356284 );
buf ( n356286 , n8597 );
and ( n8599 , n8595 , n356286 );
or ( n8600 , n8594 , n8599 );
buf ( n356289 , n355409 );
not ( n8602 , n356289 );
nor ( n8603 , n4625 , n352312 );
buf ( n8604 , n8603 );
buf ( n356293 , n8604 );
not ( n8606 , n356293 );
or ( n8607 , n8602 , n8606 );
buf ( n356296 , n352295 );
buf ( n356297 , n554 );
buf ( n356298 , n562 );
xor ( n8611 , n356297 , n356298 );
buf ( n356300 , n8611 );
buf ( n356301 , n356300 );
nand ( n8614 , n356296 , n356301 );
buf ( n356303 , n8614 );
buf ( n356304 , n356303 );
nand ( n8617 , n8607 , n356304 );
buf ( n356306 , n8617 );
buf ( n356307 , n355440 );
not ( n8620 , n356307 );
buf ( n356309 , n351330 );
not ( n8622 , n356309 );
or ( n8623 , n8620 , n8622 );
buf ( n356312 , n3650 );
buf ( n356313 , n552 );
buf ( n356314 , n564 );
xor ( n8627 , n356313 , n356314 );
buf ( n356316 , n8627 );
buf ( n356317 , n356316 );
nand ( n8630 , n356312 , n356317 );
buf ( n356319 , n8630 );
buf ( n356320 , n356319 );
nand ( n8633 , n8623 , n356320 );
buf ( n356322 , n8633 );
xor ( n8635 , n356306 , n356322 );
buf ( n356324 , n7787 );
not ( n8637 , n356324 );
buf ( n356326 , n2236 );
not ( n8639 , n356326 );
or ( n8640 , n8637 , n8639 );
buf ( n356329 , n349933 );
buf ( n356330 , n548 );
buf ( n356331 , n568 );
xor ( n8644 , n356330 , n356331 );
buf ( n356333 , n8644 );
buf ( n356334 , n356333 );
nand ( n8647 , n356329 , n356334 );
buf ( n356336 , n8647 );
buf ( n356337 , n356336 );
nand ( n8650 , n8640 , n356337 );
buf ( n356339 , n8650 );
xor ( n8652 , n8635 , n356339 );
buf ( n356341 , n355394 );
not ( n8654 , n356341 );
buf ( n356343 , n355364 );
buf ( n356344 , n355371 );
nand ( n8657 , n356343 , n356344 );
buf ( n356346 , n8657 );
buf ( n356347 , n356346 );
not ( n8660 , n356347 );
or ( n8661 , n8654 , n8660 );
buf ( n356350 , n355367 );
buf ( n356351 , n355376 );
nand ( n8664 , n356350 , n356351 );
buf ( n356353 , n8664 );
buf ( n356354 , n356353 );
nand ( n8667 , n8661 , n356354 );
buf ( n356356 , n8667 );
buf ( n356357 , n356356 );
or ( n8670 , n7725 , n355446 );
nand ( n8671 , n8670 , n355429 );
buf ( n356360 , n8671 );
nand ( n8673 , n355446 , n7725 );
buf ( n356362 , n8673 );
nand ( n8675 , n356360 , n356362 );
buf ( n356364 , n8675 );
buf ( n356365 , n356364 );
xor ( n8678 , n356357 , n356365 );
xor ( n8679 , n355468 , n355478 );
and ( n8680 , n8679 , n355496 );
and ( n8681 , n355468 , n355478 );
or ( n8682 , n8680 , n8681 );
buf ( n356371 , n8682 );
buf ( n356372 , n356371 );
xor ( n8685 , n8678 , n356372 );
buf ( n356374 , n8685 );
xor ( n8687 , n8652 , n356374 );
not ( n8688 , n355450 );
not ( n8689 , n7711 );
or ( n8690 , n8688 , n8689 );
not ( n8691 , n7712 );
not ( n8692 , n7759 );
or ( n8693 , n8691 , n8692 );
nand ( n8694 , n8693 , n355498 );
nand ( n8695 , n8690 , n8694 );
xnor ( n8696 , n8687 , n8695 );
buf ( n356385 , n8696 );
buf ( n8698 , n356385 );
buf ( n356387 , n8698 );
xor ( n8700 , n8600 , n356387 );
buf ( n356389 , n8700 );
buf ( n356390 , n355519 );
not ( n8703 , n356390 );
buf ( n356392 , n355536 );
not ( n8705 , n356392 );
or ( n8706 , n8703 , n8705 );
buf ( n356395 , n355536 );
buf ( n356396 , n355519 );
or ( n8709 , n356395 , n356396 );
buf ( n356398 , n355728 );
nand ( n8711 , n8709 , n356398 );
buf ( n356400 , n8711 );
buf ( n356401 , n356400 );
nand ( n8714 , n8706 , n356401 );
buf ( n356403 , n8714 );
buf ( n356404 , n356403 );
xor ( n8717 , n356389 , n356404 );
buf ( n356406 , n355501 );
not ( n8719 , n356406 );
buf ( n356408 , n355355 );
not ( n8721 , n356408 );
or ( n8722 , n8719 , n8721 );
buf ( n356411 , n355355 );
buf ( n356412 , n355501 );
or ( n8725 , n356411 , n356412 );
buf ( n356414 , n355350 );
nand ( n8727 , n8725 , n356414 );
buf ( n356416 , n8727 );
buf ( n356417 , n356416 );
nand ( n8730 , n8722 , n356417 );
buf ( n356419 , n8730 );
buf ( n356420 , n356419 );
xor ( n8733 , n355672 , n355678 );
and ( n8734 , n8733 , n355726 );
and ( n8735 , n355672 , n355678 );
or ( n8736 , n8734 , n8735 );
buf ( n356425 , n8736 );
buf ( n356426 , n356425 );
xor ( n8739 , n356420 , n356426 );
buf ( n356428 , n558 );
buf ( n356429 , n576 );
and ( n8742 , n356428 , n356429 );
buf ( n356431 , n8742 );
buf ( n356432 , n356431 );
buf ( n356433 , n347697 );
xor ( n8746 , n356432 , n356433 );
buf ( n356435 , n355623 );
not ( n8748 , n356435 );
buf ( n356437 , n354687 );
buf ( n356438 , n353193 );
nor ( n8751 , n356437 , n356438 );
buf ( n356440 , n8751 );
buf ( n356441 , n356440 );
not ( n8754 , n356441 );
or ( n8755 , n8748 , n8754 );
buf ( n356444 , n353193 );
buf ( n8757 , n356444 );
buf ( n356446 , n8757 );
buf ( n356447 , n356446 );
xor ( n8760 , n576 , n556 );
buf ( n356449 , n8760 );
nand ( n8762 , n356447 , n356449 );
buf ( n356451 , n8762 );
buf ( n356452 , n356451 );
nand ( n8765 , n8755 , n356452 );
buf ( n356454 , n8765 );
buf ( n356455 , n356454 );
xor ( n8768 , n8746 , n356455 );
buf ( n356457 , n8768 );
buf ( n356458 , n356457 );
buf ( n356459 , n355640 );
not ( n8772 , n356459 );
buf ( n356461 , n350699 );
not ( n8774 , n356461 );
or ( n8775 , n8772 , n8774 );
buf ( n356464 , n350705 );
xor ( n8777 , n582 , n550 );
buf ( n356466 , n8777 );
nand ( n8779 , n356464 , n356466 );
buf ( n356468 , n8779 );
buf ( n356469 , n356468 );
nand ( n8782 , n8775 , n356469 );
buf ( n356471 , n8782 );
buf ( n356472 , n356471 );
not ( n8785 , n356472 );
buf ( n356474 , n8785 );
buf ( n356475 , n355562 );
not ( n8788 , n356475 );
buf ( n356477 , n347671 );
not ( n8790 , n356477 );
or ( n8791 , n8788 , n8790 );
buf ( n356480 , n347530 );
buf ( n356481 , n546 );
buf ( n356482 , n586 );
xor ( n8795 , n356481 , n356482 );
buf ( n356484 , n8795 );
buf ( n356485 , n356484 );
nand ( n8798 , n356480 , n356485 );
buf ( n356487 , n8798 );
buf ( n356488 , n356487 );
nand ( n8801 , n8791 , n356488 );
buf ( n356490 , n8801 );
not ( n8803 , n356490 );
not ( n8804 , n355603 );
not ( n8805 , n347554 );
or ( n8806 , n8804 , n8805 );
buf ( n356495 , n544 );
buf ( n356496 , n588 );
xor ( n8809 , n356495 , n356496 );
buf ( n356498 , n8809 );
buf ( n356499 , n356498 );
buf ( n356500 , n347568 );
nand ( n8813 , n356499 , n356500 );
buf ( n356502 , n8813 );
nand ( n8815 , n8806 , n356502 );
not ( n8816 , n8815 );
not ( n8817 , n8816 );
or ( n8818 , n8803 , n8817 );
or ( n8819 , n8816 , n356490 );
nand ( n8820 , n8818 , n8819 );
xnor ( n8821 , n356474 , n8820 );
buf ( n356510 , n8821 );
xor ( n8823 , n356458 , n356510 );
xor ( n8824 , n355707 , n355712 );
and ( n8825 , n8824 , n355720 );
and ( n8826 , n355707 , n355712 );
or ( n8827 , n8825 , n8826 );
buf ( n356516 , n8827 );
buf ( n356517 , n356516 );
xor ( n8830 , n8823 , n356517 );
buf ( n356519 , n8830 );
buf ( n356520 , n356519 );
xor ( n8833 , n355685 , n355703 );
and ( n8834 , n8833 , n355723 );
and ( n8835 , n355685 , n355703 );
or ( n8836 , n8834 , n8835 );
buf ( n356525 , n8836 );
buf ( n356526 , n356525 );
xor ( n8839 , n356520 , n356526 );
buf ( n356528 , n7860 );
not ( n8841 , n356528 );
buf ( n356530 , n5162 );
not ( n8843 , n356530 );
or ( n8844 , n8841 , n8843 );
buf ( n356533 , n354788 );
xor ( n8846 , n578 , n554 );
buf ( n356535 , n8846 );
nand ( n8848 , n356533 , n356535 );
buf ( n356537 , n8848 );
buf ( n356538 , n356537 );
nand ( n8851 , n8844 , n356538 );
buf ( n356540 , n8851 );
buf ( n356541 , n356540 );
buf ( n356542 , n7884 );
not ( n8855 , n356542 );
buf ( n356544 , n3870 );
not ( n8857 , n356544 );
or ( n8858 , n8855 , n8857 );
buf ( n356547 , n351559 );
xor ( n8860 , n580 , n552 );
buf ( n356549 , n8860 );
nand ( n8862 , n356547 , n356549 );
buf ( n356551 , n8862 );
buf ( n356552 , n356551 );
nand ( n8865 , n8858 , n356552 );
buf ( n356554 , n8865 );
buf ( n356555 , n356554 );
xor ( n8868 , n356541 , n356555 );
buf ( n356557 , n355658 );
not ( n8870 , n356557 );
buf ( n356559 , n2471 );
not ( n8872 , n356559 );
or ( n8873 , n8870 , n8872 );
buf ( n356562 , n348617 );
xor ( n8875 , n584 , n548 );
buf ( n356564 , n8875 );
nand ( n8877 , n356562 , n356564 );
buf ( n356566 , n8877 );
buf ( n356567 , n356566 );
nand ( n8880 , n8873 , n356567 );
buf ( n356569 , n8880 );
buf ( n356570 , n356569 );
not ( n8883 , n356570 );
buf ( n356572 , n8883 );
buf ( n356573 , n356572 );
xor ( n8886 , n8868 , n356573 );
buf ( n356575 , n8886 );
buf ( n356576 , n356575 );
buf ( n356577 , n7923 );
not ( n8890 , n356577 );
buf ( n356579 , n355670 );
nand ( n8892 , n8890 , n356579 );
buf ( n356581 , n8892 );
buf ( n356582 , n356581 );
not ( n8895 , n7923 );
not ( n8896 , n355667 );
or ( n8897 , n8895 , n8896 );
nand ( n8898 , n8897 , n7889 );
buf ( n356587 , n8898 );
nand ( n8900 , n356582 , n356587 );
buf ( n356589 , n8900 );
buf ( n356590 , n356589 );
xor ( n8903 , n356576 , n356590 );
buf ( n356592 , n355610 );
not ( n8905 , n356592 );
buf ( n356594 , n355589 );
not ( n8907 , n356594 );
buf ( n356596 , n355593 );
nand ( n8909 , n8907 , n356596 );
buf ( n356598 , n8909 );
buf ( n356599 , n356598 );
not ( n8912 , n356599 );
or ( n8913 , n8905 , n8912 );
buf ( n356602 , n355593 );
not ( n8915 , n356602 );
buf ( n356604 , n355589 );
nand ( n8917 , n8915 , n356604 );
buf ( n356606 , n8917 );
buf ( n356607 , n356606 );
nand ( n8920 , n8913 , n356607 );
buf ( n356609 , n8920 );
buf ( n356610 , n356609 );
buf ( n356611 , n355554 );
buf ( n356612 , n7888 );
or ( n8925 , n356611 , n356612 );
buf ( n356614 , n7878 );
nand ( n8927 , n8925 , n356614 );
buf ( n356616 , n8927 );
buf ( n356617 , n356616 );
buf ( n356618 , n355554 );
buf ( n356619 , n7888 );
nand ( n8932 , n356618 , n356619 );
buf ( n356621 , n8932 );
buf ( n356622 , n356621 );
nand ( n8935 , n356617 , n356622 );
buf ( n356624 , n8935 );
buf ( n356625 , n356624 );
xor ( n8938 , n356610 , n356625 );
not ( n8939 , n355646 );
not ( n8940 , n355629 );
or ( n8941 , n8939 , n8940 );
buf ( n356630 , n355646 );
buf ( n356631 , n355629 );
nor ( n8944 , n356630 , n356631 );
buf ( n356633 , n8944 );
buf ( n356634 , n355664 );
not ( n8947 , n356634 );
buf ( n356636 , n8947 );
or ( n8949 , n356633 , n356636 );
nand ( n8950 , n8941 , n8949 );
buf ( n356639 , n8950 );
xor ( n8952 , n8938 , n356639 );
buf ( n356641 , n8952 );
buf ( n356642 , n356641 );
xor ( n8955 , n8903 , n356642 );
buf ( n356644 , n8955 );
buf ( n356645 , n356644 );
xor ( n8958 , n8839 , n356645 );
buf ( n356647 , n8958 );
buf ( n356648 , n356647 );
xor ( n8961 , n8739 , n356648 );
buf ( n356650 , n8961 );
buf ( n356651 , n356650 );
xor ( n8964 , n8717 , n356651 );
buf ( n356653 , n8964 );
not ( n8966 , n8041 );
not ( n8967 , n355509 );
nand ( n8968 , n8967 , n7815 );
not ( n8969 , n8968 );
or ( n8970 , n8966 , n8969 );
nand ( n8971 , n7814 , n355509 );
nand ( n8972 , n8970 , n8971 );
nor ( n8973 , n356653 , n8972 );
not ( n8974 , n8973 );
buf ( n356663 , n356653 );
buf ( n356664 , n8972 );
nand ( n8977 , n356663 , n356664 );
buf ( n356666 , n8977 );
nand ( n8979 , n8974 , n356666 );
xor ( n8980 , n8490 , n8979 );
not ( n8981 , n8980 );
nand ( n8982 , n8485 , n8981 );
nand ( n8983 , n8484 , n8980 );
and ( n8984 , n8982 , n8983 );
and ( n8985 , n8357 , n8984 );
not ( n8986 , n8357 );
not ( n8987 , n8984 );
and ( n8988 , n8986 , n8987 );
nor ( n8989 , n8985 , n8988 );
buf ( n8990 , n8989 );
nand ( n8991 , n8990 , n8303 );
not ( n8992 , n8991 );
nand ( n8993 , n8352 , n8992 );
nor ( n8994 , n8254 , n8258 );
nor ( n8995 , n8473 , n8994 );
not ( n8996 , n8995 );
not ( n8997 , n8272 );
or ( n8998 , n8996 , n8997 );
not ( n8999 , n8472 );
not ( n9000 , n8365 );
and ( n9001 , n8999 , n9000 );
nand ( n9002 , n8254 , n8258 );
nor ( n9003 , n9001 , n9002 );
nor ( n9004 , n9003 , n8477 );
nand ( n9005 , n8998 , n9004 );
not ( n9006 , n9005 );
xor ( n9007 , n8379 , n8390 );
and ( n9008 , n9007 , n8396 );
and ( n9009 , n8379 , n8390 );
or ( n9010 , n9008 , n9009 );
xor ( n9011 , n8402 , n8413 );
and ( n9012 , n9011 , n8418 );
and ( n9013 , n8402 , n8413 );
or ( n9014 , n9012 , n9013 );
xor ( n9015 , n9010 , n9014 );
not ( n9016 , n1916 );
not ( n9017 , n7245 );
not ( n9018 , n9017 );
not ( n9019 , n9018 );
or ( n9020 , n9016 , n9019 );
not ( n9021 , n556 );
not ( n9022 , n8184 );
or ( n9023 , n9021 , n9022 );
nand ( n9024 , n348119 , n8183 );
nand ( n9025 , n9023 , n9024 );
and ( n9026 , n9025 , n348088 );
and ( n9027 , n7246 , n1919 );
nor ( n9028 , n9026 , n9027 );
nand ( n9029 , n9020 , n9028 );
not ( n9030 , n4078 );
not ( n9031 , n8409 );
or ( n9032 , n9030 , n9031 );
and ( n9033 , n2071 , n550 );
not ( n9034 , n2071 );
and ( n9035 , n9034 , n1880 );
nor ( n9036 , n9033 , n9035 );
nand ( n9037 , n9036 , n1875 );
nand ( n9038 , n9032 , n9037 );
xor ( n9039 , n9029 , n9038 );
not ( n9040 , n1022 );
not ( n9041 , n8430 );
or ( n9042 , n9040 , n9041 );
xor ( n9043 , n554 , n6081 );
nand ( n9044 , n1925 , n9043 );
nand ( n9045 , n9042 , n9044 );
xor ( n9046 , n9039 , n9045 );
xor ( n9047 , n9015 , n9046 );
xor ( n9048 , n8456 , n8460 );
and ( n9049 , n9048 , n8465 );
and ( n9050 , n8456 , n8460 );
or ( n9051 , n9049 , n9050 );
xor ( n9052 , n9047 , n9051 );
xor ( n9053 , n8432 , n8450 );
and ( n9054 , n9053 , n8455 );
and ( n9055 , n8432 , n8450 );
or ( n9056 , n9054 , n9055 );
xor ( n9057 , n8442 , n8444 );
and ( n9058 , n9057 , n8449 );
and ( n9059 , n8442 , n8444 );
or ( n9060 , n9058 , n9059 );
not ( n9061 , n348234 );
nand ( n9062 , n9061 , n348268 );
not ( n9063 , n9062 );
not ( n9064 , n348146 );
nand ( n9065 , n9064 , n544 );
not ( n9066 , n9065 );
or ( n9067 , n9063 , n9066 );
or ( n9068 , n9065 , n9062 );
nand ( n9069 , n9067 , n9068 );
not ( n9070 , n8215 );
not ( n9071 , n966 );
xor ( n9072 , n544 , n9071 );
not ( n9073 , n9072 );
or ( n9074 , n9070 , n9073 );
nand ( n9075 , n8438 , n8223 );
nand ( n9076 , n9074 , n9075 );
xor ( n9077 , n9069 , n9076 );
xor ( n9078 , n9060 , n9077 );
not ( n9079 , n5751 );
not ( n9080 , n8377 );
or ( n9081 , n9079 , n9080 );
not ( n9082 , n548 );
not ( n9083 , n1844 );
or ( n9084 , n9082 , n9083 );
nand ( n9085 , n1843 , n351773 );
nand ( n9086 , n9084 , n9085 );
nand ( n9087 , n9086 , n2019 );
nand ( n9088 , n9081 , n9087 );
not ( n9089 , n546 );
not ( n9090 , n2002 );
or ( n9091 , n9089 , n9090 );
nand ( n9092 , n997 , n5761 );
nand ( n9093 , n9091 , n9092 );
not ( n9094 , n9093 );
not ( n9095 , n5757 );
or ( n9096 , n9094 , n9095 );
nand ( n9097 , n8388 , n8381 );
nand ( n9098 , n9096 , n9097 );
xor ( n9099 , n9088 , n9098 );
and ( n9100 , n552 , n5937 );
not ( n9101 , n552 );
and ( n9102 , n9101 , n353618 );
or ( n9103 , n9100 , n9102 );
not ( n9104 , n9103 );
not ( n9105 , n1011 );
or ( n9106 , n9104 , n9105 );
not ( n9107 , n8392 );
nand ( n9108 , n9107 , n1871 );
nand ( n9109 , n9106 , n9108 );
xor ( n9110 , n9099 , n9109 );
xor ( n9111 , n9078 , n9110 );
xor ( n9112 , n9056 , n9111 );
xor ( n9113 , n8369 , n8397 );
and ( n9114 , n9113 , n8419 );
and ( n9115 , n8369 , n8397 );
or ( n9116 , n9114 , n9115 );
xor ( n9117 , n9112 , n9116 );
xor ( n9118 , n9052 , n9117 );
xor ( n9119 , n8420 , n8466 );
and ( n9120 , n9119 , n8471 );
and ( n9121 , n8420 , n8466 );
or ( n9122 , n9120 , n9121 );
nor ( n9123 , n9118 , n9122 );
not ( n9124 , n9123 );
nand ( n9125 , n9118 , n9122 );
buf ( n9126 , n9125 );
nand ( n9127 , n9124 , n9126 );
and ( n9128 , n9006 , n9127 );
not ( n9129 , n9006 );
not ( n9130 , n9127 );
and ( n9131 , n9129 , n9130 );
nor ( n9132 , n9128 , n9131 );
not ( n9133 , n9132 );
nor ( n9134 , n8973 , n8052 );
not ( n9135 , n9134 );
not ( n9136 , n8487 );
or ( n9137 , n9135 , n9136 );
or ( n9138 , n8054 , n8973 );
nand ( n9139 , n9138 , n356666 );
buf ( n356828 , n9139 );
not ( n9141 , n356828 );
buf ( n356830 , n9141 );
nand ( n9143 , n9137 , n356830 );
buf ( n356832 , n557 );
buf ( n356833 , n560 );
and ( n9146 , n356832 , n356833 );
buf ( n356835 , n9146 );
buf ( n356836 , n356835 );
buf ( n356837 , n8559 );
not ( n9150 , n356837 );
buf ( n356839 , n2851 );
not ( n9152 , n356839 );
or ( n9153 , n9150 , n9152 );
buf ( n356842 , n2550 );
xor ( n9155 , n566 , n549 );
buf ( n356844 , n9155 );
nand ( n9157 , n356842 , n356844 );
buf ( n356846 , n9157 );
buf ( n356847 , n356846 );
nand ( n9160 , n9153 , n356847 );
buf ( n356849 , n9160 );
buf ( n356850 , n356849 );
xor ( n9163 , n356836 , n356850 );
buf ( n356852 , n356233 );
not ( n9165 , n356852 );
buf ( n356854 , n347344 );
not ( n9167 , n356854 );
or ( n9168 , n9165 , n9167 );
buf ( n356857 , n347350 );
buf ( n356858 , n545 );
buf ( n356859 , n570 );
xor ( n9172 , n356858 , n356859 );
buf ( n356861 , n9172 );
buf ( n356862 , n356861 );
nand ( n9175 , n356857 , n356862 );
buf ( n356864 , n9175 );
buf ( n356865 , n356864 );
nand ( n9178 , n9168 , n356865 );
buf ( n356867 , n9178 );
buf ( n356868 , n356867 );
xor ( n9181 , n9163 , n356868 );
buf ( n356870 , n9181 );
buf ( n356871 , n356870 );
buf ( n356872 , n356195 );
not ( n9185 , n356872 );
buf ( n9186 , n354458 );
buf ( n356875 , n9186 );
not ( n9188 , n356875 );
or ( n9189 , n9185 , n9188 );
buf ( n356878 , n5407 );
buf ( n356879 , n555 );
buf ( n356880 , n560 );
xor ( n9193 , n356879 , n356880 );
buf ( n356882 , n9193 );
buf ( n356883 , n356882 );
nand ( n9196 , n356878 , n356883 );
buf ( n356885 , n9196 );
buf ( n356886 , n356885 );
nand ( n9199 , n9189 , n356886 );
buf ( n356888 , n9199 );
buf ( n356889 , n356888 );
buf ( n356890 , n356339 );
xor ( n9203 , n356889 , n356890 );
buf ( n356892 , n356217 );
not ( n9205 , n356892 );
buf ( n356894 , n347378 );
not ( n9207 , n356894 );
or ( n9208 , n9205 , n9207 );
buf ( n356897 , n572 );
buf ( n356898 , n347382 );
nand ( n9211 , n356897 , n356898 );
buf ( n356900 , n9211 );
buf ( n356901 , n356900 );
nand ( n9214 , n9208 , n356901 );
buf ( n356903 , n9214 );
buf ( n356904 , n356903 );
not ( n9217 , n356904 );
buf ( n356906 , n9217 );
buf ( n356907 , n356906 );
xor ( n9220 , n9203 , n356907 );
buf ( n356909 , n9220 );
buf ( n356910 , n356909 );
xor ( n9223 , n356871 , n356910 );
xor ( n9224 , n356357 , n356365 );
and ( n9225 , n9224 , n356372 );
and ( n9226 , n356357 , n356365 );
or ( n9227 , n9225 , n9226 );
buf ( n356916 , n9227 );
buf ( n356917 , n356916 );
xor ( n9230 , n9223 , n356917 );
buf ( n356919 , n9230 );
buf ( n356920 , n356919 );
buf ( n356921 , n8652 );
not ( n9234 , n356921 );
buf ( n356923 , n356374 );
not ( n9236 , n356923 );
buf ( n356925 , n9236 );
buf ( n356926 , n356925 );
not ( n9239 , n356926 );
or ( n9240 , n9234 , n9239 );
buf ( n356929 , n8695 );
nand ( n9242 , n9240 , n356929 );
buf ( n356931 , n9242 );
buf ( n356932 , n356931 );
buf ( n356933 , n8652 );
not ( n9246 , n356933 );
buf ( n356935 , n356374 );
nand ( n9248 , n9246 , n356935 );
buf ( n356937 , n9248 );
buf ( n356938 , n356937 );
nand ( n9251 , n356932 , n356938 );
buf ( n356940 , n9251 );
buf ( n356941 , n356940 );
xor ( n9254 , n356920 , n356941 );
buf ( n356943 , n356322 );
buf ( n356944 , n356306 );
nor ( n9257 , n356943 , n356944 );
buf ( n356946 , n9257 );
buf ( n356947 , n356946 );
buf ( n356948 , n356339 );
or ( n9261 , n356947 , n356948 );
buf ( n356950 , n356322 );
buf ( n356951 , n356306 );
nand ( n9264 , n356950 , n356951 );
buf ( n356953 , n9264 );
buf ( n356954 , n356953 );
nand ( n9267 , n9261 , n356954 );
buf ( n356956 , n9267 );
buf ( n356957 , n356956 );
buf ( n356958 , n356188 );
buf ( n356959 , n574 );
nand ( n9272 , n356958 , n356959 );
buf ( n356961 , n9272 );
not ( n9274 , n356961 );
not ( n9275 , n8511 );
or ( n9276 , n9274 , n9275 );
or ( n9277 , n356188 , n574 );
nand ( n9278 , n9276 , n9277 );
buf ( n356967 , n9278 );
buf ( n356968 , n356239 );
not ( n9281 , n356968 );
buf ( n356970 , n356223 );
not ( n9283 , n356970 );
or ( n9284 , n9281 , n9283 );
or ( n9285 , n356239 , n356223 );
nand ( n9286 , n9285 , n356253 );
buf ( n356975 , n9286 );
nand ( n9288 , n9284 , n356975 );
buf ( n356977 , n9288 );
buf ( n356978 , n356977 );
xor ( n9291 , n356967 , n356978 );
buf ( n356980 , n356316 );
not ( n9293 , n356980 );
buf ( n356982 , n4490 );
not ( n9295 , n356982 );
or ( n9296 , n9293 , n9295 );
xor ( n9297 , n551 , n564 );
nand ( n9298 , n3650 , n9297 );
buf ( n356987 , n9298 );
nand ( n9300 , n9296 , n356987 );
buf ( n356989 , n9300 );
buf ( n356990 , n356989 );
buf ( n356991 , n356300 );
not ( n9304 , n356991 );
buf ( n356993 , n8603 );
not ( n9306 , n356993 );
or ( n9307 , n9304 , n9306 );
buf ( n356996 , n352295 );
buf ( n356997 , n553 );
buf ( n356998 , n562 );
xor ( n9311 , n356997 , n356998 );
buf ( n357000 , n9311 );
buf ( n357001 , n357000 );
nand ( n9314 , n356996 , n357001 );
buf ( n357003 , n9314 );
buf ( n357004 , n357003 );
nand ( n9317 , n9307 , n357004 );
buf ( n357006 , n9317 );
buf ( n357007 , n357006 );
xor ( n9320 , n356990 , n357007 );
buf ( n357009 , n356333 );
not ( n9322 , n357009 );
buf ( n357011 , n2236 );
not ( n9324 , n357011 );
or ( n9325 , n9322 , n9324 );
buf ( n357014 , n2579 );
buf ( n357015 , n547 );
buf ( n357016 , n568 );
xor ( n9329 , n357015 , n357016 );
buf ( n357018 , n9329 );
buf ( n357019 , n357018 );
nand ( n9332 , n357014 , n357019 );
buf ( n357021 , n9332 );
buf ( n357022 , n357021 );
nand ( n9335 , n9325 , n357022 );
buf ( n357024 , n9335 );
buf ( n357025 , n357024 );
xor ( n9338 , n9320 , n357025 );
buf ( n357027 , n9338 );
buf ( n357028 , n357027 );
xor ( n9341 , n9291 , n357028 );
buf ( n357030 , n9341 );
buf ( n357031 , n357030 );
xor ( n9344 , n356957 , n357031 );
or ( n9345 , n8583 , n356205 );
nand ( n9346 , n9345 , n8574 );
buf ( n357035 , n9346 );
buf ( n357036 , n8583 );
buf ( n357037 , n356205 );
nand ( n9350 , n357036 , n357037 );
buf ( n357039 , n9350 );
buf ( n357040 , n357039 );
nand ( n9353 , n357035 , n357040 );
buf ( n357042 , n9353 );
buf ( n357043 , n357042 );
xor ( n9356 , n9344 , n357043 );
buf ( n357045 , n9356 );
buf ( n357046 , n357045 );
xor ( n9359 , n9254 , n357046 );
buf ( n357048 , n9359 );
buf ( n357049 , n357048 );
xor ( n9362 , n356420 , n356426 );
and ( n9363 , n9362 , n356648 );
and ( n9364 , n356420 , n356426 );
or ( n9365 , n9363 , n9364 );
buf ( n357054 , n9365 );
buf ( n357055 , n357054 );
xor ( n9368 , n357049 , n357055 );
not ( n9369 , n8696 );
buf ( n357058 , n356183 );
not ( n9371 , n357058 );
buf ( n357060 , n9371 );
nand ( n9373 , n357060 , n356281 );
not ( n9374 , n9373 );
or ( n9375 , n9369 , n9374 );
nand ( n9376 , n356286 , n356183 );
nand ( n9377 , n9375 , n9376 );
buf ( n357066 , n9377 );
xor ( n9379 , n356520 , n356526 );
and ( n9380 , n9379 , n356645 );
and ( n9381 , n356520 , n356526 );
or ( n9382 , n9380 , n9381 );
buf ( n357071 , n9382 );
buf ( n357072 , n357071 );
xor ( n9385 , n357066 , n357072 );
buf ( n357074 , n356484 );
not ( n9387 , n357074 );
buf ( n357076 , n347671 );
not ( n9389 , n357076 );
or ( n9390 , n9387 , n9389 );
buf ( n357079 , n347530 );
buf ( n357080 , n545 );
buf ( n357081 , n586 );
xor ( n9394 , n357080 , n357081 );
buf ( n357083 , n9394 );
buf ( n357084 , n357083 );
nand ( n9397 , n357079 , n357084 );
buf ( n357086 , n9397 );
buf ( n357087 , n357086 );
nand ( n9400 , n9390 , n357087 );
buf ( n357089 , n9400 );
buf ( n357090 , n357089 );
buf ( n357091 , n557 );
buf ( n357092 , n576 );
nand ( n9405 , n357091 , n357092 );
buf ( n357094 , n9405 );
buf ( n357095 , n357094 );
not ( n9408 , n357095 );
buf ( n357097 , n9408 );
buf ( n357098 , n357097 );
and ( n9411 , n357090 , n357098 );
not ( n9412 , n357090 );
buf ( n357101 , n357094 );
and ( n9414 , n9412 , n357101 );
nor ( n9415 , n9411 , n9414 );
buf ( n357104 , n9415 );
buf ( n357105 , n8777 );
not ( n9418 , n357105 );
buf ( n357107 , n350699 );
not ( n9420 , n357107 );
or ( n9421 , n9418 , n9420 );
buf ( n357110 , n350377 );
xor ( n9423 , n582 , n549 );
buf ( n357112 , n9423 );
nand ( n9425 , n357110 , n357112 );
buf ( n357114 , n9425 );
buf ( n357115 , n357114 );
nand ( n9428 , n9421 , n357115 );
buf ( n357117 , n9428 );
xor ( n9430 , n357104 , n357117 );
buf ( n357119 , n9430 );
buf ( n357120 , n8760 );
not ( n9433 , n357120 );
buf ( n357122 , n356440 );
not ( n9435 , n357122 );
or ( n9436 , n9433 , n9435 );
buf ( n357125 , n356446 );
buf ( n357126 , n555 );
buf ( n357127 , n576 );
xor ( n9440 , n357126 , n357127 );
buf ( n357129 , n9440 );
buf ( n357130 , n357129 );
nand ( n9443 , n357125 , n357130 );
buf ( n357132 , n9443 );
buf ( n357133 , n357132 );
nand ( n9446 , n9436 , n357133 );
buf ( n357135 , n9446 );
buf ( n357136 , n357135 );
buf ( n357137 , n356498 );
not ( n9450 , n357137 );
buf ( n357139 , n347554 );
not ( n9452 , n357139 );
or ( n9453 , n9450 , n9452 );
buf ( n357142 , n588 );
buf ( n357143 , n347568 );
nand ( n9456 , n357142 , n357143 );
buf ( n357145 , n9456 );
buf ( n357146 , n357145 );
nand ( n9459 , n9453 , n357146 );
buf ( n357148 , n9459 );
buf ( n357149 , n357148 );
not ( n9462 , n357149 );
buf ( n357151 , n9462 );
buf ( n357152 , n357151 );
xor ( n9465 , n357136 , n357152 );
buf ( n357154 , n356569 );
xor ( n9467 , n9465 , n357154 );
buf ( n357156 , n9467 );
buf ( n357157 , n357156 );
xor ( n9470 , n357119 , n357157 );
xor ( n9471 , n356610 , n356625 );
and ( n9472 , n9471 , n356639 );
and ( n9473 , n356610 , n356625 );
or ( n9474 , n9472 , n9473 );
buf ( n357163 , n9474 );
buf ( n357164 , n357163 );
xor ( n9477 , n9470 , n357164 );
buf ( n357166 , n9477 );
buf ( n357167 , n357166 );
xor ( n9480 , n356576 , n356590 );
and ( n9481 , n9480 , n356642 );
and ( n9482 , n356576 , n356590 );
or ( n9483 , n9481 , n9482 );
buf ( n357172 , n9483 );
buf ( n357173 , n357172 );
xor ( n9486 , n357167 , n357173 );
xor ( n9487 , n356541 , n356555 );
and ( n9488 , n9487 , n356573 );
and ( n9489 , n356541 , n356555 );
or ( n9490 , n9488 , n9489 );
buf ( n357179 , n9490 );
buf ( n357180 , n357179 );
xor ( n9493 , n356432 , n356433 );
and ( n9494 , n9493 , n356455 );
and ( n9495 , n356432 , n356433 );
or ( n9496 , n9494 , n9495 );
buf ( n357185 , n9496 );
buf ( n357186 , n357185 );
buf ( n357187 , n356471 );
not ( n9500 , n357187 );
buf ( n357189 , n8815 );
not ( n9502 , n357189 );
or ( n9503 , n9500 , n9502 );
buf ( n357192 , n356474 );
not ( n9505 , n357192 );
buf ( n357194 , n8816 );
not ( n9507 , n357194 );
or ( n9508 , n9505 , n9507 );
buf ( n357197 , n356490 );
nand ( n9510 , n9508 , n357197 );
buf ( n357199 , n9510 );
buf ( n357200 , n357199 );
nand ( n9513 , n9503 , n357200 );
buf ( n357202 , n9513 );
buf ( n357203 , n357202 );
xor ( n9516 , n357186 , n357203 );
buf ( n357205 , n551 );
buf ( n357206 , n580 );
xor ( n9519 , n357205 , n357206 );
buf ( n357208 , n9519 );
not ( n9521 , n357208 );
not ( n9522 , n351038 );
or ( n9523 , n9521 , n9522 );
nand ( n9524 , n3868 , n351035 , n8860 );
nand ( n9525 , n9523 , n9524 );
buf ( n357214 , n9525 );
buf ( n357215 , n8846 );
not ( n9528 , n357215 );
buf ( n357217 , n5162 );
not ( n9530 , n357217 );
or ( n9531 , n9528 , n9530 );
buf ( n357220 , n352491 );
buf ( n357221 , n553 );
buf ( n357222 , n578 );
xor ( n9535 , n357221 , n357222 );
buf ( n357224 , n9535 );
buf ( n357225 , n357224 );
nand ( n9538 , n357220 , n357225 );
buf ( n357227 , n9538 );
buf ( n357228 , n357227 );
nand ( n9541 , n9531 , n357228 );
buf ( n357230 , n9541 );
buf ( n357231 , n357230 );
xor ( n9544 , n357214 , n357231 );
buf ( n357233 , n8875 );
not ( n9546 , n357233 );
buf ( n357235 , n2471 );
not ( n9548 , n357235 );
or ( n9549 , n9546 , n9548 );
buf ( n357238 , n348629 );
xor ( n9551 , n584 , n547 );
buf ( n357240 , n9551 );
nand ( n9553 , n357238 , n357240 );
buf ( n357242 , n9553 );
buf ( n357243 , n357242 );
nand ( n9556 , n9549 , n357243 );
buf ( n357245 , n9556 );
buf ( n357246 , n357245 );
xor ( n9559 , n9544 , n357246 );
buf ( n357248 , n9559 );
buf ( n357249 , n357248 );
xor ( n9562 , n9516 , n357249 );
buf ( n357251 , n9562 );
buf ( n357252 , n357251 );
xor ( n9565 , n357180 , n357252 );
xor ( n9566 , n356458 , n356510 );
and ( n9567 , n9566 , n356517 );
and ( n9568 , n356458 , n356510 );
or ( n9569 , n9567 , n9568 );
buf ( n357258 , n9569 );
buf ( n357259 , n357258 );
xor ( n9572 , n9565 , n357259 );
buf ( n357261 , n9572 );
buf ( n357262 , n357261 );
xor ( n9575 , n9486 , n357262 );
buf ( n357264 , n9575 );
buf ( n357265 , n357264 );
xor ( n9578 , n9385 , n357265 );
buf ( n357267 , n9578 );
buf ( n357268 , n357267 );
xor ( n9581 , n9368 , n357268 );
buf ( n357270 , n9581 );
xor ( n9583 , n356389 , n356404 );
and ( n9584 , n9583 , n356651 );
and ( n9585 , n356389 , n356404 );
or ( n9586 , n9584 , n9585 );
buf ( n357275 , n9586 );
or ( n9588 , n357270 , n357275 );
buf ( n357277 , n357270 );
buf ( n357278 , n357275 );
nand ( n9591 , n357277 , n357278 );
buf ( n357280 , n9591 );
nand ( n9593 , n9588 , n357280 );
and ( n9594 , n9143 , n9593 );
not ( n9595 , n9143 );
not ( n9596 , n9593 );
and ( n9597 , n9595 , n9596 );
nor ( n9598 , n9594 , n9597 );
not ( n9599 , n9598 );
nand ( n9600 , n9133 , n9599 );
not ( n9601 , n9600 );
not ( n9602 , n9132 );
nor ( n9603 , n9602 , n9599 );
or ( n9604 , n9601 , n9603 );
not ( n9605 , n9604 );
not ( n9606 , n8484 );
not ( n9607 , n8980 );
or ( n9608 , n9606 , n9607 );
nand ( n9609 , n9608 , n8283 );
not ( n9610 , n9609 );
nand ( n9611 , n9610 , n8354 );
not ( n9612 , n8279 );
not ( n9613 , n9612 );
not ( n9614 , n8983 );
or ( n9615 , n9613 , n9614 );
nand ( n9616 , n9615 , n8982 );
buf ( n9617 , n9616 );
not ( n9618 , n9617 );
nand ( n9619 , n9611 , n9618 );
not ( n9620 , n9619 );
or ( n9621 , n9605 , n9620 );
nor ( n9622 , n9604 , n9617 );
nand ( n9623 , n9611 , n9622 );
nand ( n9624 , n9621 , n9623 );
buf ( n9625 , n9624 );
buf ( n357314 , n9625 );
buf ( n9627 , n357314 );
buf ( n357316 , n9627 );
buf ( n9629 , n357316 );
not ( n9630 , n9629 );
and ( n9631 , n8993 , n9630 );
not ( n9632 , n8993 );
and ( n9633 , n9632 , n9629 );
nor ( n9634 , n9631 , n9633 );
buf ( n9635 , n9634 );
buf ( n9636 , n9635 );
not ( n9637 , n9636 );
buf ( n357326 , n9637 );
not ( n9639 , n357326 );
or ( n9640 , n8351 , n9639 );
buf ( n357329 , n9635 );
not ( n9642 , n606 );
buf ( n357331 , n9642 );
nand ( n9644 , n357329 , n357331 );
buf ( n357333 , n9644 );
buf ( n357334 , n357333 );
nand ( n9647 , n9640 , n357334 );
buf ( n357336 , n9647 );
buf ( n357337 , n357336 );
not ( n9650 , n357337 );
or ( n9651 , n8349 , n9650 );
buf ( n357340 , n606 );
not ( n9653 , n357340 );
not ( n9654 , n8311 );
not ( n9655 , n8321 );
or ( n9656 , n9654 , n9655 );
nand ( n9657 , n9656 , n8303 );
buf ( n357346 , n8990 );
buf ( n9659 , n357346 );
buf ( n357348 , n9659 );
or ( n9661 , n9657 , n357348 );
nand ( n9662 , n357348 , n9657 );
nand ( n9663 , n9661 , n9662 );
buf ( n9664 , n9663 );
buf ( n357353 , n9664 );
not ( n9666 , n357353 );
buf ( n357355 , n9666 );
buf ( n357356 , n357355 );
not ( n9669 , n357356 );
or ( n9670 , n9653 , n9669 );
buf ( n357359 , n9664 );
buf ( n357360 , n9642 );
nand ( n9673 , n357359 , n357360 );
buf ( n357362 , n9673 );
buf ( n357363 , n357362 );
nand ( n9676 , n9670 , n357363 );
buf ( n357365 , n9676 );
buf ( n357366 , n357365 );
buf ( n357367 , n9642 );
buf ( n357368 , n607 );
nor ( n9681 , n357367 , n357368 );
buf ( n357370 , n9681 );
buf ( n357371 , n357370 );
buf ( n9684 , n357371 );
buf ( n357373 , n9684 );
buf ( n357374 , n357373 );
buf ( n9687 , n357374 );
buf ( n357376 , n9687 );
buf ( n357377 , n357376 );
nand ( n9690 , n357366 , n357377 );
buf ( n357379 , n9690 );
buf ( n357380 , n357379 );
nand ( n9693 , n9651 , n357380 );
buf ( n357382 , n9693 );
buf ( n357383 , n357382 );
xor ( n9696 , n8347 , n357383 );
buf ( n357385 , n9696 );
buf ( n357386 , n357385 );
xor ( n9699 , n7597 , n357386 );
buf ( n357388 , n9699 );
buf ( n357389 , n357388 );
not ( n9702 , n357389 );
buf ( n357391 , n607 );
not ( n9704 , n357391 );
buf ( n357393 , n357365 );
not ( n9706 , n357393 );
or ( n9707 , n9704 , n9706 );
not ( n9708 , n8333 );
and ( n9709 , n9708 , n9642 );
not ( n9710 , n9708 );
and ( n9711 , n9710 , n606 );
nor ( n9712 , n9709 , n9711 );
buf ( n357401 , n9712 );
buf ( n357402 , n357376 );
nand ( n9715 , n357401 , n357402 );
buf ( n357404 , n9715 );
buf ( n357405 , n357404 );
nand ( n9718 , n9707 , n357405 );
buf ( n357407 , n9718 );
buf ( n357408 , n357407 );
buf ( n357409 , n4361 );
not ( n9722 , n357409 );
buf ( n357411 , n355115 );
not ( n9724 , n357411 );
or ( n9725 , n9722 , n9724 );
buf ( n357414 , n4443 );
buf ( n357415 , n598 );
not ( n9728 , n357415 );
buf ( n357417 , n4298 );
not ( n9730 , n357417 );
or ( n9731 , n9728 , n9730 );
buf ( n357420 , n348884 );
buf ( n357421 , n347312 );
nand ( n9734 , n357420 , n357421 );
buf ( n357423 , n9734 );
buf ( n357424 , n357423 );
nand ( n9737 , n9731 , n357424 );
buf ( n357426 , n9737 );
buf ( n357427 , n357426 );
nand ( n9740 , n357414 , n357427 );
buf ( n357429 , n9740 );
buf ( n357430 , n357429 );
nand ( n9743 , n9725 , n357430 );
buf ( n357432 , n9743 );
buf ( n357433 , n357432 );
xor ( n9746 , n349257 , n349282 );
xor ( n9747 , n9746 , n349386 );
buf ( n357436 , n9747 );
buf ( n357437 , n357436 );
xor ( n9750 , n357433 , n357437 );
buf ( n9751 , n1721 );
buf ( n357440 , n9751 );
not ( n9753 , n357440 );
buf ( n357442 , n355158 );
not ( n9755 , n357442 );
or ( n9756 , n9753 , n9755 );
and ( n9757 , n351952 , n600 );
not ( n9758 , n351952 );
and ( n9759 , n9758 , n4192 );
or ( n9760 , n9757 , n9759 );
buf ( n357449 , n9760 );
buf ( n357450 , n351924 );
nand ( n9763 , n357449 , n357450 );
buf ( n357452 , n9763 );
buf ( n357453 , n357452 );
nand ( n9766 , n9756 , n357453 );
buf ( n357455 , n9766 );
buf ( n357456 , n357455 );
and ( n9769 , n9750 , n357456 );
and ( n9770 , n357433 , n357437 );
or ( n9771 , n9769 , n9770 );
buf ( n357460 , n9771 );
buf ( n357461 , n357460 );
not ( n9774 , n352149 );
not ( n9775 , n355203 );
or ( n9776 , n9774 , n9775 );
buf ( n357465 , n602 );
not ( n9778 , n357465 );
buf ( n357467 , n351901 );
not ( n9780 , n357467 );
or ( n9781 , n9778 , n9780 );
buf ( n357470 , n4221 );
buf ( n357471 , n349406 );
nand ( n9784 , n357470 , n357471 );
buf ( n357473 , n9784 );
buf ( n357474 , n357473 );
nand ( n9787 , n9781 , n357474 );
buf ( n357476 , n9787 );
buf ( n357477 , n357476 );
buf ( n357478 , n354113 );
nand ( n9791 , n357477 , n357478 );
buf ( n357480 , n9791 );
nand ( n9793 , n9776 , n357480 );
buf ( n357482 , n9793 );
xor ( n9795 , n357461 , n357482 );
xor ( n9796 , n355123 , n355127 );
xor ( n9797 , n9796 , n355166 );
buf ( n357486 , n9797 );
buf ( n357487 , n357486 );
and ( n9800 , n9795 , n357487 );
and ( n9801 , n357461 , n357482 );
or ( n9802 , n9800 , n9801 );
buf ( n357491 , n9802 );
buf ( n357492 , n357491 );
buf ( n357493 , n6599 );
not ( n9806 , n357493 );
buf ( n357495 , n7372 );
not ( n9808 , n357495 );
or ( n9809 , n9806 , n9808 );
not ( n9810 , n6399 );
not ( n9811 , n354080 );
or ( n9812 , n9810 , n9811 );
nand ( n9813 , n354079 , n6398 );
nand ( n9814 , n9812 , n9813 );
buf ( n357503 , n9814 );
not ( n9816 , n357503 );
buf ( n357505 , n9816 );
and ( n9818 , n604 , n357505 );
not ( n9819 , n604 );
and ( n9820 , n9819 , n9814 );
or ( n9821 , n9818 , n9820 );
buf ( n357510 , n9821 );
buf ( n357511 , n355075 );
nand ( n9824 , n357510 , n357511 );
buf ( n357513 , n9824 );
buf ( n357514 , n357513 );
nand ( n9827 , n9809 , n357514 );
buf ( n357516 , n9827 );
buf ( n357517 , n357516 );
xor ( n9830 , n357492 , n357517 );
xor ( n9831 , n355171 , n355211 );
xor ( n9832 , n9831 , n355246 );
buf ( n357521 , n9832 );
buf ( n357522 , n357521 );
and ( n9835 , n9830 , n357522 );
and ( n9836 , n357492 , n357517 );
or ( n9837 , n9835 , n9836 );
buf ( n357526 , n9837 );
buf ( n357527 , n357526 );
xor ( n9840 , n357408 , n357527 );
xor ( n9841 , n355082 , n355251 );
xor ( n9842 , n9841 , n355279 );
buf ( n357531 , n9842 );
buf ( n357532 , n357531 );
and ( n9845 , n9840 , n357532 );
and ( n9846 , n357408 , n357527 );
or ( n9847 , n9845 , n9846 );
buf ( n357536 , n9847 );
buf ( n357537 , n357536 );
not ( n9850 , n357537 );
buf ( n357539 , n9850 );
buf ( n357540 , n357539 );
nand ( n9853 , n9702 , n357540 );
buf ( n357542 , n9853 );
not ( n9855 , n357542 );
buf ( n357544 , n607 );
not ( n9857 , n357544 );
buf ( n357546 , n606 );
not ( n9859 , n357546 );
buf ( n357548 , n7360 );
not ( n9861 , n357548 );
or ( n9862 , n9859 , n9861 );
buf ( n357551 , n7363 );
buf ( n357552 , n9642 );
nand ( n9865 , n357551 , n357552 );
buf ( n357554 , n9865 );
buf ( n357555 , n357554 );
nand ( n9868 , n9862 , n357555 );
buf ( n357557 , n9868 );
buf ( n357558 , n357557 );
not ( n9871 , n357558 );
or ( n9872 , n9857 , n9871 );
buf ( n357561 , n606 );
not ( n9874 , n357561 );
buf ( n357563 , n354056 );
not ( n9876 , n357563 );
or ( n9877 , n9874 , n9876 );
buf ( n357566 , n354053 );
buf ( n357567 , n9642 );
nand ( n9880 , n357566 , n357567 );
buf ( n357569 , n9880 );
buf ( n357570 , n357569 );
nand ( n9883 , n9877 , n357570 );
buf ( n357572 , n9883 );
buf ( n357573 , n357572 );
buf ( n357574 , n357376 );
nand ( n9887 , n357573 , n357574 );
buf ( n357576 , n9887 );
buf ( n357577 , n357576 );
nand ( n9890 , n9872 , n357577 );
buf ( n357579 , n9890 );
buf ( n357580 , n357579 );
buf ( n357581 , n9751 );
not ( n9894 , n357581 );
buf ( n357583 , n9760 );
not ( n9896 , n357583 );
or ( n9897 , n9894 , n9896 );
buf ( n357586 , n600 );
not ( n9899 , n357586 );
buf ( n357588 , n1145 );
not ( n9901 , n357588 );
buf ( n357590 , n9901 );
buf ( n357591 , n357590 );
not ( n9904 , n357591 );
or ( n9905 , n9899 , n9904 );
buf ( n357594 , n357590 );
not ( n9907 , n357594 );
buf ( n357596 , n9907 );
buf ( n357597 , n357596 );
buf ( n357598 , n4192 );
nand ( n9911 , n357597 , n357598 );
buf ( n357600 , n9911 );
buf ( n357601 , n357600 );
nand ( n9914 , n9905 , n357601 );
buf ( n357603 , n9914 );
buf ( n357604 , n357603 );
buf ( n357605 , n351924 );
nand ( n9918 , n357604 , n357605 );
buf ( n357607 , n9918 );
buf ( n357608 , n357607 );
nand ( n9921 , n9897 , n357608 );
buf ( n357610 , n9921 );
buf ( n357611 , n357610 );
buf ( n357612 , n4361 );
not ( n9925 , n357612 );
buf ( n357614 , n357426 );
not ( n9927 , n357614 );
or ( n9928 , n9925 , n9927 );
buf ( n357617 , n598 );
not ( n9930 , n357617 );
buf ( n357619 , n349232 );
not ( n9932 , n357619 );
or ( n9933 , n9930 , n9932 );
buf ( n357622 , n354213 );
buf ( n357623 , n347312 );
nand ( n9936 , n357622 , n357623 );
buf ( n357625 , n9936 );
buf ( n357626 , n357625 );
nand ( n9939 , n9933 , n357626 );
buf ( n357628 , n9939 );
buf ( n357629 , n357628 );
buf ( n357630 , n4443 );
nand ( n9943 , n357629 , n357630 );
buf ( n357632 , n9943 );
buf ( n357633 , n357632 );
nand ( n9946 , n9928 , n357633 );
buf ( n357635 , n9946 );
buf ( n357636 , n357635 );
xor ( n9949 , n349294 , n349319 );
xor ( n9950 , n9949 , n349381 );
buf ( n357639 , n9950 );
buf ( n357640 , n357639 );
xor ( n9953 , n357636 , n357640 );
xor ( n9954 , n349325 , n349363 );
xor ( n9955 , n9954 , n349377 );
buf ( n357644 , n9955 );
buf ( n357645 , n357644 );
buf ( n357646 , n4361 );
not ( n9959 , n357646 );
buf ( n357648 , n357628 );
not ( n9961 , n357648 );
or ( n9962 , n9959 , n9961 );
buf ( n357651 , n598 );
not ( n9964 , n357651 );
buf ( n357653 , n349070 );
not ( n9966 , n357653 );
or ( n9967 , n9964 , n9966 );
buf ( n357656 , n347312 );
buf ( n357657 , n1375 );
nand ( n9970 , n357656 , n357657 );
buf ( n357659 , n9970 );
buf ( n357660 , n357659 );
nand ( n9973 , n9967 , n357660 );
buf ( n357662 , n9973 );
buf ( n357663 , n357662 );
buf ( n357664 , n352124 );
nand ( n9977 , n357663 , n357664 );
buf ( n357666 , n9977 );
buf ( n357667 , n357666 );
nand ( n9980 , n9962 , n357667 );
buf ( n357669 , n9980 );
buf ( n357670 , n357669 );
xor ( n9983 , n357645 , n357670 );
buf ( n357672 , n349359 );
not ( n9985 , n357672 );
buf ( n357674 , n1654 );
not ( n9987 , n357674 );
or ( n9988 , n9985 , n9987 );
buf ( n357677 , n1654 );
buf ( n357678 , n349359 );
or ( n9991 , n357677 , n357678 );
nand ( n9992 , n9988 , n9991 );
buf ( n357681 , n9992 );
buf ( n357682 , n357681 );
buf ( n357683 , n4361 );
not ( n9996 , n357683 );
buf ( n357685 , n357662 );
not ( n9998 , n357685 );
or ( n9999 , n9996 , n9998 );
buf ( n357688 , n598 );
not ( n10001 , n357688 );
buf ( n357690 , n349106 );
not ( n10003 , n357690 );
or ( n10004 , n10001 , n10003 );
buf ( n357693 , n1305 );
buf ( n357694 , n347312 );
nand ( n10007 , n357693 , n357694 );
buf ( n357696 , n10007 );
buf ( n357697 , n357696 );
nand ( n10010 , n10004 , n357697 );
buf ( n357699 , n10010 );
buf ( n357700 , n357699 );
buf ( n357701 , n352124 );
nand ( n10014 , n357700 , n357701 );
buf ( n357703 , n10014 );
buf ( n357704 , n357703 );
nand ( n10017 , n9999 , n357704 );
buf ( n357706 , n10017 );
buf ( n357707 , n357706 );
xor ( n10020 , n357682 , n357707 );
buf ( n357709 , n1202 );
buf ( n357710 , n347319 );
not ( n10023 , n357710 );
buf ( n357712 , n10023 );
buf ( n357713 , n357712 );
nor ( n10026 , n357709 , n357713 );
buf ( n357715 , n10026 );
buf ( n357716 , n357715 );
not ( n10029 , n4361 );
not ( n10030 , n598 );
not ( n10031 , n348925 );
or ( n10032 , n10030 , n10031 );
buf ( n357721 , n1215 );
buf ( n357722 , n347312 );
nand ( n10035 , n357721 , n357722 );
buf ( n357724 , n10035 );
nand ( n10037 , n10032 , n357724 );
not ( n10038 , n10037 );
or ( n10039 , n10029 , n10038 );
buf ( n357728 , n352124 );
buf ( n357729 , n598 );
nand ( n10042 , n357728 , n357729 );
buf ( n357731 , n10042 );
buf ( n357732 , n357731 );
not ( n10045 , n357732 );
buf ( n357734 , n1256 );
not ( n10047 , n357734 );
and ( n10048 , n10045 , n10047 );
buf ( n357737 , n1256 );
buf ( n357738 , n352124 );
buf ( n357739 , n598 );
not ( n10052 , n357739 );
and ( n10053 , n357738 , n10052 );
buf ( n357742 , n10053 );
buf ( n357743 , n357742 );
and ( n10056 , n357737 , n357743 );
nor ( n10057 , n10048 , n10056 );
buf ( n357746 , n10057 );
nand ( n10059 , n10039 , n357746 );
buf ( n357748 , n10059 );
buf ( n357749 , n599 );
buf ( n357750 , n600 );
or ( n10063 , n357749 , n357750 );
buf ( n357752 , n1256 );
nand ( n10065 , n10063 , n357752 );
buf ( n357754 , n10065 );
buf ( n357755 , n357754 );
buf ( n357756 , n599 );
buf ( n357757 , n600 );
and ( n10070 , n357756 , n357757 );
buf ( n357759 , n347312 );
nor ( n10072 , n10070 , n357759 );
buf ( n357761 , n10072 );
buf ( n357762 , n357761 );
nand ( n10075 , n357755 , n357762 );
buf ( n357764 , n10075 );
buf ( n357765 , n357764 );
not ( n10078 , n357765 );
and ( n10079 , n357748 , n10078 );
buf ( n357768 , n10079 );
buf ( n357769 , n357768 );
xor ( n10082 , n357716 , n357769 );
buf ( n357771 , n4361 );
not ( n10084 , n357771 );
buf ( n357773 , n357699 );
not ( n10086 , n357773 );
or ( n10087 , n10084 , n10086 );
nand ( n10088 , n10037 , n352124 );
buf ( n357777 , n10088 );
nand ( n10090 , n10087 , n357777 );
buf ( n357779 , n10090 );
buf ( n357780 , n357779 );
and ( n10093 , n10082 , n357780 );
or ( n10095 , n10093 , C0 );
buf ( n357783 , n10095 );
buf ( n357784 , n357783 );
and ( n10098 , n10020 , n357784 );
and ( n10099 , n357682 , n357707 );
or ( n10100 , n10098 , n10099 );
buf ( n357788 , n10100 );
buf ( n357789 , n357788 );
and ( n10103 , n9983 , n357789 );
and ( n10104 , n357645 , n357670 );
or ( n10105 , n10103 , n10104 );
buf ( n357793 , n10105 );
buf ( n357794 , n357793 );
xor ( n10108 , n9953 , n357794 );
buf ( n357796 , n10108 );
buf ( n357797 , n357796 );
xor ( n10111 , n357611 , n357797 );
buf ( n357799 , n352149 );
not ( n10113 , n357799 );
buf ( n357801 , n602 );
not ( n10115 , n357801 );
buf ( n357803 , n352066 );
not ( n10117 , n357803 );
or ( n10118 , n10115 , n10117 );
buf ( n357806 , n4388 );
buf ( n357807 , n349406 );
nand ( n10121 , n357806 , n357807 );
buf ( n357809 , n10121 );
buf ( n357810 , n357809 );
nand ( n10124 , n10118 , n357810 );
buf ( n357812 , n10124 );
buf ( n357813 , n357812 );
not ( n10127 , n357813 );
or ( n10128 , n10113 , n10127 );
buf ( n357816 , n602 );
not ( n10130 , n357816 );
buf ( n357818 , n352095 );
not ( n10132 , n357818 );
or ( n10133 , n10130 , n10132 );
buf ( n357821 , n354251 );
buf ( n357822 , n349406 );
nand ( n10136 , n357821 , n357822 );
buf ( n357824 , n10136 );
buf ( n357825 , n357824 );
nand ( n10139 , n10133 , n357825 );
buf ( n357827 , n10139 );
buf ( n357828 , n357827 );
buf ( n357829 , n354113 );
nand ( n10143 , n357828 , n357829 );
buf ( n357831 , n10143 );
buf ( n357832 , n357831 );
nand ( n10146 , n10128 , n357832 );
buf ( n357834 , n10146 );
buf ( n357835 , n357834 );
and ( n10149 , n10111 , n357835 );
and ( n10150 , n357611 , n357797 );
or ( n10151 , n10149 , n10150 );
buf ( n357839 , n10151 );
buf ( n357840 , n357839 );
buf ( n357841 , n6600 );
not ( n10155 , n357841 );
buf ( n357843 , n604 );
buf ( n357844 , n6458 );
and ( n10158 , n357843 , n357844 );
not ( n10159 , n357843 );
buf ( n357847 , n355178 );
and ( n10161 , n10159 , n357847 );
nor ( n10162 , n10158 , n10161 );
buf ( n357850 , n10162 );
buf ( n357851 , n357850 );
not ( n10165 , n357851 );
or ( n10166 , n10155 , n10165 );
and ( n10167 , n604 , n4179 );
not ( n10168 , n604 );
buf ( n357856 , n4183 );
buf ( n10170 , n357856 );
buf ( n357858 , n10170 );
and ( n10172 , n10168 , n357858 );
or ( n10173 , n10167 , n10172 );
buf ( n357861 , n10173 );
buf ( n357862 , n355075 );
nand ( n10176 , n357861 , n357862 );
buf ( n357864 , n10176 );
buf ( n357865 , n357864 );
nand ( n10179 , n10166 , n357865 );
buf ( n357867 , n10179 );
buf ( n357868 , n357867 );
xor ( n10182 , n357840 , n357868 );
xor ( n10183 , n357636 , n357640 );
and ( n10184 , n10183 , n357794 );
and ( n10185 , n357636 , n357640 );
or ( n10186 , n10184 , n10185 );
buf ( n357874 , n10186 );
buf ( n357875 , n357874 );
buf ( n357876 , n352149 );
not ( n10190 , n357876 );
buf ( n357878 , n357476 );
not ( n10192 , n357878 );
or ( n10193 , n10190 , n10192 );
buf ( n357881 , n357812 );
buf ( n357882 , n354113 );
nand ( n10196 , n357881 , n357882 );
buf ( n357884 , n10196 );
buf ( n357885 , n357884 );
nand ( n10199 , n10193 , n357885 );
buf ( n357887 , n10199 );
buf ( n357888 , n357887 );
xor ( n10202 , n357875 , n357888 );
xor ( n10203 , n357433 , n357437 );
xor ( n10204 , n10203 , n357456 );
buf ( n357892 , n10204 );
buf ( n357893 , n357892 );
xor ( n10207 , n10202 , n357893 );
buf ( n357895 , n10207 );
buf ( n357896 , n357895 );
and ( n10210 , n10182 , n357896 );
and ( n10211 , n357840 , n357868 );
or ( n10212 , n10210 , n10211 );
buf ( n357900 , n10212 );
buf ( n357901 , n357900 );
xor ( n10215 , n357580 , n357901 );
xor ( n10216 , n357875 , n357888 );
and ( n10217 , n10216 , n357893 );
and ( n10218 , n357875 , n357888 );
or ( n10219 , n10217 , n10218 );
buf ( n357907 , n10219 );
buf ( n357908 , n357907 );
xor ( n10222 , n357461 , n357482 );
xor ( n10223 , n10222 , n357487 );
buf ( n357911 , n10223 );
buf ( n357912 , n357911 );
xor ( n10226 , n357908 , n357912 );
buf ( n357914 , n6599 );
not ( n10228 , n357914 );
buf ( n357916 , n9821 );
not ( n10230 , n357916 );
or ( n10231 , n10228 , n10230 );
buf ( n357919 , n357850 );
buf ( n357920 , n355075 );
nand ( n10234 , n357919 , n357920 );
buf ( n357922 , n10234 );
buf ( n357923 , n357922 );
nand ( n10237 , n10231 , n357923 );
buf ( n357925 , n10237 );
buf ( n357926 , n357925 );
xor ( n10240 , n10226 , n357926 );
buf ( n357928 , n10240 );
buf ( n357929 , n357928 );
xor ( n10243 , n10215 , n357929 );
buf ( n357931 , n10243 );
buf ( n357932 , n357931 );
buf ( n357933 , n1722 );
not ( n10247 , n357933 );
buf ( n357935 , n357603 );
not ( n10249 , n357935 );
or ( n10250 , n10247 , n10249 );
buf ( n357938 , n600 );
not ( n10252 , n357938 );
buf ( n357940 , n4298 );
not ( n10254 , n357940 );
or ( n10255 , n10252 , n10254 );
buf ( n357943 , n4192 );
buf ( n357944 , n1179 );
nand ( n10258 , n357943 , n357944 );
buf ( n357946 , n10258 );
buf ( n357947 , n357946 );
nand ( n10261 , n10255 , n357947 );
buf ( n357949 , n10261 );
buf ( n357950 , n357949 );
buf ( n357951 , n351924 );
nand ( n10265 , n357950 , n357951 );
buf ( n357953 , n10265 );
buf ( n357954 , n357953 );
nand ( n10268 , n10250 , n357954 );
buf ( n357956 , n10268 );
buf ( n357957 , n357956 );
xor ( n10271 , n357645 , n357670 );
xor ( n10272 , n10271 , n357789 );
buf ( n357960 , n10272 );
buf ( n357961 , n357960 );
xor ( n10275 , n357957 , n357961 );
buf ( n357963 , n1722 );
not ( n10277 , n357963 );
buf ( n357965 , n357949 );
not ( n10279 , n357965 );
or ( n10280 , n10277 , n10279 );
buf ( n357968 , n600 );
not ( n10282 , n357968 );
buf ( n357970 , n349049 );
not ( n10284 , n357970 );
or ( n10285 , n10282 , n10284 );
buf ( n357973 , n354213 );
buf ( n357974 , n4192 );
nand ( n10288 , n357973 , n357974 );
buf ( n357976 , n10288 );
buf ( n357977 , n357976 );
nand ( n10291 , n10285 , n357977 );
buf ( n357979 , n10291 );
buf ( n357980 , n357979 );
buf ( n357981 , n351924 );
nand ( n10295 , n357980 , n357981 );
buf ( n357983 , n10295 );
buf ( n357984 , n357983 );
nand ( n10298 , n10280 , n357984 );
buf ( n357986 , n10298 );
buf ( n357987 , n357986 );
xor ( n10301 , n357682 , n357707 );
xor ( n10302 , n10301 , n357784 );
buf ( n357990 , n10302 );
buf ( n357991 , n357990 );
xor ( n10305 , n357987 , n357991 );
xor ( n10306 , n357716 , n357769 );
xor ( n10307 , n10306 , n357780 );
buf ( n357995 , n10307 );
buf ( n357996 , n357995 );
buf ( n357997 , n1722 );
not ( n10311 , n357997 );
buf ( n357999 , n357979 );
not ( n10313 , n357999 );
or ( n10314 , n10311 , n10313 );
buf ( n358002 , n600 );
not ( n10316 , n358002 );
buf ( n358004 , n349070 );
not ( n10318 , n358004 );
or ( n10319 , n10316 , n10318 );
buf ( n358007 , n1375 );
buf ( n358008 , n4192 );
nand ( n10322 , n358007 , n358008 );
buf ( n358010 , n10322 );
buf ( n358011 , n358010 );
nand ( n10325 , n10319 , n358011 );
buf ( n358013 , n10325 );
buf ( n358014 , n358013 );
buf ( n358015 , n351924 );
nand ( n10329 , n358014 , n358015 );
buf ( n358017 , n10329 );
buf ( n358018 , n358017 );
nand ( n10332 , n10314 , n358018 );
buf ( n358020 , n10332 );
buf ( n358021 , n358020 );
xor ( n10335 , n357996 , n358021 );
buf ( n358023 , n357764 );
not ( n10337 , n358023 );
buf ( n358025 , n10059 );
not ( n10339 , n358025 );
or ( n10340 , n10337 , n10339 );
buf ( n358028 , n10059 );
buf ( n358029 , n357764 );
or ( n10343 , n358028 , n358029 );
nand ( n10344 , n10340 , n10343 );
buf ( n358032 , n10344 );
buf ( n358033 , n358032 );
buf ( n358034 , n1202 );
buf ( n358035 , n352112 );
nor ( n10349 , n358034 , n358035 );
buf ( n358037 , n10349 );
buf ( n358038 , n358037 );
buf ( n358039 , n1722 );
not ( n10353 , n358039 );
buf ( n358041 , n10353 );
not ( n10355 , n600 );
nor ( n10356 , n358041 , n10355 );
not ( n10357 , n10356 );
not ( n10358 , n348925 );
or ( n10359 , n10357 , n10358 );
buf ( n10360 , n348922 );
nor ( n10361 , n358041 , n600 );
and ( n10362 , n10360 , n10361 );
buf ( n358050 , n1256 );
buf ( n358051 , n351924 );
buf ( n358052 , n600 );
not ( n10366 , n358052 );
and ( n10367 , n358051 , n10366 );
buf ( n358055 , n10367 );
buf ( n358056 , n358055 );
and ( n10370 , n358050 , n358056 );
buf ( n358058 , n1202 );
buf ( n358059 , n351924 );
buf ( n358060 , n600 );
nand ( n10374 , n358059 , n358060 );
buf ( n358062 , n10374 );
buf ( n358063 , n358062 );
not ( n10377 , n358063 );
buf ( n358065 , n10377 );
buf ( n358066 , n358065 );
and ( n10380 , n358058 , n358066 );
nor ( n10381 , n10370 , n10380 );
buf ( n358069 , n10381 );
not ( n10383 , n358069 );
nor ( n10384 , n10362 , n10383 );
nand ( n10385 , n10359 , n10384 );
buf ( n358073 , n10385 );
not ( n10387 , n358073 );
buf ( n358075 , n601 );
buf ( n358076 , n602 );
or ( n10390 , n358075 , n358076 );
buf ( n358078 , n1256 );
nand ( n10392 , n10390 , n358078 );
buf ( n358080 , n10392 );
buf ( n358081 , n358080 );
buf ( n358082 , n601 );
buf ( n358083 , n602 );
nand ( n10397 , n358082 , n358083 );
buf ( n358085 , n10397 );
buf ( n358086 , n358085 );
buf ( n358087 , n600 );
nand ( n10401 , n358081 , n358086 , n358087 );
buf ( n358089 , n10401 );
buf ( n358090 , n358089 );
nor ( n10404 , n10387 , n358090 );
buf ( n358092 , n10404 );
buf ( n358093 , n358092 );
xor ( n10407 , n358038 , n358093 );
not ( n10408 , n1722 );
not ( n10409 , n1297 );
not ( n10413 , n600 );
and ( n10414 , C1 , n10413 );
or ( n10415 , C0 , n10414 );
and ( n10416 , n10409 , n10415 );
not ( n10417 , n10409 );
not ( n10419 , n4192 );
and ( n10420 , C1 , n10419 );
or ( n10424 , n10420 , C0 );
and ( n10425 , n10417 , n10424 );
or ( n10426 , n10416 , n10425 );
not ( n10427 , n10426 );
or ( n10428 , n10408 , n10427 );
or ( n10429 , n600 , n10360 );
or ( n10430 , n348925 , n10355 );
nand ( n10431 , n10429 , n10430 , n351924 );
nand ( n10432 , n10428 , n10431 );
buf ( n358113 , n10432 );
and ( n10434 , n10407 , n358113 );
or ( n10436 , n10434 , C0 );
buf ( n358116 , n10436 );
buf ( n358117 , n358116 );
xor ( n10439 , n358033 , n358117 );
buf ( n358119 , n1722 );
not ( n10441 , n358119 );
buf ( n358121 , n358013 );
not ( n10443 , n358121 );
or ( n10444 , n10441 , n10443 );
nand ( n10445 , n10426 , n351924 );
buf ( n358125 , n10445 );
nand ( n10447 , n10444 , n358125 );
buf ( n358127 , n10447 );
buf ( n358128 , n358127 );
and ( n10450 , n10439 , n358128 );
and ( n10451 , n358033 , n358117 );
or ( n10452 , n10450 , n10451 );
buf ( n358132 , n10452 );
buf ( n358133 , n358132 );
and ( n10455 , n10335 , n358133 );
and ( n10456 , n357996 , n358021 );
or ( n10457 , n10455 , n10456 );
buf ( n358137 , n10457 );
buf ( n358138 , n358137 );
and ( n10460 , n10305 , n358138 );
and ( n10461 , n357987 , n357991 );
or ( n10462 , n10460 , n10461 );
buf ( n358142 , n10462 );
buf ( n358143 , n358142 );
and ( n10465 , n10275 , n358143 );
and ( n10466 , n357957 , n357961 );
or ( n10467 , n10465 , n10466 );
buf ( n358147 , n10467 );
buf ( n358148 , n358147 );
buf ( n358149 , n6600 );
not ( n10471 , n358149 );
buf ( n358151 , n10173 );
not ( n10473 , n358151 );
or ( n10474 , n10471 , n10473 );
buf ( n358154 , n355075 );
and ( n10476 , n604 , n4221 );
not ( n10477 , n604 );
and ( n10478 , n10477 , n351901 );
nor ( n10479 , n10476 , n10478 );
buf ( n358159 , n10479 );
nand ( n10481 , n358154 , n358159 );
buf ( n358161 , n10481 );
buf ( n358162 , n358161 );
nand ( n10484 , n10474 , n358162 );
buf ( n358164 , n10484 );
buf ( n358165 , n358164 );
xor ( n10487 , n358148 , n358165 );
xor ( n10488 , n357611 , n357797 );
xor ( n10489 , n10488 , n357835 );
buf ( n358169 , n10489 );
buf ( n358170 , n358169 );
and ( n10492 , n10487 , n358170 );
and ( n10493 , n358148 , n358165 );
or ( n10494 , n10492 , n10493 );
buf ( n358174 , n10494 );
buf ( n358175 , n358174 );
buf ( n358176 , n607 );
not ( n10498 , n358176 );
buf ( n358178 , n357572 );
not ( n10500 , n358178 );
or ( n10501 , n10498 , n10500 );
buf ( n358181 , n606 );
not ( n10503 , n358181 );
buf ( n358183 , n354087 );
not ( n10505 , n358183 );
or ( n10506 , n10503 , n10505 );
buf ( n358186 , n354093 );
buf ( n358187 , n9642 );
nand ( n10509 , n358186 , n358187 );
buf ( n358189 , n10509 );
buf ( n358190 , n358189 );
nand ( n10512 , n10506 , n358190 );
buf ( n358192 , n10512 );
buf ( n358193 , n358192 );
buf ( n358194 , n357373 );
nand ( n10516 , n358193 , n358194 );
buf ( n358196 , n10516 );
buf ( n358197 , n358196 );
nand ( n10519 , n10501 , n358197 );
buf ( n358199 , n10519 );
buf ( n358200 , n358199 );
xor ( n10522 , n358175 , n358200 );
xor ( n10523 , n357840 , n357868 );
xor ( n10524 , n10523 , n357896 );
buf ( n358204 , n10524 );
buf ( n358205 , n358204 );
and ( n10527 , n10522 , n358205 );
and ( n10528 , n358175 , n358200 );
or ( n10529 , n10527 , n10528 );
buf ( n358209 , n10529 );
buf ( n358210 , n358209 );
nor ( n10532 , n357932 , n358210 );
buf ( n358212 , n10532 );
buf ( n358213 , n358212 );
not ( n10535 , n358213 );
buf ( n358215 , n10535 );
not ( n10537 , n358215 );
xor ( n10538 , n358175 , n358200 );
xor ( n10539 , n10538 , n358205 );
buf ( n358219 , n10539 );
buf ( n358220 , n358219 );
buf ( n358221 , n352149 );
not ( n10543 , n358221 );
buf ( n358223 , n357827 );
not ( n10545 , n358223 );
or ( n10546 , n10543 , n10545 );
buf ( n358226 , n602 );
not ( n10548 , n358226 );
buf ( n358228 , n351952 );
not ( n10550 , n358228 );
or ( n10551 , n10548 , n10550 );
buf ( n358231 , n349406 );
buf ( n358232 , n351958 );
nand ( n10554 , n358231 , n358232 );
buf ( n358234 , n10554 );
buf ( n358235 , n358234 );
nand ( n10557 , n10551 , n358235 );
buf ( n358237 , n10557 );
buf ( n358238 , n358237 );
buf ( n358239 , n354113 );
nand ( n10561 , n358238 , n358239 );
buf ( n358241 , n10561 );
buf ( n358242 , n358241 );
nand ( n10564 , n10546 , n358242 );
buf ( n358244 , n10564 );
buf ( n358245 , n358244 );
buf ( n358246 , n6600 );
not ( n10568 , n358246 );
buf ( n358248 , n10479 );
not ( n10570 , n358248 );
or ( n10571 , n10568 , n10570 );
buf ( n358251 , n604 );
not ( n10573 , n358251 );
not ( n10574 , n352065 );
buf ( n358254 , n10574 );
not ( n10576 , n358254 );
or ( n10577 , n10573 , n10576 );
buf ( n358257 , n604 );
not ( n10579 , n358257 );
buf ( n358259 , n352065 );
nand ( n10581 , n10579 , n358259 );
buf ( n358261 , n10581 );
buf ( n358262 , n358261 );
nand ( n10584 , n10577 , n358262 );
buf ( n358264 , n10584 );
buf ( n358265 , n358264 );
buf ( n358266 , n355072 );
nand ( n10588 , n358265 , n358266 );
buf ( n358268 , n10588 );
buf ( n358269 , n358268 );
nand ( n10591 , n10571 , n358269 );
buf ( n358271 , n10591 );
buf ( n358272 , n358271 );
xor ( n10594 , n358245 , n358272 );
xor ( n10595 , n357957 , n357961 );
xor ( n10596 , n10595 , n358143 );
buf ( n358276 , n10596 );
buf ( n358277 , n358276 );
and ( n10599 , n10594 , n358277 );
and ( n10600 , n358245 , n358272 );
or ( n10601 , n10599 , n10600 );
buf ( n358281 , n10601 );
buf ( n358282 , n358281 );
xor ( n10604 , n358148 , n358165 );
xor ( n10605 , n10604 , n358170 );
buf ( n358285 , n10605 );
buf ( n358286 , n358285 );
xor ( n10608 , n358282 , n358286 );
buf ( n358288 , n607 );
not ( n10610 , n358288 );
buf ( n358290 , n358192 );
not ( n10612 , n358290 );
or ( n10613 , n10610 , n10612 );
not ( n10614 , n6458 );
not ( n10615 , n9642 );
or ( n10616 , n10614 , n10615 );
not ( n10617 , n6458 );
nand ( n10618 , n10617 , n606 );
nand ( n10619 , n10616 , n10618 );
buf ( n358299 , n10619 );
buf ( n358300 , n357373 );
nand ( n10622 , n358299 , n358300 );
buf ( n358302 , n10622 );
buf ( n358303 , n358302 );
nand ( n10625 , n10613 , n358303 );
buf ( n358305 , n10625 );
buf ( n358306 , n358305 );
and ( n10628 , n10608 , n358306 );
and ( n10629 , n358282 , n358286 );
or ( n10630 , n10628 , n10629 );
buf ( n358310 , n10630 );
buf ( n358311 , n358310 );
nor ( n10633 , n358220 , n358311 );
buf ( n358313 , n10633 );
not ( n10635 , n358313 );
not ( n10636 , n10635 );
buf ( n358316 , n352149 );
not ( n10638 , n358316 );
buf ( n358318 , n602 );
not ( n10640 , n358318 );
buf ( n358320 , n4298 );
not ( n10642 , n358320 );
or ( n10643 , n10640 , n10642 );
buf ( n358323 , n349406 );
buf ( n358324 , n1179 );
nand ( n10646 , n358323 , n358324 );
buf ( n358326 , n10646 );
buf ( n358327 , n358326 );
nand ( n10649 , n10643 , n358327 );
buf ( n358329 , n10649 );
buf ( n358330 , n358329 );
not ( n10652 , n358330 );
or ( n10653 , n10638 , n10652 );
buf ( n358333 , n602 );
not ( n10655 , n358333 );
buf ( n358335 , n349232 );
not ( n10657 , n358335 );
or ( n10658 , n10655 , n10657 );
buf ( n358338 , n354213 );
buf ( n358339 , n349406 );
nand ( n10661 , n358338 , n358339 );
buf ( n358341 , n10661 );
buf ( n358342 , n358341 );
nand ( n10664 , n10658 , n358342 );
buf ( n358344 , n10664 );
buf ( n358345 , n358344 );
buf ( n358346 , n354113 );
nand ( n10668 , n358345 , n358346 );
buf ( n358348 , n10668 );
buf ( n358349 , n358348 );
nand ( n10671 , n10653 , n358349 );
buf ( n358351 , n10671 );
buf ( n358352 , n358351 );
xor ( n10674 , n358033 , n358117 );
xor ( n10675 , n10674 , n358128 );
buf ( n358355 , n10675 );
buf ( n358356 , n358355 );
xor ( n10678 , n358352 , n358356 );
xor ( n10679 , n358038 , n358093 );
xor ( n10680 , n10679 , n358113 );
buf ( n358360 , n10680 );
buf ( n358361 , n358360 );
buf ( n358362 , n352149 );
not ( n10684 , n358362 );
buf ( n358364 , n358344 );
not ( n10686 , n358364 );
or ( n10687 , n10684 , n10686 );
buf ( n358367 , n349406 );
not ( n10689 , n358367 );
buf ( n358369 , n1375 );
not ( n10691 , n358369 );
or ( n10692 , n10689 , n10691 );
not ( n10693 , n1375 );
nand ( n10694 , n10693 , n602 );
buf ( n358374 , n10694 );
nand ( n10696 , n10692 , n358374 );
buf ( n358376 , n10696 );
buf ( n358377 , n358376 );
buf ( n358378 , n354113 );
nand ( n10700 , n358377 , n358378 );
buf ( n358380 , n10700 );
buf ( n358381 , n358380 );
nand ( n10703 , n10687 , n358381 );
buf ( n358383 , n10703 );
buf ( n358384 , n358383 );
xor ( n10706 , n358361 , n358384 );
buf ( n358386 , n358089 );
not ( n10708 , n358386 );
buf ( n358388 , n10385 );
not ( n10710 , n358388 );
or ( n10711 , n10708 , n10710 );
buf ( n358391 , n10385 );
buf ( n358392 , n358089 );
or ( n10714 , n358391 , n358392 );
nand ( n10715 , n10711 , n10714 );
buf ( n358395 , n10715 );
buf ( n358396 , n358395 );
buf ( n358397 , n1202 );
buf ( n358398 , n358041 );
nor ( n10720 , n358397 , n358398 );
buf ( n358400 , n10720 );
buf ( n358401 , n358400 );
buf ( n358402 , n349406 );
buf ( n358403 , n1215 );
and ( n10725 , n358402 , n358403 );
not ( n10726 , n358402 );
buf ( n358406 , n348931 );
and ( n10728 , n10726 , n358406 );
nor ( n10729 , n10725 , n10728 );
buf ( n358409 , n10729 );
buf ( n358410 , n358409 );
buf ( n358411 , n4464 );
or ( n10733 , n358410 , n358411 );
buf ( n358413 , n1256 );
buf ( n358414 , n354113 );
buf ( n358415 , n349406 );
and ( n10737 , n358414 , n358415 );
buf ( n358417 , n10737 );
buf ( n358418 , n358417 );
and ( n10740 , n358413 , n358418 );
buf ( n358420 , n1202 );
buf ( n358421 , n354113 );
buf ( n358422 , n602 );
and ( n10744 , n358421 , n358422 );
buf ( n358424 , n10744 );
buf ( n358425 , n358424 );
and ( n10747 , n358420 , n358425 );
nor ( n10748 , n10740 , n10747 );
buf ( n358428 , n10748 );
buf ( n358429 , n358428 );
nand ( n10751 , n10733 , n358429 );
buf ( n358431 , n10751 );
buf ( n358432 , n358431 );
not ( n10754 , n358432 );
buf ( n358434 , n603 );
buf ( n358435 , n604 );
or ( n10757 , n358434 , n358435 );
buf ( n358437 , n1256 );
nand ( n10759 , n10757 , n358437 );
buf ( n358439 , n10759 );
buf ( n358440 , n358439 );
buf ( n358441 , n352145 );
buf ( n358442 , n602 );
nand ( n10764 , n358440 , n358441 , n358442 );
buf ( n358444 , n10764 );
buf ( n358445 , n358444 );
nor ( n10767 , n10754 , n358445 );
buf ( n358447 , n10767 );
buf ( n358448 , n358447 );
xor ( n10770 , n358401 , n358448 );
or ( n10771 , n4464 , n349406 );
nor ( n10772 , n10771 , n1305 );
not ( n10773 , n354113 );
nor ( n10774 , n10773 , n358409 );
nor ( n10775 , n10772 , n10774 );
not ( n10776 , n4464 );
nand ( n10777 , n10776 , n1305 , n349406 );
nand ( n10778 , n10775 , n10777 );
buf ( n358458 , n10778 );
and ( n10780 , n10770 , n358458 );
or ( n10782 , n10780 , C0 );
buf ( n358461 , n10782 );
buf ( n358462 , n358461 );
xor ( n10785 , n358396 , n358462 );
buf ( n358464 , n352149 );
not ( n10787 , n358464 );
buf ( n358466 , n358376 );
not ( n10789 , n358466 );
or ( n10790 , n10787 , n10789 );
xnor ( n10791 , n349406 , n1305 );
nand ( n10792 , n10791 , n354113 );
buf ( n358471 , n10792 );
nand ( n10794 , n10790 , n358471 );
buf ( n358473 , n10794 );
buf ( n358474 , n358473 );
and ( n10797 , n10785 , n358474 );
and ( n10798 , n358396 , n358462 );
or ( n10799 , n10797 , n10798 );
buf ( n358478 , n10799 );
buf ( n358479 , n358478 );
and ( n10802 , n10706 , n358479 );
and ( n10803 , n358361 , n358384 );
or ( n10804 , n10802 , n10803 );
buf ( n358483 , n10804 );
buf ( n358484 , n358483 );
and ( n10807 , n10678 , n358484 );
and ( n10808 , n358352 , n358356 );
or ( n10809 , n10807 , n10808 );
buf ( n358488 , n10809 );
buf ( n358489 , n358488 );
buf ( n358490 , n607 );
not ( n10813 , n358490 );
buf ( n358492 , n606 );
buf ( n358493 , n4221 );
and ( n10816 , n358492 , n358493 );
not ( n10817 , n358492 );
buf ( n358496 , n351901 );
and ( n10819 , n10817 , n358496 );
nor ( n10820 , n10816 , n10819 );
buf ( n358499 , n10820 );
buf ( n358500 , n358499 );
not ( n10823 , n358500 );
or ( n10824 , n10813 , n10823 );
buf ( n358503 , n606 );
not ( n10826 , n358503 );
buf ( n358505 , n10574 );
not ( n10828 , n358505 );
or ( n10829 , n10826 , n10828 );
buf ( n358508 , n9642 );
buf ( n358509 , n352065 );
nand ( n10832 , n358508 , n358509 );
buf ( n358511 , n10832 );
buf ( n358512 , n358511 );
nand ( n10835 , n10829 , n358512 );
buf ( n358514 , n10835 );
buf ( n358515 , n358514 );
buf ( n358516 , n357373 );
nand ( n10839 , n358515 , n358516 );
buf ( n358518 , n10839 );
buf ( n358519 , n358518 );
nand ( n10842 , n10824 , n358519 );
buf ( n358521 , n10842 );
buf ( n358522 , n358521 );
xor ( n10845 , n358489 , n358522 );
buf ( n358524 , n352149 );
not ( n10847 , n358524 );
buf ( n358526 , n602 );
not ( n10849 , n358526 );
buf ( n358528 , n357590 );
not ( n10851 , n358528 );
or ( n10852 , n10849 , n10851 );
buf ( n358531 , n357596 );
buf ( n358532 , n349406 );
nand ( n10855 , n358531 , n358532 );
buf ( n358534 , n10855 );
buf ( n358535 , n358534 );
nand ( n10858 , n10852 , n358535 );
buf ( n358537 , n10858 );
buf ( n358538 , n358537 );
not ( n10861 , n358538 );
or ( n10862 , n10847 , n10861 );
buf ( n358541 , n358329 );
buf ( n358542 , n354113 );
nand ( n10865 , n358541 , n358542 );
buf ( n358544 , n10865 );
buf ( n358545 , n358544 );
nand ( n10868 , n10862 , n358545 );
buf ( n358547 , n10868 );
buf ( n358548 , n358547 );
xor ( n10871 , n357996 , n358021 );
xor ( n10872 , n10871 , n358133 );
buf ( n358551 , n10872 );
buf ( n358552 , n358551 );
xor ( n10875 , n358548 , n358552 );
buf ( n358554 , n6599 );
not ( n10877 , n358554 );
buf ( n358556 , n604 );
not ( n10879 , n358556 );
buf ( n358558 , n4410 );
not ( n10881 , n358558 );
or ( n10882 , n10879 , n10881 );
buf ( n358561 , n604 );
not ( n10884 , n358561 );
buf ( n358563 , n6561 );
nand ( n10886 , n10884 , n358563 );
buf ( n358565 , n10886 );
buf ( n358566 , n358565 );
nand ( n10889 , n10882 , n358566 );
buf ( n358568 , n10889 );
buf ( n358569 , n358568 );
not ( n10892 , n358569 );
or ( n10893 , n10877 , n10892 );
not ( n10894 , n604 );
not ( n10895 , n351952 );
or ( n10896 , n10894 , n10895 );
buf ( n358575 , n604 );
not ( n10898 , n358575 );
buf ( n358577 , n4266 );
nand ( n10900 , n10898 , n358577 );
buf ( n358579 , n10900 );
nand ( n10902 , n10896 , n358579 );
buf ( n358581 , n10902 );
buf ( n358582 , n355072 );
nand ( n10905 , n358581 , n358582 );
buf ( n358584 , n10905 );
buf ( n358585 , n358584 );
nand ( n10908 , n10893 , n358585 );
buf ( n358587 , n10908 );
buf ( n358588 , n358587 );
xor ( n10911 , n10875 , n358588 );
buf ( n358590 , n10911 );
buf ( n358591 , n358590 );
xor ( n10914 , n10845 , n358591 );
buf ( n358593 , n10914 );
buf ( n358594 , n358593 );
not ( n10917 , n358594 );
not ( n10918 , n6599 );
not ( n10919 , n10902 );
or ( n10920 , n10918 , n10919 );
xor ( n10921 , n604 , n348855 );
nand ( n10922 , n10921 , n355072 );
nand ( n10923 , n10920 , n10922 );
buf ( n358602 , n10923 );
xor ( n10925 , n358352 , n358356 );
xor ( n10926 , n10925 , n358484 );
buf ( n358605 , n10926 );
buf ( n358606 , n358605 );
xor ( n10929 , n358602 , n358606 );
buf ( n358608 , n607 );
not ( n10931 , n358608 );
buf ( n358610 , n358514 );
not ( n10933 , n358610 );
or ( n10934 , n10931 , n10933 );
buf ( n358613 , n606 );
not ( n10936 , n358613 );
buf ( n358615 , n4410 );
not ( n10938 , n358615 );
or ( n10939 , n10936 , n10938 );
not ( n10940 , n4410 );
nand ( n10941 , n10940 , n9642 );
buf ( n358620 , n10941 );
nand ( n10943 , n10939 , n358620 );
buf ( n358622 , n10943 );
buf ( n358623 , n358622 );
buf ( n358624 , n357373 );
nand ( n10947 , n358623 , n358624 );
buf ( n358626 , n10947 );
buf ( n358627 , n358626 );
nand ( n10950 , n10934 , n358627 );
buf ( n358629 , n10950 );
buf ( n358630 , n358629 );
and ( n10953 , n10929 , n358630 );
and ( n10954 , n358602 , n358606 );
or ( n10955 , n10953 , n10954 );
buf ( n358634 , n10955 );
buf ( n358635 , n358634 );
not ( n10958 , n358635 );
buf ( n358637 , n10958 );
buf ( n358638 , n358637 );
nand ( n10961 , n10917 , n358638 );
buf ( n358640 , n10961 );
not ( n10963 , n358640 );
buf ( n358642 , n6599 );
not ( n10965 , n358642 );
buf ( n358644 , n10921 );
not ( n10967 , n358644 );
or ( n10968 , n10965 , n10967 );
not ( n10969 , n1179 );
and ( n10970 , n604 , n10969 );
not ( n10971 , n604 );
and ( n10972 , n10971 , n1179 );
or ( n10973 , n10970 , n10972 );
buf ( n358652 , n10973 );
buf ( n358653 , n355072 );
nand ( n10976 , n358652 , n358653 );
buf ( n358655 , n10976 );
buf ( n358656 , n358655 );
nand ( n10979 , n10968 , n358656 );
buf ( n358658 , n10979 );
buf ( n358659 , n358658 );
xor ( n10982 , n358361 , n358384 );
xor ( n10983 , n10982 , n358479 );
buf ( n358662 , n10983 );
buf ( n358663 , n358662 );
xor ( n10986 , n358659 , n358663 );
buf ( n358665 , n607 );
not ( n10988 , n358665 );
buf ( n358667 , n358622 );
not ( n10990 , n358667 );
or ( n10991 , n10988 , n10990 );
buf ( n358670 , n606 );
buf ( n358671 , n4266 );
xor ( n10994 , n358670 , n358671 );
buf ( n358673 , n10994 );
buf ( n358674 , n358673 );
buf ( n358675 , n357373 );
nand ( n10998 , n358674 , n358675 );
buf ( n358677 , n10998 );
buf ( n358678 , n358677 );
nand ( n11001 , n10991 , n358678 );
buf ( n358680 , n11001 );
buf ( n358681 , n358680 );
and ( n11004 , n10986 , n358681 );
and ( n11005 , n358659 , n358663 );
or ( n11006 , n11004 , n11005 );
buf ( n358685 , n11006 );
xor ( n11008 , n358602 , n358606 );
xor ( n11009 , n11008 , n358630 );
buf ( n358688 , n11009 );
xor ( n11011 , n358685 , n358688 );
buf ( n358690 , n6599 );
not ( n11013 , n358690 );
buf ( n358692 , n10973 );
not ( n11015 , n358692 );
or ( n11016 , n11013 , n11015 );
buf ( n358695 , n604 );
not ( n11018 , n358695 );
buf ( n358697 , n349049 );
not ( n11020 , n358697 );
or ( n11021 , n11018 , n11020 );
buf ( n358700 , n604 );
not ( n11023 , n358700 );
buf ( n358702 , n349046 );
nand ( n11025 , n11023 , n358702 );
buf ( n358704 , n11025 );
buf ( n358705 , n358704 );
nand ( n11028 , n11021 , n358705 );
buf ( n358707 , n11028 );
buf ( n358708 , n358707 );
buf ( n358709 , n355072 );
nand ( n11032 , n358708 , n358709 );
buf ( n358711 , n11032 );
buf ( n358712 , n358711 );
nand ( n11035 , n11016 , n358712 );
buf ( n358714 , n11035 );
buf ( n358715 , n358714 );
xor ( n11038 , n358396 , n358462 );
xor ( n11039 , n11038 , n358474 );
buf ( n358718 , n11039 );
buf ( n358719 , n358718 );
xor ( n11042 , n358715 , n358719 );
xor ( n11043 , n358401 , n358448 );
xor ( n11044 , n11043 , n358458 );
buf ( n358723 , n11044 );
buf ( n358724 , n358723 );
buf ( n358725 , n6599 );
not ( n11048 , n358725 );
buf ( n358727 , n358707 );
not ( n11050 , n358727 );
or ( n11051 , n11048 , n11050 );
not ( n11052 , n604 );
not ( n11053 , n10693 );
or ( n11054 , n11052 , n11053 );
or ( n11055 , n10693 , n604 );
nand ( n11056 , n11054 , n11055 );
buf ( n358735 , n11056 );
buf ( n358736 , n355072 );
nand ( n11059 , n358735 , n358736 );
buf ( n358738 , n11059 );
buf ( n358739 , n358738 );
nand ( n11062 , n11051 , n358739 );
buf ( n358741 , n11062 );
buf ( n358742 , n358741 );
xor ( n11065 , n358724 , n358742 );
buf ( n358744 , n358444 );
not ( n11067 , n358744 );
buf ( n358746 , n358431 );
not ( n11069 , n358746 );
or ( n11070 , n11067 , n11069 );
buf ( n358749 , n358431 );
buf ( n358750 , n358444 );
or ( n11073 , n358749 , n358750 );
nand ( n11074 , n11070 , n11073 );
buf ( n358753 , n11074 );
buf ( n358754 , n358753 );
buf ( n358755 , n6599 );
not ( n11078 , n358755 );
buf ( n358757 , n11056 );
not ( n11080 , n358757 );
or ( n11081 , n11078 , n11080 );
and ( n11082 , n604 , n349106 );
not ( n11083 , n604 );
and ( n11084 , n11083 , n1305 );
or ( n11085 , n11082 , n11084 );
buf ( n358764 , n11085 );
buf ( n358765 , n355072 );
nand ( n11088 , n358764 , n358765 );
buf ( n358767 , n11088 );
buf ( n358768 , n358767 );
nand ( n11091 , n11081 , n358768 );
buf ( n358770 , n11091 );
buf ( n358771 , n358770 );
xor ( n11094 , n358754 , n358771 );
buf ( n358773 , n1202 );
buf ( n358774 , n4464 );
nor ( n11097 , n358773 , n358774 );
buf ( n358776 , n11097 );
buf ( n358777 , n358776 );
buf ( n358778 , n6599 );
not ( n11101 , n358778 );
buf ( n358780 , n604 );
not ( n11103 , n358780 );
buf ( n358782 , n1214 );
not ( n11105 , n358782 );
or ( n11106 , n11103 , n11105 );
buf ( n358785 , n604 );
not ( n11108 , n358785 );
buf ( n358787 , n1215 );
nand ( n11110 , n11108 , n358787 );
buf ( n358789 , n11110 );
buf ( n358790 , n358789 );
nand ( n11113 , n11106 , n358790 );
buf ( n358792 , n11113 );
buf ( n358793 , n358792 );
not ( n11116 , n358793 );
or ( n11117 , n11101 , n11116 );
buf ( n358796 , n604 );
buf ( n358797 , n1256 );
and ( n11120 , n358796 , n358797 );
not ( n11121 , n358796 );
buf ( n358800 , n1202 );
and ( n11123 , n11121 , n358800 );
nor ( n11124 , n11120 , n11123 );
buf ( n358803 , n11124 );
buf ( n358804 , n358803 );
buf ( n358805 , n355072 );
nand ( n11128 , n358804 , n358805 );
buf ( n358807 , n11128 );
buf ( n358808 , n358807 );
nand ( n11131 , n11117 , n358808 );
buf ( n358810 , n11131 );
buf ( n358811 , n358810 );
not ( n11134 , n358811 );
buf ( n358813 , n605 );
buf ( n358814 , n606 );
or ( n11137 , n358813 , n358814 );
buf ( n358816 , n1256 );
nand ( n11139 , n11137 , n358816 );
buf ( n358818 , n11139 );
buf ( n358819 , n358818 );
buf ( n358820 , n605 );
buf ( n358821 , n606 );
and ( n11144 , n358820 , n358821 );
not ( n11145 , n604 );
buf ( n358824 , n11145 );
nor ( n11147 , n11144 , n358824 );
buf ( n358826 , n11147 );
buf ( n358827 , n358826 );
nand ( n11150 , n358819 , n358827 );
buf ( n358829 , n11150 );
buf ( n358830 , n358829 );
nor ( n11153 , n11134 , n358830 );
buf ( n358832 , n11153 );
buf ( n358833 , n358832 );
xor ( n11156 , n358777 , n358833 );
buf ( n358835 , n6599 );
not ( n11158 , n358835 );
buf ( n358837 , n11085 );
not ( n11160 , n358837 );
or ( n11161 , n11158 , n11160 );
buf ( n358840 , n358792 );
buf ( n358841 , n355072 );
nand ( n11164 , n358840 , n358841 );
buf ( n358843 , n11164 );
buf ( n358844 , n358843 );
nand ( n11167 , n11161 , n358844 );
buf ( n358846 , n11167 );
buf ( n358847 , n358846 );
and ( n11170 , n11156 , n358847 );
or ( n11172 , n11170 , C0 );
buf ( n358850 , n11172 );
buf ( n358851 , n358850 );
and ( n11175 , n11094 , n358851 );
and ( n11176 , n358754 , n358771 );
or ( n11177 , n11175 , n11176 );
buf ( n358855 , n11177 );
buf ( n358856 , n358855 );
and ( n11180 , n11065 , n358856 );
and ( n11181 , n358724 , n358742 );
or ( n11182 , n11180 , n11181 );
buf ( n358860 , n11182 );
buf ( n358861 , n358860 );
and ( n11185 , n11042 , n358861 );
and ( n11186 , n358715 , n358719 );
or ( n11187 , n11185 , n11186 );
buf ( n358865 , n11187 );
xor ( n11189 , n358659 , n358663 );
xor ( n11190 , n11189 , n358681 );
buf ( n358868 , n11190 );
xor ( n11192 , n358865 , n358868 );
xor ( n11193 , n358724 , n358742 );
xor ( n11194 , n11193 , n358856 );
buf ( n358872 , n11194 );
not ( n11196 , n358872 );
buf ( n358874 , n607 );
not ( n11198 , n358874 );
buf ( n358876 , n606 );
buf ( n358877 , n348855 );
and ( n11201 , n358876 , n358877 );
not ( n11202 , n358876 );
buf ( n358880 , n357590 );
and ( n11204 , n11202 , n358880 );
nor ( n11205 , n11201 , n11204 );
buf ( n358883 , n11205 );
buf ( n358884 , n358883 );
not ( n11208 , n358884 );
or ( n11209 , n11198 , n11208 );
not ( n11210 , n606 );
not ( n11211 , n4298 );
or ( n11212 , n11210 , n11211 );
buf ( n358890 , n1179 );
buf ( n358891 , n9642 );
nand ( n11215 , n358890 , n358891 );
buf ( n358893 , n11215 );
nand ( n11217 , n11212 , n358893 );
buf ( n358895 , n11217 );
buf ( n358896 , n357373 );
nand ( n11220 , n358895 , n358896 );
buf ( n358898 , n11220 );
buf ( n358899 , n358898 );
nand ( n11223 , n11209 , n358899 );
buf ( n358901 , n11223 );
not ( n11225 , n358901 );
nand ( n11226 , n11196 , n11225 );
not ( n11227 , n607 );
not ( n11228 , n358893 );
not ( n11229 , n11228 );
or ( n11230 , n11227 , n11229 );
and ( n11231 , n607 , n606 );
and ( n11232 , n10969 , n11231 );
and ( n11233 , n1349 , n9642 );
not ( n11234 , n1349 );
and ( n11235 , n11234 , n606 );
or ( n11236 , n11233 , n11235 );
and ( n11237 , n11236 , n357373 );
nor ( n11238 , n11232 , n11237 );
nand ( n11239 , n11230 , n11238 );
buf ( n358917 , n11239 );
xor ( n11241 , n358754 , n358771 );
xor ( n11242 , n11241 , n358851 );
buf ( n358920 , n11242 );
buf ( n358921 , n358920 );
xor ( n11245 , n358917 , n358921 );
buf ( n358923 , n358829 );
not ( n11247 , n358923 );
buf ( n358925 , n358810 );
not ( n11249 , n358925 );
or ( n11250 , n11247 , n11249 );
buf ( n358928 , n358810 );
buf ( n358929 , n358829 );
or ( n11253 , n358928 , n358929 );
nand ( n11254 , n11250 , n11253 );
buf ( n358932 , n11254 );
buf ( n358933 , n358932 );
buf ( n358934 , n1202 );
buf ( n358935 , n6599 );
not ( n11259 , n358935 );
buf ( n358937 , n11259 );
buf ( n358938 , n358937 );
nor ( n11262 , n358934 , n358938 );
buf ( n358940 , n11262 );
buf ( n358941 , n358940 );
buf ( n358942 , n606 );
not ( n11266 , n358942 );
buf ( n358944 , n1214 );
not ( n11268 , n358944 );
or ( n11269 , n11266 , n11268 );
buf ( n358947 , n1215 );
buf ( n358948 , n9642 );
nand ( n11272 , n358947 , n358948 );
buf ( n358950 , n11272 );
buf ( n358951 , n358950 );
nand ( n11275 , n11269 , n358951 );
buf ( n358953 , n11275 );
buf ( n358954 , n358953 );
buf ( n358955 , n607 );
and ( n11279 , n358954 , n358955 );
buf ( n358957 , n357370 );
not ( n11281 , n358957 );
buf ( n358959 , n1256 );
nor ( n11283 , n11281 , n358959 );
buf ( n358961 , n11283 );
buf ( n358962 , n358961 );
nor ( n11286 , n11279 , n358962 );
buf ( n358964 , n11286 );
buf ( n358965 , n358964 );
buf ( n358966 , n1202 );
buf ( n358967 , n607 );
not ( n11291 , n358967 );
buf ( n358969 , n11291 );
buf ( n358970 , n358969 );
nor ( n11294 , n358966 , n358970 );
buf ( n358972 , n11294 );
buf ( n358973 , n358972 );
buf ( n11297 , n358973 );
buf ( n358975 , n11297 );
buf ( n358976 , n358975 );
buf ( n358977 , n9642 );
or ( n11301 , n358976 , n358977 );
buf ( n358979 , n11301 );
buf ( n358980 , n358979 );
nor ( n11304 , n358965 , n358980 );
buf ( n358982 , n11304 );
buf ( n358983 , n358982 );
xor ( n11307 , n358941 , n358983 );
xor ( n11308 , n1301 , n9642 );
buf ( n358986 , n11308 );
buf ( n358987 , n358969 );
or ( n11311 , n358986 , n358987 );
buf ( n358989 , n357370 );
buf ( n358990 , n358953 );
nand ( n11314 , n358989 , n358990 );
buf ( n358992 , n11314 );
buf ( n358993 , n358992 );
nand ( n11317 , n11311 , n358993 );
buf ( n358995 , n11317 );
buf ( n358996 , n358995 );
and ( n11320 , n11307 , n358996 );
or ( n11322 , n11320 , C0 );
buf ( n358999 , n11322 );
buf ( n359000 , n358999 );
xor ( n11325 , n358933 , n359000 );
not ( n11326 , n9642 );
not ( n11327 , n10693 );
or ( n11328 , n11326 , n11327 );
nand ( n11329 , n1375 , n606 );
nand ( n11330 , n11328 , n11329 );
buf ( n359007 , n11330 );
buf ( n359008 , n358969 );
or ( n11333 , n359007 , n359008 );
buf ( n359010 , n11308 );
not ( n11335 , n359010 );
buf ( n359012 , n357373 );
nand ( n11337 , n11335 , n359012 );
buf ( n359014 , n11337 );
buf ( n359015 , n359014 );
nand ( n11340 , n11333 , n359015 );
buf ( n359017 , n11340 );
buf ( n359018 , n359017 );
and ( n11343 , n11325 , n359018 );
and ( n11344 , n358933 , n359000 );
or ( n11345 , n11343 , n11344 );
buf ( n359022 , n11345 );
not ( n11347 , n359022 );
buf ( n359024 , n607 );
not ( n11349 , n359024 );
buf ( n359026 , n11236 );
not ( n11351 , n359026 );
or ( n11352 , n11349 , n11351 );
buf ( n359029 , n11330 );
not ( n11354 , n359029 );
buf ( n359031 , n357373 );
nand ( n11356 , n11354 , n359031 );
buf ( n359033 , n11356 );
buf ( n359034 , n359033 );
nand ( n11359 , n11352 , n359034 );
buf ( n359036 , n11359 );
xor ( n11361 , n358777 , n358833 );
xor ( n11362 , n11361 , n358847 );
buf ( n359039 , n11362 );
nor ( n11364 , n359036 , n359039 );
or ( n11365 , n11347 , n11364 );
nand ( n11366 , n359039 , n359036 );
nand ( n11367 , n11365 , n11366 );
buf ( n359044 , n11367 );
and ( n11369 , n11245 , n359044 );
and ( n11370 , n358917 , n358921 );
or ( n11371 , n11369 , n11370 );
buf ( n359048 , n11371 );
and ( n11373 , n11226 , n359048 );
and ( n11374 , n358872 , n358901 );
nor ( n11375 , n11373 , n11374 );
buf ( n359052 , n11375 );
xor ( n11377 , n358715 , n358719 );
xor ( n11378 , n11377 , n358861 );
buf ( n359055 , n11378 );
buf ( n359056 , n359055 );
not ( n11381 , n358883 );
not ( n11382 , n357373 );
or ( n11383 , n11381 , n11382 );
buf ( n359060 , n358673 );
not ( n11385 , n359060 );
buf ( n359062 , n11385 );
or ( n11387 , n359062 , n358969 );
nand ( n11388 , n11383 , n11387 );
buf ( n359065 , n11388 );
nor ( n11390 , n359056 , n359065 );
buf ( n359067 , n11390 );
buf ( n359068 , n359067 );
or ( n11393 , n359052 , n359068 );
buf ( n359070 , n359055 );
buf ( n359071 , n11388 );
nand ( n11396 , n359070 , n359071 );
buf ( n359073 , n11396 );
buf ( n359074 , n359073 );
nand ( n11399 , n11393 , n359074 );
buf ( n359076 , n11399 );
and ( n11401 , n11192 , n359076 );
and ( n11402 , n358865 , n358868 );
or ( n11403 , n11401 , n11402 );
and ( n11404 , n11011 , n11403 );
and ( n11405 , n358685 , n358688 );
or ( n11406 , n11404 , n11405 );
not ( n11407 , n11406 );
or ( n11408 , n10963 , n11407 );
buf ( n359085 , n358593 );
buf ( n359086 , n358634 );
nand ( n11411 , n359085 , n359086 );
buf ( n359088 , n11411 );
nand ( n11413 , n11408 , n359088 );
buf ( n359090 , n11413 );
not ( n11415 , n359090 );
xor ( n11416 , n358489 , n358522 );
and ( n11417 , n11416 , n358591 );
and ( n11418 , n358489 , n358522 );
or ( n11419 , n11417 , n11418 );
buf ( n359096 , n11419 );
not ( n11421 , n359096 );
buf ( n359098 , n607 );
not ( n11423 , n359098 );
and ( n11424 , n606 , n4179 );
not ( n11425 , n606 );
and ( n11426 , n11425 , n4183 );
or ( n11427 , n11424 , n11426 );
buf ( n359104 , n11427 );
not ( n11429 , n359104 );
or ( n11430 , n11423 , n11429 );
buf ( n359107 , n358499 );
buf ( n359108 , n357373 );
nand ( n11433 , n359107 , n359108 );
buf ( n359110 , n11433 );
buf ( n359111 , n359110 );
nand ( n11436 , n11430 , n359111 );
buf ( n359113 , n11436 );
buf ( n359114 , n359113 );
xor ( n11439 , n358548 , n358552 );
and ( n11440 , n11439 , n358588 );
and ( n11441 , n358548 , n358552 );
or ( n11442 , n11440 , n11441 );
buf ( n359119 , n11442 );
buf ( n359120 , n359119 );
xor ( n11445 , n359114 , n359120 );
buf ( n359122 , n352149 );
not ( n11447 , n359122 );
buf ( n359124 , n358237 );
not ( n11449 , n359124 );
or ( n11450 , n11447 , n11449 );
buf ( n359127 , n358537 );
buf ( n359128 , n354113 );
nand ( n11453 , n359127 , n359128 );
buf ( n359130 , n11453 );
buf ( n359131 , n359130 );
nand ( n11456 , n11450 , n359131 );
buf ( n359133 , n11456 );
buf ( n359134 , n359133 );
xor ( n11459 , n357987 , n357991 );
xor ( n11460 , n11459 , n358138 );
buf ( n359137 , n11460 );
buf ( n359138 , n359137 );
xor ( n11463 , n359134 , n359138 );
buf ( n359140 , n6599 );
not ( n11465 , n359140 );
buf ( n359142 , n358264 );
not ( n11467 , n359142 );
or ( n11468 , n11465 , n11467 );
buf ( n359145 , n358568 );
buf ( n11470 , n359145 );
buf ( n359147 , n11470 );
buf ( n359148 , n359147 );
buf ( n359149 , n355072 );
nand ( n11474 , n359148 , n359149 );
buf ( n359151 , n11474 );
buf ( n359152 , n359151 );
nand ( n11477 , n11468 , n359152 );
buf ( n359154 , n11477 );
buf ( n359155 , n359154 );
xor ( n11480 , n11463 , n359155 );
buf ( n359157 , n11480 );
buf ( n359158 , n359157 );
xor ( n11483 , n11445 , n359158 );
buf ( n359160 , n11483 );
buf ( n359161 , n359160 );
not ( n11486 , n359161 );
buf ( n359163 , n11486 );
nand ( n11488 , n11421 , n359163 );
buf ( n359165 , n11488 );
not ( n11490 , n359165 );
or ( n11491 , n11415 , n11490 );
buf ( n359168 , n359163 );
not ( n11493 , n359168 );
buf ( n359170 , n359096 );
nand ( n11495 , n11493 , n359170 );
buf ( n359172 , n11495 );
buf ( n359173 , n359172 );
nand ( n11498 , n11491 , n359173 );
buf ( n359175 , n11498 );
buf ( n359176 , n359175 );
not ( n11501 , n359176 );
xor ( n11502 , n359134 , n359138 );
and ( n11503 , n11502 , n359155 );
and ( n11504 , n359134 , n359138 );
or ( n11505 , n11503 , n11504 );
buf ( n359182 , n11505 );
buf ( n359183 , n359182 );
xor ( n11508 , n358245 , n358272 );
xor ( n11509 , n11508 , n358277 );
buf ( n359186 , n11509 );
buf ( n359187 , n359186 );
xor ( n11512 , n359183 , n359187 );
buf ( n359189 , n607 );
not ( n11514 , n359189 );
buf ( n359191 , n10619 );
not ( n11516 , n359191 );
or ( n11517 , n11514 , n11516 );
buf ( n359194 , n11427 );
buf ( n359195 , n357373 );
nand ( n11520 , n359194 , n359195 );
buf ( n359197 , n11520 );
buf ( n359198 , n359197 );
nand ( n11523 , n11517 , n359198 );
buf ( n359200 , n11523 );
buf ( n359201 , n359200 );
xor ( n11526 , n11512 , n359201 );
buf ( n359203 , n11526 );
buf ( n359204 , n359203 );
xor ( n11529 , n359114 , n359120 );
and ( n11530 , n11529 , n359158 );
and ( n11531 , n359114 , n359120 );
or ( n11532 , n11530 , n11531 );
buf ( n359209 , n11532 );
buf ( n359210 , n359209 );
nor ( n11535 , n359204 , n359210 );
buf ( n359212 , n11535 );
buf ( n359213 , n359212 );
not ( n11538 , n359213 );
buf ( n359215 , n11538 );
buf ( n359216 , n359215 );
not ( n11541 , n359216 );
or ( n11542 , n11501 , n11541 );
buf ( n359219 , n359203 );
buf ( n359220 , n359209 );
nand ( n11545 , n359219 , n359220 );
buf ( n359222 , n11545 );
buf ( n359223 , n359222 );
nand ( n11548 , n11542 , n359223 );
buf ( n359225 , n11548 );
not ( n11550 , n359225 );
xor ( n11551 , n358282 , n358286 );
xor ( n11552 , n11551 , n358306 );
buf ( n359229 , n11552 );
buf ( n359230 , n359229 );
not ( n11555 , n359230 );
xor ( n11556 , n359183 , n359187 );
and ( n11557 , n11556 , n359201 );
and ( n11558 , n359183 , n359187 );
or ( n11559 , n11557 , n11558 );
buf ( n359236 , n11559 );
buf ( n359237 , n359236 );
not ( n11562 , n359237 );
buf ( n359239 , n11562 );
buf ( n359240 , n359239 );
nand ( n11565 , n11555 , n359240 );
buf ( n359242 , n11565 );
not ( n11567 , n359242 );
or ( n11568 , n11550 , n11567 );
buf ( n359245 , n359229 );
buf ( n359246 , n359236 );
nand ( n11571 , n359245 , n359246 );
buf ( n359248 , n11571 );
nand ( n11573 , n11568 , n359248 );
not ( n11574 , n11573 );
or ( n11575 , n10636 , n11574 );
nand ( n11576 , n358219 , n358310 );
nand ( n11577 , n11575 , n11576 );
not ( n11578 , n11577 );
or ( n11579 , n10537 , n11578 );
buf ( n359256 , n357931 );
buf ( n359257 , n358209 );
nand ( n11582 , n359256 , n359257 );
buf ( n359259 , n11582 );
nand ( n11584 , n11579 , n359259 );
buf ( n359261 , n11584 );
not ( n11586 , n359261 );
buf ( n359263 , n11586 );
xor ( n11588 , n357908 , n357912 );
and ( n11589 , n11588 , n357926 );
and ( n11590 , n357908 , n357912 );
or ( n11591 , n11589 , n11590 );
buf ( n359268 , n11591 );
buf ( n359269 , n359268 );
not ( n11594 , n607 );
not ( n11595 , n9712 );
or ( n11596 , n11594 , n11595 );
nand ( n11597 , n357557 , n357376 );
nand ( n11598 , n11596 , n11597 );
buf ( n359275 , n11598 );
xor ( n11600 , n359269 , n359275 );
xor ( n11601 , n357492 , n357517 );
xor ( n11602 , n11601 , n357522 );
buf ( n359279 , n11602 );
buf ( n359280 , n359279 );
xor ( n11605 , n11600 , n359280 );
buf ( n359282 , n11605 );
buf ( n359283 , n359282 );
xor ( n11608 , n357580 , n357901 );
and ( n11609 , n11608 , n357929 );
and ( n11610 , n357580 , n357901 );
or ( n11611 , n11609 , n11610 );
buf ( n359288 , n11611 );
buf ( n359289 , n359288 );
nor ( n11614 , n359283 , n359289 );
buf ( n359291 , n11614 );
or ( n11616 , n359263 , n359291 );
buf ( n359293 , n359282 );
buf ( n359294 , n359288 );
nand ( n11619 , n359293 , n359294 );
buf ( n359296 , n11619 );
nand ( n11621 , n11616 , n359296 );
not ( n11622 , n11621 );
xor ( n11623 , n357408 , n357527 );
xor ( n11624 , n11623 , n357532 );
buf ( n359301 , n11624 );
buf ( n359302 , n359301 );
not ( n11627 , n359302 );
xor ( n11628 , n359269 , n359275 );
and ( n11629 , n11628 , n359280 );
and ( n11630 , n359269 , n359275 );
or ( n11631 , n11629 , n11630 );
buf ( n359308 , n11631 );
buf ( n359309 , n359308 );
not ( n11634 , n359309 );
buf ( n359311 , n11634 );
buf ( n359312 , n359311 );
nand ( n11637 , n11627 , n359312 );
buf ( n359314 , n11637 );
not ( n11639 , n359314 );
or ( n11640 , n11622 , n11639 );
buf ( n359317 , n359301 );
buf ( n359318 , n359308 );
nand ( n11643 , n359317 , n359318 );
buf ( n359320 , n11643 );
nand ( n11645 , n11640 , n359320 );
not ( n11646 , n11645 );
or ( n11647 , n9855 , n11646 );
nand ( n11648 , n357388 , n357536 );
buf ( n11649 , n11648 );
nand ( n11650 , n11647 , n11649 );
xor ( n11651 , n354127 , n354149 );
and ( n11652 , n11651 , n354275 );
and ( n11653 , n354127 , n354149 );
or ( n11654 , n11652 , n11653 );
buf ( n359331 , n11654 );
buf ( n359332 , n359331 );
buf ( n359333 , n352149 );
not ( n11658 , n359333 );
buf ( n359335 , n602 );
not ( n11660 , n359335 );
buf ( n359337 , n7360 );
not ( n11662 , n359337 );
or ( n11663 , n11660 , n11662 );
buf ( n359340 , n7363 );
buf ( n359341 , n349406 );
nand ( n11666 , n359340 , n359341 );
buf ( n359343 , n11666 );
buf ( n359344 , n359343 );
nand ( n11669 , n11663 , n359344 );
buf ( n359346 , n11669 );
buf ( n359347 , n359346 );
not ( n11672 , n359347 );
or ( n11673 , n11658 , n11672 );
buf ( n359350 , n354066 );
buf ( n359351 , n354113 );
nand ( n11676 , n359350 , n359351 );
buf ( n359353 , n11676 );
buf ( n359354 , n359353 );
nand ( n11679 , n11673 , n359354 );
buf ( n359356 , n11679 );
buf ( n359357 , n359356 );
xor ( n11682 , n359332 , n359357 );
xor ( n11683 , n354156 , n354181 );
and ( n11684 , n11683 , n354272 );
and ( n11685 , n354156 , n354181 );
or ( n11686 , n11684 , n11685 );
buf ( n359363 , n11686 );
buf ( n359364 , n359363 );
buf ( n359365 , n1722 );
not ( n11690 , n359365 );
buf ( n359367 , n600 );
not ( n11692 , n359367 );
buf ( n359369 , n354087 );
not ( n11694 , n359369 );
or ( n11695 , n11692 , n11694 );
buf ( n359372 , n6460 );
buf ( n359373 , n9814 );
nand ( n11698 , n359372 , n359373 );
buf ( n359375 , n11698 );
buf ( n359376 , n359375 );
nand ( n11701 , n11695 , n359376 );
buf ( n359378 , n11701 );
buf ( n359379 , n359378 );
not ( n11704 , n359379 );
or ( n11705 , n11690 , n11704 );
nand ( n11706 , n354146 , n351924 );
buf ( n359383 , n11706 );
nand ( n11708 , n11705 , n359383 );
buf ( n359385 , n11708 );
buf ( n359386 , n359385 );
xor ( n11711 , n359364 , n359386 );
xor ( n11712 , n354199 , n354236 );
and ( n11713 , n11712 , n354269 );
and ( n11714 , n354199 , n354236 );
or ( n11715 , n11713 , n11714 );
buf ( n359392 , n11715 );
buf ( n359393 , n359392 );
not ( n11718 , n4361 );
not ( n11719 , n598 );
not ( n11720 , n351870 );
or ( n11721 , n11719 , n11720 );
buf ( n359398 , n357858 );
buf ( n359399 , n347312 );
nand ( n11724 , n359398 , n359399 );
buf ( n359401 , n11724 );
nand ( n11726 , n11721 , n359401 );
not ( n11727 , n11726 );
or ( n11728 , n11718 , n11727 );
nand ( n11729 , n354170 , n4443 );
nand ( n11730 , n11728 , n11729 );
buf ( n359407 , n11730 );
xor ( n11732 , n359393 , n359407 );
not ( n11733 , n349035 );
not ( n11734 , n351958 );
not ( n11735 , n348975 );
or ( n11736 , n11734 , n11735 );
nand ( n11737 , n594 , n351952 );
nand ( n11738 , n11736 , n11737 );
not ( n11739 , n11738 );
or ( n11740 , n11733 , n11739 );
buf ( n359417 , n6504 );
buf ( n359418 , n1397 );
nand ( n11743 , n359417 , n359418 );
buf ( n359420 , n11743 );
nand ( n11745 , n11740 , n359420 );
buf ( n359422 , n11745 );
buf ( n359423 , n349067 );
buf ( n359424 , n592 );
and ( n11749 , n359423 , n359424 );
buf ( n359426 , n11749 );
buf ( n359427 , n359426 );
buf ( n359428 , n348946 );
not ( n11753 , n359428 );
buf ( n359430 , n592 );
not ( n11755 , n4298 );
buf ( n359432 , n11755 );
xor ( n11757 , n359430 , n359432 );
buf ( n359434 , n11757 );
buf ( n359435 , n359434 );
not ( n11760 , n359435 );
or ( n11761 , n11753 , n11760 );
buf ( n359438 , n354220 );
buf ( n359439 , n1250 );
nand ( n11764 , n359438 , n359439 );
buf ( n359441 , n11764 );
buf ( n359442 , n359441 );
nand ( n11767 , n11761 , n359442 );
buf ( n359444 , n11767 );
buf ( n359445 , n359444 );
xor ( n11770 , n359427 , n359445 );
xor ( n11771 , n354204 , n354226 );
and ( n11772 , n11771 , n354233 );
and ( n11773 , n354204 , n354226 );
or ( n11774 , n11772 , n11773 );
buf ( n359451 , n11774 );
buf ( n359452 , n359451 );
xor ( n11777 , n11770 , n359452 );
buf ( n359454 , n11777 );
buf ( n359455 , n359454 );
xor ( n11780 , n359422 , n359455 );
buf ( n359457 , n347319 );
not ( n11782 , n359457 );
buf ( n359459 , n596 );
not ( n11784 , n359459 );
buf ( n359461 , n7445 );
not ( n11786 , n359461 );
or ( n11787 , n11784 , n11786 );
buf ( n359464 , n4388 );
buf ( n359465 , n348865 );
nand ( n11790 , n359464 , n359465 );
buf ( n359467 , n11790 );
buf ( n359468 , n359467 );
nand ( n11793 , n11787 , n359468 );
buf ( n359470 , n11793 );
buf ( n359471 , n359470 );
not ( n11796 , n359471 );
or ( n11797 , n11782 , n11796 );
buf ( n359474 , n354258 );
buf ( n359475 , n348898 );
nand ( n11800 , n359474 , n359475 );
buf ( n359477 , n11800 );
buf ( n359478 , n359477 );
nand ( n11803 , n11797 , n359478 );
buf ( n359480 , n11803 );
buf ( n359481 , n359480 );
xor ( n11806 , n11780 , n359481 );
buf ( n359483 , n11806 );
buf ( n359484 , n359483 );
xor ( n11809 , n11732 , n359484 );
buf ( n359486 , n11809 );
buf ( n359487 , n359486 );
xor ( n11812 , n11711 , n359487 );
buf ( n359489 , n11812 );
buf ( n359490 , n359489 );
xor ( n11815 , n11682 , n359490 );
buf ( n359492 , n11815 );
buf ( n359493 , n359492 );
xor ( n11818 , n355291 , n356034 );
and ( n11819 , n11818 , n357383 );
and ( n11820 , n355291 , n356034 );
or ( n11821 , n11819 , n11820 );
buf ( n359498 , n11821 );
buf ( n359499 , n359498 );
xor ( n11824 , n359493 , n359499 );
xor ( n11825 , n352140 , n354120 );
and ( n11826 , n11825 , n354278 );
and ( n11827 , n352140 , n354120 );
or ( n11828 , n11826 , n11827 );
buf ( n359505 , n11828 );
buf ( n359506 , n359505 );
buf ( n359507 , n6600 );
not ( n11832 , n359507 );
and ( n11833 , n604 , n357355 );
not ( n11834 , n604 );
and ( n11835 , n11834 , n9664 );
or ( n11836 , n11833 , n11835 );
buf ( n359513 , n11836 );
not ( n11838 , n359513 );
or ( n11839 , n11832 , n11838 );
buf ( n359516 , n8335 );
buf ( n359517 , n355075 );
nand ( n11842 , n359516 , n359517 );
buf ( n359519 , n11842 );
buf ( n359520 , n359519 );
nand ( n11845 , n11839 , n359520 );
buf ( n359522 , n11845 );
buf ( n359523 , n359522 );
xor ( n11848 , n359506 , n359523 );
buf ( n359525 , n607 );
not ( n11850 , n359525 );
buf ( n359527 , n606 );
not ( n11852 , n359527 );
nor ( n11853 , n9609 , n9603 );
not ( n11854 , n11853 );
not ( n11855 , n8297 );
or ( n11856 , n11854 , n11855 );
not ( n11857 , n8485 );
not ( n11858 , n8981 );
and ( n11859 , n11857 , n11858 );
nor ( n11860 , n11859 , n9603 );
nand ( n11861 , n8982 , n8279 );
and ( n11862 , n11860 , n11861 );
nor ( n11863 , n11862 , n9601 );
nand ( n11864 , n11856 , n11863 );
xor ( n11865 , n356889 , n356890 );
and ( n11866 , n11865 , n356907 );
and ( n11867 , n356889 , n356890 );
or ( n11868 , n11866 , n11867 );
buf ( n359545 , n11868 );
buf ( n359546 , n359545 );
buf ( n359547 , n556 );
buf ( n359548 , n560 );
and ( n11873 , n359547 , n359548 );
buf ( n359550 , n11873 );
buf ( n359551 , n359550 );
buf ( n359552 , n9297 );
not ( n11877 , n359552 );
buf ( n359554 , n351330 );
not ( n11879 , n359554 );
or ( n11880 , n11877 , n11879 );
buf ( n359557 , n3650 );
buf ( n359558 , n550 );
buf ( n359559 , n564 );
xor ( n11884 , n359558 , n359559 );
buf ( n359561 , n11884 );
buf ( n359562 , n359561 );
nand ( n11887 , n359557 , n359562 );
buf ( n359564 , n11887 );
buf ( n359565 , n359564 );
nand ( n11890 , n11880 , n359565 );
buf ( n359567 , n11890 );
buf ( n359568 , n359567 );
xor ( n11893 , n359551 , n359568 );
buf ( n359570 , n357018 );
not ( n11895 , n359570 );
buf ( n359572 , n2236 );
not ( n11897 , n359572 );
or ( n11898 , n11895 , n11897 );
buf ( n359575 , n349933 );
xor ( n11900 , n568 , n546 );
buf ( n359577 , n11900 );
nand ( n11902 , n359575 , n359577 );
buf ( n359579 , n11902 );
buf ( n359580 , n359579 );
nand ( n11905 , n11898 , n359580 );
buf ( n359582 , n11905 );
buf ( n359583 , n359582 );
xor ( n11908 , n11893 , n359583 );
buf ( n359585 , n11908 );
buf ( n359586 , n359585 );
xor ( n11911 , n359546 , n359586 );
not ( n11912 , n357000 );
not ( n11913 , n8604 );
or ( n11914 , n11912 , n11913 );
buf ( n359591 , n352295 );
buf ( n359592 , n552 );
buf ( n359593 , n562 );
xor ( n11918 , n359592 , n359593 );
buf ( n359595 , n11918 );
buf ( n359596 , n359595 );
nand ( n11921 , n359591 , n359596 );
buf ( n359598 , n11921 );
nand ( n11923 , n11914 , n359598 );
not ( n11924 , n11923 );
buf ( n359601 , n356882 );
not ( n11926 , n359601 );
buf ( n359603 , n9186 );
not ( n11928 , n359603 );
or ( n11929 , n11926 , n11928 );
buf ( n359606 , n5407 );
buf ( n359607 , n554 );
buf ( n359608 , n560 );
xor ( n11933 , n359607 , n359608 );
buf ( n359610 , n11933 );
buf ( n359611 , n359610 );
nand ( n11936 , n359606 , n359611 );
buf ( n359613 , n11936 );
buf ( n359614 , n359613 );
nand ( n11939 , n11929 , n359614 );
buf ( n359616 , n11939 );
and ( n11941 , n11924 , n359616 );
not ( n11942 , n11924 );
not ( n11943 , n359616 );
and ( n11944 , n11942 , n11943 );
nor ( n11945 , n11941 , n11944 );
and ( n11946 , n11945 , n356906 );
not ( n11947 , n11945 );
and ( n11948 , n11947 , n356903 );
nor ( n11949 , n11946 , n11948 );
buf ( n359626 , n11949 );
xor ( n11951 , n11911 , n359626 );
buf ( n359628 , n11951 );
buf ( n359629 , n359628 );
xor ( n11954 , n356957 , n357031 );
and ( n11955 , n11954 , n357043 );
and ( n11956 , n356957 , n357031 );
or ( n11957 , n11955 , n11956 );
buf ( n359634 , n11957 );
buf ( n359635 , n359634 );
xor ( n11960 , n359629 , n359635 );
xor ( n11961 , n356967 , n356978 );
and ( n11962 , n11961 , n357028 );
and ( n11963 , n356967 , n356978 );
or ( n11964 , n11962 , n11963 );
buf ( n359641 , n11964 );
buf ( n359642 , n359641 );
xor ( n11967 , n356836 , n356850 );
and ( n11968 , n11967 , n356868 );
and ( n11969 , n356836 , n356850 );
or ( n11970 , n11968 , n11969 );
buf ( n359647 , n11970 );
buf ( n359648 , n359647 );
xor ( n11973 , n356990 , n357007 );
and ( n11974 , n11973 , n357025 );
and ( n11975 , n356990 , n357007 );
or ( n11976 , n11974 , n11975 );
buf ( n359653 , n11976 );
buf ( n359654 , n359653 );
xor ( n11979 , n359648 , n359654 );
buf ( n359656 , n356861 );
not ( n11981 , n359656 );
buf ( n359658 , n354366 );
not ( n11983 , n359658 );
or ( n11984 , n11981 , n11983 );
buf ( n359661 , n348473 );
buf ( n359662 , n544 );
buf ( n359663 , n570 );
xor ( n11988 , n359662 , n359663 );
buf ( n359665 , n11988 );
buf ( n359666 , n359665 );
nand ( n11991 , n359661 , n359666 );
buf ( n359668 , n11991 );
buf ( n359669 , n359668 );
nand ( n11994 , n11984 , n359669 );
buf ( n359671 , n11994 );
buf ( n359672 , n359671 );
or ( n11997 , n347382 , n3241 );
nand ( n11998 , n11997 , n572 );
buf ( n359675 , n11998 );
xor ( n12000 , n359672 , n359675 );
buf ( n359677 , n9155 );
not ( n12002 , n359677 );
buf ( n359679 , n350874 );
not ( n12004 , n359679 );
or ( n12005 , n12002 , n12004 );
buf ( n359682 , n2550 );
buf ( n359683 , n548 );
buf ( n359684 , n566 );
xor ( n12009 , n359683 , n359684 );
buf ( n359686 , n12009 );
buf ( n359687 , n359686 );
nand ( n12012 , n359682 , n359687 );
buf ( n359689 , n12012 );
buf ( n359690 , n359689 );
nand ( n12015 , n12005 , n359690 );
buf ( n359692 , n12015 );
buf ( n359693 , n359692 );
xor ( n12018 , n12000 , n359693 );
buf ( n359695 , n12018 );
buf ( n359696 , n359695 );
xor ( n12021 , n11979 , n359696 );
buf ( n359698 , n12021 );
buf ( n359699 , n359698 );
xor ( n12024 , n359642 , n359699 );
xor ( n12025 , n356871 , n356910 );
and ( n12026 , n12025 , n356917 );
and ( n12027 , n356871 , n356910 );
or ( n12028 , n12026 , n12027 );
buf ( n359705 , n12028 );
buf ( n359706 , n359705 );
xor ( n12031 , n12024 , n359706 );
buf ( n359708 , n12031 );
buf ( n359709 , n359708 );
xor ( n12034 , n11960 , n359709 );
buf ( n359711 , n12034 );
buf ( n359712 , n359711 );
xor ( n12037 , n357066 , n357072 );
and ( n12038 , n12037 , n357265 );
and ( n12039 , n357066 , n357072 );
or ( n12040 , n12038 , n12039 );
buf ( n359717 , n12040 );
buf ( n359718 , n359717 );
xor ( n12043 , n359712 , n359718 );
xor ( n12044 , n356920 , n356941 );
and ( n12045 , n12044 , n357046 );
and ( n12046 , n356920 , n356941 );
or ( n12047 , n12045 , n12046 );
buf ( n359724 , n12047 );
buf ( n359725 , n359724 );
xor ( n12050 , n357167 , n357173 );
and ( n12051 , n12050 , n357262 );
and ( n12052 , n357167 , n357173 );
or ( n12053 , n12051 , n12052 );
buf ( n359730 , n12053 );
buf ( n359731 , n359730 );
xor ( n12056 , n359725 , n359731 );
xor ( n12057 , n357136 , n357152 );
and ( n12058 , n12057 , n357154 );
and ( n12059 , n357136 , n357152 );
or ( n12060 , n12058 , n12059 );
buf ( n359737 , n12060 );
buf ( n359738 , n359737 );
buf ( n359739 , n556 );
buf ( n359740 , n576 );
and ( n12065 , n359739 , n359740 );
buf ( n359742 , n12065 );
buf ( n359743 , n359742 );
not ( n12068 , n357208 );
not ( n12069 , n3869 );
not ( n12070 , n12069 );
or ( n12071 , n12068 , n12070 );
not ( n12072 , n550 );
not ( n12073 , n6052 );
or ( n12074 , n12072 , n12073 );
nand ( n12075 , n5123 , n580 );
nand ( n12076 , n12074 , n12075 );
nand ( n12077 , n3345 , n12076 );
nand ( n12078 , n12071 , n12077 );
buf ( n359755 , n12078 );
xor ( n12080 , n359743 , n359755 );
buf ( n359757 , n9551 );
not ( n12082 , n359757 );
buf ( n359759 , n2471 );
not ( n12084 , n359759 );
or ( n12085 , n12082 , n12084 );
buf ( n359762 , n348617 );
xor ( n12087 , n584 , n546 );
buf ( n359764 , n12087 );
nand ( n12089 , n359762 , n359764 );
buf ( n359766 , n12089 );
buf ( n359767 , n359766 );
nand ( n12092 , n12085 , n359767 );
buf ( n359769 , n12092 );
buf ( n359770 , n359769 );
xor ( n12095 , n12080 , n359770 );
buf ( n359772 , n12095 );
buf ( n359773 , n359772 );
xor ( n12098 , n359738 , n359773 );
buf ( n359775 , n357129 );
not ( n12100 , n359775 );
buf ( n359777 , n356440 );
not ( n12102 , n359777 );
or ( n12103 , n12100 , n12102 );
buf ( n359780 , n356446 );
buf ( n359781 , n554 );
buf ( n359782 , n576 );
xor ( n12107 , n359781 , n359782 );
buf ( n359784 , n12107 );
buf ( n359785 , n359784 );
nand ( n12110 , n359780 , n359785 );
buf ( n359787 , n12110 );
buf ( n359788 , n359787 );
nand ( n12113 , n12103 , n359788 );
buf ( n359790 , n12113 );
buf ( n359791 , n359790 );
buf ( n359792 , n357224 );
not ( n12117 , n359792 );
buf ( n359794 , n355543 );
not ( n12119 , n359794 );
or ( n12120 , n12117 , n12119 );
buf ( n359797 , n352491 );
xor ( n12122 , n578 , n552 );
buf ( n359799 , n12122 );
nand ( n12124 , n359797 , n359799 );
buf ( n359801 , n12124 );
buf ( n359802 , n359801 );
nand ( n12127 , n12120 , n359802 );
buf ( n359804 , n12127 );
buf ( n359805 , n359804 );
xor ( n12130 , n359791 , n359805 );
buf ( n359807 , n12130 );
buf ( n359808 , n359807 );
buf ( n359809 , n357148 );
xor ( n12134 , n359808 , n359809 );
buf ( n359811 , n12134 );
buf ( n359812 , n359811 );
xor ( n12137 , n12098 , n359812 );
buf ( n359814 , n12137 );
buf ( n359815 , n359814 );
xor ( n12140 , n357180 , n357252 );
and ( n12141 , n12140 , n357259 );
and ( n12142 , n357180 , n357252 );
or ( n12143 , n12141 , n12142 );
buf ( n359820 , n12143 );
buf ( n359821 , n359820 );
xor ( n12146 , n359815 , n359821 );
xor ( n12147 , n357186 , n357203 );
and ( n12148 , n12147 , n357249 );
and ( n12149 , n357186 , n357203 );
or ( n12150 , n12148 , n12149 );
buf ( n359827 , n12150 );
buf ( n359828 , n359827 );
buf ( n359829 , n357117 );
buf ( n359830 , n357097 );
or ( n12155 , n359829 , n359830 );
buf ( n359832 , n357089 );
nand ( n12157 , n12155 , n359832 );
buf ( n359834 , n12157 );
buf ( n359835 , n359834 );
buf ( n359836 , n357117 );
buf ( n359837 , n357097 );
nand ( n12162 , n359836 , n359837 );
buf ( n359839 , n12162 );
buf ( n359840 , n359839 );
nand ( n12165 , n359835 , n359840 );
buf ( n359842 , n12165 );
buf ( n359843 , n359842 );
xor ( n12168 , n357214 , n357231 );
and ( n12169 , n12168 , n357246 );
and ( n12170 , n357214 , n357231 );
or ( n12171 , n12169 , n12170 );
buf ( n359848 , n12171 );
buf ( n359849 , n359848 );
xor ( n12174 , n359843 , n359849 );
buf ( n359851 , n9423 );
not ( n12176 , n359851 );
buf ( n359853 , n350699 );
not ( n12178 , n359853 );
or ( n12179 , n12176 , n12178 );
buf ( n359856 , n350705 );
buf ( n359857 , n548 );
buf ( n359858 , n582 );
xor ( n12183 , n359857 , n359858 );
buf ( n359860 , n12183 );
buf ( n359861 , n359860 );
nand ( n12186 , n359856 , n359861 );
buf ( n359863 , n12186 );
buf ( n359864 , n359863 );
nand ( n12189 , n12179 , n359864 );
buf ( n359866 , n12189 );
buf ( n359867 , n357083 );
not ( n12192 , n359867 );
buf ( n359869 , n350110 );
not ( n12194 , n359869 );
or ( n12195 , n12192 , n12194 );
buf ( n359872 , n347530 );
buf ( n359873 , n544 );
buf ( n359874 , n586 );
xor ( n12199 , n359873 , n359874 );
buf ( n359876 , n12199 );
buf ( n359877 , n359876 );
nand ( n12202 , n359872 , n359877 );
buf ( n359879 , n12202 );
buf ( n359880 , n359879 );
nand ( n12205 , n12195 , n359880 );
buf ( n359882 , n12205 );
xor ( n12207 , n359866 , n359882 );
not ( n12208 , n347565 );
buf ( n359885 , n12208 );
not ( n12210 , n359885 );
buf ( n359887 , n350130 );
not ( n12212 , n359887 );
or ( n12213 , n12210 , n12212 );
buf ( n359890 , n588 );
nand ( n12215 , n12213 , n359890 );
buf ( n359892 , n12215 );
xor ( n12217 , n12207 , n359892 );
buf ( n359894 , n12217 );
xor ( n12219 , n12174 , n359894 );
buf ( n359896 , n12219 );
buf ( n359897 , n359896 );
xor ( n12222 , n359828 , n359897 );
xor ( n12223 , n357119 , n357157 );
and ( n12224 , n12223 , n357164 );
and ( n12225 , n357119 , n357157 );
or ( n12226 , n12224 , n12225 );
buf ( n359903 , n12226 );
buf ( n359904 , n359903 );
xor ( n12229 , n12222 , n359904 );
buf ( n359906 , n12229 );
buf ( n359907 , n359906 );
xor ( n12232 , n12146 , n359907 );
buf ( n359909 , n12232 );
buf ( n359910 , n359909 );
xor ( n12235 , n12056 , n359910 );
buf ( n359912 , n12235 );
buf ( n359913 , n359912 );
xor ( n12238 , n12043 , n359913 );
buf ( n359915 , n12238 );
xor ( n12240 , n357049 , n357055 );
and ( n12241 , n12240 , n357268 );
and ( n12242 , n357049 , n357055 );
or ( n12243 , n12241 , n12242 );
buf ( n359920 , n12243 );
nor ( n12245 , n359915 , n359920 );
buf ( n12246 , n12245 );
buf ( n359923 , n359915 );
buf ( n359924 , n359920 );
and ( n12249 , n359923 , n359924 );
buf ( n359926 , n12249 );
nor ( n12251 , n12246 , n359926 );
not ( n12252 , n12251 );
not ( n12253 , n12252 );
buf ( n359930 , n9139 );
not ( n12255 , n359930 );
buf ( n359932 , n9588 );
not ( n12257 , n359932 );
or ( n12258 , n12255 , n12257 );
buf ( n359935 , n357280 );
nand ( n12260 , n12258 , n359935 );
buf ( n359937 , n12260 );
buf ( n359938 , n359937 );
not ( n12263 , n359938 );
buf ( n359940 , n12263 );
and ( n12265 , n9588 , n9134 );
nand ( n12266 , n12265 , n8487 );
nand ( n12267 , n359940 , n12266 );
not ( n12268 , n12267 );
or ( n12269 , n12253 , n12268 );
nand ( n12270 , n359940 , n12266 , n12251 );
nand ( n12271 , n12269 , n12270 );
not ( n12272 , n12271 );
not ( n12273 , n9124 );
not ( n12274 , n9005 );
or ( n12275 , n12273 , n12274 );
nand ( n12276 , n12275 , n9126 );
xor ( n12277 , n9047 , n9051 );
and ( n12278 , n12277 , n9117 );
and ( n12279 , n9047 , n9051 );
or ( n12280 , n12278 , n12279 );
not ( n12281 , n12280 );
not ( n12282 , n7272 );
not ( n12283 , n9093 );
or ( n12284 , n12282 , n12283 );
not ( n12285 , n5990 );
and ( n12286 , n1788 , n5761 );
not ( n12287 , n1788 );
and ( n12288 , n12287 , n546 );
or ( n12289 , n12286 , n12288 );
nand ( n12290 , n12285 , n12289 );
nand ( n12291 , n12284 , n12290 );
not ( n12292 , n8215 );
not ( n12293 , n1751 );
nand ( n12294 , n12293 , n7283 );
nand ( n12295 , n4114 , n544 );
nand ( n12296 , n12294 , n12295 );
not ( n12297 , n12296 );
or ( n12298 , n12292 , n12297 );
nand ( n12299 , n9072 , n8223 );
nand ( n12300 , n12298 , n12299 );
xor ( n12301 , n12291 , n12300 );
not ( n12302 , n1875 );
not ( n12303 , n1880 );
not ( n12304 , n353641 );
or ( n12305 , n12303 , n12304 );
nand ( n12306 , n550 , n4057 );
nand ( n12307 , n12305 , n12306 );
not ( n12308 , n12307 );
or ( n12309 , n12302 , n12308 );
nand ( n12310 , n9036 , n4078 );
nand ( n12311 , n12309 , n12310 );
xor ( n12312 , n12301 , n12311 );
xor ( n12313 , n9088 , n9098 );
and ( n12314 , n12313 , n9109 );
and ( n12315 , n9088 , n9098 );
or ( n12316 , n12314 , n12315 );
xor ( n12317 , n12312 , n12316 );
not ( n12318 , n1925 );
not ( n12319 , n554 );
not ( n12320 , n7245 );
or ( n12321 , n12319 , n12320 );
not ( n12322 , n7245 );
nand ( n12323 , n12322 , n348175 );
nand ( n12324 , n12321 , n12323 );
not ( n12325 , n12324 );
or ( n12326 , n12318 , n12325 );
nand ( n12327 , n9043 , n1022 );
nand ( n12328 , n12326 , n12327 );
not ( n12329 , n5735 );
not ( n12330 , n548 );
not ( n12331 , n1975 );
or ( n12332 , n12330 , n12331 );
nand ( n12333 , n1974 , n351773 );
nand ( n12334 , n12332 , n12333 );
not ( n12335 , n12334 );
or ( n12336 , n12329 , n12335 );
nand ( n12337 , n9086 , n5751 );
nand ( n12338 , n12336 , n12337 );
xor ( n12339 , n12328 , n12338 );
not ( n12340 , n1871 );
not ( n12341 , n9103 );
or ( n12342 , n12340 , n12341 );
and ( n12343 , n552 , n6035 );
not ( n12344 , n552 );
and ( n12345 , n12344 , n6034 );
or ( n12346 , n12343 , n12345 );
nand ( n12347 , n12346 , n1011 );
nand ( n12348 , n12342 , n12347 );
xor ( n12349 , n12339 , n12348 );
xor ( n12350 , n12317 , n12349 );
and ( n12351 , n9076 , n9069 );
not ( n12352 , n348153 );
not ( n12353 , n9025 );
or ( n12354 , n12352 , n12353 );
nand ( n12355 , n12354 , n6011 );
not ( n12356 , n544 );
not ( n12357 , n9064 );
or ( n12358 , n12356 , n12357 );
nand ( n12359 , n12358 , n9062 );
xor ( n12360 , n12355 , n12359 );
not ( n12361 , n1856 );
nand ( n12362 , n12361 , n544 );
xor ( n12363 , n12360 , n12362 );
xor ( n12364 , n12351 , n12363 );
xor ( n12365 , n9029 , n9038 );
and ( n12366 , n12365 , n9045 );
and ( n12367 , n9029 , n9038 );
or ( n12368 , n12366 , n12367 );
xor ( n12369 , n12364 , n12368 );
xor ( n12370 , n9060 , n9077 );
and ( n12371 , n12370 , n9110 );
and ( n12372 , n9060 , n9077 );
or ( n12373 , n12371 , n12372 );
xor ( n12374 , n12369 , n12373 );
xor ( n12375 , n9010 , n9014 );
and ( n12376 , n12375 , n9046 );
and ( n12377 , n9010 , n9014 );
or ( n12378 , n12376 , n12377 );
xor ( n12379 , n12374 , n12378 );
xor ( n12380 , n12350 , n12379 );
xor ( n12381 , n9056 , n9111 );
and ( n12382 , n12381 , n9116 );
and ( n12383 , n9056 , n9111 );
or ( n12384 , n12382 , n12383 );
xor ( n12385 , n12380 , n12384 );
buf ( n12386 , n12385 );
not ( n12387 , n12386 );
or ( n12388 , n12281 , n12387 );
nor ( n12389 , n12385 , n12280 );
not ( n12390 , n12389 );
nand ( n12391 , n12388 , n12390 );
not ( n12392 , n12391 );
and ( n12393 , n12276 , n12392 );
not ( n12394 , n12276 );
and ( n12395 , n12394 , n12391 );
nor ( n12396 , n12393 , n12395 );
nor ( n12397 , n12272 , n12396 );
not ( n12398 , n12397 );
nand ( n12399 , n12396 , n12272 );
buf ( n12400 , n12399 );
nand ( n12401 , n12398 , n12400 );
and ( n12402 , n11864 , n12401 );
not ( n12403 , n11864 );
not ( n12404 , n12401 );
and ( n12405 , n12403 , n12404 );
nor ( n12406 , n12402 , n12405 );
not ( n12407 , n12406 );
buf ( n360084 , n12407 );
buf ( n12409 , n360084 );
buf ( n360086 , n12409 );
not ( n12411 , n360086 );
not ( n12412 , n357316 );
nor ( n12413 , n12412 , n8991 );
nand ( n12414 , n8323 , n12413 );
not ( n12415 , n12414 );
or ( n12416 , n12411 , n12415 );
not ( n12417 , n12414 );
not ( n12418 , n360086 );
nand ( n12419 , n12417 , n12418 );
nand ( n12420 , n12416 , n12419 );
buf ( n360097 , n12420 );
not ( n12422 , n360097 );
buf ( n360099 , n12422 );
buf ( n360100 , n360099 );
not ( n12425 , n360100 );
or ( n12426 , n11852 , n12425 );
buf ( n360103 , n12420 );
buf ( n12428 , n360103 );
buf ( n360105 , n12428 );
buf ( n360106 , n360105 );
buf ( n360107 , n9642 );
nand ( n12432 , n360106 , n360107 );
buf ( n360109 , n12432 );
buf ( n360110 , n360109 );
nand ( n12435 , n12426 , n360110 );
buf ( n360112 , n12435 );
buf ( n360113 , n360112 );
not ( n12438 , n360113 );
or ( n12439 , n11850 , n12438 );
buf ( n360116 , n357336 );
buf ( n360117 , n357376 );
nand ( n12442 , n360116 , n360117 );
buf ( n360119 , n12442 );
buf ( n360120 , n360119 );
nand ( n12445 , n12439 , n360120 );
buf ( n360122 , n12445 );
buf ( n360123 , n360122 );
xor ( n12448 , n11848 , n360123 );
buf ( n360125 , n12448 );
buf ( n360126 , n360125 );
xor ( n12451 , n11824 , n360126 );
buf ( n360128 , n12451 );
xor ( n12453 , n354281 , n355284 );
and ( n12454 , n12453 , n357386 );
and ( n12455 , n354281 , n355284 );
or ( n12456 , n12454 , n12455 );
buf ( n360133 , n12456 );
or ( n12458 , n360128 , n360133 );
buf ( n360135 , n12458 );
buf ( n360136 , n360128 );
buf ( n360137 , n360133 );
nand ( n12462 , n360136 , n360137 );
buf ( n360139 , n12462 );
buf ( n360140 , n360139 );
buf ( n12465 , n360140 );
buf ( n360142 , n12465 );
buf ( n360143 , n360142 );
nand ( n12468 , n360135 , n360143 );
buf ( n360145 , n12468 );
xnor ( n12470 , n11650 , n360145 );
buf ( n12471 , n12470 );
not ( n12472 , n359301 );
not ( n12473 , n359308 );
or ( n12474 , n12472 , n12473 );
nand ( n12475 , n12474 , n359314 );
buf ( n360152 , n11621 );
buf ( n12477 , n360152 );
buf ( n360154 , n12477 );
xnor ( n12479 , n12475 , n360154 );
buf ( n12480 , n12479 );
not ( n12481 , n4370 );
buf ( n12482 , n1060 );
buf ( n12483 , n3603 );
buf ( n12484 , n1129 );
buf ( n12485 , n920 );
buf ( n12486 , n352888 );
buf ( n12487 , n352640 );
buf ( n12488 , n351640 );
buf ( n12489 , n351089 );
buf ( n12490 , n350495 );
buf ( n12491 , n354581 );
buf ( n12492 , n4751 );
buf ( n12493 , n347580 );
buf ( n12494 , n2323 );
buf ( n12495 , n348532 );
buf ( n12496 , n347428 );
buf ( n12497 , n354608 );
buf ( n12498 , n347718 );
buf ( n12499 , n350178 );
buf ( n12500 , n4992 );
buf ( n12501 , n352439 );
buf ( n12502 , n350971 );
buf ( n12503 , n350808 );
buf ( n12504 , n357264 );
not ( n12505 , n9616 );
nand ( n12506 , n9598 , n9132 );
and ( n12507 , n12399 , n12506 );
not ( n12508 , n12507 );
or ( n12509 , n12505 , n12508 );
not ( n12510 , n12271 );
nand ( n12511 , n12510 , n12396 );
and ( n12512 , n12511 , n9601 );
nor ( n12513 , n12512 , n12397 );
nand ( n12514 , n12509 , n12513 );
not ( n12515 , n12514 );
nand ( n12516 , n9610 , n12507 );
not ( n12517 , n12516 );
nand ( n12518 , n12517 , n8354 );
nand ( n12519 , n12515 , n12518 );
nor ( n12520 , n12389 , n9123 );
not ( n12521 , n12520 );
not ( n12522 , n9005 );
or ( n12523 , n12521 , n12522 );
not ( n12524 , n12280 );
not ( n12525 , n12385 );
or ( n12526 , n12524 , n12525 );
nand ( n12527 , n12526 , n9125 );
nand ( n12528 , n12527 , n12390 );
nand ( n12529 , n12523 , n12528 );
buf ( n12530 , n12529 );
xor ( n12531 , n12328 , n12338 );
and ( n12532 , n12531 , n12348 );
and ( n12533 , n12328 , n12338 );
or ( n12534 , n12532 , n12533 );
xor ( n12535 , n12291 , n12300 );
and ( n12536 , n12535 , n12311 );
and ( n12537 , n12291 , n12300 );
or ( n12538 , n12536 , n12537 );
xor ( n12539 , n12534 , n12538 );
not ( n12540 , n1022 );
not ( n12541 , n12324 );
or ( n12542 , n12540 , n12541 );
buf ( n12543 , n8185 );
and ( n12544 , n554 , n12543 );
not ( n12545 , n554 );
not ( n12546 , n8185 );
and ( n12547 , n12545 , n12546 );
nor ( n12548 , n12544 , n12547 );
nand ( n12549 , n12548 , n1925 );
nand ( n12550 , n12542 , n12549 );
not ( n12551 , n5751 );
not ( n12552 , n12334 );
or ( n12553 , n12551 , n12552 );
and ( n12554 , n2071 , n548 );
not ( n12555 , n2071 );
and ( n12556 , n12555 , n351773 );
nor ( n12557 , n12554 , n12556 );
buf ( n12558 , n12557 );
nand ( n12559 , n12558 , n8133 );
nand ( n12560 , n12553 , n12559 );
xor ( n12561 , n12550 , n12560 );
not ( n12562 , n1871 );
not ( n12563 , n12346 );
or ( n12564 , n12562 , n12563 );
and ( n12565 , n552 , n6082 );
not ( n12566 , n552 );
and ( n12567 , n12566 , n6081 );
or ( n12568 , n12565 , n12567 );
nand ( n12569 , n12568 , n4109 );
nand ( n12570 , n12564 , n12569 );
xor ( n12571 , n12561 , n12570 );
xor ( n12572 , n12539 , n12571 );
xor ( n12573 , n12351 , n12363 );
and ( n12574 , n12573 , n12368 );
and ( n12575 , n12351 , n12363 );
or ( n12576 , n12574 , n12575 );
xor ( n12577 , n12355 , n12359 );
and ( n12578 , n12577 , n12362 );
and ( n12579 , n12355 , n12359 );
or ( n12580 , n12578 , n12579 );
not ( n12581 , n348089 );
not ( n12582 , n348152 );
or ( n12583 , n12581 , n12582 );
nand ( n12584 , n12583 , n556 );
and ( n12585 , n544 , n9071 );
xor ( n12586 , n12584 , n12585 );
not ( n12587 , n12362 );
xor ( n12588 , n12586 , n12587 );
xor ( n12589 , n12580 , n12588 );
not ( n12590 , n5757 );
not ( n12591 , n546 );
not ( n12592 , n5827 );
or ( n12593 , n12591 , n12592 );
nand ( n12594 , n5761 , n1843 );
nand ( n12595 , n12593 , n12594 );
not ( n12596 , n12595 );
or ( n12597 , n12590 , n12596 );
nand ( n12598 , n12289 , n8381 );
nand ( n12599 , n12597 , n12598 );
not ( n12600 , n8215 );
xor ( n12601 , n544 , n997 );
not ( n12602 , n12601 );
or ( n12603 , n12600 , n12602 );
not ( n12604 , n12294 );
not ( n12605 , n12295 );
or ( n12606 , n12604 , n12605 );
nand ( n12607 , n12606 , n8223 );
nand ( n12608 , n12603 , n12607 );
xor ( n12609 , n12599 , n12608 );
not ( n12610 , n1875 );
not ( n12611 , n550 );
not ( n12612 , n5937 );
or ( n12613 , n12611 , n12612 );
nand ( n12614 , n353618 , n1880 );
nand ( n12615 , n12613 , n12614 );
not ( n12616 , n12615 );
or ( n12617 , n12610 , n12616 );
nand ( n12618 , n12307 , n4078 );
nand ( n12619 , n12617 , n12618 );
xor ( n12620 , n12609 , n12619 );
xor ( n12621 , n12589 , n12620 );
xor ( n12622 , n12576 , n12621 );
xor ( n12623 , n12312 , n12316 );
and ( n12624 , n12623 , n12349 );
and ( n12625 , n12312 , n12316 );
or ( n12626 , n12624 , n12625 );
xor ( n12627 , n12622 , n12626 );
xor ( n12628 , n12572 , n12627 );
xor ( n12629 , n12369 , n12373 );
and ( n12630 , n12629 , n12378 );
and ( n12631 , n12369 , n12373 );
or ( n12632 , n12630 , n12631 );
xor ( n12633 , n12628 , n12632 );
xor ( n12634 , n12350 , n12379 );
and ( n12635 , n12634 , n12384 );
and ( n12636 , n12350 , n12379 );
or ( n12637 , n12635 , n12636 );
nor ( n12638 , n12633 , n12637 );
buf ( n12639 , n12638 );
not ( n12640 , n12639 );
nand ( n12641 , n12633 , n12637 );
nand ( n12642 , n12640 , n12641 );
not ( n12643 , n12642 );
and ( n12644 , n12530 , n12643 );
not ( n12645 , n12530 );
and ( n12646 , n12645 , n12642 );
nor ( n12647 , n12644 , n12646 );
xor ( n12648 , n359546 , n359586 );
and ( n12649 , n12648 , n359626 );
and ( n12650 , n359546 , n359586 );
or ( n12651 , n12649 , n12650 );
buf ( n360328 , n12651 );
buf ( n360329 , n360328 );
xor ( n12654 , n359642 , n359699 );
and ( n12655 , n12654 , n359706 );
and ( n12656 , n359642 , n359699 );
or ( n12657 , n12655 , n12656 );
buf ( n360334 , n12657 );
buf ( n360335 , n360334 );
xor ( n12660 , n360329 , n360335 );
xor ( n12661 , n359648 , n359654 );
and ( n12662 , n12661 , n359696 );
and ( n12663 , n359648 , n359654 );
or ( n12664 , n12662 , n12663 );
buf ( n360341 , n12664 );
buf ( n360342 , n360341 );
buf ( n360343 , n359665 );
not ( n12668 , n360343 );
buf ( n360345 , n347344 );
not ( n12670 , n360345 );
or ( n12671 , n12668 , n12670 );
buf ( n360348 , n570 );
buf ( n360349 , n347350 );
nand ( n12674 , n360348 , n360349 );
buf ( n360351 , n12674 );
buf ( n360352 , n360351 );
nand ( n12677 , n12671 , n360352 );
buf ( n360354 , n12677 );
buf ( n360355 , n360354 );
not ( n12680 , n360355 );
buf ( n360357 , n12680 );
buf ( n360358 , n360357 );
xor ( n12683 , n359551 , n359568 );
and ( n12684 , n12683 , n359583 );
and ( n12685 , n359551 , n359568 );
or ( n12686 , n12684 , n12685 );
buf ( n360363 , n12686 );
buf ( n360364 , n360363 );
xor ( n12689 , n360358 , n360364 );
xor ( n12690 , n359672 , n359675 );
and ( n12691 , n12690 , n359693 );
and ( n12692 , n359672 , n359675 );
or ( n12693 , n12691 , n12692 );
buf ( n360370 , n12693 );
buf ( n360371 , n360370 );
xor ( n12696 , n12689 , n360371 );
buf ( n360373 , n12696 );
buf ( n360374 , n360373 );
xor ( n12699 , n360342 , n360374 );
buf ( n360376 , n11943 );
not ( n12701 , n360376 );
buf ( n360378 , n11924 );
not ( n12703 , n360378 );
or ( n12704 , n12701 , n12703 );
buf ( n360381 , n356903 );
nand ( n12706 , n12704 , n360381 );
buf ( n360383 , n12706 );
buf ( n360384 , n360383 );
buf ( n360385 , n11923 );
buf ( n360386 , n359616 );
nand ( n12711 , n360385 , n360386 );
buf ( n360388 , n12711 );
buf ( n360389 , n360388 );
nand ( n12714 , n360384 , n360389 );
buf ( n360391 , n12714 );
buf ( n360392 , n360391 );
buf ( n360393 , n555 );
buf ( n360394 , n560 );
and ( n12719 , n360393 , n360394 );
buf ( n360396 , n12719 );
buf ( n360397 , n360396 );
buf ( n360398 , n359610 );
not ( n12723 , n360398 );
buf ( n360400 , n9186 );
not ( n12725 , n360400 );
or ( n12726 , n12723 , n12725 );
buf ( n360403 , n5407 );
buf ( n360404 , n553 );
buf ( n360405 , n560 );
xor ( n12730 , n360404 , n360405 );
buf ( n360407 , n12730 );
buf ( n360408 , n360407 );
nand ( n12733 , n360403 , n360408 );
buf ( n360410 , n12733 );
buf ( n360411 , n360410 );
nand ( n12736 , n12726 , n360411 );
buf ( n360413 , n12736 );
buf ( n360414 , n360413 );
xor ( n12739 , n360397 , n360414 );
buf ( n360416 , n359686 );
not ( n12741 , n360416 );
buf ( n360418 , n350874 );
buf ( n12743 , n360418 );
buf ( n360420 , n12743 );
buf ( n360421 , n360420 );
not ( n12746 , n360421 );
or ( n12747 , n12741 , n12746 );
buf ( n360424 , n2550 );
buf ( n360425 , n547 );
buf ( n360426 , n566 );
xor ( n12751 , n360425 , n360426 );
buf ( n360428 , n12751 );
buf ( n360429 , n360428 );
nand ( n12754 , n360424 , n360429 );
buf ( n360431 , n12754 );
buf ( n360432 , n360431 );
nand ( n12757 , n12747 , n360432 );
buf ( n360434 , n12757 );
buf ( n360435 , n360434 );
xor ( n12760 , n12739 , n360435 );
buf ( n360437 , n12760 );
buf ( n360438 , n360437 );
xor ( n12763 , n360392 , n360438 );
buf ( n360440 , n359561 );
not ( n12765 , n360440 );
buf ( n360442 , n351330 );
not ( n12767 , n360442 );
or ( n12768 , n12765 , n12767 );
buf ( n360445 , n3650 );
buf ( n360446 , n549 );
buf ( n360447 , n564 );
xor ( n12772 , n360446 , n360447 );
buf ( n360449 , n12772 );
buf ( n360450 , n360449 );
nand ( n12775 , n360445 , n360450 );
buf ( n360452 , n12775 );
buf ( n360453 , n360452 );
nand ( n12778 , n12768 , n360453 );
buf ( n360455 , n12778 );
buf ( n360456 , n360455 );
buf ( n360457 , n359595 );
not ( n12782 , n360457 );
buf ( n360459 , n8604 );
not ( n12784 , n360459 );
or ( n12785 , n12782 , n12784 );
buf ( n360462 , n352295 );
buf ( n360463 , n551 );
buf ( n360464 , n562 );
xor ( n12789 , n360463 , n360464 );
buf ( n360466 , n12789 );
buf ( n360467 , n360466 );
nand ( n12792 , n360462 , n360467 );
buf ( n360469 , n12792 );
buf ( n360470 , n360469 );
nand ( n12795 , n12785 , n360470 );
buf ( n360472 , n12795 );
buf ( n360473 , n360472 );
xor ( n12798 , n360456 , n360473 );
buf ( n360475 , n11900 );
not ( n12800 , n360475 );
buf ( n360477 , n2236 );
not ( n12802 , n360477 );
or ( n12803 , n12800 , n12802 );
buf ( n360480 , n349933 );
buf ( n360481 , n545 );
buf ( n360482 , n568 );
xor ( n12807 , n360481 , n360482 );
buf ( n360484 , n12807 );
buf ( n360485 , n360484 );
nand ( n12810 , n360480 , n360485 );
buf ( n360487 , n12810 );
buf ( n360488 , n360487 );
nand ( n12813 , n12803 , n360488 );
buf ( n360490 , n12813 );
buf ( n360491 , n360490 );
xor ( n12816 , n12798 , n360491 );
buf ( n360493 , n12816 );
buf ( n360494 , n360493 );
xor ( n12819 , n12763 , n360494 );
buf ( n360496 , n12819 );
buf ( n360497 , n360496 );
xor ( n12822 , n12699 , n360497 );
buf ( n360499 , n12822 );
buf ( n360500 , n360499 );
xor ( n12825 , n12660 , n360500 );
buf ( n360502 , n12825 );
buf ( n360503 , n360502 );
xor ( n12828 , n359725 , n359731 );
and ( n12829 , n12828 , n359910 );
and ( n12830 , n359725 , n359731 );
or ( n12831 , n12829 , n12830 );
buf ( n360508 , n12831 );
buf ( n360509 , n360508 );
xor ( n12834 , n360503 , n360509 );
xor ( n12835 , n359629 , n359635 );
and ( n12836 , n12835 , n359709 );
and ( n12837 , n359629 , n359635 );
or ( n12838 , n12836 , n12837 );
buf ( n360515 , n12838 );
buf ( n360516 , n360515 );
xor ( n12841 , n359815 , n359821 );
and ( n12842 , n12841 , n359907 );
and ( n12843 , n359815 , n359821 );
or ( n12844 , n12842 , n12843 );
buf ( n360521 , n12844 );
buf ( n360522 , n360521 );
xor ( n12847 , n360516 , n360522 );
xor ( n12848 , n359738 , n359773 );
and ( n12849 , n12848 , n359812 );
and ( n12850 , n359738 , n359773 );
or ( n12851 , n12849 , n12850 );
buf ( n360528 , n12851 );
buf ( n360529 , n360528 );
buf ( n360530 , n359876 );
not ( n12855 , n360530 );
buf ( n360532 , n347671 );
not ( n12857 , n360532 );
or ( n12858 , n12855 , n12857 );
buf ( n360535 , n347530 );
buf ( n360536 , n586 );
nand ( n12861 , n360535 , n360536 );
buf ( n360538 , n12861 );
buf ( n360539 , n360538 );
nand ( n12864 , n12858 , n360539 );
buf ( n360541 , n12864 );
buf ( n360542 , n360541 );
not ( n12867 , n360542 );
buf ( n360544 , n12867 );
buf ( n360545 , n360544 );
xor ( n12870 , n359743 , n359755 );
and ( n12871 , n12870 , n359770 );
and ( n12872 , n359743 , n359755 );
or ( n12873 , n12871 , n12872 );
buf ( n360550 , n12873 );
buf ( n360551 , n360550 );
xor ( n12876 , n360545 , n360551 );
buf ( n360553 , n359892 );
buf ( n360554 , n359882 );
or ( n12879 , n360553 , n360554 );
buf ( n360556 , n359866 );
nand ( n12881 , n12879 , n360556 );
buf ( n360558 , n12881 );
buf ( n360559 , n360558 );
buf ( n360560 , n359892 );
buf ( n360561 , n359882 );
nand ( n12886 , n360560 , n360561 );
buf ( n360563 , n12886 );
buf ( n360564 , n360563 );
nand ( n12889 , n360559 , n360564 );
buf ( n360566 , n12889 );
buf ( n360567 , n360566 );
xor ( n12892 , n12876 , n360567 );
buf ( n360569 , n12892 );
buf ( n360570 , n360569 );
xor ( n12895 , n359843 , n359849 );
and ( n12896 , n12895 , n359894 );
and ( n12897 , n359843 , n359849 );
or ( n12898 , n12896 , n12897 );
buf ( n360575 , n12898 );
buf ( n360576 , n360575 );
xor ( n12901 , n360570 , n360576 );
buf ( n360578 , n359804 );
not ( n12903 , n360578 );
buf ( n360580 , n357148 );
not ( n12905 , n360580 );
or ( n12906 , n12903 , n12905 );
buf ( n360583 , n357148 );
buf ( n360584 , n359804 );
or ( n12909 , n360583 , n360584 );
buf ( n360586 , n359790 );
nand ( n12911 , n12909 , n360586 );
buf ( n360588 , n12911 );
buf ( n360589 , n360588 );
nand ( n12914 , n12906 , n360589 );
buf ( n360591 , n12914 );
buf ( n360592 , n360591 );
nand ( n12917 , n555 , n576 );
not ( n12918 , n356440 );
not ( n12919 , n359784 );
or ( n12920 , n12918 , n12919 );
buf ( n360597 , n353193 );
buf ( n360598 , n553 );
buf ( n360599 , n576 );
xor ( n12924 , n360598 , n360599 );
buf ( n360601 , n12924 );
buf ( n360602 , n360601 );
nand ( n12927 , n360597 , n360602 );
buf ( n360604 , n12927 );
nand ( n12929 , n12920 , n360604 );
xor ( n12930 , n12917 , n12929 );
not ( n12931 , n359860 );
not ( n12932 , n350699 );
or ( n12933 , n12931 , n12932 );
buf ( n360610 , n350705 );
buf ( n360611 , n547 );
buf ( n360612 , n582 );
xor ( n12937 , n360611 , n360612 );
buf ( n360614 , n12937 );
buf ( n360615 , n360614 );
nand ( n12940 , n360610 , n360615 );
buf ( n360617 , n12940 );
nand ( n12942 , n12933 , n360617 );
xnor ( n12943 , n12930 , n12942 );
buf ( n360620 , n12943 );
xor ( n12945 , n360592 , n360620 );
not ( n12946 , n12122 );
not ( n12947 , n355543 );
or ( n12948 , n12946 , n12947 );
buf ( n360625 , n352491 );
buf ( n360626 , n551 );
buf ( n360627 , n578 );
xor ( n12952 , n360626 , n360627 );
buf ( n360629 , n12952 );
buf ( n360630 , n360629 );
nand ( n12955 , n360625 , n360630 );
buf ( n360632 , n12955 );
nand ( n12957 , n12948 , n360632 );
buf ( n360634 , n12087 );
not ( n12959 , n360634 );
buf ( n360636 , n5570 );
not ( n12961 , n360636 );
or ( n12962 , n12959 , n12961 );
buf ( n360639 , n348617 );
xor ( n12964 , n584 , n545 );
buf ( n360641 , n12964 );
nand ( n12966 , n360639 , n360641 );
buf ( n360643 , n12966 );
buf ( n360644 , n360643 );
nand ( n12969 , n12962 , n360644 );
buf ( n360646 , n12969 );
xor ( n12971 , n12957 , n360646 );
buf ( n360648 , n549 );
buf ( n360649 , n580 );
xor ( n12974 , n360648 , n360649 );
buf ( n360651 , n12974 );
not ( n12976 , n360651 );
not ( n12977 , n351559 );
or ( n12978 , n12976 , n12977 );
nand ( n12979 , n12076 , n3870 );
nand ( n12980 , n12978 , n12979 );
xor ( n12981 , n12971 , n12980 );
buf ( n360658 , n12981 );
xor ( n12983 , n12945 , n360658 );
buf ( n360660 , n12983 );
buf ( n360661 , n360660 );
xor ( n12986 , n12901 , n360661 );
buf ( n360663 , n12986 );
buf ( n360664 , n360663 );
xor ( n12989 , n360529 , n360664 );
xor ( n12990 , n359828 , n359897 );
and ( n12991 , n12990 , n359904 );
and ( n12992 , n359828 , n359897 );
or ( n12993 , n12991 , n12992 );
buf ( n360670 , n12993 );
buf ( n360671 , n360670 );
xor ( n12996 , n12989 , n360671 );
buf ( n360673 , n12996 );
buf ( n360674 , n360673 );
xor ( n12999 , n12847 , n360674 );
buf ( n360676 , n12999 );
buf ( n360677 , n360676 );
xor ( n13002 , n12834 , n360677 );
buf ( n360679 , n13002 );
buf ( n360680 , n360679 );
not ( n13005 , n360680 );
buf ( n360682 , n13005 );
buf ( n360683 , n360682 );
xor ( n13008 , n359712 , n359718 );
and ( n13009 , n13008 , n359913 );
and ( n13010 , n359712 , n359718 );
or ( n13011 , n13009 , n13010 );
buf ( n360688 , n13011 );
buf ( n360689 , n360688 );
not ( n13014 , n360689 );
buf ( n360691 , n13014 );
buf ( n360692 , n360691 );
nand ( n13017 , n360683 , n360692 );
buf ( n360694 , n13017 );
buf ( n360695 , n360694 );
buf ( n13020 , n360695 );
buf ( n360697 , n13020 );
not ( n13022 , n360691 );
nand ( n13023 , n13022 , n360679 );
and ( n13024 , n360697 , n13023 );
not ( n13025 , n12245 );
not ( n13026 , n8973 );
nand ( n13027 , n13025 , n13026 , n9588 , n8053 );
buf ( n360704 , n13027 );
not ( n13029 , n360704 );
buf ( n360706 , n13029 );
not ( n13031 , n360706 );
not ( n13032 , n355795 );
or ( n13033 , n13031 , n13032 );
not ( n13034 , n357270 );
not ( n13035 , n357275 );
and ( n13036 , n13034 , n13035 );
nor ( n13037 , n13036 , n12245 );
not ( n13038 , n13037 );
not ( n13039 , n9139 );
or ( n13040 , n13038 , n13039 );
buf ( n360717 , n12245 );
not ( n13042 , n360717 );
buf ( n360719 , n357280 );
not ( n13044 , n360719 );
and ( n13045 , n13042 , n13044 );
buf ( n360722 , n359926 );
nor ( n13047 , n13045 , n360722 );
buf ( n360724 , n13047 );
nand ( n13049 , n13040 , n360724 );
buf ( n360726 , n13049 );
not ( n13051 , n360726 );
buf ( n360728 , n13051 );
nand ( n13053 , n13033 , n360728 );
and ( n13054 , n13024 , n13053 );
not ( n13055 , n13024 );
not ( n13056 , n360728 );
nor ( n13057 , n355792 , n13027 );
nor ( n13058 , n13056 , n13057 );
and ( n13059 , n13055 , n13058 );
nor ( n13060 , n13054 , n13059 );
not ( n13061 , n13060 );
nor ( n13062 , n12647 , n13061 );
not ( n13063 , n13062 );
not ( n13064 , n13060 );
nand ( n13065 , n13064 , n12647 );
buf ( n13066 , n13065 );
and ( n13067 , n13063 , n13066 );
and ( n13068 , n12519 , n13067 );
not ( n13069 , n12519 );
not ( n13070 , n13067 );
and ( n13071 , n13069 , n13070 );
nor ( n13072 , n13068 , n13071 );
nand ( n13073 , n13072 , n9625 , n12407 );
nand ( n13074 , n8990 , n8303 );
nor ( n13075 , n13073 , n13074 );
not ( n13076 , n12640 );
not ( n13077 , n12529 );
or ( n13078 , n13076 , n13077 );
buf ( n13079 , n12641 );
nand ( n13080 , n13078 , n13079 );
not ( n13081 , n8215 );
not ( n13082 , n544 );
not ( n13083 , n3996 );
or ( n13084 , n13082 , n13083 );
nand ( n13085 , n1788 , n7283 );
nand ( n13086 , n13084 , n13085 );
not ( n13087 , n13086 );
or ( n13088 , n13081 , n13087 );
nand ( n13089 , n12601 , n8223 );
nand ( n13090 , n13088 , n13089 );
buf ( n13091 , n348266 );
and ( n13092 , n13091 , n544 );
xor ( n13093 , n13090 , n13092 );
not ( n13094 , n4109 );
and ( n13095 , n552 , n7247 );
not ( n13096 , n552 );
and ( n13097 , n13096 , n9017 );
or ( n13098 , n13095 , n13097 );
not ( n13099 , n13098 );
or ( n13100 , n13094 , n13099 );
nand ( n13101 , n12568 , n1871 );
nand ( n13102 , n13100 , n13101 );
xor ( n13103 , n13093 , n13102 );
xor ( n13104 , n12550 , n12560 );
and ( n13105 , n13104 , n12570 );
and ( n13106 , n12550 , n12560 );
or ( n13107 , n13105 , n13106 );
xor ( n13108 , n13103 , n13107 );
not ( n13109 , n2019 );
not ( n13110 , n548 );
not ( n13111 , n4057 );
or ( n13112 , n13110 , n13111 );
nand ( n13113 , n351734 , n4031 );
not ( n13114 , n13113 );
not ( n13115 , n351739 );
or ( n13116 , n13114 , n13115 );
nand ( n13117 , n13116 , n351773 );
nand ( n13118 , n13112 , n13117 );
not ( n13119 , n13118 );
or ( n13120 , n13109 , n13119 );
nand ( n13121 , n12557 , n5751 );
nand ( n13122 , n13120 , n13121 );
not ( n13123 , n5757 );
not ( n13124 , n546 );
not ( n13125 , n4011 );
or ( n13126 , n13124 , n13125 );
nand ( n13127 , n1974 , n5761 );
nand ( n13128 , n13126 , n13127 );
not ( n13129 , n13128 );
or ( n13130 , n13123 , n13129 );
nand ( n13131 , n12595 , n8381 );
nand ( n13132 , n13130 , n13131 );
xor ( n13133 , n13122 , n13132 );
not ( n13134 , n1875 );
not ( n13135 , n550 );
not ( n13136 , n6035 );
or ( n13137 , n13135 , n13136 );
nand ( n13138 , n6034 , n1880 );
nand ( n13139 , n13137 , n13138 );
not ( n13140 , n13139 );
or ( n13141 , n13134 , n13140 );
nand ( n13142 , n12615 , n4078 );
nand ( n13143 , n13141 , n13142 );
xor ( n13144 , n13133 , n13143 );
xor ( n13145 , n13108 , n13144 );
xor ( n13146 , n12580 , n12588 );
and ( n13147 , n13146 , n12620 );
and ( n13148 , n12580 , n12588 );
or ( n13149 , n13147 , n13148 );
buf ( n13150 , n12548 );
and ( n13151 , n13150 , n5718 );
nor ( n13152 , n8424 , n348175 );
nor ( n13153 , n13151 , n13152 );
xor ( n13154 , n12584 , n12585 );
and ( n13155 , n13154 , n12587 );
and ( n13156 , n12584 , n12585 );
or ( n13157 , n13155 , n13156 );
xor ( n13158 , n13153 , n13157 );
xor ( n13159 , n12599 , n12608 );
and ( n13160 , n13159 , n12619 );
and ( n13161 , n12599 , n12608 );
or ( n13162 , n13160 , n13161 );
xor ( n13163 , n13158 , n13162 );
xor ( n13164 , n13149 , n13163 );
xor ( n13165 , n12534 , n12538 );
and ( n13166 , n13165 , n12571 );
and ( n13167 , n12534 , n12538 );
or ( n13168 , n13166 , n13167 );
xor ( n13169 , n13164 , n13168 );
xor ( n13170 , n13145 , n13169 );
xor ( n13171 , n12576 , n12621 );
and ( n13172 , n13171 , n12626 );
and ( n13173 , n12576 , n12621 );
or ( n13174 , n13172 , n13173 );
xor ( n13175 , n13170 , n13174 );
xor ( n13176 , n12572 , n12627 );
and ( n13177 , n13176 , n12632 );
and ( n13178 , n12572 , n12627 );
or ( n13179 , n13177 , n13178 );
nand ( n13180 , n13175 , n13179 );
not ( n13181 , n13175 );
not ( n13182 , n13179 );
nand ( n13183 , n13181 , n13182 );
nand ( n13184 , n13180 , n13183 );
not ( n13185 , n13184 );
and ( n13186 , n13080 , n13185 );
not ( n13187 , n13080 );
and ( n13188 , n13187 , n13184 );
nor ( n13189 , n13186 , n13188 );
buf ( n360866 , n355795 );
not ( n13191 , n360866 );
buf ( n360868 , n360697 );
not ( n13193 , n360868 );
buf ( n360870 , n13027 );
nor ( n13195 , n13193 , n360870 );
buf ( n360872 , n13195 );
buf ( n360873 , n360872 );
not ( n13198 , n360873 );
or ( n13199 , n13191 , n13198 );
not ( n13200 , n360697 );
not ( n13201 , n13049 );
or ( n13202 , n13200 , n13201 );
nand ( n13203 , n13202 , n13023 );
buf ( n360880 , n13203 );
not ( n13205 , n360880 );
buf ( n360882 , n13205 );
buf ( n360883 , n360882 );
nand ( n13208 , n13199 , n360883 );
buf ( n360885 , n13208 );
xor ( n13210 , n360397 , n360414 );
and ( n13211 , n13210 , n360435 );
and ( n13212 , n360397 , n360414 );
or ( n13213 , n13211 , n13212 );
buf ( n360890 , n13213 );
buf ( n360891 , n360890 );
buf ( n360892 , n360484 );
not ( n13217 , n360892 );
buf ( n360894 , n2236 );
not ( n13219 , n360894 );
or ( n13220 , n13217 , n13219 );
buf ( n360897 , n349933 );
buf ( n360898 , n544 );
buf ( n360899 , n568 );
xor ( n13224 , n360898 , n360899 );
buf ( n360901 , n13224 );
buf ( n360902 , n360901 );
nand ( n13227 , n360897 , n360902 );
buf ( n360904 , n13227 );
buf ( n360905 , n360904 );
nand ( n13230 , n13220 , n360905 );
buf ( n360907 , n13230 );
buf ( n360908 , n360907 );
buf ( n360909 , n360449 );
not ( n13234 , n360909 );
buf ( n360911 , n351330 );
buf ( n13236 , n360911 );
buf ( n360913 , n13236 );
buf ( n360914 , n360913 );
not ( n13239 , n360914 );
or ( n13240 , n13234 , n13239 );
buf ( n360917 , n3650 );
buf ( n360918 , n548 );
buf ( n360919 , n564 );
xor ( n13244 , n360918 , n360919 );
buf ( n360921 , n13244 );
buf ( n360922 , n360921 );
nand ( n13247 , n360917 , n360922 );
buf ( n360924 , n13247 );
buf ( n360925 , n360924 );
nand ( n13250 , n13240 , n360925 );
buf ( n360927 , n13250 );
buf ( n360928 , n360927 );
xor ( n13253 , n360908 , n360928 );
buf ( n360930 , n347350 );
buf ( n360931 , n347344 );
or ( n13256 , n360930 , n360931 );
buf ( n360933 , n570 );
nand ( n13258 , n13256 , n360933 );
buf ( n360935 , n13258 );
buf ( n360936 , n360935 );
xor ( n13261 , n13253 , n360936 );
buf ( n360938 , n13261 );
buf ( n360939 , n360938 );
xor ( n13264 , n360891 , n360939 );
buf ( n360941 , n360407 );
not ( n13266 , n360941 );
buf ( n360943 , n9186 );
not ( n13268 , n360943 );
or ( n13269 , n13266 , n13268 );
buf ( n360946 , n5407 );
buf ( n360947 , n552 );
buf ( n360948 , n560 );
xor ( n13273 , n360947 , n360948 );
buf ( n360950 , n13273 );
buf ( n360951 , n360950 );
nand ( n13276 , n360946 , n360951 );
buf ( n360953 , n13276 );
buf ( n360954 , n360953 );
nand ( n13279 , n13269 , n360954 );
buf ( n360956 , n13279 );
buf ( n360957 , n360956 );
buf ( n360958 , n360466 );
not ( n13283 , n360958 );
buf ( n360960 , n8604 );
not ( n13285 , n360960 );
or ( n13286 , n13283 , n13285 );
buf ( n360963 , n352295 );
buf ( n360964 , n550 );
buf ( n360965 , n562 );
xor ( n13290 , n360964 , n360965 );
buf ( n360967 , n13290 );
buf ( n360968 , n360967 );
nand ( n13293 , n360963 , n360968 );
buf ( n360970 , n13293 );
buf ( n360971 , n360970 );
nand ( n13296 , n13286 , n360971 );
buf ( n360973 , n13296 );
buf ( n360974 , n360973 );
xor ( n13299 , n360957 , n360974 );
buf ( n360976 , n360428 );
not ( n13301 , n360976 );
buf ( n360978 , n360420 );
not ( n13303 , n360978 );
or ( n13304 , n13301 , n13303 );
buf ( n360981 , n2550 );
buf ( n360982 , n546 );
buf ( n360983 , n566 );
xor ( n13308 , n360982 , n360983 );
buf ( n360985 , n13308 );
buf ( n360986 , n360985 );
nand ( n13311 , n360981 , n360986 );
buf ( n360988 , n13311 );
buf ( n360989 , n360988 );
nand ( n13314 , n13304 , n360989 );
buf ( n360991 , n13314 );
buf ( n360992 , n360991 );
xor ( n13317 , n13299 , n360992 );
buf ( n360994 , n13317 );
buf ( n360995 , n360994 );
xor ( n13320 , n13264 , n360995 );
buf ( n360997 , n13320 );
buf ( n360998 , n360997 );
xor ( n13323 , n360342 , n360374 );
and ( n13324 , n13323 , n360497 );
and ( n13325 , n360342 , n360374 );
or ( n13326 , n13324 , n13325 );
buf ( n361003 , n13326 );
buf ( n361004 , n361003 );
xor ( n13329 , n360998 , n361004 );
buf ( n361006 , n554 );
buf ( n361007 , n560 );
and ( n13332 , n361006 , n361007 );
buf ( n361009 , n13332 );
buf ( n361010 , n361009 );
buf ( n361011 , n360354 );
xor ( n13336 , n361010 , n361011 );
xor ( n13337 , n360456 , n360473 );
and ( n13338 , n13337 , n360491 );
and ( n13339 , n360456 , n360473 );
or ( n13340 , n13338 , n13339 );
buf ( n361017 , n13340 );
buf ( n361018 , n361017 );
xor ( n13343 , n13336 , n361018 );
buf ( n361020 , n13343 );
buf ( n361021 , n361020 );
xor ( n13346 , n360358 , n360364 );
and ( n13347 , n13346 , n360371 );
and ( n13348 , n360358 , n360364 );
or ( n13349 , n13347 , n13348 );
buf ( n361026 , n13349 );
buf ( n361027 , n361026 );
xor ( n13352 , n361021 , n361027 );
xor ( n13353 , n360392 , n360438 );
and ( n13354 , n13353 , n360494 );
and ( n13355 , n360392 , n360438 );
or ( n13356 , n13354 , n13355 );
buf ( n361033 , n13356 );
buf ( n361034 , n361033 );
xor ( n13359 , n13352 , n361034 );
buf ( n361036 , n13359 );
buf ( n361037 , n361036 );
xor ( n13362 , n13329 , n361037 );
buf ( n361039 , n13362 );
not ( n13364 , n12917 );
not ( n13365 , n12929 );
not ( n13366 , n13365 );
or ( n13367 , n13364 , n13366 );
nand ( n13368 , n13367 , n12942 );
not ( n13369 , n12917 );
nand ( n13370 , n13369 , n12929 );
nand ( n13371 , n13368 , n13370 );
buf ( n361048 , n13371 );
buf ( n361049 , n347530 );
buf ( n361050 , n350110 );
or ( n13375 , n361049 , n361050 );
buf ( n361052 , n586 );
nand ( n13377 , n13375 , n361052 );
buf ( n361054 , n13377 );
buf ( n361055 , n361054 );
buf ( n361056 , n12964 );
not ( n13381 , n361056 );
buf ( n361058 , n5570 );
not ( n13383 , n361058 );
or ( n13384 , n13381 , n13383 );
xor ( n13385 , n584 , n544 );
nand ( n13386 , n348617 , n13385 );
buf ( n361063 , n13386 );
nand ( n13388 , n13384 , n361063 );
buf ( n361065 , n13388 );
buf ( n361066 , n361065 );
xor ( n13391 , n361055 , n361066 );
buf ( n361068 , n360651 );
not ( n13393 , n361068 );
buf ( n361070 , n3870 );
not ( n13395 , n361070 );
or ( n13396 , n13393 , n13395 );
buf ( n361073 , n351559 );
buf ( n361074 , n548 );
buf ( n361075 , n580 );
xor ( n13400 , n361074 , n361075 );
buf ( n361077 , n13400 );
buf ( n361078 , n361077 );
nand ( n13403 , n361073 , n361078 );
buf ( n361080 , n13403 );
buf ( n361081 , n361080 );
nand ( n13406 , n13396 , n361081 );
buf ( n361083 , n13406 );
buf ( n361084 , n361083 );
xor ( n13409 , n13391 , n361084 );
buf ( n361086 , n13409 );
buf ( n361087 , n361086 );
xor ( n13412 , n361048 , n361087 );
buf ( n361089 , n360614 );
not ( n13414 , n361089 );
buf ( n361091 , n350699 );
not ( n13416 , n361091 );
or ( n13417 , n13414 , n13416 );
buf ( n361094 , n350705 );
buf ( n361095 , n546 );
buf ( n361096 , n582 );
xor ( n13421 , n361095 , n361096 );
buf ( n361098 , n13421 );
buf ( n361099 , n361098 );
nand ( n13424 , n361094 , n361099 );
buf ( n361101 , n13424 );
buf ( n361102 , n361101 );
nand ( n13427 , n13417 , n361102 );
buf ( n361104 , n13427 );
buf ( n361105 , n361104 );
buf ( n361106 , n360601 );
not ( n13431 , n361106 );
buf ( n361108 , n356440 );
buf ( n13433 , n361108 );
buf ( n361110 , n13433 );
buf ( n361111 , n361110 );
not ( n13436 , n361111 );
or ( n13437 , n13431 , n13436 );
buf ( n361114 , n356446 );
buf ( n361115 , n552 );
buf ( n361116 , n576 );
xor ( n13441 , n361115 , n361116 );
buf ( n361118 , n13441 );
buf ( n361119 , n361118 );
nand ( n13444 , n361114 , n361119 );
buf ( n361121 , n13444 );
buf ( n361122 , n361121 );
nand ( n13447 , n13437 , n361122 );
buf ( n361124 , n13447 );
buf ( n361125 , n361124 );
xor ( n13450 , n361105 , n361125 );
buf ( n361127 , n360629 );
not ( n13452 , n361127 );
buf ( n361129 , n5162 );
buf ( n13454 , n361129 );
buf ( n361131 , n13454 );
buf ( n361132 , n361131 );
not ( n13457 , n361132 );
or ( n13458 , n13452 , n13457 );
buf ( n361135 , n354788 );
buf ( n361136 , n550 );
buf ( n361137 , n578 );
xor ( n13462 , n361136 , n361137 );
buf ( n361139 , n13462 );
buf ( n361140 , n361139 );
nand ( n13465 , n361135 , n361140 );
buf ( n361142 , n13465 );
buf ( n361143 , n361142 );
nand ( n13468 , n13458 , n361143 );
buf ( n361145 , n13468 );
buf ( n361146 , n361145 );
xor ( n13471 , n13450 , n361146 );
buf ( n361148 , n13471 );
buf ( n361149 , n361148 );
xor ( n13474 , n13412 , n361149 );
buf ( n361151 , n13474 );
buf ( n361152 , n361151 );
buf ( n361153 , n554 );
buf ( n361154 , n576 );
nand ( n13479 , n361153 , n361154 );
buf ( n361156 , n13479 );
xor ( n13481 , n360541 , n361156 );
not ( n13482 , n12957 );
not ( n13483 , n360646 );
or ( n13484 , n13482 , n13483 );
or ( n13485 , n12957 , n360646 );
nand ( n13486 , n13485 , n12980 );
nand ( n13487 , n13484 , n13486 );
xnor ( n13488 , n13481 , n13487 );
buf ( n361165 , n13488 );
xor ( n13490 , n360545 , n360551 );
and ( n13491 , n13490 , n360567 );
and ( n13492 , n360545 , n360551 );
or ( n13493 , n13491 , n13492 );
buf ( n361170 , n13493 );
buf ( n361171 , n361170 );
xor ( n13496 , n361165 , n361171 );
xor ( n13497 , n360592 , n360620 );
and ( n13498 , n13497 , n360658 );
and ( n13499 , n360592 , n360620 );
or ( n13500 , n13498 , n13499 );
buf ( n361177 , n13500 );
buf ( n361178 , n361177 );
xor ( n13503 , n13496 , n361178 );
buf ( n361180 , n13503 );
buf ( n361181 , n361180 );
xor ( n13506 , n361152 , n361181 );
xor ( n13507 , n360570 , n360576 );
and ( n13508 , n13507 , n360661 );
and ( n13509 , n360570 , n360576 );
or ( n13510 , n13508 , n13509 );
buf ( n361187 , n13510 );
buf ( n361188 , n361187 );
xor ( n13513 , n13506 , n361188 );
buf ( n361190 , n13513 );
xor ( n13515 , n360329 , n360335 );
and ( n13516 , n13515 , n360500 );
and ( n13517 , n360329 , n360335 );
or ( n13518 , n13516 , n13517 );
buf ( n361195 , n13518 );
xor ( n13520 , n361190 , n361195 );
xor ( n13521 , n360529 , n360664 );
and ( n13522 , n13521 , n360671 );
and ( n13523 , n360529 , n360664 );
or ( n13524 , n13522 , n13523 );
buf ( n361201 , n13524 );
xor ( n13526 , n13520 , n361201 );
xor ( n13527 , n361039 , n13526 );
xor ( n13528 , n360516 , n360522 );
and ( n13529 , n13528 , n360674 );
and ( n13530 , n360516 , n360522 );
or ( n13531 , n13529 , n13530 );
buf ( n361208 , n13531 );
xor ( n13533 , n13527 , n361208 );
buf ( n361210 , n13533 );
not ( n13535 , n361210 );
buf ( n361212 , n13535 );
buf ( n361213 , n361212 );
xor ( n13538 , n360503 , n360509 );
and ( n13539 , n13538 , n360677 );
and ( n13540 , n360503 , n360509 );
or ( n13541 , n13539 , n13540 );
buf ( n361218 , n13541 );
buf ( n361219 , n361218 );
not ( n13544 , n361219 );
buf ( n361221 , n13544 );
buf ( n361222 , n361221 );
nand ( n13547 , n361213 , n361222 );
buf ( n361224 , n13547 );
buf ( n361225 , n361224 );
buf ( n13550 , n361225 );
buf ( n361227 , n13550 );
not ( n13552 , n361212 );
nand ( n13553 , n13552 , n361218 );
buf ( n361230 , n13553 );
buf ( n13555 , n361230 );
buf ( n361232 , n13555 );
nand ( n13557 , n361227 , n361232 );
and ( n13558 , n360885 , n13557 );
not ( n13559 , n360885 );
and ( n13560 , n361227 , n361232 );
and ( n13561 , n13559 , n13560 );
nor ( n13562 , n13558 , n13561 );
nand ( n13563 , n13189 , n13562 );
nand ( n13564 , n13563 , n13065 );
not ( n13565 , n13564 );
not ( n13566 , n13565 );
not ( n13567 , n13566 );
buf ( n361244 , n355789 );
not ( n13569 , n361244 );
buf ( n361246 , n13569 );
nand ( n13571 , n361246 , n360706 );
buf ( n361248 , n361224 );
buf ( n361249 , n360694 );
and ( n13574 , n361248 , n361249 );
buf ( n361251 , n13574 );
buf ( n361252 , n361251 );
buf ( n13577 , n361252 );
buf ( n361254 , n13577 );
not ( n13579 , n361254 );
or ( n13580 , n13571 , n13579 );
buf ( n361257 , n361251 );
not ( n13582 , n361257 );
buf ( n361259 , n13049 );
not ( n13584 , n361259 );
or ( n13585 , n13582 , n13584 );
nand ( n13586 , n13553 , n13023 );
buf ( n361263 , n13586 );
buf ( n361264 , n361227 );
nand ( n13589 , n361263 , n361264 );
buf ( n361266 , n13589 );
buf ( n361267 , n361266 );
nand ( n13592 , n13585 , n361267 );
buf ( n361269 , n13592 );
not ( n13594 , n361269 );
nand ( n13595 , n13580 , n13594 );
not ( n13596 , n13595 );
xor ( n13597 , n361039 , n13526 );
and ( n13598 , n13597 , n361208 );
and ( n13599 , n361039 , n13526 );
or ( n13600 , n13598 , n13599 );
buf ( n361277 , n553 );
buf ( n361278 , n560 );
and ( n13603 , n361277 , n361278 );
buf ( n361280 , n13603 );
buf ( n361281 , n361280 );
buf ( n361282 , n360921 );
not ( n13607 , n361282 );
buf ( n361284 , n360913 );
not ( n13609 , n361284 );
or ( n13610 , n13607 , n13609 );
buf ( n361287 , n3650 );
buf ( n361288 , n547 );
buf ( n361289 , n564 );
xor ( n13614 , n361288 , n361289 );
buf ( n361291 , n13614 );
buf ( n361292 , n361291 );
nand ( n13617 , n361287 , n361292 );
buf ( n361294 , n13617 );
buf ( n361295 , n361294 );
nand ( n13620 , n13610 , n361295 );
buf ( n361297 , n13620 );
buf ( n361298 , n361297 );
xor ( n13623 , n361281 , n361298 );
buf ( n361300 , n360420 );
buf ( n361301 , n360985 );
and ( n13626 , n361300 , n361301 );
buf ( n361303 , n2550 );
buf ( n361304 , n545 );
buf ( n361305 , n566 );
xor ( n13630 , n361304 , n361305 );
buf ( n361307 , n13630 );
buf ( n361308 , n361307 );
and ( n13633 , n361303 , n361308 );
nor ( n13634 , n13626 , n13633 );
buf ( n361311 , n13634 );
buf ( n361312 , n361311 );
xor ( n13637 , n13623 , n361312 );
buf ( n361314 , n13637 );
buf ( n361315 , n361314 );
xor ( n13640 , n361010 , n361011 );
and ( n13641 , n13640 , n361018 );
and ( n13642 , n361010 , n361011 );
or ( n13643 , n13641 , n13642 );
buf ( n361320 , n13643 );
buf ( n361321 , n361320 );
xor ( n13646 , n361315 , n361321 );
xor ( n13647 , n360891 , n360939 );
and ( n13648 , n13647 , n360995 );
and ( n13649 , n360891 , n360939 );
or ( n13650 , n13648 , n13649 );
buf ( n361327 , n13650 );
buf ( n361328 , n361327 );
xor ( n13653 , n13646 , n361328 );
buf ( n361330 , n13653 );
xor ( n13655 , n360957 , n360974 );
and ( n13656 , n13655 , n360992 );
and ( n13657 , n360957 , n360974 );
or ( n13658 , n13656 , n13657 );
buf ( n361335 , n13658 );
buf ( n361336 , n361335 );
buf ( n361337 , n360901 );
not ( n13662 , n361337 );
buf ( n361339 , n2236 );
not ( n13664 , n361339 );
or ( n13665 , n13662 , n13664 );
buf ( n361342 , n349933 );
buf ( n361343 , n568 );
nand ( n13668 , n361342 , n361343 );
buf ( n361345 , n13668 );
buf ( n361346 , n361345 );
nand ( n13671 , n13665 , n361346 );
buf ( n361348 , n13671 );
buf ( n361349 , n360967 );
not ( n13674 , n361349 );
buf ( n361351 , n8604 );
not ( n13676 , n361351 );
or ( n13677 , n13674 , n13676 );
buf ( n361354 , n352295 );
xor ( n13679 , n549 , n562 );
buf ( n361356 , n13679 );
nand ( n13681 , n361354 , n361356 );
buf ( n361358 , n13681 );
buf ( n361359 , n361358 );
nand ( n13684 , n13677 , n361359 );
buf ( n361361 , n13684 );
xor ( n13686 , n361348 , n361361 );
buf ( n361363 , n360950 );
not ( n13688 , n361363 );
buf ( n361365 , n9186 );
not ( n13690 , n361365 );
or ( n13691 , n13688 , n13690 );
buf ( n361368 , n5407 );
buf ( n361369 , n551 );
buf ( n361370 , n560 );
xor ( n13695 , n361369 , n361370 );
buf ( n361372 , n13695 );
buf ( n361373 , n361372 );
nand ( n13698 , n361368 , n361373 );
buf ( n361375 , n13698 );
buf ( n361376 , n361375 );
nand ( n13701 , n13691 , n361376 );
buf ( n361378 , n13701 );
xor ( n13703 , n13686 , n361378 );
buf ( n361380 , n13703 );
xor ( n13705 , n361336 , n361380 );
xor ( n13706 , n360908 , n360928 );
and ( n13707 , n13706 , n360936 );
and ( n13708 , n360908 , n360928 );
or ( n13709 , n13707 , n13708 );
buf ( n361386 , n13709 );
buf ( n361387 , n361386 );
xor ( n13712 , n13705 , n361387 );
buf ( n361389 , n13712 );
buf ( n13714 , n361389 );
xor ( n13715 , n361021 , n361027 );
and ( n13716 , n13715 , n361034 );
and ( n13717 , n361021 , n361027 );
or ( n13718 , n13716 , n13717 );
buf ( n361395 , n13718 );
nand ( n13720 , n361330 , n13714 , n361395 );
not ( n13721 , n361330 );
not ( n13722 , n13714 );
nand ( n13723 , n13721 , n361395 , n13722 );
not ( n13724 , n361395 );
nand ( n13725 , n13724 , n361330 , n13722 );
not ( n13726 , n361330 );
nand ( n13727 , n13726 , n13724 , n13714 );
nand ( n13728 , n13720 , n13723 , n13725 , n13727 );
xor ( n13729 , n361190 , n361195 );
and ( n13730 , n13729 , n361201 );
and ( n13731 , n361190 , n361195 );
or ( n13732 , n13730 , n13731 );
xor ( n13733 , n13728 , n13732 );
xor ( n13734 , n361152 , n361181 );
and ( n13735 , n13734 , n361188 );
and ( n13736 , n361152 , n361181 );
or ( n13737 , n13735 , n13736 );
buf ( n361414 , n13737 );
xor ( n13739 , n361105 , n361125 );
and ( n13740 , n13739 , n361146 );
and ( n13741 , n361105 , n361125 );
or ( n13742 , n13740 , n13741 );
buf ( n361419 , n13742 );
buf ( n361420 , n361419 );
xor ( n13745 , n361055 , n361066 );
and ( n13746 , n13745 , n361084 );
and ( n13747 , n361055 , n361066 );
or ( n13748 , n13746 , n13747 );
buf ( n361425 , n13748 );
buf ( n361426 , n361425 );
xor ( n13751 , n361420 , n361426 );
not ( n13752 , n13385 );
not ( n13753 , n2471 );
or ( n13754 , n13752 , n13753 );
nand ( n13755 , n350726 , n584 );
nand ( n13756 , n13754 , n13755 );
not ( n13757 , n13756 );
buf ( n361434 , n361118 );
not ( n13759 , n361434 );
buf ( n361436 , n361110 );
not ( n13761 , n361436 );
or ( n13762 , n13759 , n13761 );
buf ( n361439 , n356446 );
buf ( n361440 , n551 );
buf ( n361441 , n576 );
xor ( n13766 , n361440 , n361441 );
buf ( n361443 , n13766 );
buf ( n361444 , n361443 );
nand ( n13769 , n361439 , n361444 );
buf ( n361446 , n13769 );
buf ( n361447 , n361446 );
nand ( n13772 , n13762 , n361447 );
buf ( n361449 , n13772 );
not ( n13774 , n361449 );
not ( n13775 , n13774 );
or ( n13776 , n13757 , n13775 );
not ( n13777 , n13756 );
nand ( n13778 , n13777 , n361449 );
nand ( n13779 , n13776 , n13778 );
buf ( n361456 , n361139 );
not ( n13781 , n361456 );
buf ( n361458 , n361131 );
not ( n13783 , n361458 );
or ( n13784 , n13781 , n13783 );
buf ( n361461 , n354788 );
buf ( n361462 , n549 );
buf ( n361463 , n578 );
xor ( n13788 , n361462 , n361463 );
buf ( n361465 , n13788 );
buf ( n361466 , n361465 );
nand ( n13791 , n361461 , n361466 );
buf ( n361468 , n13791 );
buf ( n361469 , n361468 );
nand ( n13794 , n13784 , n361469 );
buf ( n361471 , n13794 );
and ( n13796 , n13779 , n361471 );
not ( n13797 , n13779 );
not ( n13798 , n361471 );
and ( n13799 , n13797 , n13798 );
nor ( n13800 , n13796 , n13799 );
buf ( n361477 , n13800 );
xor ( n13802 , n13751 , n361477 );
buf ( n361479 , n13802 );
buf ( n361480 , n361479 );
buf ( n361481 , n553 );
buf ( n361482 , n576 );
and ( n13807 , n361481 , n361482 );
buf ( n361484 , n13807 );
buf ( n361485 , n361484 );
buf ( n361486 , n361077 );
not ( n13811 , n361486 );
buf ( n361488 , n3870 );
not ( n13813 , n361488 );
or ( n13814 , n13811 , n13813 );
buf ( n361491 , n351559 );
buf ( n361492 , n547 );
buf ( n361493 , n580 );
xor ( n13818 , n361492 , n361493 );
buf ( n361495 , n13818 );
buf ( n361496 , n361495 );
nand ( n13821 , n361491 , n361496 );
buf ( n361498 , n13821 );
buf ( n361499 , n361498 );
nand ( n13824 , n13814 , n361499 );
buf ( n361501 , n13824 );
buf ( n361502 , n361501 );
xor ( n13827 , n361485 , n361502 );
not ( n13828 , n361098 );
not ( n13829 , n350699 );
or ( n13830 , n13828 , n13829 );
buf ( n361507 , n350705 );
buf ( n361508 , n545 );
buf ( n361509 , n582 );
xor ( n13834 , n361508 , n361509 );
buf ( n361511 , n13834 );
buf ( n361512 , n361511 );
nand ( n13837 , n361507 , n361512 );
buf ( n361514 , n13837 );
nand ( n13839 , n13830 , n361514 );
buf ( n361516 , n13839 );
not ( n13841 , n361516 );
buf ( n361518 , n13841 );
buf ( n361519 , n361518 );
xor ( n13844 , n13827 , n361519 );
buf ( n361521 , n13844 );
buf ( n361522 , n361521 );
buf ( n361523 , n360544 );
buf ( n361524 , n361156 );
nand ( n13849 , n361523 , n361524 );
buf ( n361526 , n13849 );
buf ( n361527 , n361526 );
not ( n13852 , n361527 );
buf ( n361529 , n13487 );
not ( n13854 , n361529 );
or ( n13855 , n13852 , n13854 );
buf ( n361532 , n361156 );
not ( n13857 , n361532 );
buf ( n361534 , n360541 );
nand ( n13859 , n13857 , n361534 );
buf ( n361536 , n13859 );
buf ( n361537 , n361536 );
nand ( n13862 , n13855 , n361537 );
buf ( n361539 , n13862 );
buf ( n361540 , n361539 );
xor ( n13865 , n361522 , n361540 );
xor ( n13866 , n361048 , n361087 );
and ( n13867 , n13866 , n361149 );
and ( n13868 , n361048 , n361087 );
or ( n13869 , n13867 , n13868 );
buf ( n361546 , n13869 );
buf ( n361547 , n361546 );
xor ( n13872 , n13865 , n361547 );
buf ( n361549 , n13872 );
buf ( n361550 , n361549 );
xor ( n13875 , n361480 , n361550 );
xor ( n13876 , n361165 , n361171 );
and ( n13877 , n13876 , n361178 );
and ( n13878 , n361165 , n361171 );
or ( n13879 , n13877 , n13878 );
buf ( n361556 , n13879 );
buf ( n361557 , n361556 );
xor ( n13882 , n13875 , n361557 );
buf ( n361559 , n13882 );
xor ( n13884 , n361414 , n361559 );
xor ( n13885 , n360998 , n361004 );
and ( n13886 , n13885 , n361037 );
and ( n13887 , n360998 , n361004 );
or ( n13888 , n13886 , n13887 );
buf ( n361565 , n13888 );
xor ( n13890 , n13884 , n361565 );
xor ( n13891 , n13733 , n13890 );
nor ( n13892 , n13600 , n13891 );
buf ( n361569 , n13892 );
not ( n13894 , n361569 );
buf ( n361571 , n13894 );
nand ( n13896 , n13891 , n13600 );
nand ( n13897 , n361571 , n13896 );
buf ( n13898 , n13897 );
not ( n13899 , n13898 );
and ( n13900 , n13596 , n13899 );
and ( n13901 , n13595 , n13898 );
nor ( n13902 , n13900 , n13901 );
nor ( n13903 , n13175 , n13179 );
nor ( n13904 , n12637 , n12633 );
nor ( n13905 , n13903 , n13904 );
nand ( n13906 , n13905 , n12520 );
not ( n13907 , n13906 );
not ( n13908 , n13907 );
not ( n13909 , n9005 );
or ( n13910 , n13908 , n13909 );
not ( n13911 , n12527 );
nor ( n13912 , n12385 , n12280 );
nor ( n13913 , n12638 , n13912 );
not ( n13914 , n13913 );
or ( n13915 , n13911 , n13914 );
nand ( n13916 , n12633 , n12637 );
and ( n13917 , n13180 , n13916 );
nand ( n13918 , n13915 , n13917 );
buf ( n13919 , n13183 );
nand ( n13920 , n13918 , n13919 );
nand ( n13921 , n13910 , n13920 );
buf ( n13922 , n13921 );
xor ( n13923 , n13122 , n13132 );
and ( n13924 , n13923 , n13143 );
and ( n13925 , n13122 , n13132 );
or ( n13926 , n13924 , n13925 );
not ( n13927 , n8424 );
not ( n13928 , n5717 );
or ( n13929 , n13927 , n13928 );
nand ( n13930 , n13929 , n554 );
not ( n13931 , n8223 );
not ( n13932 , n13086 );
or ( n13933 , n13931 , n13932 );
not ( n13934 , n544 );
not ( n13935 , n1843 );
not ( n13936 , n13935 );
or ( n13937 , n13934 , n13936 );
nand ( n13938 , n1843 , n7283 );
nand ( n13939 , n13937 , n13938 );
nand ( n13940 , n13939 , n8215 );
nand ( n13941 , n13933 , n13940 );
xor ( n13942 , n13930 , n13941 );
and ( n13943 , n544 , n997 );
xor ( n13944 , n13942 , n13943 );
xor ( n13945 , n13926 , n13944 );
not ( n13946 , n1871 );
not ( n13947 , n13098 );
or ( n13948 , n13946 , n13947 );
and ( n13949 , n552 , n12546 );
not ( n13950 , n552 );
and ( n13951 , n13950 , n12543 );
or ( n13952 , n13949 , n13951 );
nand ( n13953 , n13952 , n4109 );
nand ( n13954 , n13948 , n13953 );
not ( n13955 , n8133 );
not ( n13956 , n548 );
not ( n13957 , n5937 );
or ( n13958 , n13956 , n13957 );
nand ( n13959 , n353618 , n351773 );
nand ( n13960 , n13958 , n13959 );
not ( n13961 , n13960 );
or ( n13962 , n13955 , n13961 );
nand ( n13963 , n13118 , n5751 );
nand ( n13964 , n13962 , n13963 );
xor ( n13965 , n13954 , n13964 );
not ( n13966 , n13153 );
xor ( n13967 , n13965 , n13966 );
xor ( n13968 , n13945 , n13967 );
xor ( n13969 , n13153 , n13157 );
and ( n13970 , n13969 , n13162 );
and ( n13971 , n13153 , n13157 );
or ( n13972 , n13970 , n13971 );
not ( n13973 , n8381 );
not ( n13974 , n13128 );
or ( n13975 , n13973 , n13974 );
and ( n13976 , n5730 , n5761 );
not ( n13977 , n5730 );
and ( n13978 , n13977 , n546 );
or ( n13979 , n13976 , n13978 );
nand ( n13980 , n13979 , n5757 );
nand ( n13981 , n13975 , n13980 );
not ( n13982 , n4078 );
not ( n13983 , n13139 );
or ( n13984 , n13982 , n13983 );
not ( n13985 , n550 );
not ( n13986 , n6082 );
or ( n13987 , n13985 , n13986 );
nand ( n13988 , n6081 , n1880 );
nand ( n13989 , n13987 , n13988 );
nand ( n13990 , n13989 , n1875 );
nand ( n13991 , n13984 , n13990 );
xor ( n13992 , n13981 , n13991 );
xor ( n13993 , n13090 , n13092 );
and ( n13994 , n13993 , n13102 );
and ( n13995 , n13090 , n13092 );
or ( n13996 , n13994 , n13995 );
xor ( n13997 , n13992 , n13996 );
xor ( n13998 , n13972 , n13997 );
xor ( n13999 , n13103 , n13107 );
and ( n14000 , n13999 , n13144 );
and ( n14001 , n13103 , n13107 );
or ( n14002 , n14000 , n14001 );
xor ( n14003 , n13998 , n14002 );
xor ( n14004 , n13968 , n14003 );
xor ( n14005 , n13149 , n13163 );
and ( n14006 , n14005 , n13168 );
and ( n14007 , n13149 , n13163 );
or ( n14008 , n14006 , n14007 );
xor ( n14009 , n14004 , n14008 );
buf ( n14010 , n14009 );
not ( n14011 , n14010 );
xor ( n14012 , n13145 , n13169 );
and ( n14013 , n14012 , n13174 );
and ( n14014 , n13145 , n13169 );
or ( n14015 , n14013 , n14014 );
not ( n14016 , n14015 );
nand ( n14017 , n14011 , n14016 );
nand ( n14018 , n14009 , n14015 );
nand ( n14019 , n14017 , n14018 );
not ( n14020 , n14019 );
and ( n14021 , n13922 , n14020 );
not ( n14022 , n13922 );
and ( n14023 , n14022 , n14019 );
nor ( n14024 , n14021 , n14023 );
nand ( n14025 , n13902 , n14024 );
and ( n14026 , n12517 , n14025 );
nand ( n14027 , n13567 , n14026 , n8298 );
and ( n14028 , n13565 , n14025 );
not ( n14029 , n12514 );
not ( n14030 , n14029 );
and ( n14031 , n14028 , n14030 );
not ( n14032 , n14025 );
not ( n14033 , n13563 );
not ( n14034 , n13062 );
or ( n14035 , n14033 , n14034 );
not ( n14036 , n13189 );
not ( n14037 , n13562 );
nand ( n14038 , n14036 , n14037 );
nand ( n14039 , n14035 , n14038 );
not ( n14040 , n14039 );
or ( n14041 , n14032 , n14040 );
nor ( n14042 , n13902 , n14024 );
not ( n14043 , n14042 );
nand ( n14044 , n14041 , n14043 );
nor ( n14045 , n14031 , n14044 );
nand ( n14046 , n14027 , n14045 );
not ( n14047 , n14017 );
not ( n14048 , n13921 );
or ( n14049 , n14047 , n14048 );
buf ( n14050 , n14018 );
nand ( n14051 , n14049 , n14050 );
xor ( n14052 , n13930 , n13941 );
and ( n14053 , n14052 , n13943 );
and ( n14054 , n13930 , n13941 );
or ( n14055 , n14053 , n14054 );
xor ( n14056 , n13954 , n13964 );
and ( n14057 , n14056 , n13966 );
and ( n14058 , n13954 , n13964 );
or ( n14059 , n14057 , n14058 );
xor ( n14060 , n14055 , n14059 );
not ( n14061 , n8215 );
xor ( n14062 , n544 , n5720 );
not ( n14063 , n14062 );
or ( n14064 , n14061 , n14063 );
nand ( n14065 , n13939 , n8223 );
nand ( n14066 , n14064 , n14065 );
not ( n14067 , n5751 );
not ( n14068 , n13960 );
or ( n14069 , n14067 , n14068 );
not ( n14070 , n548 );
not ( n14071 , n6035 );
or ( n14072 , n14070 , n14071 );
nand ( n14073 , n6034 , n351773 );
nand ( n14074 , n14072 , n14073 );
nand ( n14075 , n14074 , n8133 );
nand ( n14076 , n14069 , n14075 );
xor ( n14077 , n14066 , n14076 );
and ( n14078 , n13952 , n1871 );
nor ( n14079 , n14078 , n7214 );
xor ( n14080 , n14077 , n14079 );
xor ( n14081 , n14060 , n14080 );
not ( n14082 , n544 );
buf ( n14083 , n1789 );
nor ( n14084 , n14082 , n14083 );
not ( n14085 , n1875 );
not ( n14086 , n550 );
buf ( n14087 , n7246 );
not ( n14088 , n14087 );
not ( n14089 , n14088 );
or ( n14090 , n14086 , n14089 );
nand ( n14091 , n14087 , n1880 );
nand ( n14092 , n14090 , n14091 );
not ( n14093 , n14092 );
or ( n14094 , n14085 , n14093 );
nand ( n14095 , n13989 , n4078 );
nand ( n14096 , n14094 , n14095 );
xor ( n14097 , n14084 , n14096 );
not ( n14098 , n8381 );
not ( n14099 , n13979 );
or ( n14100 , n14098 , n14099 );
not ( n14101 , n546 );
not ( n14102 , n5962 );
or ( n14103 , n14101 , n14102 );
nand ( n14104 , n353641 , n5761 );
nand ( n14105 , n14103 , n14104 );
nand ( n14106 , n14105 , n353673 );
nand ( n14107 , n14100 , n14106 );
xor ( n14108 , n14097 , n14107 );
xor ( n14109 , n13981 , n13991 );
and ( n14110 , n14109 , n13996 );
and ( n14111 , n13981 , n13991 );
or ( n14112 , n14110 , n14111 );
xor ( n14113 , n14108 , n14112 );
xor ( n14114 , n13926 , n13944 );
and ( n14115 , n14114 , n13967 );
and ( n14116 , n13926 , n13944 );
or ( n14117 , n14115 , n14116 );
xor ( n14118 , n14113 , n14117 );
xor ( n14119 , n14081 , n14118 );
xor ( n14120 , n13972 , n13997 );
and ( n14121 , n14120 , n14002 );
and ( n14122 , n13972 , n13997 );
or ( n14123 , n14121 , n14122 );
xor ( n14124 , n14119 , n14123 );
xor ( n14125 , n13968 , n14003 );
and ( n14126 , n14125 , n14008 );
and ( n14127 , n13968 , n14003 );
or ( n14128 , n14126 , n14127 );
nor ( n14129 , n14124 , n14128 );
not ( n14130 , n14129 );
buf ( n14131 , n14124 );
nand ( n14132 , n14131 , n14128 );
nand ( n14133 , n14130 , n14132 );
not ( n14134 , n14133 );
and ( n14135 , n14051 , n14134 );
not ( n14136 , n14051 );
and ( n14137 , n14136 , n14133 );
nor ( n14138 , n14135 , n14137 );
buf ( n361815 , n361251 );
buf ( n361816 , n361571 );
and ( n14141 , n361815 , n361816 );
buf ( n361818 , n14141 );
not ( n14143 , n361818 );
not ( n14144 , n360706 );
not ( n14145 , n361246 );
or ( n14146 , n14144 , n14145 );
nand ( n14147 , n14146 , n360728 );
not ( n14148 , n14147 );
or ( n14149 , n14143 , n14148 );
nand ( n14150 , n13586 , n361571 , n361227 );
nand ( n14151 , n14150 , n13896 );
xor ( n14152 , n13728 , n13732 );
and ( n14153 , n14152 , n13890 );
and ( n14154 , n13728 , n13732 );
or ( n14155 , n14153 , n14154 );
buf ( n361832 , n14155 );
xor ( n14157 , n361336 , n361380 );
and ( n14158 , n14157 , n361387 );
and ( n14159 , n361336 , n361380 );
or ( n14160 , n14158 , n14159 );
buf ( n361837 , n14160 );
buf ( n361838 , n361837 );
buf ( n361839 , n361311 );
not ( n14164 , n361839 );
buf ( n361841 , n14164 );
buf ( n361842 , n361841 );
buf ( n361843 , n361378 );
not ( n14168 , n361843 );
buf ( n361845 , n361348 );
not ( n14170 , n361845 );
or ( n14171 , n14168 , n14170 );
buf ( n361848 , n361348 );
buf ( n361849 , n361378 );
or ( n14174 , n361848 , n361849 );
buf ( n361851 , n361361 );
nand ( n14176 , n14174 , n361851 );
buf ( n361853 , n14176 );
buf ( n361854 , n361853 );
nand ( n14179 , n14171 , n361854 );
buf ( n361856 , n14179 );
buf ( n361857 , n361856 );
xor ( n14182 , n361842 , n361857 );
buf ( n361859 , n552 );
buf ( n361860 , n560 );
and ( n14185 , n361859 , n361860 );
buf ( n361862 , n14185 );
buf ( n361863 , n361862 );
buf ( n361864 , n361372 );
not ( n14189 , n361864 );
buf ( n361866 , n9186 );
not ( n14191 , n361866 );
or ( n14192 , n14189 , n14191 );
buf ( n361869 , n5407 );
buf ( n361870 , n550 );
buf ( n361871 , n560 );
xor ( n14196 , n361870 , n361871 );
buf ( n361873 , n14196 );
buf ( n361874 , n361873 );
nand ( n14199 , n361869 , n361874 );
buf ( n361876 , n14199 );
buf ( n361877 , n361876 );
nand ( n14202 , n14192 , n361877 );
buf ( n361879 , n14202 );
buf ( n361880 , n361879 );
xor ( n14205 , n361863 , n361880 );
buf ( n361882 , n361291 );
not ( n14207 , n361882 );
buf ( n361884 , n360913 );
not ( n14209 , n361884 );
or ( n14210 , n14207 , n14209 );
buf ( n361887 , n3650 );
buf ( n361888 , n546 );
buf ( n361889 , n564 );
xor ( n14214 , n361888 , n361889 );
buf ( n361891 , n14214 );
buf ( n361892 , n361891 );
nand ( n14217 , n361887 , n361892 );
buf ( n361894 , n14217 );
buf ( n361895 , n361894 );
nand ( n14220 , n14210 , n361895 );
buf ( n361897 , n14220 );
buf ( n361898 , n361897 );
xor ( n14223 , n14205 , n361898 );
buf ( n361900 , n14223 );
buf ( n361901 , n361900 );
xor ( n14226 , n14182 , n361901 );
buf ( n361903 , n14226 );
buf ( n361904 , n361307 );
not ( n14229 , n361904 );
buf ( n361906 , n360420 );
not ( n14231 , n361906 );
or ( n14232 , n14229 , n14231 );
buf ( n361909 , n2550 );
buf ( n361910 , n544 );
buf ( n361911 , n566 );
xor ( n14236 , n361910 , n361911 );
buf ( n361913 , n14236 );
buf ( n361914 , n361913 );
nand ( n14239 , n361909 , n361914 );
buf ( n361916 , n14239 );
buf ( n361917 , n361916 );
nand ( n14242 , n14232 , n361917 );
buf ( n361919 , n14242 );
buf ( n361920 , n361919 );
not ( n14245 , n361920 );
buf ( n361922 , n2236 );
buf ( n361923 , n349933 );
or ( n14248 , n361922 , n361923 );
buf ( n361925 , n568 );
nand ( n14250 , n14248 , n361925 );
buf ( n361927 , n14250 );
buf ( n361928 , n361927 );
not ( n14253 , n361928 );
buf ( n361930 , n14253 );
buf ( n361931 , n361930 );
not ( n14256 , n361931 );
or ( n14257 , n14245 , n14256 );
buf ( n361934 , n361919 );
buf ( n361935 , n361930 );
or ( n14260 , n361934 , n361935 );
nand ( n14261 , n14257 , n14260 );
buf ( n361938 , n14261 );
buf ( n361939 , n361938 );
buf ( n361940 , n548 );
buf ( n361941 , n562 );
xor ( n14266 , n361940 , n361941 );
buf ( n361943 , n14266 );
and ( n14268 , n352295 , n361943 );
nand ( n14269 , n13679 , n8603 );
not ( n14270 , n14269 );
nor ( n14271 , n14268 , n14270 );
buf ( n361948 , n14271 );
and ( n14273 , n361939 , n361948 );
not ( n14274 , n361939 );
not ( n14275 , n361943 );
not ( n14276 , n352295 );
or ( n14277 , n14275 , n14276 );
nand ( n14278 , n14277 , n14269 );
buf ( n361955 , n14278 );
and ( n14280 , n14274 , n361955 );
nor ( n14281 , n14273 , n14280 );
buf ( n361958 , n14281 );
buf ( n361959 , n361958 );
not ( n14284 , n361959 );
buf ( n361961 , n14284 );
xor ( n14286 , n361281 , n361298 );
and ( n14287 , n14286 , n361312 );
and ( n14288 , n361281 , n361298 );
or ( n14289 , n14287 , n14288 );
buf ( n361966 , n14289 );
buf ( n361967 , n361966 );
not ( n14292 , n361967 );
buf ( n361969 , n14292 );
xor ( n14294 , n361961 , n361969 );
xnor ( n14295 , n361903 , n14294 );
buf ( n361972 , n14295 );
xor ( n14297 , n361838 , n361972 );
xor ( n14298 , n361315 , n361321 );
and ( n14299 , n14298 , n361328 );
and ( n14300 , n361315 , n361321 );
or ( n14301 , n14299 , n14300 );
buf ( n361978 , n14301 );
buf ( n361979 , n361978 );
xor ( n14304 , n14297 , n361979 );
buf ( n361981 , n14304 );
buf ( n361982 , n361981 );
xor ( n14307 , n361414 , n361559 );
and ( n14308 , n14307 , n361565 );
and ( n14309 , n361414 , n361559 );
or ( n14310 , n14308 , n14309 );
buf ( n361987 , n14310 );
xor ( n14312 , n361982 , n361987 );
xor ( n14313 , n361480 , n361550 );
and ( n14314 , n14313 , n361557 );
and ( n14315 , n361480 , n361550 );
or ( n14316 , n14314 , n14315 );
buf ( n361993 , n14316 );
buf ( n361994 , n361993 );
xor ( n14319 , n361420 , n361426 );
and ( n14320 , n14319 , n361477 );
and ( n14321 , n361420 , n361426 );
or ( n14322 , n14320 , n14321 );
buf ( n361999 , n14322 );
buf ( n362000 , n361999 );
xor ( n14325 , n361522 , n361540 );
and ( n14326 , n14325 , n361547 );
and ( n14327 , n361522 , n361540 );
or ( n14328 , n14326 , n14327 );
buf ( n362005 , n14328 );
buf ( n362006 , n362005 );
xor ( n14331 , n362000 , n362006 );
xor ( n14332 , n361485 , n361502 );
and ( n14333 , n14332 , n361519 );
and ( n14334 , n361485 , n361502 );
or ( n14335 , n14333 , n14334 );
buf ( n362012 , n14335 );
buf ( n362013 , n362012 );
buf ( n362014 , n361511 );
not ( n14339 , n362014 );
buf ( n362016 , n350699 );
not ( n14341 , n362016 );
or ( n14342 , n14339 , n14341 );
buf ( n362019 , n350705 );
buf ( n362020 , n544 );
buf ( n362021 , n582 );
xor ( n14346 , n362020 , n362021 );
buf ( n362023 , n14346 );
buf ( n362024 , n362023 );
nand ( n14349 , n362019 , n362024 );
buf ( n362026 , n14349 );
buf ( n362027 , n362026 );
nand ( n14352 , n14342 , n362027 );
buf ( n362029 , n14352 );
buf ( n362030 , n362029 );
not ( n14355 , n348626 );
not ( n14356 , n2470 );
or ( n14357 , n14355 , n14356 );
nand ( n14358 , n14357 , n584 );
buf ( n362035 , n14358 );
xor ( n14360 , n362030 , n362035 );
buf ( n362037 , n361465 );
not ( n14362 , n362037 );
buf ( n362039 , n361131 );
not ( n14364 , n362039 );
or ( n14365 , n14362 , n14364 );
buf ( n362042 , n354788 );
buf ( n362043 , n548 );
buf ( n362044 , n578 );
xor ( n14369 , n362043 , n362044 );
buf ( n362046 , n14369 );
buf ( n362047 , n362046 );
nand ( n14372 , n362042 , n362047 );
buf ( n362049 , n14372 );
buf ( n362050 , n362049 );
nand ( n14375 , n14365 , n362050 );
buf ( n362052 , n14375 );
buf ( n362053 , n362052 );
xor ( n14378 , n14360 , n362053 );
buf ( n362055 , n14378 );
buf ( n362056 , n362055 );
xor ( n14381 , n362013 , n362056 );
not ( n14382 , n361449 );
not ( n14383 , n361471 );
or ( n14384 , n14382 , n14383 );
or ( n14385 , n361471 , n361449 );
nand ( n14386 , n14385 , n13756 );
nand ( n14387 , n14384 , n14386 );
xor ( n14388 , n13839 , n14387 );
buf ( n362065 , n552 );
buf ( n362066 , n576 );
and ( n14391 , n362065 , n362066 );
buf ( n362068 , n14391 );
buf ( n362069 , n361495 );
not ( n14394 , n362069 );
buf ( n362071 , n3870 );
not ( n14396 , n362071 );
or ( n14397 , n14394 , n14396 );
buf ( n362074 , n351559 );
buf ( n362075 , n546 );
buf ( n362076 , n580 );
xor ( n14401 , n362075 , n362076 );
buf ( n362078 , n14401 );
buf ( n362079 , n362078 );
nand ( n14404 , n362074 , n362079 );
buf ( n362081 , n14404 );
buf ( n362082 , n362081 );
nand ( n14407 , n14397 , n362082 );
buf ( n362084 , n14407 );
xor ( n14409 , n362068 , n362084 );
buf ( n362086 , n361443 );
not ( n14411 , n362086 );
buf ( n362088 , n361110 );
not ( n14413 , n362088 );
or ( n14414 , n14411 , n14413 );
buf ( n362091 , n356446 );
buf ( n362092 , n550 );
buf ( n362093 , n576 );
xor ( n14418 , n362092 , n362093 );
buf ( n362095 , n14418 );
buf ( n362096 , n362095 );
nand ( n14421 , n362091 , n362096 );
buf ( n362098 , n14421 );
buf ( n362099 , n362098 );
nand ( n14424 , n14414 , n362099 );
buf ( n362101 , n14424 );
xor ( n14426 , n14409 , n362101 );
xor ( n14427 , n14388 , n14426 );
buf ( n362104 , n14427 );
xor ( n14429 , n14381 , n362104 );
buf ( n362106 , n14429 );
buf ( n362107 , n362106 );
xor ( n14432 , n14331 , n362107 );
buf ( n362109 , n14432 );
buf ( n362110 , n362109 );
xor ( n14435 , n361994 , n362110 );
not ( n14436 , n361330 );
not ( n14437 , n13714 );
or ( n14438 , n14436 , n14437 );
or ( n14439 , n361330 , n13714 );
nand ( n14440 , n14439 , n361395 );
nand ( n14441 , n14438 , n14440 );
buf ( n362118 , n14441 );
xor ( n14443 , n14435 , n362118 );
buf ( n362120 , n14443 );
buf ( n362121 , n362120 );
xor ( n14446 , n14312 , n362121 );
buf ( n362123 , n14446 );
buf ( n362124 , n362123 );
nor ( n14449 , n361832 , n362124 );
buf ( n362126 , n14449 );
buf ( n362127 , n362126 );
buf ( n14452 , n362127 );
buf ( n362129 , n14452 );
not ( n14454 , n362129 );
buf ( n362131 , n14155 );
buf ( n362132 , n362123 );
nand ( n14457 , n362131 , n362132 );
buf ( n362134 , n14457 );
nand ( n14459 , n14454 , n362134 );
nor ( n14460 , n14151 , n14459 );
nand ( n14461 , n14149 , n14460 );
nand ( n14462 , n14151 , n14459 );
nand ( n14463 , n14147 , n14459 , n361818 );
nand ( n14464 , n14461 , n14462 , n14463 );
not ( n14465 , n14464 );
nand ( n14466 , n14138 , n14465 );
buf ( n14467 , n14466 );
not ( n14468 , n14138 );
buf ( n14469 , n14464 );
nand ( n14470 , n14468 , n14469 );
buf ( n14471 , n14470 );
nand ( n14472 , n14467 , n14471 );
xnor ( n14473 , n14046 , n14472 );
nand ( n14474 , n14043 , n14025 );
not ( n14475 , n14474 );
not ( n14476 , n14475 );
nand ( n14477 , n12514 , n13565 );
not ( n14478 , n14039 );
nand ( n14479 , n13565 , n12517 , n8298 );
nand ( n14480 , n14477 , n14478 , n14479 );
not ( n14481 , n14480 );
not ( n14482 , n14481 );
or ( n14483 , n14476 , n14482 );
nand ( n14484 , n14480 , n14474 );
nand ( n14485 , n14483 , n14484 );
and ( n14486 , n14038 , n13563 );
not ( n14487 , n11863 );
and ( n14488 , n13065 , n12400 );
and ( n14489 , n14487 , n14488 );
not ( n14490 , n12397 );
not ( n14491 , n13065 );
or ( n14492 , n14490 , n14491 );
nand ( n14493 , n14492 , n13063 );
nor ( n14494 , n14489 , n14493 );
nand ( n14495 , n13066 , n8298 , n12517 );
nand ( n14496 , n14494 , n14495 );
xor ( n14497 , n14486 , n14496 );
buf ( n14498 , n14497 );
nand ( n14499 , n13075 , n14473 , n14485 , n14498 );
not ( n14500 , n14499 );
not ( n14501 , n14500 );
not ( n14502 , n14501 );
not ( n14503 , n13902 );
not ( n14504 , n14024 );
or ( n14505 , n14503 , n14504 );
nand ( n14506 , n14505 , n14466 );
not ( n14507 , n14506 );
and ( n14508 , n13563 , n13065 );
nand ( n14509 , n14507 , n14508 );
not ( n14510 , n14509 );
buf ( n14511 , n14510 );
not ( n14512 , n14029 );
and ( n14513 , n14511 , n14512 );
not ( n14514 , n14507 );
not ( n14515 , n14039 );
or ( n14516 , n14514 , n14515 );
not ( n14517 , n14042 );
not ( n14518 , n14466 );
or ( n14519 , n14517 , n14518 );
nand ( n14520 , n14519 , n14470 );
not ( n14521 , n14520 );
nand ( n14522 , n14516 , n14521 );
nor ( n14523 , n14513 , n14522 );
nand ( n14524 , n14510 , n12517 );
not ( n14525 , n14524 );
nand ( n14526 , n8298 , n14525 );
nand ( n14527 , n14523 , n14526 );
not ( n14528 , n14527 );
xor ( n14529 , n14081 , n14118 );
and ( n14530 , n14529 , n14123 );
and ( n14531 , n14081 , n14118 );
or ( n14532 , n14530 , n14531 );
not ( n14533 , n14532 );
xor ( n14534 , n14055 , n14059 );
and ( n14535 , n14534 , n14080 );
and ( n14536 , n14055 , n14059 );
or ( n14537 , n14535 , n14536 );
not ( n14538 , n8393 );
not ( n14539 , n353522 );
or ( n14540 , n14538 , n14539 );
nand ( n14541 , n14540 , n552 );
not ( n14542 , n544 );
nor ( n14543 , n14542 , n13935 );
xor ( n14544 , n14541 , n14543 );
not ( n14545 , n4078 );
not ( n14546 , n14092 );
or ( n14547 , n14545 , n14546 );
not ( n14548 , n1880 );
buf ( n14549 , n12543 );
not ( n14550 , n14549 );
or ( n14551 , n14548 , n14550 );
not ( n14552 , n14549 );
nand ( n14553 , n14552 , n550 );
nand ( n14554 , n14551 , n14553 );
nand ( n14555 , n14554 , n1875 );
nand ( n14556 , n14547 , n14555 );
xor ( n14557 , n14544 , n14556 );
not ( n14558 , n8381 );
not ( n14559 , n14105 );
or ( n14560 , n14558 , n14559 );
not ( n14561 , n546 );
not ( n14562 , n5937 );
or ( n14563 , n14561 , n14562 );
nand ( n14564 , n353618 , n5761 );
nand ( n14565 , n14563 , n14564 );
nand ( n14566 , n14565 , n353673 );
nand ( n14567 , n14560 , n14566 );
not ( n14568 , n8223 );
not ( n14569 , n14062 );
or ( n14570 , n14568 , n14569 );
xor ( n14571 , n544 , n5730 );
nand ( n14572 , n14571 , n8215 );
nand ( n14573 , n14570 , n14572 );
xor ( n14574 , n14567 , n14573 );
not ( n14575 , n5751 );
not ( n14576 , n14074 );
or ( n14577 , n14575 , n14576 );
not ( n14578 , n548 );
not ( n14579 , n6082 );
or ( n14580 , n14578 , n14579 );
not ( n14581 , n6082 );
nand ( n14582 , n14581 , n351773 );
nand ( n14583 , n14580 , n14582 );
nand ( n14584 , n14583 , n8133 );
nand ( n14585 , n14577 , n14584 );
xor ( n14586 , n14574 , n14585 );
xor ( n14587 , n14557 , n14586 );
not ( n14588 , n14079 );
xor ( n14589 , n14084 , n14096 );
and ( n14590 , n14589 , n14107 );
and ( n14591 , n14084 , n14096 );
or ( n14592 , n14590 , n14591 );
xor ( n14593 , n14588 , n14592 );
xor ( n14594 , n14066 , n14076 );
and ( n14595 , n14594 , n14079 );
and ( n14596 , n14066 , n14076 );
or ( n14597 , n14595 , n14596 );
xor ( n14598 , n14593 , n14597 );
xor ( n14599 , n14587 , n14598 );
xor ( n14600 , n14537 , n14599 );
xor ( n14601 , n14108 , n14112 );
and ( n14602 , n14601 , n14117 );
and ( n14603 , n14108 , n14112 );
or ( n14604 , n14602 , n14603 );
xor ( n14605 , n14600 , n14604 );
not ( n14606 , n14605 );
nand ( n14607 , n14533 , n14606 );
nand ( n14608 , n14532 , n14605 );
nand ( n14609 , n14607 , n14608 );
not ( n14610 , n14609 );
not ( n14611 , n14610 );
nor ( n14612 , n14010 , n14015 );
nor ( n14613 , n14129 , n14612 );
not ( n14614 , n14613 );
not ( n14615 , n13922 );
or ( n14616 , n14614 , n14615 );
nor ( n14617 , n14128 , n14124 );
or ( n14618 , n14617 , n14018 );
nand ( n14619 , n14124 , n14128 );
nand ( n14620 , n14618 , n14619 );
buf ( n14621 , n14620 );
not ( n14622 , n14621 );
nand ( n14623 , n14616 , n14622 );
not ( n14624 , n14623 );
not ( n14625 , n14624 );
or ( n14626 , n14611 , n14625 );
nand ( n14627 , n14623 , n14609 );
nand ( n14628 , n14626 , n14627 );
xor ( n14629 , n361838 , n361972 );
and ( n14630 , n14629 , n361979 );
and ( n14631 , n361838 , n361972 );
or ( n14632 , n14630 , n14631 );
buf ( n362309 , n14632 );
buf ( n362310 , n362309 );
xor ( n14635 , n13839 , n14387 );
and ( n14636 , n14635 , n14426 );
and ( n14637 , n13839 , n14387 );
or ( n14638 , n14636 , n14637 );
buf ( n362315 , n14638 );
buf ( n362316 , n551 );
buf ( n362317 , n576 );
and ( n14642 , n362316 , n362317 );
buf ( n362319 , n14642 );
not ( n14644 , n362023 );
not ( n14645 , n350699 );
or ( n14646 , n14644 , n14645 );
buf ( n362323 , n350705 );
buf ( n362324 , n582 );
nand ( n14649 , n362323 , n362324 );
buf ( n362326 , n14649 );
nand ( n14651 , n14646 , n362326 );
xor ( n14652 , n362319 , n14651 );
buf ( n362329 , n362095 );
not ( n14654 , n362329 );
buf ( n362331 , n361110 );
not ( n14656 , n362331 );
or ( n14657 , n14654 , n14656 );
buf ( n362334 , n356446 );
buf ( n362335 , n549 );
buf ( n362336 , n576 );
xor ( n14661 , n362335 , n362336 );
buf ( n362338 , n14661 );
buf ( n362339 , n362338 );
nand ( n14664 , n362334 , n362339 );
buf ( n362341 , n14664 );
buf ( n362342 , n362341 );
nand ( n14667 , n14657 , n362342 );
buf ( n362344 , n14667 );
xor ( n14669 , n14652 , n362344 );
buf ( n362346 , n14669 );
xor ( n14671 , n362030 , n362035 );
and ( n14672 , n14671 , n362053 );
and ( n14673 , n362030 , n362035 );
or ( n14674 , n14672 , n14673 );
buf ( n362351 , n14674 );
buf ( n362352 , n362351 );
xor ( n14677 , n362346 , n362352 );
buf ( n362354 , n362046 );
not ( n14679 , n362354 );
buf ( n362356 , n361131 );
not ( n14681 , n362356 );
or ( n14682 , n14679 , n14681 );
buf ( n362359 , n354788 );
buf ( n362360 , n547 );
buf ( n362361 , n578 );
xor ( n14686 , n362360 , n362361 );
buf ( n362363 , n14686 );
buf ( n362364 , n362363 );
nand ( n14689 , n362359 , n362364 );
buf ( n362366 , n14689 );
buf ( n362367 , n362366 );
nand ( n14692 , n14682 , n362367 );
buf ( n362369 , n14692 );
buf ( n362370 , n362369 );
buf ( n362371 , n362078 );
not ( n14696 , n362371 );
buf ( n362373 , n3870 );
buf ( n14698 , n362373 );
buf ( n362375 , n14698 );
buf ( n362376 , n362375 );
not ( n14701 , n362376 );
or ( n14702 , n14696 , n14701 );
buf ( n362379 , n351559 );
buf ( n362380 , n545 );
buf ( n362381 , n580 );
xor ( n14706 , n362380 , n362381 );
buf ( n362383 , n14706 );
buf ( n362384 , n362383 );
nand ( n14709 , n362379 , n362384 );
buf ( n362386 , n14709 );
buf ( n362387 , n362386 );
nand ( n14712 , n14702 , n362387 );
buf ( n362389 , n14712 );
buf ( n362390 , n362389 );
not ( n14715 , n362390 );
buf ( n362392 , n14715 );
buf ( n362393 , n362392 );
xor ( n14718 , n362370 , n362393 );
not ( n14719 , n362101 );
or ( n14720 , n362084 , n362068 );
not ( n14721 , n14720 );
or ( n14722 , n14719 , n14721 );
nand ( n14723 , n362084 , n362068 );
nand ( n14724 , n14722 , n14723 );
buf ( n362401 , n14724 );
xor ( n14726 , n14718 , n362401 );
buf ( n362403 , n14726 );
buf ( n362404 , n362403 );
xor ( n14729 , n14677 , n362404 );
buf ( n362406 , n14729 );
buf ( n362407 , n362406 );
xor ( n14732 , n362315 , n362407 );
xor ( n14733 , n362013 , n362056 );
and ( n14734 , n14733 , n362104 );
and ( n14735 , n362013 , n362056 );
or ( n14736 , n14734 , n14735 );
buf ( n362413 , n14736 );
buf ( n362414 , n362413 );
xor ( n14739 , n14732 , n362414 );
buf ( n362416 , n14739 );
buf ( n362417 , n362416 );
not ( n14742 , n362417 );
buf ( n362419 , n14742 );
buf ( n362420 , n362419 );
and ( n14745 , n362310 , n362420 );
not ( n14746 , n362310 );
buf ( n362423 , n362416 );
and ( n14748 , n14746 , n362423 );
nor ( n14749 , n14745 , n14748 );
buf ( n362426 , n14749 );
xor ( n14751 , n362000 , n362006 );
and ( n14752 , n14751 , n362107 );
and ( n14753 , n362000 , n362006 );
or ( n14754 , n14752 , n14753 );
buf ( n362431 , n14754 );
not ( n14756 , n362431 );
and ( n14757 , n362426 , n14756 );
not ( n14758 , n362426 );
and ( n14759 , n14758 , n362431 );
nor ( n14760 , n14757 , n14759 );
not ( n14761 , n14760 );
not ( n14762 , n14761 );
xor ( n14763 , n361994 , n362110 );
and ( n14764 , n14763 , n362118 );
and ( n14765 , n361994 , n362110 );
or ( n14766 , n14764 , n14765 );
buf ( n362443 , n14766 );
xor ( n14768 , n361842 , n361857 );
and ( n14769 , n14768 , n361901 );
and ( n14770 , n361842 , n361857 );
or ( n14771 , n14769 , n14770 );
buf ( n362448 , n14771 );
buf ( n362449 , n362448 );
buf ( n362450 , n551 );
buf ( n362451 , n560 );
and ( n14776 , n362450 , n362451 );
buf ( n362453 , n14776 );
buf ( n362454 , n362453 );
buf ( n362455 , n361873 );
not ( n14780 , n362455 );
buf ( n362457 , n9186 );
not ( n14782 , n362457 );
or ( n14783 , n14780 , n14782 );
buf ( n362460 , n5407 );
buf ( n362461 , n549 );
buf ( n362462 , n560 );
xor ( n14787 , n362461 , n362462 );
buf ( n362464 , n14787 );
buf ( n362465 , n362464 );
nand ( n14790 , n362460 , n362465 );
buf ( n362467 , n14790 );
buf ( n362468 , n362467 );
nand ( n14793 , n14783 , n362468 );
buf ( n362470 , n14793 );
buf ( n362471 , n362470 );
xor ( n14796 , n362454 , n362471 );
buf ( n362473 , n361913 );
not ( n14798 , n362473 );
buf ( n362475 , n360420 );
not ( n14800 , n362475 );
or ( n14801 , n14798 , n14800 );
buf ( n362478 , n2550 );
buf ( n362479 , n566 );
nand ( n14804 , n362478 , n362479 );
buf ( n362481 , n14804 );
buf ( n362482 , n362481 );
nand ( n14807 , n14801 , n362482 );
buf ( n362484 , n14807 );
buf ( n362485 , n362484 );
xor ( n14810 , n14796 , n362485 );
buf ( n362487 , n14810 );
buf ( n362488 , n362487 );
buf ( n362489 , n14271 );
not ( n14814 , n362489 );
buf ( n362491 , n361930 );
not ( n14816 , n362491 );
or ( n14817 , n14814 , n14816 );
buf ( n362494 , n361919 );
nand ( n14819 , n14817 , n362494 );
buf ( n362496 , n14819 );
buf ( n362497 , n362496 );
buf ( n362498 , n361927 );
buf ( n362499 , n14278 );
nand ( n14824 , n362498 , n362499 );
buf ( n362501 , n14824 );
buf ( n362502 , n362501 );
nand ( n14827 , n362497 , n362502 );
buf ( n362504 , n14827 );
buf ( n362505 , n362504 );
xor ( n14830 , n362488 , n362505 );
buf ( n362507 , n361943 );
not ( n14832 , n362507 );
buf ( n362509 , n8604 );
not ( n14834 , n362509 );
or ( n14835 , n14832 , n14834 );
buf ( n362512 , n352295 );
buf ( n362513 , n547 );
buf ( n362514 , n562 );
xor ( n14839 , n362513 , n362514 );
buf ( n362516 , n14839 );
buf ( n362517 , n362516 );
nand ( n14842 , n362512 , n362517 );
buf ( n362519 , n14842 );
buf ( n362520 , n362519 );
nand ( n14845 , n14835 , n362520 );
buf ( n362522 , n14845 );
buf ( n362523 , n362522 );
buf ( n362524 , n361891 );
not ( n14849 , n362524 );
buf ( n362526 , n360913 );
not ( n14851 , n362526 );
or ( n14852 , n14849 , n14851 );
buf ( n362529 , n3650 );
buf ( n362530 , n545 );
buf ( n362531 , n564 );
xor ( n14856 , n362530 , n362531 );
buf ( n362533 , n14856 );
buf ( n362534 , n362533 );
nand ( n14859 , n362529 , n362534 );
buf ( n362536 , n14859 );
buf ( n362537 , n362536 );
nand ( n14862 , n14852 , n362537 );
buf ( n362539 , n14862 );
buf ( n362540 , n362539 );
not ( n14865 , n362540 );
buf ( n362542 , n14865 );
buf ( n362543 , n362542 );
xor ( n14868 , n362523 , n362543 );
xor ( n14869 , n361863 , n361880 );
and ( n14870 , n14869 , n361898 );
and ( n14871 , n361863 , n361880 );
or ( n14872 , n14870 , n14871 );
buf ( n362549 , n14872 );
buf ( n362550 , n362549 );
xor ( n14875 , n14868 , n362550 );
buf ( n362552 , n14875 );
buf ( n362553 , n362552 );
xor ( n14878 , n14830 , n362553 );
buf ( n362555 , n14878 );
buf ( n362556 , n362555 );
xor ( n14881 , n362449 , n362556 );
buf ( n362558 , n361958 );
buf ( n362559 , n361969 );
nand ( n14884 , n362558 , n362559 );
buf ( n362561 , n14884 );
buf ( n362562 , n362561 );
not ( n14887 , n362562 );
buf ( n362564 , n361903 );
not ( n14889 , n362564 );
or ( n14890 , n14887 , n14889 );
buf ( n362567 , n361961 );
buf ( n362568 , n361966 );
nand ( n14893 , n362567 , n362568 );
buf ( n362570 , n14893 );
buf ( n362571 , n362570 );
nand ( n14896 , n14890 , n362571 );
buf ( n362573 , n14896 );
buf ( n362574 , n362573 );
xor ( n14899 , n14881 , n362574 );
buf ( n362576 , n14899 );
buf ( n362577 , n362576 );
not ( n14902 , n362577 );
buf ( n362579 , n14902 );
and ( n14904 , n362443 , n362579 );
not ( n14905 , n362443 );
and ( n14906 , n14905 , n362576 );
nor ( n14907 , n14904 , n14906 );
not ( n14908 , n14907 );
not ( n14909 , n14908 );
or ( n14910 , n14762 , n14909 );
nand ( n14911 , n14907 , n14760 );
nand ( n14912 , n14910 , n14911 );
buf ( n362589 , n14912 );
xor ( n14914 , n361982 , n361987 );
and ( n14915 , n14914 , n362121 );
and ( n14916 , n361982 , n361987 );
or ( n14917 , n14915 , n14916 );
buf ( n362594 , n14917 );
buf ( n362595 , n362594 );
nor ( n14920 , n362589 , n362595 );
buf ( n362597 , n14920 );
buf ( n362598 , n362597 );
not ( n14923 , n362598 );
buf ( n362600 , n14923 );
buf ( n362601 , n362600 );
buf ( n362602 , n14912 );
buf ( n362603 , n362594 );
nand ( n14928 , n362602 , n362603 );
buf ( n362605 , n14928 );
buf ( n362606 , n362605 );
nand ( n14931 , n362601 , n362606 );
buf ( n362608 , n14931 );
not ( n14933 , n362608 );
buf ( n362610 , n355792 );
not ( n14935 , n362610 );
buf ( n362612 , n14935 );
not ( n14937 , n362612 );
buf ( n362614 , n361251 );
buf ( n362615 , n13892 );
buf ( n362616 , n362126 );
nor ( n14941 , n362615 , n362616 );
buf ( n362618 , n14941 );
buf ( n362619 , n362618 );
and ( n14944 , n362614 , n362619 );
buf ( n362621 , n14944 );
nand ( n14946 , n362621 , n360706 );
not ( n14947 , n14946 );
not ( n14948 , n14947 );
or ( n14949 , n14937 , n14948 );
not ( n14950 , n13049 );
not ( n14951 , n362621 );
or ( n14952 , n14950 , n14951 );
and ( n14953 , n13896 , n362134 );
not ( n14954 , n14953 );
not ( n14955 , n14150 );
or ( n14956 , n14954 , n14955 );
buf ( n362633 , n362129 );
not ( n14958 , n362633 );
buf ( n362635 , n14958 );
nand ( n14960 , n14956 , n362635 );
nand ( n14961 , n14952 , n14960 );
not ( n14962 , n14961 );
nand ( n14963 , n14949 , n14962 );
not ( n14964 , n14963 );
not ( n14965 , n14964 );
or ( n14966 , n14933 , n14965 );
buf ( n362643 , n362608 );
not ( n14968 , n362643 );
buf ( n362645 , n14968 );
not ( n14970 , n362645 );
or ( n14971 , n14970 , n14964 );
nand ( n14972 , n14966 , n14971 );
nand ( n14973 , n14628 , n14972 );
not ( n14974 , n13053 );
not ( n14975 , n361254 );
buf ( n362652 , n362618 );
buf ( n362653 , n362600 );
nand ( n14978 , n362652 , n362653 );
buf ( n362655 , n14978 );
nor ( n14980 , n14975 , n362655 );
not ( n14981 , n14980 );
or ( n14982 , n14974 , n14981 );
not ( n14983 , n362655 );
not ( n14984 , n361266 );
and ( n14985 , n14983 , n14984 );
not ( n14986 , n362134 );
nor ( n14987 , n362129 , n13896 );
nor ( n14988 , n14986 , n14987 );
buf ( n362665 , n14988 );
buf ( n362666 , n362597 );
or ( n14991 , n362665 , n362666 );
buf ( n362668 , n362605 );
nand ( n14993 , n14991 , n362668 );
buf ( n362670 , n14993 );
nor ( n14995 , n14985 , n362670 );
nand ( n14996 , n14982 , n14995 );
buf ( n362673 , n14761 );
buf ( n362674 , n362579 );
nand ( n14999 , n362673 , n362674 );
buf ( n362676 , n14999 );
buf ( n362677 , n362676 );
buf ( n15002 , n362443 );
buf ( n362679 , n15002 );
and ( n15004 , n362677 , n362679 );
buf ( n362681 , n14761 );
buf ( n362682 , n362579 );
nor ( n15007 , n362681 , n362682 );
buf ( n362684 , n15007 );
buf ( n362685 , n362684 );
nor ( n15010 , n15004 , n362685 );
buf ( n362687 , n15010 );
buf ( n362688 , n362687 );
not ( n15013 , n362688 );
buf ( n362690 , n15013 );
buf ( n362691 , n362690 );
xor ( n15016 , n362449 , n362556 );
and ( n15017 , n15016 , n362574 );
and ( n15018 , n362449 , n362556 );
or ( n15019 , n15017 , n15018 );
buf ( n362696 , n15019 );
buf ( n362697 , n362696 );
xor ( n15022 , n362370 , n362393 );
and ( n15023 , n15022 , n362401 );
and ( n15024 , n362370 , n362393 );
or ( n15025 , n15023 , n15024 );
buf ( n362702 , n15025 );
buf ( n362703 , n362702 );
xor ( n15028 , n362319 , n14651 );
and ( n15029 , n15028 , n362344 );
and ( n15030 , n362319 , n14651 );
or ( n15031 , n15029 , n15030 );
not ( n15032 , n15031 );
buf ( n362709 , n550 );
buf ( n362710 , n576 );
and ( n15035 , n362709 , n362710 );
buf ( n362712 , n15035 );
buf ( n362713 , n362712 );
buf ( n362714 , n362389 );
xor ( n15039 , n362713 , n362714 );
buf ( n362716 , n362363 );
not ( n15041 , n362716 );
buf ( n362718 , n361131 );
not ( n15043 , n362718 );
or ( n15044 , n15041 , n15043 );
buf ( n362721 , n354788 );
buf ( n362722 , n546 );
buf ( n362723 , n578 );
xor ( n15048 , n362722 , n362723 );
buf ( n362725 , n15048 );
buf ( n362726 , n362725 );
nand ( n15051 , n362721 , n362726 );
buf ( n362728 , n15051 );
buf ( n362729 , n362728 );
nand ( n15054 , n15044 , n362729 );
buf ( n362731 , n15054 );
buf ( n362732 , n362731 );
xor ( n15057 , n15039 , n362732 );
buf ( n362734 , n15057 );
not ( n15059 , n362734 );
and ( n15060 , n15032 , n15059 );
not ( n15061 , n15032 );
not ( n15062 , n15059 );
and ( n15063 , n15061 , n15062 );
nor ( n15064 , n15060 , n15063 );
buf ( n362741 , n350705 );
not ( n15066 , n362741 );
buf ( n362743 , n15066 );
buf ( n362744 , n362743 );
not ( n15069 , n362744 );
buf ( n362746 , n3009 );
not ( n15071 , n362746 );
or ( n15072 , n15069 , n15071 );
buf ( n362749 , n582 );
nand ( n15074 , n15072 , n362749 );
buf ( n362751 , n15074 );
buf ( n362752 , n362338 );
not ( n15077 , n362752 );
buf ( n362754 , n361110 );
not ( n15079 , n362754 );
or ( n15080 , n15077 , n15079 );
buf ( n362757 , n356446 );
buf ( n362758 , n548 );
buf ( n362759 , n576 );
xor ( n15084 , n362758 , n362759 );
buf ( n362761 , n15084 );
buf ( n362762 , n362761 );
nand ( n15087 , n362757 , n362762 );
buf ( n362764 , n15087 );
buf ( n362765 , n362764 );
nand ( n15090 , n15080 , n362765 );
buf ( n362767 , n15090 );
not ( n15092 , n362767 );
and ( n15093 , n362751 , n15092 );
not ( n15094 , n362751 );
not ( n15095 , n15092 );
and ( n15096 , n15094 , n15095 );
or ( n15097 , n15093 , n15096 );
buf ( n362774 , n362383 );
not ( n15099 , n362774 );
buf ( n362776 , n362375 );
not ( n15101 , n362776 );
or ( n15102 , n15099 , n15101 );
buf ( n362779 , n351559 );
buf ( n362780 , n544 );
buf ( n362781 , n580 );
xor ( n15106 , n362780 , n362781 );
buf ( n362783 , n15106 );
buf ( n362784 , n362783 );
nand ( n15109 , n362779 , n362784 );
buf ( n362786 , n15109 );
buf ( n362787 , n362786 );
nand ( n15112 , n15102 , n362787 );
buf ( n362789 , n15112 );
not ( n15114 , n362789 );
not ( n15115 , n15114 );
xor ( n15116 , n15097 , n15115 );
and ( n15117 , n15064 , n15116 );
not ( n15118 , n15064 );
not ( n15119 , n15116 );
and ( n15120 , n15118 , n15119 );
nor ( n15121 , n15117 , n15120 );
buf ( n362798 , n15121 );
xor ( n15123 , n362703 , n362798 );
xor ( n15124 , n362346 , n362352 );
and ( n15125 , n15124 , n362404 );
and ( n15126 , n362346 , n362352 );
or ( n15127 , n15125 , n15126 );
buf ( n362804 , n15127 );
buf ( n362805 , n362804 );
xor ( n15130 , n15123 , n362805 );
buf ( n362807 , n15130 );
buf ( n362808 , n362807 );
xor ( n15133 , n362315 , n362407 );
and ( n15134 , n15133 , n362414 );
and ( n15135 , n362315 , n362407 );
or ( n15136 , n15134 , n15135 );
buf ( n362813 , n15136 );
buf ( n362814 , n362813 );
xor ( n15139 , n362808 , n362814 );
xor ( n15140 , n362523 , n362543 );
and ( n15141 , n15140 , n362550 );
and ( n15142 , n362523 , n362543 );
or ( n15143 , n15141 , n15142 );
buf ( n362820 , n15143 );
buf ( n362821 , n362820 );
xor ( n15146 , n362454 , n362471 );
and ( n15147 , n15146 , n362485 );
and ( n15148 , n362454 , n362471 );
or ( n15149 , n15147 , n15148 );
buf ( n362826 , n15149 );
buf ( n362827 , n362826 );
buf ( n362828 , n550 );
buf ( n362829 , n560 );
and ( n15154 , n362828 , n362829 );
buf ( n362831 , n15154 );
buf ( n362832 , n362831 );
buf ( n362833 , n362539 );
xor ( n15158 , n362832 , n362833 );
buf ( n362835 , n362516 );
not ( n15160 , n362835 );
buf ( n362837 , n8604 );
not ( n15162 , n362837 );
or ( n15163 , n15160 , n15162 );
buf ( n362840 , n352295 );
buf ( n362841 , n546 );
buf ( n362842 , n562 );
xor ( n15167 , n362841 , n362842 );
buf ( n362844 , n15167 );
buf ( n362845 , n362844 );
nand ( n15170 , n362840 , n362845 );
buf ( n362847 , n15170 );
buf ( n362848 , n362847 );
nand ( n15173 , n15163 , n362848 );
buf ( n362850 , n15173 );
buf ( n362851 , n362850 );
xor ( n15176 , n15158 , n362851 );
buf ( n362853 , n15176 );
buf ( n362854 , n362853 );
xor ( n15179 , n362827 , n362854 );
buf ( n362856 , n362464 );
not ( n15181 , n362856 );
buf ( n362858 , n9186 );
not ( n15183 , n362858 );
or ( n15184 , n15181 , n15183 );
buf ( n362861 , n5407 );
buf ( n362862 , n548 );
buf ( n362863 , n560 );
xor ( n15188 , n362862 , n362863 );
buf ( n362865 , n15188 );
buf ( n362866 , n362865 );
nand ( n15191 , n362861 , n362866 );
buf ( n362868 , n15191 );
buf ( n362869 , n362868 );
nand ( n15194 , n15184 , n362869 );
buf ( n362871 , n15194 );
buf ( n362872 , n362871 );
buf ( n362873 , n362533 );
not ( n15198 , n362873 );
buf ( n362875 , n360913 );
not ( n15200 , n362875 );
or ( n15201 , n15198 , n15200 );
buf ( n362878 , n3650 );
xor ( n15203 , n564 , n544 );
buf ( n362880 , n15203 );
nand ( n15205 , n362878 , n362880 );
buf ( n362882 , n15205 );
buf ( n362883 , n362882 );
nand ( n15208 , n15201 , n362883 );
buf ( n362885 , n15208 );
buf ( n362886 , n362885 );
xor ( n15211 , n362872 , n362886 );
buf ( n362888 , n2550 );
buf ( n362889 , n360420 );
or ( n15214 , n362888 , n362889 );
buf ( n362891 , n566 );
nand ( n15216 , n15214 , n362891 );
buf ( n362893 , n15216 );
buf ( n362894 , n362893 );
xor ( n15219 , n15211 , n362894 );
buf ( n362896 , n15219 );
buf ( n362897 , n362896 );
xor ( n15222 , n15179 , n362897 );
buf ( n362899 , n15222 );
buf ( n362900 , n362899 );
xor ( n15225 , n362821 , n362900 );
xor ( n15226 , n362488 , n362505 );
and ( n15227 , n15226 , n362553 );
and ( n15228 , n362488 , n362505 );
or ( n15229 , n15227 , n15228 );
buf ( n362906 , n15229 );
buf ( n362907 , n362906 );
xor ( n15232 , n15225 , n362907 );
buf ( n362909 , n15232 );
buf ( n362910 , n362909 );
xor ( n15235 , n15139 , n362910 );
buf ( n362912 , n15235 );
buf ( n362913 , n362912 );
xor ( n15238 , n362697 , n362913 );
buf ( n362915 , n362431 );
not ( n15240 , n362915 );
buf ( n362917 , n362309 );
not ( n15242 , n362917 );
or ( n15243 , n15240 , n15242 );
buf ( n362920 , n362309 );
buf ( n362921 , n362431 );
or ( n15246 , n362920 , n362921 );
buf ( n362923 , n362416 );
nand ( n15248 , n15246 , n362923 );
buf ( n362925 , n15248 );
buf ( n362926 , n362925 );
nand ( n15251 , n15243 , n362926 );
buf ( n362928 , n15251 );
buf ( n362929 , n362928 );
xor ( n15254 , n15238 , n362929 );
buf ( n362931 , n15254 );
buf ( n362932 , n362931 );
nor ( n15257 , n362691 , n362932 );
buf ( n362934 , n15257 );
not ( n15259 , n362934 );
buf ( n362936 , n362931 );
buf ( n362937 , n362690 );
nand ( n15262 , n362936 , n362937 );
buf ( n362939 , n15262 );
nand ( n15264 , n15259 , n362939 );
and ( n15265 , n14996 , n15264 );
not ( n15266 , n14996 );
not ( n15267 , n15264 );
and ( n15268 , n15266 , n15267 );
nor ( n15269 , n15265 , n15268 );
nand ( n15270 , n14613 , n14607 );
not ( n15271 , n15270 );
nand ( n15272 , n13922 , n15271 );
not ( n15273 , n15272 );
not ( n15274 , n14532 );
nand ( n15275 , n15274 , n14606 );
not ( n15276 , n15275 );
not ( n15277 , n14620 );
or ( n15278 , n15276 , n15277 );
nand ( n15279 , n15278 , n14608 );
not ( n15280 , n15279 );
buf ( n15281 , n15280 );
not ( n15282 , n15281 );
or ( n15283 , n15273 , n15282 );
and ( n15284 , n544 , n5720 );
not ( n15285 , n5757 );
not ( n15286 , n546 );
buf ( n15287 , n6035 );
not ( n15288 , n15287 );
or ( n15289 , n15286 , n15288 );
not ( n15290 , n15287 );
nand ( n15291 , n15290 , n5761 );
nand ( n15292 , n15289 , n15291 );
not ( n15293 , n15292 );
or ( n15294 , n15285 , n15293 );
nand ( n15295 , n14565 , n8381 );
nand ( n15296 , n15294 , n15295 );
xor ( n15297 , n15284 , n15296 );
xor ( n15298 , n14567 , n14573 );
and ( n15299 , n15298 , n14585 );
and ( n15300 , n14567 , n14573 );
or ( n15301 , n15299 , n15300 );
xor ( n15302 , n15297 , n15301 );
xor ( n15303 , n14541 , n14543 );
and ( n15304 , n15303 , n14556 );
and ( n15305 , n14541 , n14543 );
or ( n15306 , n15304 , n15305 );
not ( n15307 , n8133 );
not ( n15308 , n548 );
not ( n15309 , n14088 );
or ( n15310 , n15308 , n15309 );
nand ( n15311 , n14087 , n351773 );
nand ( n15312 , n15310 , n15311 );
not ( n15313 , n15312 );
or ( n15314 , n15307 , n15313 );
nand ( n15315 , n14583 , n5751 );
nand ( n15316 , n15314 , n15315 );
not ( n15317 , n14554 );
not ( n15318 , n15317 );
not ( n15319 , n4078 );
not ( n15320 , n15319 );
and ( n15321 , n15318 , n15320 );
and ( n15322 , n1875 , n550 );
nor ( n15323 , n15321 , n15322 );
xor ( n15324 , n15316 , n15323 );
not ( n15325 , n8215 );
xor ( n15326 , n544 , n353641 );
not ( n15327 , n15326 );
or ( n15328 , n15325 , n15327 );
nand ( n15329 , n14571 , n8223 );
nand ( n15330 , n15328 , n15329 );
xor ( n15331 , n15324 , n15330 );
xor ( n15332 , n15306 , n15331 );
xor ( n15333 , n14588 , n14592 );
and ( n15334 , n15333 , n14597 );
and ( n15335 , n14588 , n14592 );
or ( n15336 , n15334 , n15335 );
xor ( n15337 , n15332 , n15336 );
xor ( n15338 , n15302 , n15337 );
xor ( n15339 , n14557 , n14586 );
and ( n15340 , n15339 , n14598 );
and ( n15341 , n14557 , n14586 );
or ( n15342 , n15340 , n15341 );
xor ( n15343 , n15338 , n15342 );
xor ( n15344 , n14537 , n14599 );
and ( n15345 , n15344 , n14604 );
and ( n15346 , n14537 , n14599 );
or ( n15347 , n15345 , n15346 );
xor ( n15348 , n15343 , n15347 );
nand ( n15349 , n15283 , n15348 );
nor ( n15350 , n15347 , n15343 );
not ( n15351 , n15350 );
nand ( n15352 , n15347 , n15343 );
nand ( n15353 , n15351 , n15352 );
nand ( n15354 , n15272 , n15281 , n15353 );
nand ( n15355 , n15269 , n15349 , n15354 );
and ( n15356 , n14973 , n15355 );
xor ( n15357 , n362821 , n362900 );
and ( n15358 , n15357 , n362907 );
and ( n15359 , n362821 , n362900 );
or ( n15360 , n15358 , n15359 );
buf ( n363037 , n15360 );
buf ( n363038 , n363037 );
xor ( n15363 , n362808 , n362814 );
and ( n15364 , n15363 , n362910 );
and ( n15365 , n362808 , n362814 );
or ( n15366 , n15364 , n15365 );
buf ( n363043 , n15366 );
buf ( n363044 , n363043 );
xor ( n15369 , n363038 , n363044 );
xor ( n15370 , n362832 , n362833 );
and ( n15371 , n15370 , n362851 );
and ( n15372 , n362832 , n362833 );
or ( n15373 , n15371 , n15372 );
buf ( n363050 , n15373 );
buf ( n363051 , n363050 );
buf ( n363052 , n15203 );
not ( n15377 , n363052 );
buf ( n363054 , n360913 );
not ( n15379 , n363054 );
or ( n15380 , n15377 , n15379 );
buf ( n363057 , n3650 );
buf ( n363058 , n564 );
nand ( n15383 , n363057 , n363058 );
buf ( n363060 , n15383 );
buf ( n363061 , n363060 );
nand ( n15386 , n15380 , n363061 );
buf ( n363063 , n15386 );
buf ( n363064 , n363063 );
not ( n15389 , n363064 );
buf ( n363066 , n15389 );
buf ( n363067 , n363066 );
xor ( n15392 , n362872 , n362886 );
and ( n15393 , n15392 , n362894 );
and ( n15394 , n362872 , n362886 );
or ( n15395 , n15393 , n15394 );
buf ( n363072 , n15395 );
buf ( n363073 , n363072 );
xor ( n15398 , n363067 , n363073 );
buf ( n363075 , n549 );
buf ( n363076 , n560 );
and ( n15401 , n363075 , n363076 );
buf ( n363078 , n15401 );
buf ( n363079 , n363078 );
buf ( n363080 , n362865 );
not ( n15405 , n363080 );
buf ( n363082 , n9186 );
not ( n15407 , n363082 );
or ( n15408 , n15405 , n15407 );
buf ( n363085 , n5407 );
xor ( n15410 , n560 , n547 );
buf ( n363087 , n15410 );
nand ( n15412 , n363085 , n363087 );
buf ( n363089 , n15412 );
buf ( n363090 , n363089 );
nand ( n15415 , n15408 , n363090 );
buf ( n363092 , n15415 );
buf ( n363093 , n363092 );
xor ( n15418 , n363079 , n363093 );
buf ( n363095 , n362844 );
not ( n15420 , n363095 );
buf ( n363097 , n8604 );
not ( n15422 , n363097 );
or ( n15423 , n15420 , n15422 );
buf ( n363100 , n352295 );
buf ( n363101 , n545 );
buf ( n363102 , n562 );
xor ( n15427 , n363101 , n363102 );
buf ( n363104 , n15427 );
buf ( n363105 , n363104 );
nand ( n15430 , n363100 , n363105 );
buf ( n363107 , n15430 );
buf ( n363108 , n363107 );
nand ( n15433 , n15423 , n363108 );
buf ( n363110 , n15433 );
buf ( n363111 , n363110 );
xor ( n15436 , n15418 , n363111 );
buf ( n363113 , n15436 );
buf ( n363114 , n363113 );
xor ( n15439 , n15398 , n363114 );
buf ( n363116 , n15439 );
buf ( n363117 , n363116 );
xor ( n15442 , n363051 , n363117 );
xor ( n15443 , n362827 , n362854 );
and ( n15444 , n15443 , n362897 );
and ( n15445 , n362827 , n362854 );
or ( n15446 , n15444 , n15445 );
buf ( n363123 , n15446 );
buf ( n363124 , n363123 );
xor ( n15449 , n15442 , n363124 );
buf ( n363126 , n15449 );
buf ( n363127 , n363126 );
xor ( n15452 , n362713 , n362714 );
and ( n15453 , n15452 , n362732 );
and ( n15454 , n362713 , n362714 );
or ( n15455 , n15453 , n15454 );
buf ( n363132 , n15455 );
not ( n15457 , n15032 );
not ( n15458 , n15059 );
or ( n15459 , n15457 , n15458 );
nand ( n15460 , n15459 , n15116 );
not ( n15461 , n15032 );
nand ( n15462 , n15461 , n15062 );
nand ( n15463 , n15460 , n15462 );
xor ( n15464 , n363132 , n15463 );
not ( n15465 , n362783 );
not ( n15466 , n362375 );
or ( n15467 , n15465 , n15466 );
buf ( n363144 , n351559 );
buf ( n363145 , n580 );
nand ( n15470 , n363144 , n363145 );
buf ( n363147 , n15470 );
nand ( n15472 , n15467 , n363147 );
not ( n15473 , n15472 );
not ( n15474 , n15114 );
nand ( n15475 , n15474 , n15095 );
not ( n15476 , n15092 );
not ( n15477 , n15114 );
or ( n15478 , n15476 , n15477 );
nand ( n15479 , n15478 , n362751 );
nand ( n15480 , n15475 , n15479 );
xor ( n15481 , n15473 , n15480 );
buf ( n363158 , n549 );
buf ( n363159 , n576 );
and ( n15484 , n363158 , n363159 );
buf ( n363161 , n15484 );
buf ( n363162 , n362725 );
not ( n15487 , n363162 );
buf ( n363164 , n361131 );
not ( n15489 , n363164 );
or ( n15490 , n15487 , n15489 );
buf ( n363167 , n354788 );
buf ( n363168 , n545 );
buf ( n363169 , n578 );
xor ( n15494 , n363168 , n363169 );
buf ( n363171 , n15494 );
buf ( n363172 , n363171 );
nand ( n15497 , n363167 , n363172 );
buf ( n363174 , n15497 );
buf ( n363175 , n363174 );
nand ( n15500 , n15490 , n363175 );
buf ( n363177 , n15500 );
xor ( n15502 , n363161 , n363177 );
buf ( n363179 , n362761 );
not ( n15504 , n363179 );
buf ( n363181 , n361110 );
not ( n15506 , n363181 );
or ( n15507 , n15504 , n15506 );
buf ( n363184 , n356446 );
buf ( n363185 , n576 );
buf ( n363186 , n547 );
xor ( n15511 , n363185 , n363186 );
buf ( n363188 , n15511 );
buf ( n363189 , n363188 );
nand ( n15514 , n363184 , n363189 );
buf ( n363191 , n15514 );
buf ( n363192 , n363191 );
nand ( n15517 , n15507 , n363192 );
buf ( n363194 , n15517 );
xor ( n15519 , n15502 , n363194 );
xor ( n15520 , n15481 , n15519 );
xor ( n15521 , n15464 , n15520 );
buf ( n363198 , n15521 );
xor ( n15523 , n363127 , n363198 );
xor ( n15524 , n362703 , n362798 );
and ( n15525 , n15524 , n362805 );
and ( n15526 , n362703 , n362798 );
or ( n15527 , n15525 , n15526 );
buf ( n363204 , n15527 );
buf ( n363205 , n363204 );
xor ( n15530 , n15523 , n363205 );
buf ( n363207 , n15530 );
buf ( n363208 , n363207 );
xor ( n15533 , n15369 , n363208 );
buf ( n363210 , n15533 );
buf ( n363211 , n363210 );
xor ( n15536 , n362697 , n362913 );
and ( n15537 , n15536 , n362929 );
and ( n15538 , n362697 , n362913 );
or ( n15539 , n15537 , n15538 );
buf ( n363216 , n15539 );
buf ( n363217 , n363216 );
and ( n15542 , n363211 , n363217 );
buf ( n363219 , n15542 );
buf ( n363220 , n363219 );
not ( n15545 , n363220 );
buf ( n363222 , n15545 );
buf ( n363223 , n363216 );
buf ( n363224 , n363210 );
nor ( n15549 , n363223 , n363224 );
buf ( n363226 , n15549 );
buf ( n363227 , n363226 );
not ( n15552 , n363227 );
buf ( n363229 , n15552 );
nand ( n15554 , n363222 , n363229 );
not ( n15555 , n15554 );
buf ( n15556 , n362621 );
buf ( n363233 , n362597 );
buf ( n363234 , n362934 );
nor ( n15559 , n363233 , n363234 );
buf ( n363236 , n15559 );
buf ( n363237 , n363236 );
buf ( n15562 , n363237 );
buf ( n363239 , n15562 );
nand ( n15564 , n362612 , n360706 , n15556 , n363239 );
nand ( n15565 , n14961 , n363239 );
buf ( n363242 , n362934 );
buf ( n363243 , n362605 );
or ( n15568 , n363242 , n363243 );
buf ( n363245 , n362939 );
nand ( n15570 , n15568 , n363245 );
buf ( n363247 , n15570 );
buf ( n15572 , n363247 );
not ( n15573 , n15572 );
nand ( n15574 , n15564 , n15565 , n15573 );
not ( n15575 , n15574 );
or ( n15576 , n15555 , n15575 );
nor ( n15577 , n15572 , n15554 );
nand ( n15578 , n15565 , n15577 , n15564 );
nand ( n15579 , n15576 , n15578 );
not ( n15580 , n15579 );
not ( n15581 , n15580 );
or ( n15582 , n15347 , n15343 );
not ( n15583 , n15582 );
not ( n15584 , n15279 );
or ( n15585 , n15583 , n15584 );
nand ( n15586 , n15585 , n15352 );
not ( n15587 , n15586 );
not ( n15588 , n13920 );
nand ( n15589 , n9005 , n13907 );
not ( n15590 , n15589 );
or ( n15591 , n15588 , n15590 );
nor ( n15592 , n15270 , n15350 );
nand ( n15593 , n15591 , n15592 );
nand ( n15594 , n15587 , n15593 );
buf ( n15595 , n15594 );
xor ( n15596 , n15302 , n15337 );
and ( n15597 , n15596 , n15342 );
and ( n15598 , n15302 , n15337 );
or ( n15599 , n15597 , n15598 );
xor ( n15600 , n15284 , n15296 );
and ( n15601 , n15600 , n15301 );
and ( n15602 , n15284 , n15296 );
or ( n15603 , n15601 , n15602 );
xor ( n15604 , n15316 , n15323 );
and ( n15605 , n15604 , n15330 );
and ( n15606 , n15316 , n15323 );
or ( n15607 , n15605 , n15606 );
not ( n15608 , n8411 );
not ( n15609 , n15319 );
or ( n15610 , n15608 , n15609 );
nand ( n15611 , n15610 , n550 );
not ( n15612 , n5751 );
not ( n15613 , n15312 );
or ( n15614 , n15612 , n15613 );
not ( n15615 , n548 );
not ( n15616 , n14552 );
or ( n15617 , n15615 , n15616 );
nand ( n15618 , n14549 , n351773 );
nand ( n15619 , n15617 , n15618 );
nand ( n15620 , n15619 , n8133 );
nand ( n15621 , n15614 , n15620 );
xor ( n15622 , n15611 , n15621 );
not ( n15623 , n8223 );
not ( n15624 , n15326 );
or ( n15625 , n15623 , n15624 );
buf ( n15626 , n353618 );
xor ( n15627 , n544 , n15626 );
nand ( n15628 , n15627 , n8215 );
nand ( n15629 , n15625 , n15628 );
xor ( n15630 , n15622 , n15629 );
xor ( n15631 , n15607 , n15630 );
and ( n15632 , n544 , n5730 );
not ( n15633 , n8381 );
not ( n15634 , n15292 );
or ( n15635 , n15633 , n15634 );
not ( n15636 , n546 );
not ( n15637 , n6082 );
or ( n15638 , n15636 , n15637 );
nand ( n15639 , n14581 , n5761 );
nand ( n15640 , n15638 , n15639 );
nand ( n15641 , n15640 , n353673 );
nand ( n15642 , n15635 , n15641 );
xor ( n15643 , n15632 , n15642 );
not ( n15644 , n15323 );
xor ( n15645 , n15643 , n15644 );
xor ( n15646 , n15631 , n15645 );
xor ( n15647 , n15603 , n15646 );
xor ( n15648 , n15306 , n15331 );
and ( n15649 , n15648 , n15336 );
and ( n15650 , n15306 , n15331 );
or ( n15651 , n15649 , n15650 );
xor ( n15652 , n15647 , n15651 );
not ( n15653 , n15652 );
not ( n15654 , n15653 );
and ( n15655 , n15599 , n15654 );
not ( n15656 , n15599 );
and ( n15657 , n15656 , n15653 );
nor ( n15658 , n15655 , n15657 );
and ( n15659 , n15595 , n15658 );
not ( n15660 , n15595 );
not ( n15661 , n15658 );
and ( n15662 , n15660 , n15661 );
nor ( n15663 , n15659 , n15662 );
not ( n15664 , n15663 );
or ( n15665 , n15581 , n15664 );
not ( n15666 , n15599 );
nand ( n15667 , n15666 , n15653 );
not ( n15668 , n15667 );
not ( n15669 , n15594 );
or ( n15670 , n15668 , n15669 );
nand ( n15671 , n15599 , n15654 );
nand ( n15672 , n15670 , n15671 );
not ( n15673 , n15672 );
xor ( n15674 , n15603 , n15646 );
and ( n15675 , n15674 , n15651 );
and ( n15676 , n15603 , n15646 );
or ( n15677 , n15675 , n15676 );
not ( n15678 , n15677 );
not ( n15679 , n15678 );
and ( n15680 , n544 , n353641 );
not ( n15681 , n5757 );
not ( n15682 , n546 );
not ( n15683 , n14088 );
or ( n15684 , n15682 , n15683 );
nand ( n15685 , n14087 , n5761 );
nand ( n15686 , n15684 , n15685 );
not ( n15687 , n15686 );
or ( n15688 , n15681 , n15687 );
nand ( n15689 , n15640 , n8381 );
nand ( n15690 , n15688 , n15689 );
xor ( n15691 , n15680 , n15690 );
and ( n15692 , n15619 , n5751 );
not ( n15693 , n8133 );
nor ( n15694 , n15693 , n351773 );
nor ( n15695 , n15692 , n15694 );
xor ( n15696 , n15691 , n15695 );
not ( n15697 , n8215 );
xor ( n15698 , n544 , n15290 );
not ( n15699 , n15698 );
or ( n15700 , n15697 , n15699 );
nand ( n15701 , n15627 , n8223 );
nand ( n15702 , n15700 , n15701 );
xor ( n15703 , n15632 , n15642 );
and ( n15704 , n15703 , n15644 );
and ( n15705 , n15632 , n15642 );
or ( n15706 , n15704 , n15705 );
xor ( n15707 , n15702 , n15706 );
xor ( n15708 , n15611 , n15621 );
and ( n15709 , n15708 , n15629 );
and ( n15710 , n15611 , n15621 );
or ( n15711 , n15709 , n15710 );
xor ( n15712 , n15707 , n15711 );
xor ( n15713 , n15696 , n15712 );
xor ( n15714 , n15607 , n15630 );
and ( n15715 , n15714 , n15645 );
and ( n15716 , n15607 , n15630 );
or ( n15717 , n15715 , n15716 );
xor ( n15718 , n15713 , n15717 );
not ( n15719 , n15718 );
not ( n15720 , n15719 );
or ( n15721 , n15679 , n15720 );
nand ( n15722 , n15677 , n15718 );
nand ( n15723 , n15721 , n15722 );
nand ( n15724 , n15673 , n15723 );
xor ( n15725 , n363038 , n363044 );
and ( n15726 , n15725 , n363208 );
and ( n15727 , n363038 , n363044 );
or ( n15728 , n15726 , n15727 );
buf ( n363405 , n15728 );
buf ( n363406 , n363405 );
xor ( n15731 , n363051 , n363117 );
and ( n15732 , n15731 , n363124 );
and ( n15733 , n363051 , n363117 );
or ( n15734 , n15732 , n15733 );
buf ( n363411 , n15734 );
buf ( n363412 , n363411 );
buf ( n363413 , n548 );
buf ( n363414 , n560 );
and ( n15739 , n363413 , n363414 );
buf ( n363416 , n15739 );
buf ( n363417 , n363416 );
buf ( n363418 , n363104 );
not ( n15743 , n363418 );
buf ( n363420 , n8604 );
not ( n15745 , n363420 );
or ( n15746 , n15743 , n15745 );
buf ( n363423 , n352295 );
and ( n15748 , n562 , n544 );
not ( n15749 , n562 );
and ( n15750 , n15749 , n7283 );
nor ( n15751 , n15748 , n15750 );
buf ( n363428 , n15751 );
nand ( n15753 , n363423 , n363428 );
buf ( n363430 , n15753 );
buf ( n363431 , n363430 );
nand ( n15756 , n15746 , n363431 );
buf ( n363433 , n15756 );
buf ( n363434 , n363433 );
xor ( n15759 , n363417 , n363434 );
buf ( n363436 , n3650 );
buf ( n363437 , n360913 );
or ( n15762 , n363436 , n363437 );
buf ( n363439 , n564 );
nand ( n15764 , n15762 , n363439 );
buf ( n363441 , n15764 );
buf ( n363442 , n363441 );
xor ( n15767 , n15759 , n363442 );
buf ( n363444 , n15767 );
buf ( n363445 , n363444 );
buf ( n363446 , n363063 );
buf ( n363447 , n15410 );
not ( n15772 , n363447 );
buf ( n363449 , n9186 );
not ( n15774 , n363449 );
or ( n15775 , n15772 , n15774 );
buf ( n363452 , n5407 );
buf ( n363453 , n560 );
buf ( n363454 , n546 );
xor ( n15779 , n363453 , n363454 );
buf ( n363456 , n15779 );
buf ( n363457 , n363456 );
nand ( n15782 , n363452 , n363457 );
buf ( n363459 , n15782 );
buf ( n363460 , n363459 );
nand ( n15785 , n15775 , n363460 );
buf ( n363462 , n15785 );
buf ( n363463 , n363462 );
xor ( n15788 , n363446 , n363463 );
xor ( n15789 , n363079 , n363093 );
and ( n15790 , n15789 , n363111 );
and ( n15791 , n363079 , n363093 );
or ( n15792 , n15790 , n15791 );
buf ( n363469 , n15792 );
buf ( n363470 , n363469 );
xor ( n15795 , n15788 , n363470 );
buf ( n363472 , n15795 );
buf ( n363473 , n363472 );
xor ( n15798 , n363445 , n363473 );
xor ( n15799 , n363067 , n363073 );
and ( n15800 , n15799 , n363114 );
and ( n15801 , n363067 , n363073 );
or ( n15802 , n15800 , n15801 );
buf ( n363479 , n15802 );
buf ( n363480 , n363479 );
xor ( n15805 , n15798 , n363480 );
buf ( n363482 , n15805 );
buf ( n363483 , n363482 );
or ( n15808 , n363161 , n363194 );
nand ( n15809 , n15808 , n363177 );
nand ( n15810 , n363194 , n363161 );
nand ( n15811 , n15809 , n15810 );
buf ( n363488 , n363188 );
not ( n15813 , n363488 );
buf ( n363490 , n361110 );
not ( n15815 , n363490 );
or ( n15816 , n15813 , n15815 );
buf ( n363493 , n356446 );
buf ( n363494 , n576 );
buf ( n363495 , n546 );
xor ( n15820 , n363494 , n363495 );
buf ( n363497 , n15820 );
buf ( n363498 , n363497 );
nand ( n15823 , n363493 , n363498 );
buf ( n363500 , n15823 );
buf ( n363501 , n363500 );
nand ( n15826 , n15816 , n363501 );
buf ( n363503 , n15826 );
and ( n15828 , n15472 , n363503 );
not ( n15829 , n15472 );
not ( n15830 , n363503 );
and ( n15831 , n15829 , n15830 );
nor ( n15832 , n15828 , n15831 );
xor ( n15833 , n15811 , n15832 );
xor ( n15834 , n15473 , n15480 );
and ( n15835 , n15834 , n15519 );
and ( n15836 , n15473 , n15480 );
or ( n15837 , n15835 , n15836 );
xor ( n15838 , n15833 , n15837 );
buf ( n363515 , n548 );
buf ( n363516 , n576 );
and ( n15841 , n363515 , n363516 );
buf ( n363518 , n15841 );
buf ( n363519 , n363518 );
buf ( n363520 , n363171 );
not ( n15845 , n363520 );
buf ( n363522 , n361131 );
not ( n15847 , n363522 );
or ( n15848 , n15845 , n15847 );
buf ( n363525 , n354788 );
buf ( n363526 , n544 );
buf ( n363527 , n578 );
xor ( n15852 , n363526 , n363527 );
buf ( n363529 , n15852 );
buf ( n363530 , n363529 );
nand ( n15855 , n363525 , n363530 );
buf ( n363532 , n15855 );
buf ( n363533 , n363532 );
nand ( n15858 , n15848 , n363533 );
buf ( n363535 , n15858 );
buf ( n363536 , n363535 );
xor ( n15861 , n363519 , n363536 );
buf ( n363538 , n351559 );
buf ( n363539 , n362375 );
or ( n15864 , n363538 , n363539 );
buf ( n363541 , n580 );
nand ( n15866 , n15864 , n363541 );
buf ( n363543 , n15866 );
buf ( n363544 , n363543 );
xor ( n15869 , n15861 , n363544 );
buf ( n363546 , n15869 );
xor ( n15871 , n15838 , n363546 );
buf ( n363548 , n15871 );
xor ( n15873 , n363483 , n363548 );
xor ( n15874 , n363132 , n15463 );
and ( n15875 , n15874 , n15520 );
and ( n15876 , n363132 , n15463 );
or ( n15877 , n15875 , n15876 );
buf ( n363554 , n15877 );
xor ( n15879 , n15873 , n363554 );
buf ( n363556 , n15879 );
buf ( n363557 , n363556 );
xor ( n15882 , n363412 , n363557 );
xor ( n15883 , n363127 , n363198 );
and ( n15884 , n15883 , n363205 );
and ( n15885 , n363127 , n363198 );
or ( n15886 , n15884 , n15885 );
buf ( n363563 , n15886 );
buf ( n363564 , n363563 );
xor ( n15889 , n15882 , n363564 );
buf ( n363566 , n15889 );
buf ( n363567 , n363566 );
and ( n15892 , n363406 , n363567 );
buf ( n363569 , n15892 );
buf ( n363570 , n363405 );
buf ( n363571 , n363566 );
nor ( n15896 , n363570 , n363571 );
buf ( n363573 , n15896 );
nor ( n15898 , n363569 , n363573 );
not ( n15899 , n15898 );
and ( n15900 , n363236 , n363229 );
nand ( n15901 , n14961 , n15900 );
nand ( n15902 , n14947 , n15900 , n362612 );
buf ( n363579 , n363229 );
not ( n15904 , n363579 );
buf ( n363581 , n363247 );
not ( n15906 , n363581 );
or ( n15907 , n15904 , n15906 );
buf ( n363584 , n363222 );
nand ( n15909 , n15907 , n363584 );
buf ( n363586 , n15909 );
not ( n15911 , n363586 );
nand ( n15912 , n15901 , n15902 , n15911 );
not ( n15913 , n15912 );
or ( n15914 , n15899 , n15913 );
not ( n15915 , n363569 );
buf ( n363592 , n363573 );
not ( n15917 , n363592 );
buf ( n363594 , n15917 );
nand ( n15919 , n15915 , n363594 );
nand ( n15920 , n15901 , n15902 , n15911 , n15919 );
nand ( n15921 , n15914 , n15920 );
not ( n15922 , n15723 );
nand ( n15923 , n15922 , n15672 );
nand ( n15924 , n15724 , n15921 , n15923 );
nand ( n15925 , n15665 , n15924 );
not ( n15926 , n15925 );
nand ( n15927 , n15356 , n15926 );
xor ( n15928 , n15696 , n15712 );
and ( n15929 , n15928 , n15717 );
and ( n15930 , n15696 , n15712 );
or ( n15931 , n15929 , n15930 );
or ( n15932 , n5751 , n8133 );
nand ( n15933 , n15932 , n548 );
not ( n15934 , n8381 );
not ( n15935 , n15686 );
or ( n15936 , n15934 , n15935 );
not ( n15937 , n5761 );
not ( n15938 , n14549 );
or ( n15939 , n15937 , n15938 );
nand ( n15940 , n14552 , n546 );
nand ( n15941 , n15939 , n15940 );
nand ( n15942 , n15941 , n353673 );
nand ( n15943 , n15936 , n15942 );
xor ( n15944 , n15933 , n15943 );
and ( n15945 , n544 , n15626 );
xor ( n15946 , n15944 , n15945 );
not ( n15947 , n15695 );
not ( n15948 , n8223 );
not ( n15949 , n15698 );
or ( n15950 , n15948 , n15949 );
xor ( n15951 , n544 , n14581 );
nand ( n15952 , n15951 , n8215 );
nand ( n15953 , n15950 , n15952 );
xor ( n15954 , n15947 , n15953 );
xor ( n15955 , n15680 , n15690 );
and ( n15956 , n15955 , n15695 );
and ( n15957 , n15680 , n15690 );
or ( n15958 , n15956 , n15957 );
xor ( n15959 , n15954 , n15958 );
xor ( n15960 , n15946 , n15959 );
xor ( n15961 , n15702 , n15706 );
and ( n15962 , n15961 , n15711 );
and ( n15963 , n15702 , n15706 );
or ( n15964 , n15962 , n15963 );
xor ( n15965 , n15960 , n15964 );
nor ( n15966 , n15931 , n15965 );
not ( n15967 , n15966 );
nand ( n15968 , n15931 , n15965 );
nand ( n15969 , n15967 , n15968 );
not ( n15970 , n15969 );
not ( n15971 , n15667 );
not ( n15972 , n15594 );
or ( n15973 , n15971 , n15972 );
nand ( n15974 , n15973 , n15671 );
nand ( n15975 , n15678 , n15719 );
nand ( n15976 , n15974 , n15975 );
buf ( n15977 , n15722 );
nand ( n15978 , n15976 , n15977 );
not ( n15979 , n15978 );
or ( n15980 , n15970 , n15979 );
not ( n15981 , n15977 );
nor ( n15982 , n15981 , n15969 );
nand ( n15983 , n15982 , n15976 );
nand ( n15984 , n15980 , n15983 );
not ( n15985 , n15984 );
buf ( n363662 , n363226 );
buf ( n363663 , n363573 );
nor ( n15988 , n363662 , n363663 );
buf ( n363665 , n15988 );
buf ( n363666 , n363665 );
not ( n15991 , n363666 );
buf ( n363668 , n363247 );
not ( n15993 , n363668 );
or ( n15994 , n15991 , n15993 );
buf ( n363671 , n363594 );
buf ( n363672 , n363219 );
and ( n15997 , n363671 , n363672 );
buf ( n363674 , n363569 );
nor ( n15999 , n15997 , n363674 );
buf ( n363676 , n15999 );
buf ( n363677 , n363676 );
nand ( n16002 , n15994 , n363677 );
buf ( n363679 , n16002 );
not ( n16004 , n363679 );
buf ( n363681 , n363236 );
buf ( n363682 , n363665 );
and ( n16007 , n363681 , n363682 );
buf ( n363684 , n16007 );
nand ( n16009 , n363684 , n14961 );
buf ( n363686 , n14947 );
buf ( n363687 , n362612 );
buf ( n16012 , n363687 );
buf ( n363689 , n16012 );
buf ( n363690 , n363689 );
buf ( n363691 , n363684 );
nand ( n16016 , n363686 , n363690 , n363691 );
buf ( n363693 , n16016 );
nand ( n16018 , n16004 , n16009 , n363693 );
xor ( n16019 , n363412 , n363557 );
and ( n16020 , n16019 , n363564 );
and ( n16021 , n363412 , n363557 );
or ( n16022 , n16020 , n16021 );
buf ( n363699 , n16022 );
buf ( n363700 , n363699 );
not ( n16025 , n363700 );
xor ( n16026 , n363445 , n363473 );
and ( n16027 , n16026 , n363480 );
and ( n16028 , n363445 , n363473 );
or ( n16029 , n16027 , n16028 );
buf ( n363706 , n16029 );
buf ( n363707 , n363706 );
xor ( n16032 , n363519 , n363536 );
and ( n16033 , n16032 , n363544 );
and ( n16034 , n363519 , n363536 );
or ( n16035 , n16033 , n16034 );
buf ( n363712 , n16035 );
buf ( n363713 , n363712 );
and ( n16038 , n363185 , n363186 );
buf ( n363715 , n16038 );
buf ( n363716 , n363715 );
buf ( n363717 , n363497 );
not ( n16042 , n363717 );
buf ( n363719 , n361110 );
not ( n16044 , n363719 );
or ( n16045 , n16042 , n16044 );
buf ( n363722 , n356446 );
buf ( n363723 , n545 );
buf ( n363724 , n576 );
xor ( n16049 , n363723 , n363724 );
buf ( n363726 , n16049 );
buf ( n363727 , n363726 );
nand ( n16052 , n363722 , n363727 );
buf ( n363729 , n16052 );
buf ( n363730 , n363729 );
nand ( n16055 , n16045 , n363730 );
buf ( n363732 , n16055 );
buf ( n363733 , n363732 );
xor ( n16058 , n363716 , n363733 );
buf ( n363735 , n363529 );
not ( n16060 , n363735 );
buf ( n363737 , n361131 );
not ( n16062 , n363737 );
or ( n16063 , n16060 , n16062 );
buf ( n363740 , n354788 );
buf ( n363741 , n578 );
nand ( n16066 , n363740 , n363741 );
buf ( n363743 , n16066 );
buf ( n363744 , n363743 );
nand ( n16069 , n16063 , n363744 );
buf ( n363746 , n16069 );
buf ( n363747 , n363746 );
not ( n16072 , n363747 );
buf ( n363749 , n16072 );
buf ( n363750 , n363749 );
xor ( n16075 , n16058 , n363750 );
buf ( n363752 , n16075 );
buf ( n363753 , n363752 );
xor ( n16078 , n363713 , n363753 );
not ( n16079 , n15473 );
not ( n16080 , n15830 );
or ( n16081 , n16079 , n16080 );
nand ( n16082 , n16081 , n15811 );
nand ( n16083 , n363503 , n15472 );
nand ( n16084 , n16082 , n16083 );
buf ( n363761 , n16084 );
xor ( n16086 , n16078 , n363761 );
buf ( n363763 , n16086 );
buf ( n363764 , n363763 );
xor ( n16089 , n363417 , n363434 );
and ( n16090 , n16089 , n363442 );
and ( n16091 , n363417 , n363434 );
or ( n16092 , n16090 , n16091 );
buf ( n363769 , n16092 );
buf ( n363770 , n363769 );
not ( n16095 , n363456 );
not ( n16096 , n9186 );
or ( n16097 , n16095 , n16096 );
buf ( n363774 , n5407 );
buf ( n363775 , n560 );
buf ( n363776 , n545 );
xor ( n16101 , n363775 , n363776 );
buf ( n363778 , n16101 );
buf ( n363779 , n363778 );
nand ( n16104 , n363774 , n363779 );
buf ( n363781 , n16104 );
nand ( n16106 , n16097 , n363781 );
nand ( n16107 , n560 , n547 );
not ( n16108 , n16107 );
and ( n16109 , n16106 , n16108 );
not ( n16110 , n16106 );
and ( n16111 , n16110 , n16107 );
nor ( n16112 , n16109 , n16111 );
not ( n16113 , n562 );
not ( n16114 , n352295 );
or ( n16115 , n16113 , n16114 );
nand ( n16116 , n8604 , n15751 );
nand ( n16117 , n16115 , n16116 );
and ( n16118 , n16112 , n16117 );
not ( n16119 , n16112 );
not ( n16120 , n16117 );
and ( n16121 , n16119 , n16120 );
or ( n16122 , n16118 , n16121 );
buf ( n363799 , n16122 );
xor ( n16124 , n363770 , n363799 );
xor ( n16125 , n363446 , n363463 );
and ( n16126 , n16125 , n363470 );
and ( n16127 , n363446 , n363463 );
or ( n16128 , n16126 , n16127 );
buf ( n363805 , n16128 );
buf ( n363806 , n363805 );
xor ( n16131 , n16124 , n363806 );
buf ( n363808 , n16131 );
buf ( n363809 , n363808 );
xor ( n16134 , n363764 , n363809 );
xor ( n16135 , n15833 , n15837 );
and ( n16136 , n16135 , n363546 );
and ( n16137 , n15833 , n15837 );
or ( n16138 , n16136 , n16137 );
buf ( n363815 , n16138 );
xor ( n16140 , n16134 , n363815 );
buf ( n363817 , n16140 );
buf ( n363818 , n363817 );
xor ( n16143 , n363707 , n363818 );
xor ( n16144 , n363483 , n363548 );
and ( n16145 , n16144 , n363554 );
and ( n16146 , n363483 , n363548 );
or ( n16147 , n16145 , n16146 );
buf ( n363824 , n16147 );
buf ( n363825 , n363824 );
xor ( n16150 , n16143 , n363825 );
buf ( n363827 , n16150 );
buf ( n363828 , n363827 );
not ( n16153 , n363828 );
buf ( n363830 , n16153 );
buf ( n363831 , n363830 );
nand ( n16156 , n16025 , n363831 );
buf ( n363833 , n16156 );
buf ( n363834 , n363830 );
not ( n16159 , n363834 );
buf ( n363836 , n363699 );
nand ( n16161 , n16159 , n363836 );
buf ( n363838 , n16161 );
nand ( n16163 , n363833 , n363838 );
xor ( n16164 , n16018 , n16163 );
not ( n16165 , n16164 );
or ( n16166 , n15985 , n16165 );
not ( n16167 , n15975 );
nor ( n16168 , n16167 , n15966 );
not ( n16169 , n16168 );
not ( n16170 , n15667 );
not ( n16171 , n15594 );
or ( n16172 , n16170 , n16171 );
not ( n16173 , n15653 );
nand ( n16174 , n16173 , n15599 );
nand ( n16175 , n16172 , n16174 );
not ( n16176 , n16175 );
or ( n16177 , n16169 , n16176 );
not ( n16178 , n15977 );
not ( n16179 , n15966 );
and ( n16180 , n16178 , n16179 );
and ( n16181 , n15931 , n15965 );
nor ( n16182 , n16180 , n16181 );
nand ( n16183 , n16177 , n16182 );
xor ( n16184 , n15933 , n15943 );
and ( n16185 , n16184 , n15945 );
and ( n16186 , n15933 , n15943 );
or ( n16187 , n16185 , n16186 );
not ( n16188 , n8223 );
not ( n16189 , n15951 );
or ( n16190 , n16188 , n16189 );
xor ( n16191 , n544 , n14087 );
nand ( n16192 , n16191 , n8215 );
nand ( n16193 , n16190 , n16192 );
and ( n16194 , n15941 , n8381 );
and ( n16195 , n5757 , n546 );
nor ( n16196 , n16194 , n16195 );
xor ( n16197 , n16193 , n16196 );
and ( n16198 , n544 , n15290 );
xor ( n16199 , n16197 , n16198 );
xor ( n16200 , n16187 , n16199 );
xor ( n16201 , n15947 , n15953 );
and ( n16202 , n16201 , n15958 );
and ( n16203 , n15947 , n15953 );
or ( n16204 , n16202 , n16203 );
xor ( n16205 , n16200 , n16204 );
not ( n16206 , n16205 );
xor ( n16207 , n15946 , n15959 );
and ( n16208 , n16207 , n15964 );
and ( n16209 , n15946 , n15959 );
or ( n16210 , n16208 , n16209 );
not ( n16211 , n16210 );
nand ( n16212 , n16206 , n16211 );
or ( n16213 , n16206 , n16211 );
and ( n16214 , n16212 , n16213 );
xor ( n16215 , n16183 , n16214 );
nand ( n16216 , n363684 , n363833 );
not ( n16217 , n16216 );
not ( n16218 , n16217 );
buf ( n16219 , n14961 );
not ( n16220 , n16219 );
or ( n16221 , n16218 , n16220 );
not ( n16222 , n14947 );
nor ( n16223 , n16222 , n16216 );
and ( n16224 , n16223 , n363689 );
not ( n16225 , n363833 );
not ( n16226 , n363679 );
or ( n16227 , n16225 , n16226 );
nand ( n16228 , n16227 , n363838 );
nor ( n16229 , n16224 , n16228 );
nand ( n16230 , n16221 , n16229 );
xor ( n16231 , n363707 , n363818 );
and ( n16232 , n16231 , n363825 );
and ( n16233 , n363707 , n363818 );
or ( n16234 , n16232 , n16233 );
buf ( n363911 , n16234 );
buf ( n363912 , n363911 );
not ( n16237 , n363912 );
xor ( n16238 , n363770 , n363799 );
and ( n16239 , n16238 , n363806 );
and ( n16240 , n363770 , n363799 );
or ( n16241 , n16239 , n16240 );
buf ( n363918 , n16241 );
buf ( n363919 , n363918 );
buf ( n363920 , n16117 );
not ( n16245 , n16108 );
not ( n16246 , n16106 );
or ( n16247 , n16245 , n16246 );
not ( n16248 , n16106 );
nand ( n16249 , n16248 , n16107 );
nand ( n16250 , n16120 , n16249 );
nand ( n16251 , n16247 , n16250 );
buf ( n363928 , n16251 );
xor ( n16253 , n363920 , n363928 );
and ( n16254 , n363453 , n363454 );
buf ( n363931 , n16254 );
buf ( n363932 , n363931 );
or ( n16257 , n352295 , n8604 );
nand ( n16258 , n16257 , n562 );
buf ( n363935 , n16258 );
xor ( n16260 , n363932 , n363935 );
buf ( n363937 , n363778 );
not ( n16262 , n363937 );
buf ( n363939 , n9186 );
not ( n16264 , n363939 );
or ( n16265 , n16262 , n16264 );
buf ( n363942 , n560 );
buf ( n363943 , n544 );
xnor ( n16268 , n363942 , n363943 );
buf ( n363945 , n16268 );
buf ( n363946 , n363945 );
not ( n16271 , n363946 );
buf ( n363948 , n5407 );
nand ( n16273 , n16271 , n363948 );
buf ( n363950 , n16273 );
buf ( n363951 , n363950 );
nand ( n16276 , n16265 , n363951 );
buf ( n363953 , n16276 );
buf ( n363954 , n363953 );
xor ( n16279 , n16260 , n363954 );
buf ( n363956 , n16279 );
buf ( n363957 , n363956 );
xor ( n16282 , n16253 , n363957 );
buf ( n363959 , n16282 );
buf ( n363960 , n363959 );
buf ( n363961 , n363746 );
xor ( n16286 , n363716 , n363733 );
and ( n16287 , n16286 , n363750 );
and ( n16288 , n363716 , n363733 );
or ( n16289 , n16287 , n16288 );
buf ( n363966 , n16289 );
buf ( n363967 , n363966 );
xor ( n16292 , n363961 , n363967 );
and ( n16293 , n363494 , n363495 );
buf ( n363970 , n16293 );
buf ( n363971 , n363970 );
buf ( n363972 , n363726 );
not ( n16297 , n363972 );
buf ( n363974 , n361110 );
not ( n16299 , n363974 );
or ( n16300 , n16297 , n16299 );
buf ( n363977 , n576 );
buf ( n363978 , n544 );
xnor ( n16303 , n363977 , n363978 );
buf ( n363980 , n16303 );
buf ( n363981 , n363980 );
not ( n16306 , n363981 );
buf ( n363983 , n356446 );
nand ( n16308 , n16306 , n363983 );
buf ( n363985 , n16308 );
buf ( n363986 , n363985 );
nand ( n16311 , n16300 , n363986 );
buf ( n363988 , n16311 );
buf ( n363989 , n363988 );
xor ( n16314 , n363971 , n363989 );
buf ( n363991 , n354788 );
buf ( n363992 , n361131 );
or ( n16317 , n363991 , n363992 );
buf ( n363994 , n578 );
nand ( n16319 , n16317 , n363994 );
buf ( n363996 , n16319 );
buf ( n363997 , n363996 );
xor ( n16322 , n16314 , n363997 );
buf ( n363999 , n16322 );
buf ( n364000 , n363999 );
xor ( n16325 , n16292 , n364000 );
buf ( n364002 , n16325 );
buf ( n364003 , n364002 );
xor ( n16328 , n363960 , n364003 );
xor ( n16329 , n363713 , n363753 );
and ( n16330 , n16329 , n363761 );
and ( n16331 , n363713 , n363753 );
or ( n16332 , n16330 , n16331 );
buf ( n364009 , n16332 );
buf ( n364010 , n364009 );
xor ( n16335 , n16328 , n364010 );
buf ( n364012 , n16335 );
buf ( n364013 , n364012 );
xor ( n16338 , n363919 , n364013 );
xor ( n16339 , n363764 , n363809 );
and ( n16340 , n16339 , n363815 );
and ( n16341 , n363764 , n363809 );
or ( n16342 , n16340 , n16341 );
buf ( n364019 , n16342 );
buf ( n364020 , n364019 );
xor ( n16345 , n16338 , n364020 );
buf ( n364022 , n16345 );
buf ( n364023 , n364022 );
not ( n16348 , n364023 );
buf ( n364025 , n16348 );
buf ( n364026 , n364025 );
nand ( n16351 , n16237 , n364026 );
buf ( n364028 , n16351 );
buf ( n364029 , n364028 );
buf ( n364030 , n364025 );
not ( n16355 , n364030 );
buf ( n364032 , n363911 );
nand ( n16357 , n16355 , n364032 );
buf ( n364034 , n16357 );
buf ( n364035 , n364034 );
and ( n16360 , n364029 , n364035 );
buf ( n364037 , n16360 );
xnor ( n16362 , n16230 , n364037 );
nand ( n16363 , n16215 , n16362 );
nand ( n16364 , n16166 , n16363 );
not ( n16365 , n16364 );
buf ( n364042 , n363833 );
buf ( n364043 , n364028 );
and ( n16368 , n364042 , n364043 );
buf ( n364045 , n16368 );
buf ( n364046 , n364045 );
not ( n16371 , n364046 );
buf ( n364048 , n363679 );
not ( n16373 , n364048 );
or ( n16374 , n16371 , n16373 );
buf ( n364051 , n363838 );
not ( n16376 , n364051 );
buf ( n364053 , n364028 );
not ( n16378 , n364053 );
buf ( n364055 , n16378 );
buf ( n364056 , n364055 );
not ( n16381 , n364056 );
and ( n16382 , n16376 , n16381 );
buf ( n364059 , n364034 );
not ( n16384 , n364059 );
buf ( n364061 , n16384 );
buf ( n364062 , n364061 );
nor ( n16387 , n16382 , n364062 );
buf ( n364064 , n16387 );
buf ( n364065 , n364064 );
nand ( n16390 , n16374 , n364065 );
buf ( n364067 , n16390 );
buf ( n364068 , n364067 );
not ( n16393 , n364068 );
buf ( n364070 , n16219 );
buf ( n364071 , n363684 );
buf ( n364072 , n364045 );
and ( n16397 , n364071 , n364072 );
buf ( n364074 , n16397 );
buf ( n364075 , n364074 );
nand ( n16400 , n364070 , n364075 );
buf ( n364077 , n16400 );
buf ( n364078 , n364077 );
buf ( n364079 , n14947 );
buf ( n364080 , n363689 );
buf ( n364081 , n364074 );
nand ( n16406 , n364079 , n364080 , n364081 );
buf ( n364083 , n16406 );
buf ( n364084 , n364083 );
nand ( n16409 , n16393 , n364078 , n364084 );
buf ( n364086 , n16409 );
xor ( n16411 , n363919 , n364013 );
and ( n16412 , n16411 , n364020 );
and ( n16413 , n363919 , n364013 );
or ( n16414 , n16412 , n16413 );
buf ( n364091 , n16414 );
buf ( n364092 , n364091 );
xor ( n16417 , n363920 , n363928 );
and ( n16418 , n16417 , n363957 );
and ( n16419 , n363920 , n363928 );
or ( n16420 , n16418 , n16419 );
buf ( n364097 , n16420 );
buf ( n364098 , n364097 );
buf ( n364099 , n545 );
buf ( n364100 , n560 );
nand ( n16425 , n364099 , n364100 );
buf ( n364102 , n16425 );
buf ( n364103 , n364102 );
buf ( n364104 , n9186 );
not ( n16429 , n364104 );
buf ( n364106 , n16429 );
buf ( n364107 , n364106 );
buf ( n364108 , n363945 );
or ( n16433 , n364107 , n364108 );
buf ( n364110 , n5407 );
not ( n16435 , n364110 );
buf ( n364112 , n16435 );
buf ( n364113 , n364112 );
buf ( n364114 , n6768 );
or ( n16439 , n364113 , n364114 );
nand ( n16440 , n16433 , n16439 );
buf ( n364117 , n16440 );
buf ( n364118 , n364117 );
xor ( n16443 , n364103 , n364118 );
xor ( n16444 , n363932 , n363935 );
and ( n16445 , n16444 , n363954 );
and ( n16446 , n363932 , n363935 );
or ( n16447 , n16445 , n16446 );
buf ( n364124 , n16447 );
buf ( n364125 , n364124 );
xor ( n16450 , n16443 , n364125 );
buf ( n364127 , n16450 );
buf ( n364128 , n364127 );
buf ( n364129 , n545 );
buf ( n364130 , n576 );
nand ( n16455 , n364129 , n364130 );
buf ( n364132 , n16455 );
buf ( n364133 , n364132 );
buf ( n364134 , n361110 );
not ( n16459 , n364134 );
buf ( n364136 , n16459 );
buf ( n364137 , n364136 );
buf ( n364138 , n363980 );
or ( n16463 , n364137 , n364138 );
buf ( n364140 , n356446 );
not ( n16465 , n364140 );
buf ( n364142 , n16465 );
buf ( n364143 , n364142 );
buf ( n364144 , n354303 );
or ( n16469 , n364143 , n364144 );
nand ( n16470 , n16463 , n16469 );
buf ( n364147 , n16470 );
buf ( n364148 , n364147 );
xor ( n16473 , n364133 , n364148 );
xor ( n16474 , n363971 , n363989 );
and ( n16475 , n16474 , n363997 );
and ( n16476 , n363971 , n363989 );
or ( n16477 , n16475 , n16476 );
buf ( n364154 , n16477 );
buf ( n364155 , n364154 );
xor ( n16480 , n16473 , n364155 );
buf ( n364157 , n16480 );
buf ( n364158 , n364157 );
xor ( n16483 , n364128 , n364158 );
xor ( n16484 , n363961 , n363967 );
and ( n16485 , n16484 , n364000 );
and ( n16486 , n363961 , n363967 );
or ( n16487 , n16485 , n16486 );
buf ( n364164 , n16487 );
buf ( n364165 , n364164 );
xor ( n16490 , n16483 , n364165 );
buf ( n364167 , n16490 );
buf ( n364168 , n364167 );
xor ( n16493 , n364098 , n364168 );
xor ( n16494 , n363960 , n364003 );
and ( n16495 , n16494 , n364010 );
and ( n16496 , n363960 , n364003 );
or ( n16497 , n16495 , n16496 );
buf ( n364174 , n16497 );
buf ( n364175 , n364174 );
xor ( n16500 , n16493 , n364175 );
buf ( n364177 , n16500 );
buf ( n364178 , n364177 );
and ( n16503 , n364092 , n364178 );
buf ( n364180 , n16503 );
buf ( n364181 , n364180 );
buf ( n364182 , n364091 );
buf ( n364183 , n364177 );
nor ( n16508 , n364182 , n364183 );
buf ( n364185 , n16508 );
buf ( n364186 , n364185 );
nor ( n16511 , n364181 , n364186 );
buf ( n364188 , n16511 );
not ( n16513 , n364188 );
and ( n16514 , n364086 , n16513 );
not ( n16515 , n364086 );
and ( n16516 , n16515 , n364188 );
or ( n16517 , n16514 , n16516 );
not ( n16518 , n16517 );
nand ( n16519 , n16183 , n16212 );
not ( n16520 , n16519 );
xor ( n16521 , n16187 , n16199 );
and ( n16522 , n16521 , n16204 );
and ( n16523 , n16187 , n16199 );
or ( n16524 , n16522 , n16523 );
not ( n16525 , n16524 );
and ( n16526 , n544 , n14581 );
xor ( n16527 , n16193 , n16196 );
and ( n16528 , n16527 , n16198 );
and ( n16529 , n16193 , n16196 );
or ( n16530 , n16528 , n16529 );
xor ( n16531 , n16526 , n16530 );
or ( n16532 , n8381 , n5757 );
nand ( n16533 , n16532 , n546 );
not ( n16534 , n16191 );
not ( n16535 , n8223 );
or ( n16536 , n16534 , n16535 );
and ( n16537 , n14552 , n544 );
and ( n16538 , n14549 , n7283 );
nor ( n16539 , n16537 , n16538 );
not ( n16540 , n8215 );
or ( n16541 , n16539 , n16540 );
nand ( n16542 , n16536 , n16541 );
xor ( n16543 , n16533 , n16542 );
not ( n16544 , n16196 );
xor ( n16545 , n16543 , n16544 );
xor ( n16546 , n16531 , n16545 );
not ( n16547 , n16546 );
nand ( n16548 , n16525 , n16547 );
not ( n16549 , n16548 );
nor ( n16550 , n16547 , n16525 );
nor ( n16551 , n16549 , n16550 );
and ( n16552 , n16551 , n16213 );
not ( n16553 , n16552 );
or ( n16554 , n16520 , n16553 );
not ( n16555 , n16213 );
not ( n16556 , n16519 );
or ( n16557 , n16555 , n16556 );
not ( n16558 , n16551 );
nand ( n16559 , n16557 , n16558 );
nand ( n16560 , n16554 , n16559 );
nand ( n16561 , n16518 , n16560 );
nand ( n16562 , n16365 , n16561 );
nor ( n16563 , n15927 , n16562 );
not ( n16564 , n16563 );
or ( n16565 , n14528 , n16564 );
not ( n16566 , n16562 );
nand ( n16567 , n15349 , n15354 );
not ( n16568 , n16567 );
not ( n16569 , n15269 );
not ( n16570 , n16569 );
or ( n16571 , n16568 , n16570 );
and ( n16572 , n14623 , n14609 );
not ( n16573 , n14623 );
and ( n16574 , n16573 , n14610 );
nor ( n16575 , n16572 , n16574 );
and ( n16576 , n14963 , n362645 );
not ( n16577 , n14963 );
and ( n16578 , n16577 , n362608 );
nor ( n16579 , n16576 , n16578 );
nand ( n16580 , n16575 , n16579 );
nand ( n16581 , n16571 , n16580 );
buf ( n16582 , n15355 );
nand ( n16583 , n16581 , n15926 , n16582 );
not ( n16584 , n15921 );
not ( n16585 , n16584 );
not ( n16586 , n15922 );
not ( n16587 , n15673 );
or ( n16588 , n16586 , n16587 );
nand ( n16589 , n15672 , n15723 );
nand ( n16590 , n16588 , n16589 );
nand ( n16591 , n16585 , n16590 );
not ( n16592 , n15579 );
nor ( n16593 , n16592 , n15663 );
and ( n16594 , n16591 , n16593 );
nor ( n16595 , n16590 , n15921 );
nor ( n16596 , n16594 , n16595 );
nand ( n16597 , n16583 , n16596 );
buf ( n16598 , n16597 );
and ( n16599 , n16566 , n16598 );
not ( n16600 , n16561 );
nor ( n16601 , n16164 , n15984 );
not ( n16602 , n16601 );
not ( n16603 , n16363 );
or ( n16604 , n16602 , n16603 );
or ( n16605 , n16215 , n16362 );
nand ( n16606 , n16604 , n16605 );
not ( n16607 , n16606 );
or ( n16608 , n16600 , n16607 );
not ( n16609 , n16560 );
nand ( n16610 , n16609 , n16517 );
nand ( n16611 , n16608 , n16610 );
nor ( n16612 , n16599 , n16611 );
nand ( n16613 , n16565 , n16612 );
nand ( n16614 , n16212 , n16548 );
nor ( n16615 , n15966 , n16614 );
not ( n16616 , n16615 );
not ( n16617 , n15978 );
or ( n16618 , n16616 , n16617 );
not ( n16619 , n16212 );
not ( n16620 , n16181 );
or ( n16621 , n16619 , n16620 );
nand ( n16622 , n16621 , n16213 );
and ( n16623 , n16622 , n16548 );
nor ( n16624 , n16623 , n16550 );
nand ( n16625 , n16618 , n16624 );
xor ( n16626 , n16526 , n16530 );
and ( n16627 , n16626 , n16545 );
and ( n16628 , n16526 , n16530 );
or ( n16629 , n16627 , n16628 );
not ( n16630 , n16629 );
and ( n16631 , n544 , n14087 );
not ( n16632 , n16539 );
and ( n16633 , n16632 , n8223 );
and ( n16634 , n8215 , n544 );
nor ( n16635 , n16633 , n16634 );
xor ( n16636 , n16631 , n16635 );
xor ( n16637 , n16533 , n16542 );
and ( n16638 , n16637 , n16544 );
and ( n16639 , n16533 , n16542 );
or ( n16640 , n16638 , n16639 );
xor ( n16641 , n16636 , n16640 );
not ( n16642 , n16641 );
and ( n16643 , n16630 , n16642 );
and ( n16644 , n16629 , n16641 );
nor ( n16645 , n16643 , n16644 );
and ( n16646 , n16625 , n16645 );
not ( n16647 , n16625 );
not ( n16648 , n16645 );
and ( n16649 , n16647 , n16648 );
nor ( n16650 , n16646 , n16649 );
buf ( n364327 , n364045 );
not ( n16652 , n364327 );
buf ( n364329 , n364185 );
nor ( n16654 , n16652 , n364329 );
buf ( n364331 , n16654 );
buf ( n364332 , n364331 );
not ( n16657 , n364332 );
buf ( n364334 , n363679 );
not ( n16659 , n364334 );
or ( n16660 , n16657 , n16659 );
buf ( n364337 , n364064 );
not ( n16662 , n364337 );
buf ( n364339 , n364185 );
not ( n16664 , n364339 );
and ( n16665 , n16662 , n16664 );
buf ( n364342 , n364180 );
nor ( n16667 , n16665 , n364342 );
buf ( n364344 , n16667 );
buf ( n364345 , n364344 );
nand ( n16670 , n16660 , n364345 );
buf ( n364347 , n16670 );
buf ( n364348 , n364347 );
not ( n16673 , n364348 );
buf ( n364350 , n16219 );
buf ( n364351 , n363684 );
buf ( n364352 , n364331 );
and ( n16677 , n364351 , n364352 );
buf ( n364354 , n16677 );
buf ( n364355 , n364354 );
nand ( n16680 , n364350 , n364355 );
buf ( n364357 , n16680 );
buf ( n364358 , n364357 );
buf ( n364359 , n14947 );
buf ( n364360 , n363689 );
buf ( n364361 , n364354 );
nand ( n16686 , n364359 , n364360 , n364361 );
buf ( n364363 , n16686 );
buf ( n364364 , n364363 );
nand ( n16689 , n16673 , n364358 , n364364 );
buf ( n364366 , n16689 );
buf ( n364367 , n544 );
buf ( n364368 , n576 );
nand ( n16693 , n364367 , n364368 );
buf ( n364370 , n16693 );
buf ( n364371 , n364370 );
not ( n16696 , n364371 );
buf ( n364373 , n361110 );
buf ( n364374 , n356446 );
or ( n16699 , n364373 , n364374 );
buf ( n364376 , n576 );
nand ( n16701 , n16699 , n364376 );
buf ( n364378 , n16701 );
buf ( n364379 , n364378 );
not ( n16704 , n364379 );
or ( n16705 , n16696 , n16704 );
buf ( n364382 , n364378 );
buf ( n364383 , n364370 );
or ( n16708 , n364382 , n364383 );
nand ( n16709 , n16705 , n16708 );
buf ( n364386 , n16709 );
buf ( n364387 , n364386 );
buf ( n364388 , n364132 );
xnor ( n16713 , n364387 , n364388 );
buf ( n364390 , n16713 );
buf ( n364391 , n364390 );
not ( n16716 , n364391 );
xor ( n16717 , n364133 , n364148 );
and ( n16718 , n16717 , n364155 );
and ( n16719 , n364133 , n364148 );
or ( n16720 , n16718 , n16719 );
buf ( n364397 , n16720 );
buf ( n364398 , n364397 );
buf ( n364399 , n544 );
buf ( n364400 , n560 );
nand ( n16725 , n364399 , n364400 );
buf ( n364402 , n16725 );
buf ( n364403 , n364402 );
not ( n16728 , n364403 );
buf ( n364405 , n9186 );
buf ( n364406 , n5407 );
or ( n16731 , n364405 , n364406 );
buf ( n364408 , n560 );
nand ( n16733 , n16731 , n364408 );
buf ( n364410 , n16733 );
buf ( n364411 , n364410 );
not ( n16736 , n364411 );
or ( n16737 , n16728 , n16736 );
buf ( n364414 , n364410 );
buf ( n364415 , n364402 );
or ( n16740 , n364414 , n364415 );
nand ( n16741 , n16737 , n16740 );
buf ( n364418 , n16741 );
buf ( n364419 , n364418 );
buf ( n364420 , n364102 );
xnor ( n16745 , n364419 , n364420 );
buf ( n364422 , n16745 );
buf ( n364423 , n364422 );
xnor ( n16748 , n364398 , n364423 );
buf ( n364425 , n16748 );
buf ( n364426 , n364425 );
not ( n16751 , n364426 );
or ( n16752 , n16716 , n16751 );
buf ( n364429 , n364425 );
buf ( n364430 , n364390 );
or ( n16755 , n364429 , n364430 );
nand ( n16756 , n16752 , n16755 );
buf ( n364433 , n16756 );
buf ( n364434 , n364433 );
xor ( n16759 , n364128 , n364158 );
and ( n16760 , n16759 , n364165 );
and ( n16761 , n364128 , n364158 );
or ( n16762 , n16760 , n16761 );
buf ( n364439 , n16762 );
buf ( n364440 , n364439 );
xor ( n16765 , n364103 , n364118 );
and ( n16766 , n16765 , n364125 );
and ( n16767 , n364103 , n364118 );
or ( n16768 , n16766 , n16767 );
buf ( n364445 , n16768 );
buf ( n364446 , n364445 );
xnor ( n16771 , n364440 , n364446 );
buf ( n364448 , n16771 );
buf ( n364449 , n364448 );
xnor ( n16774 , n364434 , n364449 );
buf ( n364451 , n16774 );
buf ( n364452 , n364451 );
not ( n16777 , n364452 );
xor ( n16778 , n364098 , n364168 );
and ( n16779 , n16778 , n364175 );
and ( n16780 , n364098 , n364168 );
or ( n16781 , n16779 , n16780 );
buf ( n364458 , n16781 );
buf ( n364459 , n364458 );
not ( n16784 , n364459 );
or ( n16785 , n16777 , n16784 );
buf ( n364462 , n364458 );
buf ( n364463 , n364451 );
or ( n16788 , n364462 , n364463 );
nand ( n16789 , n16785 , n16788 );
buf ( n364466 , n16789 );
xor ( n16791 , n364366 , n364466 );
nand ( n16792 , n16650 , n16791 );
or ( n16793 , n16650 , n16791 );
nand ( n16794 , n16792 , n16793 );
not ( n16795 , n16794 );
and ( n16796 , n16613 , n16795 );
not ( n16797 , n16613 );
and ( n16798 , n16797 , n16794 );
nor ( n16799 , n16796 , n16798 );
nor ( n16800 , n15927 , n16364 );
not ( n16801 , n16800 );
not ( n16802 , n14527 );
or ( n16803 , n16801 , n16802 );
and ( n16804 , n16597 , n16365 );
nor ( n16805 , n16804 , n16606 );
nand ( n16806 , n16803 , n16805 );
not ( n16807 , n16517 );
nand ( n16808 , n16807 , n16560 );
nand ( n16809 , n16610 , n16808 );
and ( n16810 , n16806 , n16809 );
not ( n16811 , n16806 );
not ( n16812 , n16809 );
and ( n16813 , n16811 , n16812 );
nor ( n16814 , n16810 , n16813 );
not ( n16815 , n16814 );
nand ( n16816 , n16605 , n16363 );
not ( n16817 , n16816 );
nand ( n16818 , n16583 , n16596 );
nand ( n16819 , n15984 , n16164 );
buf ( n16820 , n16819 );
nand ( n16821 , n16818 , n16820 );
buf ( n16822 , n8298 );
and ( n16823 , n14525 , n16822 );
nand ( n16824 , n15663 , n15580 );
and ( n16825 , n15356 , n16819 , n16591 , n16824 );
nand ( n16826 , n16823 , n16825 );
not ( n16827 , n14512 );
not ( n16828 , n14510 );
or ( n16829 , n16827 , n16828 );
not ( n16830 , n14522 );
nand ( n16831 , n16829 , n16830 );
and ( n16832 , n16825 , n16831 );
or ( n16833 , n15984 , n16164 );
not ( n16834 , n16833 );
nor ( n16835 , n16832 , n16834 );
nand ( n16836 , n16821 , n16826 , n16835 );
not ( n16837 , n16836 );
or ( n16838 , n16817 , n16837 );
not ( n16839 , n16816 );
nand ( n16840 , n16821 , n16826 , n16835 , n16839 );
nand ( n16841 , n16838 , n16840 );
and ( n16842 , n16820 , n16833 );
nand ( n16843 , n16583 , n16596 );
not ( n16844 , n16843 );
not ( n16845 , n14512 );
not ( n16846 , n14510 );
or ( n16847 , n16845 , n16846 );
nand ( n16848 , n16847 , n16830 );
not ( n16849 , n15927 );
nand ( n16850 , n16848 , n16849 );
not ( n16851 , n15927 );
nand ( n16852 , n16851 , n14525 , n16822 );
nand ( n16853 , n16844 , n16850 , n16852 );
xor ( n16854 , n16842 , n16853 );
nand ( n16855 , n16841 , n16854 );
not ( n16856 , n16855 );
nand ( n16857 , n14502 , n16799 , n16815 , n16856 );
and ( n16858 , n16824 , n15356 );
nand ( n16859 , n16858 , n16848 );
not ( n16860 , n14507 );
or ( n16861 , n16575 , n16579 );
nand ( n16862 , n16861 , n8298 );
nor ( n16863 , n16860 , n16862 );
not ( n16864 , n16863 );
not ( n16865 , n12517 );
nor ( n16866 , n16865 , n13566 );
not ( n16867 , n16866 );
or ( n16868 , n16864 , n16867 );
not ( n16869 , n16581 );
nand ( n16870 , n16868 , n16869 );
and ( n16871 , n16582 , n16824 );
and ( n16872 , n16870 , n16871 );
nor ( n16873 , n16872 , n16593 );
nand ( n16874 , n16859 , n16873 );
not ( n16875 , n16874 );
not ( n16876 , n16590 );
or ( n16877 , n16584 , n16876 );
not ( n16878 , n16595 );
nand ( n16879 , n16877 , n16878 );
not ( n16880 , n16879 );
not ( n16881 , n16880 );
or ( n16882 , n16875 , n16881 );
nand ( n16883 , n16859 , n16873 , n16879 );
nand ( n16884 , n16882 , n16883 );
not ( n16885 , n16884 );
not ( n16886 , n8298 );
not ( n16887 , n14525 );
or ( n16888 , n16886 , n16887 );
nand ( n16889 , n16888 , n14523 );
buf ( n16890 , n16580 );
buf ( n16891 , n14972 );
buf ( n16892 , n14628 );
nand ( n16893 , n16891 , n16892 );
nand ( n16894 , n16890 , n16893 );
not ( n16895 , n16894 );
and ( n16896 , n16889 , n16895 );
not ( n16897 , n16889 );
and ( n16898 , n16897 , n16894 );
nor ( n16899 , n16896 , n16898 );
buf ( n16900 , n16899 );
nand ( n16901 , n16860 , n14521 );
not ( n16902 , n16901 );
not ( n16903 , n13565 );
not ( n16904 , n12514 );
or ( n16905 , n16903 , n16904 );
nor ( n16906 , n14039 , n14520 );
nand ( n16907 , n16905 , n16906 );
not ( n16908 , n16907 );
or ( n16909 , n16902 , n16908 );
not ( n16910 , n14510 );
not ( n16911 , n16910 );
not ( n16912 , n12518 );
and ( n16913 , n16911 , n16912 );
nor ( n16914 , n16913 , n16581 );
nand ( n16915 , n16909 , n16914 );
not ( n16916 , n16893 );
and ( n16917 , n16869 , n16916 );
not ( n16918 , n16582 );
nor ( n16919 , n16917 , n16918 );
nand ( n16920 , n16915 , n16919 );
not ( n16921 , n16593 );
not ( n16922 , n16824 );
not ( n16923 , n16922 );
nand ( n16924 , n16921 , n16923 );
and ( n16925 , n16920 , n16924 );
not ( n16926 , n16920 );
not ( n16927 , n16924 );
and ( n16928 , n16926 , n16927 );
nor ( n16929 , n16925 , n16928 );
nand ( n16930 , n16907 , n16901 , n16893 );
not ( n16931 , n16569 );
not ( n16932 , n16567 );
or ( n16933 , n16931 , n16932 );
or ( n16934 , n16569 , n16567 );
nand ( n16935 , n16933 , n16934 );
not ( n16936 , n16935 );
nor ( n16937 , n16930 , n16936 );
not ( n16938 , n16937 );
not ( n16939 , n14525 );
nand ( n16940 , n16936 , n16890 );
not ( n16941 , n16940 );
nand ( n16942 , n16939 , n16930 , n16941 );
not ( n16943 , n16862 );
not ( n16944 , n16943 );
nand ( n16945 , n16930 , n16941 , n16944 );
not ( n16946 , n14524 );
nand ( n16947 , n16935 , n16943 );
not ( n16948 , n16947 );
and ( n16949 , n16946 , n16948 );
not ( n16950 , n16890 );
not ( n16951 , n16936 );
and ( n16952 , n16950 , n16951 );
nor ( n16953 , n16949 , n16952 );
nand ( n16954 , n16938 , n16942 , n16945 , n16953 );
buf ( n16955 , n16954 );
nand ( n16956 , n16885 , n16900 , n16929 , n16955 );
not ( n16957 , n16956 );
buf ( n16958 , n8323 );
nand ( n16959 , n16957 , n16958 );
nor ( n16960 , n16857 , n16959 );
not ( n16961 , n16818 );
and ( n16962 , n16808 , n16792 , n16365 );
not ( n16963 , n16962 );
or ( n16964 , n16961 , n16963 );
and ( n16965 , n16606 , n16792 , n16808 );
nand ( n16966 , n16650 , n16791 );
not ( n16967 , n16966 );
not ( n16968 , n16610 );
not ( n16969 , n16968 );
or ( n16970 , n16967 , n16969 );
nand ( n16971 , n16970 , n16793 );
nor ( n16972 , n16965 , n16971 );
nand ( n16973 , n16964 , n16972 );
not ( n16974 , n16973 );
not ( n16975 , n16822 );
not ( n16976 , n14525 );
or ( n16977 , n16975 , n16976 );
not ( n16978 , n16831 );
nand ( n16979 , n16977 , n16978 );
nand ( n16980 , n16962 , n16849 , n16979 );
nand ( n16981 , n16974 , n16980 );
not ( n16982 , n16981 );
buf ( n364659 , n16982 );
buf ( n16984 , n364659 );
buf ( n364661 , n16984 );
buf ( n364662 , n364661 );
not ( n16987 , n364662 );
buf ( n364664 , n16987 );
nor ( n16989 , n16960 , n364664 );
not ( n16990 , n16989 );
nand ( n16991 , n364664 , n16960 );
nand ( n16992 , n16990 , n16991 );
buf ( n16993 , n16992 );
not ( n16994 , n16989 );
not ( n16995 , n16994 );
nand ( n16996 , n14500 , n16900 , n16955 , n16958 );
not ( n16997 , n16927 );
nand ( n16998 , n16915 , n16919 );
not ( n16999 , n16998 );
or ( n17000 , n16997 , n16999 );
nand ( n17001 , n16915 , n16924 , n16919 );
nand ( n17002 , n17000 , n17001 );
buf ( n17003 , n17002 );
not ( n17004 , n17003 );
and ( n17005 , n16996 , n17004 );
not ( n17006 , n16996 );
and ( n17007 , n17006 , n17003 );
nor ( n17008 , n17005 , n17007 );
buf ( n17009 , n17008 );
not ( n17010 , n14499 );
nand ( n17011 , n17010 , n8327 );
not ( n17012 , n17011 );
buf ( n17013 , n16854 );
nand ( n17014 , n16957 , n17012 , n17013 );
not ( n17015 , n17014 );
not ( n17016 , n13074 );
and ( n17017 , n9625 , n12407 );
nand ( n17018 , n17016 , n17017 );
not ( n17019 , n17018 );
nand ( n17020 , n17019 , n8327 );
buf ( n17021 , n13072 );
buf ( n17022 , n17021 );
nand ( n17023 , n17019 , n17022 , n8327 );
buf ( n17024 , n14473 );
not ( n17025 , n14485 );
not ( n17026 , n17025 );
nand ( n17027 , n17024 , n17026 );
nand ( n17028 , n14498 , n17021 );
nor ( n17029 , n17027 , n17028 );
and ( n17030 , n16955 , n17029 );
nand ( n17031 , n14498 , n17021 );
buf ( n364708 , n363808 );
buf ( n364709 , n363706 );
nand ( n17034 , n5655 , n579 );
nand ( n17035 , n6388 , n580 );
nand ( n17036 , n17034 , n17035 );
buf ( n17037 , n17036 );
buf ( n364714 , n17037 );
not ( n17039 , n364714 );
buf ( n364716 , n578 );
not ( n17041 , n364716 );
buf ( n364718 , n8990 );
not ( n17043 , n364718 );
buf ( n364720 , n17043 );
buf ( n364721 , n364720 );
not ( n17046 , n364721 );
or ( n17047 , n17041 , n17046 );
buf ( n364724 , n357348 );
buf ( n364725 , n578 );
not ( n17050 , n364725 );
buf ( n364727 , n17050 );
buf ( n364728 , n364727 );
nand ( n17053 , n364724 , n364728 );
buf ( n364730 , n17053 );
buf ( n364731 , n364730 );
nand ( n17056 , n17047 , n364731 );
buf ( n364733 , n17056 );
buf ( n364734 , n364733 );
not ( n17059 , n364734 );
or ( n17060 , n17039 , n17059 );
buf ( n364737 , n578 );
not ( n17062 , n364737 );
buf ( n364739 , n8304 );
not ( n17064 , n364739 );
or ( n17065 , n17062 , n17064 );
buf ( n364742 , n8303 );
buf ( n364743 , n364727 );
nand ( n17068 , n364742 , n364743 );
buf ( n364745 , n17068 );
buf ( n364746 , n364745 );
nand ( n17071 , n17065 , n364746 );
buf ( n364748 , n17071 );
buf ( n364749 , n364748 );
buf ( n364750 , n578 );
buf ( n364751 , n579 );
nor ( n17076 , n364750 , n364751 );
buf ( n364753 , n17076 );
not ( n17078 , n364753 );
and ( n17079 , n578 , n579 );
nor ( n17080 , n17079 , n17037 );
nand ( n17081 , n17078 , n17080 );
not ( n17082 , n17081 );
buf ( n364759 , n17082 );
nand ( n17084 , n364749 , n364759 );
buf ( n364761 , n17084 );
buf ( n364762 , n364761 );
nand ( n17087 , n17060 , n364762 );
buf ( n364764 , n17087 );
buf ( n364765 , n364764 );
buf ( n364766 , n351277 );
buf ( n364767 , n584 );
or ( n17092 , n364766 , n364767 );
buf ( n364769 , n584 );
not ( n17094 , n364769 );
buf ( n364771 , n17094 );
buf ( n364772 , n364771 );
buf ( n364773 , n583 );
or ( n17098 , n364772 , n364773 );
nand ( n17099 , n17092 , n17098 );
buf ( n364776 , n17099 );
buf ( n364777 , n364776 );
buf ( n17102 , n364777 );
buf ( n364779 , n17102 );
buf ( n364780 , n364779 );
not ( n17105 , n364780 );
xor ( n17106 , n582 , n14498 );
buf ( n364783 , n17106 );
not ( n17108 , n364783 );
or ( n17109 , n17105 , n17108 );
buf ( n364786 , n582 );
not ( n17111 , n364786 );
buf ( n364788 , n17021 );
not ( n17113 , n364788 );
buf ( n364790 , n17113 );
buf ( n364791 , n364790 );
not ( n17116 , n364791 );
or ( n17117 , n17111 , n17116 );
buf ( n364794 , n17021 );
buf ( n364795 , n582 );
not ( n17120 , n364795 );
buf ( n364797 , n17120 );
buf ( n364798 , n364797 );
nand ( n17123 , n364794 , n364798 );
buf ( n364800 , n17123 );
buf ( n364801 , n364800 );
nand ( n17126 , n17117 , n364801 );
buf ( n364803 , n17126 );
buf ( n364804 , n364803 );
not ( n17129 , n364776 );
and ( n17130 , n582 , n583 );
and ( n17131 , n364797 , n351277 );
nor ( n17132 , n17130 , n17131 );
nand ( n364809 , n17129 , n17132 );
not ( n17133 , n364809 );
buf ( n364811 , n17133 );
nand ( n17135 , n364804 , n364811 );
buf ( n364813 , n17135 );
buf ( n364814 , n364813 );
nand ( n17138 , n17109 , n364814 );
buf ( n364816 , n17138 );
buf ( n364817 , n364816 );
xor ( n17141 , n364765 , n364817 );
buf ( n364819 , n576 );
nand ( n17143 , n6356 , n6359 );
buf ( n364821 , n17143 );
not ( n17145 , n364821 );
buf ( n364823 , n17145 );
buf ( n364824 , n364823 );
not ( n17148 , n364824 );
buf ( n364826 , n17148 );
buf ( n364827 , n364826 );
and ( n17151 , n364819 , n364827 );
buf ( n364829 , n17151 );
buf ( n364830 , n364829 );
buf ( n364831 , n577 );
buf ( n364832 , n578 );
xor ( n17156 , n364831 , n364832 );
buf ( n364834 , n17156 );
buf ( n364835 , n364834 );
not ( n17159 , n364835 );
buf ( n364837 , n576 );
buf ( n17161 , n7348 );
buf ( n364839 , n17161 );
xor ( n17163 , n364837 , n364839 );
buf ( n364841 , n17163 );
buf ( n364842 , n364841 );
not ( n17166 , n364842 );
or ( n17167 , n17159 , n17166 );
buf ( n364845 , n576 );
not ( n17169 , n353869 );
not ( n17170 , n353961 );
or ( n17171 , n17169 , n17170 );
nand ( n17172 , n17171 , n353965 );
not ( n17173 , n17172 );
not ( n17174 , n17173 );
buf ( n364852 , n17174 );
xor ( n17176 , n364845 , n364852 );
buf ( n364854 , n17176 );
buf ( n364855 , n364854 );
and ( n17179 , n576 , n577 );
nor ( n17180 , n17179 , n364834 );
or ( n17181 , n576 , n577 );
and ( n17182 , n17180 , n17181 );
buf ( n364860 , n17182 );
nand ( n17184 , n364855 , n364860 );
buf ( n364862 , n17184 );
buf ( n364863 , n364862 );
nand ( n17187 , n17167 , n364863 );
buf ( n364865 , n17187 );
buf ( n364866 , n364865 );
xor ( n17190 , n364830 , n364866 );
buf ( n364868 , n580 );
buf ( n364869 , n581 );
and ( n17193 , n364868 , n364869 );
and ( n17194 , n581 , n582 );
not ( n17195 , n581 );
and ( n17196 , n17195 , n364797 );
nor ( n17197 , n17194 , n17196 );
buf ( n364875 , n17197 );
buf ( n364876 , n580 );
buf ( n364877 , n581 );
nor ( n17201 , n364876 , n364877 );
buf ( n364879 , n17201 );
buf ( n364880 , n364879 );
nor ( n17204 , n17193 , n364875 , n364880 );
buf ( n364882 , n17204 );
buf ( n364883 , n364882 );
buf ( n17207 , n364883 );
buf ( n364885 , n17207 );
buf ( n17209 , n364885 );
not ( n17210 , n17209 );
not ( n17211 , n580 );
buf ( n364889 , n9625 );
not ( n17213 , n364889 );
buf ( n364891 , n17213 );
not ( n17215 , n364891 );
or ( n17216 , n17211 , n17215 );
buf ( n364894 , n580 );
not ( n17218 , n364894 );
buf ( n364896 , n17218 );
nand ( n17220 , n364896 , n9625 );
nand ( n364898 , n17216 , n17220 );
not ( n364899 , n364898 );
or ( n364900 , n17210 , n364899 );
buf ( n364901 , n12407 );
not ( n17221 , n364901 );
buf ( n364903 , n17221 );
nand ( n364904 , n364903 , n580 );
not ( n17223 , n364904 );
buf ( n364906 , n360086 );
buf ( n364907 , n364896 );
nand ( n17226 , n364906 , n364907 );
buf ( n364909 , n17226 );
not ( n17228 , n364909 );
or ( n17229 , n17223 , n17228 );
buf ( n17230 , n17197 );
nand ( n17231 , n17229 , n17230 );
nand ( n17232 , n364900 , n17231 );
buf ( n364915 , n17232 );
xor ( n17234 , n17190 , n364915 );
buf ( n364917 , n17234 );
buf ( n364918 , n364917 );
xor ( n17237 , n17141 , n364918 );
buf ( n364920 , n17237 );
buf ( n364921 , n364920 );
buf ( n364922 , n585 );
buf ( n364923 , n586 );
xor ( n17242 , n364922 , n364923 );
buf ( n364925 , n17242 );
buf ( n364926 , n364925 );
not ( n17245 , n364926 );
buf ( n364928 , n584 );
not ( n17247 , n364928 );
not ( n17248 , n14475 );
not ( n17249 , n14481 );
or ( n17250 , n17248 , n17249 );
nand ( n17251 , n17250 , n14484 );
buf ( n364934 , n17251 );
not ( n17253 , n364934 );
buf ( n364936 , n17253 );
buf ( n364937 , n364936 );
not ( n17256 , n364937 );
or ( n17257 , n17247 , n17256 );
nand ( n17258 , n14485 , n364771 );
buf ( n364941 , n17258 );
nand ( n17260 , n17257 , n364941 );
buf ( n364943 , n17260 );
buf ( n364944 , n364943 );
not ( n17263 , n364944 );
or ( n17264 , n17245 , n17263 );
buf ( n364947 , n584 );
not ( n17266 , n364947 );
buf ( n364949 , n14498 );
not ( n17268 , n364949 );
buf ( n364951 , n17268 );
buf ( n364952 , n364951 );
not ( n17271 , n364952 );
or ( n17272 , n17266 , n17271 );
buf ( n364955 , n14498 );
buf ( n364956 , n364771 );
nand ( n17275 , n364955 , n364956 );
buf ( n364958 , n17275 );
buf ( n364959 , n364958 );
nand ( n17278 , n17272 , n364959 );
buf ( n364961 , n17278 );
buf ( n364962 , n364961 );
buf ( n364963 , n584 );
buf ( n364964 , n585 );
and ( n17283 , n364963 , n364964 );
buf ( n364966 , n364925 );
buf ( n364967 , n584 );
buf ( n364968 , n585 );
nor ( n17287 , n364967 , n364968 );
buf ( n364970 , n17287 );
buf ( n364971 , n364970 );
nor ( n17290 , n17283 , n364966 , n364971 );
buf ( n364973 , n17290 );
buf ( n364974 , n364973 );
nand ( n17293 , n364962 , n364974 );
buf ( n364976 , n17293 );
buf ( n364977 , n364976 );
nand ( n17296 , n17264 , n364977 );
buf ( n364979 , n17296 );
buf ( n364980 , n364979 );
buf ( n364981 , n576 );
not ( n17300 , n364981 );
buf ( n17301 , n6351 );
buf ( n364984 , n17301 );
not ( n17303 , n364984 );
buf ( n364986 , n17303 );
buf ( n364987 , n364986 );
buf ( n364988 , n364987 );
nor ( n364989 , n17300 , n364988 );
buf ( n364990 , n364989 );
buf ( n364991 , n364990 );
buf ( n364992 , n364834 );
not ( n17306 , n364992 );
buf ( n364994 , n364854 );
not ( n17307 , n364994 );
or ( n17308 , n17306 , n17307 );
xor ( n17309 , n364819 , n364827 );
buf ( n364998 , n17309 );
buf ( n364999 , n364998 );
buf ( n365000 , n17182 );
nand ( n17313 , n364999 , n365000 );
buf ( n365002 , n17313 );
buf ( n365003 , n365002 );
nand ( n17316 , n17308 , n365003 );
buf ( n365005 , n17316 );
buf ( n365006 , n365005 );
xor ( n17319 , n364991 , n365006 );
buf ( n365008 , n17209 );
not ( n17321 , n365008 );
and ( n17322 , n8990 , n364896 );
not ( n17323 , n8990 );
and ( n17324 , n17323 , n580 );
or ( n17325 , n17322 , n17324 );
buf ( n365014 , n17325 );
not ( n17327 , n365014 );
or ( n17328 , n17321 , n17327 );
buf ( n365017 , n17197 );
not ( n17330 , n365017 );
buf ( n365019 , n17330 );
not ( n17332 , n365019 );
nand ( n17333 , n17332 , n364898 );
buf ( n365022 , n17333 );
nand ( n17335 , n17328 , n365022 );
buf ( n365024 , n17335 );
buf ( n365025 , n365024 );
xor ( n17338 , n17319 , n365025 );
buf ( n365027 , n17338 );
buf ( n365028 , n365027 );
xor ( n17341 , n364980 , n365028 );
buf ( n365030 , n12483 );
not ( n17343 , n365030 );
buf ( n365032 , n17343 );
buf ( n365033 , n365032 );
not ( n17346 , n365033 );
buf ( n365035 , n17346 );
buf ( n365036 , n365035 );
buf ( n365037 , n576 );
and ( n17350 , n365036 , n365037 );
buf ( n365039 , n17350 );
buf ( n365040 , n365039 );
buf ( n365041 , n364834 );
not ( n17354 , n365041 );
buf ( n365043 , n576 );
not ( n17356 , n365043 );
buf ( n365045 , n364986 );
not ( n17358 , n365045 );
or ( n17359 , n17356 , n17358 );
buf ( n365048 , n17301 );
buf ( n365049 , n354303 );
nand ( n17362 , n365048 , n365049 );
buf ( n365051 , n17362 );
buf ( n365052 , n365051 );
nand ( n17365 , n17359 , n365052 );
buf ( n365054 , n17365 );
buf ( n365055 , n365054 );
not ( n17368 , n365055 );
or ( n17369 , n17354 , n17368 );
buf ( n365058 , n576 );
not ( n17371 , n365058 );
buf ( n17372 , n4173 );
buf ( n365061 , n17372 );
not ( n17374 , n365061 );
buf ( n365063 , n17374 );
buf ( n365064 , n365063 );
not ( n17377 , n365064 );
or ( n17378 , n17371 , n17377 );
buf ( n365067 , n17372 );
buf ( n365068 , n354303 );
nand ( n17381 , n365067 , n365068 );
buf ( n365070 , n17381 );
buf ( n365071 , n365070 );
nand ( n365072 , n17378 , n365071 );
buf ( n365073 , n365072 );
buf ( n365074 , n365073 );
buf ( n365075 , n17182 );
nand ( n17383 , n365074 , n365075 );
buf ( n365077 , n17383 );
buf ( n365078 , n365077 );
nand ( n17385 , n17369 , n365078 );
buf ( n365080 , n17385 );
buf ( n365081 , n365080 );
xor ( n17388 , n365040 , n365081 );
buf ( n365083 , n17037 );
not ( n17390 , n365083 );
xor ( n17391 , n578 , n17172 );
buf ( n365086 , n17391 );
not ( n17393 , n365086 );
or ( n17394 , n17390 , n17393 );
buf ( n365089 , n578 );
not ( n17396 , n365089 );
buf ( n365091 , n17143 );
not ( n17398 , n365091 );
buf ( n365093 , n17398 );
buf ( n365094 , n365093 );
not ( n17401 , n365094 );
or ( n17402 , n17396 , n17401 );
buf ( n365097 , n365093 );
not ( n17404 , n365097 );
buf ( n365099 , n17404 );
buf ( n365100 , n365099 );
buf ( n365101 , n364727 );
nand ( n17408 , n365100 , n365101 );
buf ( n365103 , n17408 );
buf ( n365104 , n365103 );
nand ( n17411 , n17402 , n365104 );
buf ( n365106 , n17411 );
buf ( n365107 , n365106 );
buf ( n365108 , n17082 );
nand ( n17415 , n365107 , n365108 );
buf ( n365110 , n17415 );
buf ( n365111 , n365110 );
nand ( n17418 , n17394 , n365111 );
buf ( n365113 , n17418 );
buf ( n365114 , n365113 );
and ( n17421 , n17388 , n365114 );
and ( n17422 , n365040 , n365081 );
or ( n17423 , n17421 , n17422 );
buf ( n365118 , n17423 );
buf ( n365119 , n365118 );
buf ( n365120 , n17230 );
not ( n17427 , n365120 );
buf ( n365122 , n17325 );
not ( n17429 , n365122 );
or ( n17430 , n17427 , n17429 );
buf ( n365125 , n580 );
not ( n17432 , n365125 );
buf ( n365127 , n8303 );
not ( n17434 , n365127 );
buf ( n365129 , n17434 );
buf ( n365130 , n365129 );
not ( n17437 , n365130 );
or ( n17438 , n17432 , n17437 );
buf ( n365133 , n8303 );
buf ( n365134 , n364896 );
nand ( n17441 , n365133 , n365134 );
buf ( n365136 , n17441 );
buf ( n365137 , n365136 );
nand ( n17444 , n17438 , n365137 );
buf ( n365139 , n17444 );
buf ( n365140 , n365139 );
buf ( n365141 , n17209 );
nand ( n17448 , n365140 , n365141 );
buf ( n365143 , n17448 );
buf ( n365144 , n365143 );
nand ( n17451 , n17430 , n365144 );
buf ( n365146 , n17451 );
buf ( n365147 , n365146 );
xor ( n17454 , n365119 , n365147 );
buf ( n365149 , n364779 );
buf ( n365150 , n365149 );
buf ( n365151 , n365150 );
buf ( n365152 , n365151 );
not ( n365153 , n365152 );
buf ( n365154 , n582 );
not ( n17456 , n365154 );
buf ( n365156 , n12418 );
not ( n17457 , n365156 );
or ( n17458 , n17456 , n17457 );
buf ( n365159 , n364903 );
not ( n17460 , n365159 );
buf ( n365161 , n17460 );
buf ( n365162 , n365161 );
buf ( n365163 , n364797 );
nand ( n17464 , n365162 , n365163 );
buf ( n365165 , n17464 );
buf ( n365166 , n365165 );
nand ( n17467 , n17458 , n365166 );
buf ( n365168 , n17467 );
buf ( n365169 , n365168 );
not ( n17470 , n365169 );
or ( n17471 , n365153 , n17470 );
buf ( n365172 , n582 );
not ( n17473 , n365172 );
buf ( n365174 , n9625 );
not ( n17475 , n365174 );
buf ( n365176 , n17475 );
buf ( n365177 , n365176 );
not ( n17478 , n365177 );
or ( n17479 , n17473 , n17478 );
nand ( n17480 , n9625 , n364797 );
buf ( n365181 , n17480 );
nand ( n17482 , n17479 , n365181 );
buf ( n365183 , n17482 );
buf ( n365184 , n365183 );
buf ( n365185 , n17133 );
nand ( n17486 , n365184 , n365185 );
buf ( n365187 , n17486 );
buf ( n365188 , n365187 );
nand ( n17489 , n17471 , n365188 );
buf ( n365190 , n17489 );
buf ( n365191 , n365190 );
and ( n17492 , n17454 , n365191 );
and ( n17493 , n365119 , n365147 );
or ( n17494 , n17492 , n17493 );
buf ( n365195 , n17494 );
buf ( n365196 , n365195 );
and ( n17497 , n17341 , n365196 );
and ( n17498 , n364980 , n365028 );
or ( n17499 , n17497 , n17498 );
buf ( n365200 , n17499 );
buf ( n365201 , n365200 );
xor ( n17502 , n364921 , n365201 );
xor ( n17503 , n364991 , n365006 );
and ( n17504 , n17503 , n365025 );
and ( n17505 , n364991 , n365006 );
or ( n17506 , n17504 , n17505 );
buf ( n365207 , n17506 );
buf ( n365208 , n365207 );
buf ( n365209 , n364925 );
not ( n17510 , n365209 );
buf ( n365211 , n584 );
not ( n17512 , n365211 );
nand ( n17513 , n14027 , n14045 );
not ( n17514 , n14472 );
and ( n17515 , n17513 , n17514 );
not ( n17516 , n17513 );
and ( n17517 , n17516 , n14472 );
nor ( n17518 , n17515 , n17517 );
buf ( n17519 , n17518 );
not ( n17520 , n17519 );
buf ( n365221 , n17520 );
not ( n365222 , n365221 );
or ( n365223 , n17512 , n365222 );
buf ( n365224 , n17519 );
buf ( n365225 , n364771 );
nand ( n17521 , n365224 , n365225 );
buf ( n365227 , n17521 );
buf ( n365228 , n365227 );
nand ( n17523 , n365223 , n365228 );
buf ( n365230 , n17523 );
buf ( n365231 , n365230 );
not ( n17526 , n365231 );
or ( n17527 , n17510 , n17526 );
buf ( n365234 , n364943 );
buf ( n365235 , n364973 );
nand ( n17530 , n365234 , n365235 );
buf ( n365237 , n17530 );
buf ( n365238 , n365237 );
nand ( n17533 , n17527 , n365238 );
buf ( n365240 , n17533 );
buf ( n365241 , n365240 );
xor ( n17536 , n365208 , n365241 );
buf ( n365243 , n17037 );
not ( n17538 , n365243 );
buf ( n365245 , n364748 );
not ( n17540 , n365245 );
or ( n17541 , n17538 , n17540 );
buf ( n365248 , n578 );
not ( n17543 , n365248 );
buf ( n365250 , n7349 );
not ( n17545 , n365250 );
or ( n17546 , n17543 , n17545 );
not ( n17547 , n7349 );
buf ( n365254 , n17547 );
buf ( n365255 , n364727 );
nand ( n17550 , n365254 , n365255 );
buf ( n365257 , n17550 );
buf ( n365258 , n365257 );
nand ( n17553 , n17546 , n365258 );
buf ( n365260 , n17553 );
buf ( n365261 , n365260 );
buf ( n365262 , n17082 );
nand ( n17557 , n365261 , n365262 );
buf ( n365264 , n17557 );
buf ( n365265 , n365264 );
nand ( n17560 , n17541 , n365265 );
buf ( n365267 , n17560 );
buf ( n365268 , n365267 );
buf ( n365269 , n364779 );
not ( n17564 , n365269 );
buf ( n365271 , n364803 );
not ( n17566 , n365271 );
or ( n17567 , n17564 , n17566 );
buf ( n365274 , n365168 );
buf ( n365275 , n17133 );
nand ( n17570 , n365274 , n365275 );
buf ( n365277 , n17570 );
buf ( n365278 , n365277 );
nand ( n17573 , n17567 , n365278 );
buf ( n365280 , n17573 );
buf ( n365281 , n365280 );
xor ( n17576 , n365268 , n365281 );
buf ( n365283 , n17372 );
buf ( n365284 , n576 );
and ( n17579 , n365283 , n365284 );
buf ( n365286 , n17579 );
buf ( n365287 , n365286 );
buf ( n365288 , n364834 );
not ( n365289 , n365288 );
buf ( n365290 , n364998 );
not ( n365291 , n365290 );
or ( n17581 , n365289 , n365291 );
buf ( n365293 , n365054 );
buf ( n365294 , n17182 );
nand ( n17583 , n365293 , n365294 );
buf ( n365296 , n17583 );
buf ( n365297 , n365296 );
nand ( n17586 , n17581 , n365297 );
buf ( n365299 , n17586 );
buf ( n365300 , n365299 );
xor ( n17589 , n365287 , n365300 );
buf ( n365302 , n17037 );
not ( n17591 , n365302 );
buf ( n365304 , n365260 );
not ( n17593 , n365304 );
or ( n17594 , n17591 , n17593 );
buf ( n365307 , n17391 );
buf ( n365308 , n17082 );
nand ( n17597 , n365307 , n365308 );
buf ( n365310 , n17597 );
buf ( n365311 , n365310 );
nand ( n17600 , n17594 , n365311 );
buf ( n365313 , n17600 );
buf ( n365314 , n365313 );
and ( n17603 , n17589 , n365314 );
and ( n17604 , n365287 , n365300 );
or ( n17605 , n17603 , n17604 );
buf ( n365318 , n17605 );
buf ( n365319 , n365318 );
and ( n17608 , n17576 , n365319 );
and ( n17609 , n365268 , n365281 );
or ( n17610 , n17608 , n17609 );
buf ( n365323 , n17610 );
buf ( n365324 , n365323 );
xor ( n17613 , n17536 , n365324 );
buf ( n365326 , n17613 );
buf ( n365327 , n365326 );
xor ( n17616 , n17502 , n365327 );
buf ( n365329 , n17616 );
buf ( n365330 , n365329 );
buf ( n365331 , n17519 );
buf ( n365332 , n586 );
not ( n17621 , n365332 );
buf ( n365334 , n17621 );
buf ( n365335 , n365334 );
nand ( n17624 , n365331 , n365335 );
buf ( n365337 , n17624 );
not ( n17626 , n365337 );
not ( n17627 , n17519 );
nand ( n17628 , n17627 , n586 );
not ( n17629 , n17628 );
or ( n17630 , n17626 , n17629 );
not ( n17631 , n588 );
and ( n17632 , n587 , n17631 );
not ( n17633 , n587 );
and ( n17634 , n17633 , n588 );
or ( n365347 , n17632 , n17634 );
buf ( n365348 , n365347 );
not ( n365349 , n365348 );
buf ( n365350 , n365349 );
not ( n365351 , n365350 );
nand ( n17635 , n17630 , n365351 );
buf ( n365353 , n364936 );
not ( n365354 , n365353 );
buf ( n365355 , n365354 );
buf ( n365356 , n365355 );
buf ( n365357 , n365334 );
nand ( n17640 , n365356 , n365357 );
buf ( n365359 , n17640 );
buf ( n365360 , n17251 );
not ( n17643 , n365360 );
buf ( n365362 , n17643 );
nand ( n17645 , n365362 , n586 );
nand ( n17646 , n365359 , n17645 );
buf ( n365365 , n586 );
buf ( n365366 , n587 );
and ( n17649 , n365365 , n365366 );
buf ( n365368 , n365347 );
buf ( n365369 , n586 );
buf ( n365370 , n587 );
nor ( n17653 , n365369 , n365370 );
buf ( n365372 , n17653 );
buf ( n365373 , n365372 );
nor ( n17656 , n17649 , n365368 , n365373 );
buf ( n365375 , n17656 );
buf ( n17658 , n365375 );
nand ( n17659 , n17646 , n17658 );
nand ( n17660 , n17635 , n17659 );
buf ( n365379 , n17660 );
buf ( n365380 , n365151 );
not ( n17663 , n365380 );
buf ( n365382 , n365183 );
not ( n17665 , n365382 );
or ( n17666 , n17663 , n17665 );
not ( n17667 , n582 );
buf ( n365386 , n8990 );
not ( n17669 , n365386 );
buf ( n365388 , n17669 );
not ( n17671 , n365388 );
or ( n17672 , n17667 , n17671 );
buf ( n365391 , n8990 );
buf ( n365392 , n364797 );
nand ( n17675 , n365391 , n365392 );
buf ( n365394 , n17675 );
nand ( n17677 , n17672 , n365394 );
nand ( n17678 , n17677 , n17133 );
buf ( n365397 , n17678 );
nand ( n17680 , n17666 , n365397 );
buf ( n365399 , n17680 );
buf ( n365400 , n365399 );
buf ( n365401 , n17021 );
buf ( n365402 , n365401 );
buf ( n365403 , n365402 );
buf ( n365404 , n364925 );
not ( n365405 , n365404 );
buf ( n365406 , n365405 );
buf ( n365407 , n365406 );
buf ( n365408 , n364771 );
nor ( n17685 , n365407 , n365408 );
buf ( n365410 , n17685 );
not ( n17687 , n365410 );
nor ( n17688 , n365403 , n17687 );
not ( n17689 , n17688 );
buf ( n365414 , n584 );
not ( n17691 , n365414 );
buf ( n365416 , n364903 );
not ( n17693 , n365416 );
or ( n17694 , n17691 , n17693 );
buf ( n365419 , n360086 );
buf ( n365420 , n364771 );
nand ( n17697 , n365419 , n365420 );
buf ( n365422 , n17697 );
buf ( n365423 , n365422 );
nand ( n17700 , n17694 , n365423 );
buf ( n365425 , n17700 );
nand ( n17702 , n365425 , n364973 );
buf ( n365427 , n365406 );
buf ( n365428 , n584 );
nor ( n17705 , n365427 , n365428 );
buf ( n365430 , n17705 );
nand ( n17707 , n365403 , n365430 );
nand ( n17708 , n17689 , n17702 , n17707 );
buf ( n365433 , n17708 );
xor ( n17710 , n365400 , n365433 );
buf ( n365435 , n17230 );
not ( n17712 , n365435 );
buf ( n365437 , n580 );
not ( n17714 , n365437 );
buf ( n365439 , n7349 );
not ( n17716 , n365439 );
or ( n17717 , n17714 , n17716 );
buf ( n365442 , n7348 );
buf ( n365443 , n364896 );
nand ( n17720 , n365442 , n365443 );
buf ( n365445 , n17720 );
buf ( n365446 , n365445 );
nand ( n17723 , n17717 , n365446 );
buf ( n365448 , n17723 );
buf ( n365449 , n365448 );
not ( n365450 , n365449 );
or ( n365451 , n17712 , n365450 );
buf ( n365452 , n580 );
not ( n365453 , n365452 );
not ( n17725 , n17172 );
buf ( n365455 , n17725 );
not ( n365456 , n365455 );
or ( n17727 , n365453 , n365456 );
buf ( n365458 , n17174 );
buf ( n365459 , n364896 );
nand ( n17730 , n365458 , n365459 );
buf ( n365461 , n17730 );
buf ( n365462 , n365461 );
nand ( n17733 , n17727 , n365462 );
buf ( n365464 , n17733 );
buf ( n365465 , n365464 );
buf ( n365466 , n364885 );
nand ( n17737 , n365465 , n365466 );
buf ( n365468 , n17737 );
buf ( n365469 , n365468 );
nand ( n17740 , n365451 , n365469 );
buf ( n365471 , n17740 );
buf ( n365472 , n365471 );
buf ( n365473 , n12481 );
not ( n17744 , n365473 );
buf ( n365475 , n17744 );
buf ( n365476 , n365475 );
buf ( n365477 , n354303 );
nor ( n17748 , n365476 , n365477 );
buf ( n365479 , n17748 );
buf ( n365480 , n365479 );
buf ( n365481 , n364834 );
not ( n17752 , n365481 );
and ( n17753 , n365035 , n354303 );
not ( n17754 , n365035 );
and ( n17755 , n17754 , n576 );
or ( n17756 , n17753 , n17755 );
buf ( n365487 , n17756 );
not ( n17758 , n365487 );
or ( n17759 , n17752 , n17758 );
buf ( n365490 , n576 );
nand ( n365491 , n3585 , n3586 );
buf ( n365492 , n365491 );
not ( n365493 , n365492 );
buf ( n365494 , n365493 );
buf ( n365495 , n365494 );
not ( n17761 , n365495 );
buf ( n365497 , n17761 );
buf ( n365498 , n365497 );
xor ( n17763 , n365490 , n365498 );
buf ( n365500 , n17763 );
buf ( n365501 , n365500 );
buf ( n365502 , n17182 );
nand ( n17767 , n365501 , n365502 );
buf ( n365504 , n17767 );
buf ( n365505 , n365504 );
nand ( n17770 , n17759 , n365505 );
buf ( n365507 , n17770 );
buf ( n365508 , n365507 );
xor ( n17773 , n365480 , n365508 );
buf ( n365510 , n17037 );
not ( n17775 , n365510 );
buf ( n365512 , n578 );
not ( n17777 , n365512 );
buf ( n365514 , n17301 );
not ( n17779 , n365514 );
buf ( n365516 , n17779 );
buf ( n365517 , n365516 );
not ( n17782 , n365517 );
or ( n17783 , n17777 , n17782 );
buf ( n365520 , n364986 );
not ( n17785 , n365520 );
buf ( n365522 , n364727 );
nand ( n17787 , n17785 , n365522 );
buf ( n365524 , n17787 );
buf ( n365525 , n365524 );
nand ( n17790 , n17783 , n365525 );
buf ( n365527 , n17790 );
buf ( n365528 , n365527 );
not ( n365529 , n365528 );
or ( n365530 , n17775 , n365529 );
buf ( n365531 , n578 );
not ( n17791 , n365531 );
buf ( n365533 , n365063 );
not ( n365534 , n365533 );
or ( n17793 , n17791 , n365534 );
buf ( n365536 , n17372 );
buf ( n365537 , n364727 );
nand ( n17796 , n365536 , n365537 );
buf ( n365539 , n17796 );
buf ( n365540 , n365539 );
nand ( n17799 , n17793 , n365540 );
buf ( n365542 , n17799 );
buf ( n365543 , n365542 );
buf ( n365544 , n17082 );
nand ( n17803 , n365543 , n365544 );
buf ( n365546 , n17803 );
buf ( n365547 , n365546 );
nand ( n17806 , n365530 , n365547 );
buf ( n365549 , n17806 );
buf ( n365550 , n365549 );
and ( n17809 , n17773 , n365550 );
and ( n17810 , n365480 , n365508 );
or ( n17811 , n17809 , n17810 );
buf ( n365554 , n17811 );
buf ( n365555 , n365554 );
xor ( n17814 , n365472 , n365555 );
and ( n365557 , n365490 , n365498 );
buf ( n365558 , n365557 );
buf ( n365559 , n365558 );
buf ( n365560 , n364834 );
not ( n365561 , n365560 );
buf ( n365562 , n365073 );
not ( n17816 , n365562 );
or ( n365564 , n365561 , n17816 );
buf ( n365565 , n17756 );
buf ( n365566 , n17182 );
nand ( n17819 , n365565 , n365566 );
buf ( n365568 , n17819 );
buf ( n365569 , n365568 );
nand ( n17822 , n365564 , n365569 );
buf ( n365571 , n17822 );
buf ( n365572 , n365571 );
xor ( n17825 , n365559 , n365572 );
buf ( n365574 , n17037 );
not ( n17827 , n365574 );
buf ( n365576 , n365106 );
not ( n17829 , n365576 );
or ( n17830 , n17827 , n17829 );
buf ( n365579 , n365527 );
buf ( n365580 , n17082 );
nand ( n365581 , n365579 , n365580 );
buf ( n365582 , n365581 );
buf ( n365583 , n365582 );
nand ( n365584 , n17830 , n365583 );
buf ( n365585 , n365584 );
buf ( n365586 , n365585 );
xor ( n17834 , n17825 , n365586 );
buf ( n365588 , n17834 );
buf ( n365589 , n365588 );
and ( n17836 , n17814 , n365589 );
and ( n17837 , n365472 , n365555 );
or ( n17838 , n17836 , n17837 );
buf ( n365593 , n17838 );
buf ( n365594 , n365593 );
and ( n17841 , n17710 , n365594 );
and ( n17842 , n365400 , n365433 );
or ( n17843 , n17841 , n17842 );
buf ( n365598 , n17843 );
buf ( n365599 , n365598 );
xor ( n365600 , n365379 , n365599 );
xor ( n365601 , n365119 , n365147 );
xor ( n365602 , n365601 , n365191 );
buf ( n365603 , n365602 );
buf ( n365604 , n365603 );
and ( n17846 , n365600 , n365604 );
and ( n365606 , n365379 , n365599 );
or ( n17847 , n17846 , n365606 );
buf ( n365608 , n17847 );
buf ( n365609 , n365608 );
not ( n17850 , n365337 );
not ( n365611 , n17628 );
or ( n365612 , n17850 , n365611 );
nand ( n365613 , n365612 , n365375 );
buf ( n365614 , n16900 );
not ( n365615 , n365614 );
buf ( n365616 , n365350 );
buf ( n365617 , n365334 );
nor ( n365618 , n365616 , n365617 );
buf ( n365619 , n365618 );
buf ( n365620 , n365619 );
nand ( n365621 , n365615 , n365620 );
buf ( n365622 , n365621 );
buf ( n365623 , n16900 );
buf ( n365624 , n365350 );
buf ( n365625 , n586 );
nor ( n365626 , n365624 , n365625 );
buf ( n365627 , n365626 );
buf ( n365628 , n365627 );
nand ( n17859 , n365623 , n365628 );
buf ( n365630 , n17859 );
nand ( n17861 , n365613 , n365622 , n365630 );
buf ( n365632 , n17861 );
and ( n17863 , n589 , n347697 );
not ( n365634 , n589 );
and ( n17865 , n365634 , n590 );
or ( n365636 , n17863 , n17865 );
buf ( n17867 , n365636 );
not ( n365638 , n17867 );
and ( n17869 , n588 , n589 );
buf ( n365640 , n588 );
buf ( n365641 , n589 );
nor ( n365642 , n365640 , n365641 );
buf ( n365643 , n365642 );
nor ( n365644 , n17869 , n365643 );
nand ( n17875 , n365638 , n365644 );
not ( n365646 , n17875 );
buf ( n365647 , n365646 );
not ( n365648 , n365647 );
buf ( n365649 , n588 );
not ( n365650 , n365649 );
buf ( n365651 , n16955 );
not ( n365652 , n365651 );
buf ( n365653 , n365652 );
buf ( n365654 , n365653 );
not ( n17885 , n365654 );
or ( n365656 , n365650 , n17885 );
buf ( n365657 , n588 );
not ( n365658 , n365657 );
buf ( n365659 , n365653 );
not ( n365660 , n365659 );
buf ( n365661 , n365660 );
buf ( n365662 , n365661 );
nand ( n17893 , n365658 , n365662 );
buf ( n365664 , n17893 );
buf ( n365665 , n365664 );
nand ( n365666 , n365656 , n365665 );
buf ( n365667 , n365666 );
buf ( n365668 , n365667 );
not ( n17899 , n365668 );
or ( n365670 , n365648 , n17899 );
not ( n17901 , n17631 );
not ( n365672 , n16927 );
not ( n17903 , n16998 );
or ( n365674 , n365672 , n17903 );
nand ( n17905 , n365674 , n17001 );
not ( n365676 , n17905 );
or ( n17907 , n17901 , n365676 );
or ( n365678 , n17002 , n17631 );
nand ( n17909 , n17907 , n365678 );
buf ( n365680 , n17909 );
buf ( n365681 , n17867 );
nand ( n365682 , n365680 , n365681 );
buf ( n365683 , n365682 );
buf ( n365684 , n365683 );
nand ( n17915 , n365670 , n365684 );
buf ( n365686 , n17915 );
buf ( n365687 , n365686 );
xor ( n365688 , n365632 , n365687 );
xor ( n17919 , n365268 , n365281 );
xor ( n365690 , n17919 , n365319 );
buf ( n365691 , n365690 );
buf ( n365692 , n365691 );
xor ( n17923 , n365688 , n365692 );
buf ( n365694 , n17923 );
buf ( n365695 , n365694 );
xor ( n365696 , n365609 , n365695 );
buf ( n365697 , n591 );
not ( n365698 , n365697 );
not ( n17929 , n16880 );
not ( n365700 , n16874 );
or ( n17931 , n17929 , n365700 );
nand ( n365702 , n17931 , n16883 );
not ( n17933 , n365702 );
xor ( n365704 , n590 , n17933 );
buf ( n365705 , n365704 );
not ( n365706 , n365705 );
or ( n17937 , n365698 , n365706 );
buf ( n365708 , n590 );
not ( n17939 , n365708 );
buf ( n365710 , n17002 );
not ( n17941 , n365710 );
buf ( n365712 , n17941 );
buf ( n365713 , n365712 );
not ( n365714 , n365713 );
or ( n17945 , n17939 , n365714 );
buf ( n365716 , n590 );
not ( n17947 , n365716 );
buf ( n365718 , n17905 );
nand ( n17949 , n17947 , n365718 );
buf ( n365720 , n17949 );
buf ( n365721 , n365720 );
nand ( n365722 , n17945 , n365721 );
buf ( n365723 , n365722 );
buf ( n365724 , n365723 );
buf ( n365725 , n590 );
not ( n365726 , n365725 );
buf ( n365727 , n591 );
nor ( n365728 , n365726 , n365727 );
buf ( n365729 , n365728 );
buf ( n365730 , n365729 );
buf ( n17961 , n365730 );
buf ( n365732 , n17961 );
buf ( n365733 , n365732 );
buf ( n365734 , n365733 );
buf ( n365735 , n365734 );
buf ( n365736 , n365735 );
buf ( n17967 , n365736 );
buf ( n365738 , n17967 );
buf ( n365739 , n365738 );
nand ( n365740 , n365724 , n365739 );
buf ( n365741 , n365740 );
buf ( n365742 , n365741 );
nand ( n17973 , n17937 , n365742 );
buf ( n365744 , n17973 );
buf ( n365745 , n365744 );
buf ( n365746 , n365646 );
not ( n17977 , n365746 );
not ( n365748 , n16900 );
and ( n17979 , n588 , n365748 );
not ( n365750 , n588 );
and ( n17981 , n365750 , n16900 );
or ( n365752 , n17979 , n17981 );
buf ( n365753 , n365752 );
not ( n365754 , n365753 );
or ( n17985 , n17977 , n365754 );
buf ( n365756 , n365667 );
buf ( n365757 , n17867 );
nand ( n365758 , n365756 , n365757 );
buf ( n365759 , n365758 );
buf ( n365760 , n365759 );
nand ( n17991 , n17985 , n365760 );
buf ( n365762 , n17991 );
buf ( n365763 , n365762 );
xor ( n365764 , n365745 , n365763 );
xor ( n17995 , n365287 , n365300 );
xor ( n365766 , n17995 , n365314 );
buf ( n365767 , n365766 );
buf ( n365768 , n365767 );
buf ( n365769 , n364925 );
not ( n365770 , n365769 );
buf ( n365771 , n364961 );
not ( n365772 , n365771 );
or ( n18003 , n365770 , n365772 );
buf ( n365774 , n365403 );
not ( n18005 , n365774 );
buf ( n365776 , n18005 );
buf ( n365777 , n365776 );
buf ( n365778 , n584 );
nand ( n18009 , n365777 , n365778 );
buf ( n365780 , n18009 );
buf ( n365781 , n365780 );
not ( n365782 , n365781 );
buf ( n365783 , n365403 );
buf ( n365784 , n364771 );
nand ( n18015 , n365783 , n365784 );
buf ( n365786 , n18015 );
buf ( n365787 , n365786 );
not ( n365788 , n365787 );
or ( n18019 , n365782 , n365788 );
buf ( n365790 , n364973 );
nand ( n18021 , n18019 , n365790 );
buf ( n365792 , n18021 );
buf ( n365793 , n365792 );
nand ( n365794 , n18003 , n365793 );
buf ( n365795 , n365794 );
buf ( n365796 , n365795 );
xor ( n18027 , n365768 , n365796 );
xor ( n365798 , n365559 , n365572 );
and ( n18029 , n365798 , n365586 );
and ( n365800 , n365559 , n365572 );
or ( n18031 , n18029 , n365800 );
buf ( n365802 , n18031 );
buf ( n365803 , n365802 );
xor ( n365804 , n365040 , n365081 );
xor ( n18035 , n365804 , n365114 );
buf ( n365806 , n18035 );
buf ( n365807 , n365806 );
xor ( n365808 , n365803 , n365807 );
buf ( n365809 , n17230 );
not ( n365810 , n365809 );
buf ( n365811 , n365139 );
not ( n365812 , n365811 );
or ( n18043 , n365810 , n365812 );
buf ( n365814 , n365448 );
buf ( n365815 , n17209 );
nand ( n365816 , n365814 , n365815 );
buf ( n365817 , n365816 );
buf ( n365818 , n365817 );
nand ( n18049 , n18043 , n365818 );
buf ( n365820 , n18049 );
buf ( n365821 , n365820 );
and ( n365822 , n365808 , n365821 );
and ( n18053 , n365803 , n365807 );
or ( n365824 , n365822 , n18053 );
buf ( n365825 , n365824 );
buf ( n365826 , n365825 );
xor ( n18057 , n18027 , n365826 );
buf ( n365828 , n18057 );
buf ( n365829 , n365828 );
and ( n365830 , n365764 , n365829 );
and ( n18061 , n365745 , n365763 );
or ( n365832 , n365830 , n18061 );
buf ( n365833 , n365832 );
buf ( n365834 , n365833 );
and ( n18065 , n365696 , n365834 );
and ( n365836 , n365609 , n365695 );
or ( n18067 , n18065 , n365836 );
buf ( n365838 , n18067 );
buf ( n365839 , n365838 );
xor ( n365840 , n365330 , n365839 );
xor ( n18071 , n365632 , n365687 );
and ( n365842 , n18071 , n365692 );
and ( n18073 , n365632 , n365687 );
or ( n365844 , n365842 , n18073 );
buf ( n365845 , n365844 );
buf ( n365846 , n365845 );
buf ( n365847 , n365375 );
not ( n365848 , n365847 );
and ( n18079 , n16900 , n365334 );
not ( n365850 , n16900 );
and ( n18081 , n365850 , n586 );
or ( n365852 , n18079 , n18081 );
buf ( n365853 , n365852 );
not ( n365854 , n365853 );
or ( n18085 , n365848 , n365854 );
buf ( n365856 , n365334 );
not ( n18087 , n365856 );
buf ( n365858 , n16955 );
not ( n18089 , n365858 );
or ( n365860 , n18087 , n18089 );
buf ( n365861 , n365653 );
buf ( n365862 , n586 );
nand ( n18093 , n365861 , n365862 );
buf ( n365864 , n18093 );
buf ( n365865 , n365864 );
nand ( n365866 , n365860 , n365865 );
buf ( n365867 , n365866 );
buf ( n365868 , n365867 );
buf ( n365869 , n365351 );
nand ( n365870 , n365868 , n365869 );
buf ( n365871 , n365870 );
buf ( n365872 , n365871 );
nand ( n18103 , n18085 , n365872 );
buf ( n365874 , n18103 );
buf ( n365875 , n365874 );
not ( n365876 , n17867 );
not ( n365877 , n16884 );
not ( n365878 , n365877 );
and ( n365879 , n588 , n365878 );
not ( n365880 , n588 );
not ( n365881 , n365702 );
and ( n365882 , n365880 , n365881 );
or ( n365883 , n365879 , n365882 );
not ( n365884 , n365883 );
or ( n365885 , n365876 , n365884 );
nand ( n365886 , n17909 , n365646 );
nand ( n365887 , n365885 , n365886 );
buf ( n365888 , n365887 );
xor ( n365889 , n365875 , n365888 );
buf ( n365890 , n591 );
not ( n365891 , n365890 );
buf ( n365892 , n16841 );
xor ( n365893 , n590 , n365892 );
buf ( n365894 , n365893 );
not ( n365895 , n365894 );
or ( n365896 , n365891 , n365895 );
buf ( n365897 , n16854 );
and ( n365898 , n365897 , n590 );
not ( n365899 , n365897 );
and ( n365900 , n365899 , n348597 );
nor ( n365901 , n365898 , n365900 );
buf ( n365902 , n365901 );
buf ( n365903 , n365738 );
nand ( n365904 , n365902 , n365903 );
buf ( n365905 , n365904 );
buf ( n365906 , n365905 );
nand ( n18130 , n365896 , n365906 );
buf ( n365908 , n18130 );
buf ( n365909 , n365908 );
xor ( n18133 , n365889 , n365909 );
buf ( n365911 , n18133 );
buf ( n365912 , n365911 );
xor ( n365913 , n365846 , n365912 );
not ( n18137 , n591 );
not ( n18138 , n365901 );
or ( n365916 , n18137 , n18138 );
buf ( n365917 , n365704 );
buf ( n365918 , n365738 );
nand ( n18142 , n365917 , n365918 );
buf ( n365920 , n18142 );
nand ( n365921 , n365916 , n365920 );
buf ( n365922 , n365921 );
xor ( n18146 , n365768 , n365796 );
and ( n365924 , n18146 , n365826 );
and ( n365925 , n365768 , n365796 );
or ( n18149 , n365924 , n365925 );
buf ( n365927 , n18149 );
buf ( n365928 , n365927 );
xor ( n365929 , n365922 , n365928 );
xor ( n18153 , n364980 , n365028 );
xor ( n18154 , n18153 , n365196 );
buf ( n365932 , n18154 );
buf ( n365933 , n365932 );
and ( n18157 , n365929 , n365933 );
and ( n18158 , n365922 , n365928 );
or ( n365936 , n18157 , n18158 );
buf ( n365937 , n365936 );
buf ( n365938 , n365937 );
xor ( n18162 , n365913 , n365938 );
buf ( n365940 , n18162 );
buf ( n365941 , n365940 );
xor ( n18165 , n365840 , n365941 );
buf ( n365943 , n18165 );
buf ( n365944 , n365943 );
buf ( n365945 , n365944 );
buf ( n365946 , n365945 );
not ( n18170 , n365946 );
xor ( n365948 , n365922 , n365928 );
xor ( n365949 , n365948 , n365933 );
buf ( n365950 , n365949 );
buf ( n365951 , n365950 );
not ( n365952 , n17658 );
buf ( n365953 , n586 );
not ( n18177 , n365953 );
buf ( n365955 , n364951 );
not ( n365956 , n365955 );
or ( n365957 , n18177 , n365956 );
buf ( n365958 , n14498 );
buf ( n365959 , n365334 );
nand ( n365960 , n365958 , n365959 );
buf ( n365961 , n365960 );
buf ( n365962 , n365961 );
nand ( n18186 , n365957 , n365962 );
buf ( n365964 , n18186 );
not ( n365965 , n365964 );
or ( n18189 , n365952 , n365965 );
not ( n18190 , n17645 );
not ( n365968 , n365359 );
or ( n365969 , n18190 , n365968 );
nand ( n18193 , n365969 , n365351 );
nand ( n18194 , n18189 , n18193 );
buf ( n365972 , n18194 );
xor ( n365973 , n365803 , n365807 );
xor ( n18197 , n365973 , n365821 );
buf ( n365975 , n18197 );
buf ( n365976 , n365975 );
xor ( n365977 , n365972 , n365976 );
buf ( n365978 , n364973 );
not ( n18202 , n365978 );
buf ( n365980 , n584 );
not ( n365981 , n365980 );
buf ( n365982 , n364891 );
not ( n18206 , n365982 );
or ( n365984 , n365981 , n18206 );
buf ( n365985 , n9625 );
buf ( n365986 , n364771 );
nand ( n18210 , n365985 , n365986 );
buf ( n365988 , n18210 );
buf ( n365989 , n365988 );
nand ( n18213 , n365984 , n365989 );
buf ( n365991 , n18213 );
buf ( n365992 , n365991 );
not ( n365993 , n365992 );
or ( n18217 , n18202 , n365993 );
buf ( n365995 , n365425 );
buf ( n365996 , n364925 );
nand ( n365997 , n365995 , n365996 );
buf ( n365998 , n365997 );
buf ( n365999 , n365998 );
nand ( n366000 , n18217 , n365999 );
buf ( n366001 , n366000 );
buf ( n366002 , n366001 );
not ( n18226 , n364779 );
not ( n366004 , n17677 );
or ( n366005 , n18226 , n366004 );
buf ( n366006 , n582 );
not ( n18230 , n366006 );
buf ( n366008 , n365129 );
not ( n366009 , n366008 );
or ( n18233 , n18230 , n366009 );
buf ( n366011 , n8303 );
buf ( n366012 , n364797 );
nand ( n366013 , n366011 , n366012 );
buf ( n366014 , n366013 );
buf ( n366015 , n366014 );
nand ( n366016 , n18233 , n366015 );
buf ( n366017 , n366016 );
buf ( n366018 , n366017 );
buf ( n366019 , n17133 );
nand ( n366020 , n366018 , n366019 );
buf ( n366021 , n366020 );
nand ( n18245 , n366005 , n366021 );
buf ( n366023 , n18245 );
xor ( n18247 , n366002 , n366023 );
buf ( n18248 , n3560 );
buf ( n366026 , n18248 );
buf ( n18250 , n366026 );
buf ( n366028 , n18250 );
buf ( n366029 , n366028 );
buf ( n366030 , n576 );
and ( n18254 , n366029 , n366030 );
buf ( n366032 , n18254 );
buf ( n366033 , n366032 );
buf ( n366034 , n364834 );
not ( n18258 , n366034 );
buf ( n366036 , n365500 );
not ( n18260 , n366036 );
or ( n18261 , n18258 , n18260 );
buf ( n366039 , n576 );
not ( n18263 , n366039 );
buf ( n366041 , n12481 );
not ( n18265 , n366041 );
buf ( n366043 , n18265 );
buf ( n366044 , n366043 );
not ( n18268 , n366044 );
or ( n18269 , n18263 , n18268 );
buf ( n366047 , n366043 );
not ( n18271 , n366047 );
buf ( n366049 , n18271 );
buf ( n366050 , n366049 );
buf ( n366051 , n354303 );
nand ( n18275 , n366050 , n366051 );
buf ( n366053 , n18275 );
buf ( n366054 , n366053 );
nand ( n18278 , n18269 , n366054 );
buf ( n366056 , n18278 );
buf ( n366057 , n366056 );
buf ( n366058 , n17182 );
nand ( n18282 , n366057 , n366058 );
buf ( n366060 , n18282 );
buf ( n366061 , n366060 );
nand ( n18285 , n18261 , n366061 );
buf ( n366063 , n18285 );
buf ( n366064 , n366063 );
xor ( n18288 , n366033 , n366064 );
buf ( n366066 , n17037 );
not ( n18290 , n366066 );
buf ( n366068 , n365542 );
not ( n18292 , n366068 );
or ( n18293 , n18290 , n18292 );
buf ( n366071 , n578 );
not ( n18295 , n366071 );
buf ( n366073 , n365032 );
not ( n18297 , n366073 );
or ( n18298 , n18295 , n18297 );
buf ( n366076 , n12483 );
buf ( n366077 , n364727 );
nand ( n18301 , n366076 , n366077 );
buf ( n366079 , n18301 );
buf ( n366080 , n366079 );
nand ( n18304 , n18298 , n366080 );
buf ( n366082 , n18304 );
buf ( n366083 , n366082 );
buf ( n366084 , n17082 );
nand ( n18308 , n366083 , n366084 );
buf ( n366086 , n18308 );
buf ( n366087 , n366086 );
nand ( n18311 , n18293 , n366087 );
buf ( n366089 , n18311 );
buf ( n366090 , n366089 );
and ( n18314 , n18288 , n366090 );
and ( n18315 , n366033 , n366064 );
or ( n18316 , n18314 , n18315 );
buf ( n366094 , n18316 );
buf ( n366095 , n366094 );
buf ( n366096 , n17230 );
not ( n18320 , n366096 );
buf ( n366098 , n365464 );
not ( n18322 , n366098 );
or ( n18323 , n18320 , n18322 );
buf ( n366101 , n580 );
not ( n18325 , n366101 );
buf ( n366103 , n365093 );
not ( n18327 , n366103 );
or ( n18328 , n18325 , n18327 );
buf ( n366106 , n17143 );
buf ( n366107 , n364896 );
nand ( n18331 , n366106 , n366107 );
buf ( n366109 , n18331 );
buf ( n366110 , n366109 );
nand ( n18334 , n18328 , n366110 );
buf ( n366112 , n18334 );
buf ( n366113 , n366112 );
buf ( n366114 , n364885 );
nand ( n18338 , n366113 , n366114 );
buf ( n366116 , n18338 );
buf ( n366117 , n366116 );
nand ( n366118 , n18323 , n366117 );
buf ( n366119 , n366118 );
buf ( n366120 , n366119 );
xor ( n366121 , n366095 , n366120 );
buf ( n366122 , n12482 );
not ( n366123 , n366122 );
buf ( n366124 , n366123 );
buf ( n366125 , n366124 );
buf ( n366126 , n366125 );
buf ( n366127 , n366126 );
buf ( n366128 , n366127 );
not ( n366129 , n366128 );
buf ( n366130 , n366129 );
buf ( n366131 , n366130 );
buf ( n366132 , n576 );
and ( n366133 , n366131 , n366132 );
buf ( n366134 , n366133 );
buf ( n366135 , n366134 );
buf ( n366136 , n364834 );
not ( n366137 , n366136 );
buf ( n366138 , n366056 );
not ( n366139 , n366138 );
or ( n366140 , n366137 , n366139 );
buf ( n366141 , n576 );
not ( n366142 , n366141 );
buf ( n366143 , n366028 );
not ( n366144 , n366143 );
buf ( n366145 , n366144 );
buf ( n366146 , n366145 );
not ( n366147 , n366146 );
or ( n366148 , n366142 , n366147 );
buf ( n366149 , n366028 );
buf ( n366150 , n354303 );
nand ( n366151 , n366149 , n366150 );
buf ( n366152 , n366151 );
buf ( n366153 , n366152 );
nand ( n366154 , n366148 , n366153 );
buf ( n366155 , n366154 );
buf ( n366156 , n366155 );
buf ( n366157 , n17182 );
nand ( n366158 , n366156 , n366157 );
buf ( n366159 , n366158 );
buf ( n366160 , n366159 );
nand ( n366161 , n366140 , n366160 );
buf ( n366162 , n366161 );
buf ( n366163 , n366162 );
xor ( n366164 , n366135 , n366163 );
buf ( n366165 , n17037 );
not ( n366166 , n366165 );
buf ( n366167 , n366082 );
not ( n366168 , n366167 );
or ( n366169 , n366166 , n366168 );
buf ( n366170 , n578 );
not ( n366171 , n366170 );
buf ( n366172 , n365494 );
not ( n366173 , n366172 );
or ( n366174 , n366171 , n366173 );
buf ( n366175 , n365491 );
buf ( n366176 , n364727 );
nand ( n366177 , n366175 , n366176 );
buf ( n366178 , n366177 );
buf ( n366179 , n366178 );
nand ( n366180 , n366174 , n366179 );
buf ( n366181 , n366180 );
buf ( n366182 , n366181 );
buf ( n366183 , n17082 );
nand ( n366184 , n366182 , n366183 );
buf ( n366185 , n366184 );
buf ( n366186 , n366185 );
nand ( n366187 , n366169 , n366186 );
buf ( n366188 , n366187 );
buf ( n366189 , n366188 );
and ( n366190 , n366164 , n366189 );
and ( n366191 , n366135 , n366163 );
or ( n366192 , n366190 , n366191 );
buf ( n366193 , n366192 );
buf ( n366194 , n366193 );
buf ( n366195 , n17230 );
not ( n366196 , n366195 );
buf ( n366197 , n366112 );
not ( n366198 , n366197 );
or ( n366199 , n366196 , n366198 );
buf ( n366200 , n580 );
not ( n366201 , n366200 );
buf ( n366202 , n365516 );
not ( n366203 , n366202 );
or ( n366204 , n366201 , n366203 );
buf ( n366205 , n17301 );
buf ( n366206 , n364896 );
nand ( n366207 , n366205 , n366206 );
buf ( n366208 , n366207 );
buf ( n366209 , n366208 );
nand ( n366210 , n366204 , n366209 );
buf ( n366211 , n366210 );
buf ( n366212 , n366211 );
buf ( n366213 , n364885 );
nand ( n366214 , n366212 , n366213 );
buf ( n366215 , n366214 );
buf ( n366216 , n366215 );
nand ( n366217 , n366199 , n366216 );
buf ( n366218 , n366217 );
buf ( n366219 , n366218 );
xor ( n366220 , n366194 , n366219 );
xor ( n366221 , n366033 , n366064 );
xor ( n366222 , n366221 , n366090 );
buf ( n366223 , n366222 );
buf ( n366224 , n366223 );
and ( n366225 , n366220 , n366224 );
and ( n366226 , n366194 , n366219 );
or ( n366227 , n366225 , n366226 );
buf ( n366228 , n366227 );
buf ( n366229 , n366228 );
and ( n366230 , n366121 , n366229 );
and ( n366231 , n366095 , n366120 );
or ( n366232 , n366230 , n366231 );
buf ( n366233 , n366232 );
buf ( n366234 , n366233 );
and ( n366235 , n18247 , n366234 );
and ( n366236 , n366002 , n366023 );
or ( n366237 , n366235 , n366236 );
buf ( n366238 , n366237 );
buf ( n366239 , n366238 );
and ( n366240 , n365977 , n366239 );
and ( n366241 , n365972 , n365976 );
or ( n366242 , n366240 , n366241 );
buf ( n366243 , n366242 );
buf ( n366244 , n366243 );
xor ( n366245 , n365379 , n365599 );
xor ( n366246 , n366245 , n365604 );
buf ( n366247 , n366246 );
buf ( n366248 , n366247 );
xor ( n366249 , n366244 , n366248 );
buf ( n366250 , n17867 );
not ( n366251 , n366250 );
buf ( n366252 , n365752 );
not ( n366253 , n366252 );
or ( n366254 , n366251 , n366253 );
not ( n366255 , n17519 );
and ( n366256 , n588 , n366255 );
not ( n366257 , n588 );
and ( n366258 , n366257 , n17519 );
or ( n366259 , n366256 , n366258 );
buf ( n366260 , n366259 );
buf ( n366261 , n365646 );
nand ( n366262 , n366260 , n366261 );
buf ( n366263 , n366262 );
buf ( n366264 , n366263 );
nand ( n366265 , n366254 , n366264 );
buf ( n366266 , n366265 );
buf ( n366267 , n366266 );
xor ( n366268 , n365400 , n365433 );
xor ( n366269 , n366268 , n365594 );
buf ( n366270 , n366269 );
buf ( n366271 , n366270 );
xor ( n366272 , n366267 , n366271 );
buf ( n366273 , n365738 );
not ( n366274 , n366273 );
buf ( n366275 , n365653 );
not ( n366276 , n366275 );
buf ( n366277 , n366276 );
xor ( n366278 , n590 , n366277 );
buf ( n366279 , n366278 );
not ( n366280 , n366279 );
or ( n366281 , n366274 , n366280 );
buf ( n366282 , n365723 );
buf ( n366283 , n591 );
nand ( n366284 , n366282 , n366283 );
buf ( n366285 , n366284 );
buf ( n366286 , n366285 );
nand ( n366287 , n366281 , n366286 );
buf ( n366288 , n366287 );
buf ( n366289 , n366288 );
and ( n366290 , n366272 , n366289 );
and ( n366291 , n366267 , n366271 );
or ( n366292 , n366290 , n366291 );
buf ( n366293 , n366292 );
buf ( n366294 , n366293 );
and ( n366295 , n366249 , n366294 );
and ( n366296 , n366244 , n366248 );
or ( n366297 , n366295 , n366296 );
buf ( n366298 , n366297 );
buf ( n366299 , n366298 );
xor ( n366300 , n365951 , n366299 );
xor ( n366301 , n365609 , n365695 );
xor ( n366302 , n366301 , n365834 );
buf ( n366303 , n366302 );
buf ( n366304 , n366303 );
and ( n366305 , n366300 , n366304 );
and ( n366306 , n365951 , n366299 );
or ( n366307 , n366305 , n366306 );
buf ( n366308 , n366307 );
not ( n366309 , n366308 );
nand ( n18533 , n18170 , n366309 );
buf ( n366311 , n365946 );
buf ( n366312 , n366308 );
nand ( n366313 , n366311 , n366312 );
buf ( n366314 , n366313 );
nand ( n18538 , n18533 , n366314 );
not ( n366316 , n18538 );
not ( n366317 , n366316 );
xor ( n18541 , n365951 , n366299 );
xor ( n18542 , n18541 , n366304 );
buf ( n366320 , n18542 );
xor ( n366321 , n365745 , n365763 );
xor ( n18545 , n366321 , n365829 );
buf ( n366323 , n18545 );
buf ( n366324 , n366323 );
buf ( n366325 , n365351 );
not ( n18549 , n366325 );
buf ( n366327 , n365964 );
not ( n366328 , n366327 );
or ( n366329 , n18549 , n366328 );
and ( n18553 , n17021 , n365334 );
not ( n18554 , n17021 );
and ( n366332 , n18554 , n586 );
or ( n366333 , n18553 , n366332 );
buf ( n366334 , n366333 );
buf ( n366335 , n365375 );
nand ( n366336 , n366334 , n366335 );
buf ( n366337 , n366336 );
buf ( n366338 , n366337 );
nand ( n18562 , n366329 , n366338 );
buf ( n366340 , n18562 );
buf ( n366341 , n366340 );
xor ( n18565 , n365472 , n365555 );
xor ( n18566 , n18565 , n365589 );
buf ( n366344 , n18566 );
buf ( n366345 , n366344 );
xor ( n18569 , n366341 , n366345 );
xor ( n18570 , n365480 , n365508 );
xor ( n366348 , n18570 , n365550 );
buf ( n366349 , n366348 );
buf ( n366350 , n366349 );
buf ( n366351 , n365151 );
not ( n366352 , n366351 );
buf ( n366353 , n366017 );
not ( n18577 , n366353 );
or ( n18578 , n366352 , n18577 );
buf ( n366356 , n582 );
not ( n366357 , n366356 );
buf ( n366358 , n7349 );
not ( n18582 , n366358 );
or ( n366360 , n366357 , n18582 );
buf ( n366361 , n17547 );
buf ( n366362 , n364797 );
nand ( n18586 , n366361 , n366362 );
buf ( n366364 , n18586 );
buf ( n366365 , n366364 );
nand ( n18589 , n366360 , n366365 );
buf ( n366367 , n18589 );
buf ( n366368 , n366367 );
buf ( n366369 , n17133 );
nand ( n18593 , n366368 , n366369 );
buf ( n366371 , n18593 );
buf ( n366372 , n366371 );
nand ( n366373 , n18578 , n366372 );
buf ( n366374 , n366373 );
buf ( n366375 , n366374 );
xor ( n366376 , n366350 , n366375 );
buf ( n366377 , n364973 );
not ( n18601 , n366377 );
and ( n18602 , n357348 , n364771 );
not ( n366380 , n357348 );
and ( n366381 , n366380 , n584 );
or ( n18605 , n18602 , n366381 );
buf ( n366383 , n18605 );
not ( n366384 , n366383 );
or ( n366385 , n18601 , n366384 );
buf ( n366386 , n365991 );
buf ( n366387 , n364925 );
nand ( n366388 , n366386 , n366387 );
buf ( n366389 , n366388 );
buf ( n366390 , n366389 );
nand ( n18614 , n366385 , n366390 );
buf ( n366392 , n18614 );
buf ( n366393 , n366392 );
and ( n18617 , n366376 , n366393 );
and ( n18618 , n366350 , n366375 );
or ( n366396 , n18617 , n18618 );
buf ( n366397 , n366396 );
buf ( n366398 , n366397 );
and ( n18622 , n18569 , n366398 );
and ( n366400 , n366341 , n366345 );
or ( n366401 , n18622 , n366400 );
buf ( n366402 , n366401 );
buf ( n366403 , n366402 );
xor ( n366404 , n365972 , n365976 );
xor ( n366405 , n366404 , n366239 );
buf ( n366406 , n366405 );
buf ( n366407 , n366406 );
xor ( n366408 , n366403 , n366407 );
buf ( n366409 , n17867 );
not ( n18633 , n366409 );
buf ( n366411 , n366259 );
not ( n366412 , n366411 );
or ( n366413 , n18633 , n366412 );
and ( n18637 , n588 , n365362 );
not ( n18638 , n588 );
and ( n366416 , n18638 , n365355 );
or ( n366417 , n18637 , n366416 );
buf ( n366418 , n366417 );
buf ( n366419 , n365646 );
nand ( n366420 , n366418 , n366419 );
buf ( n366421 , n366420 );
buf ( n366422 , n366421 );
nand ( n18646 , n366413 , n366422 );
buf ( n366424 , n18646 );
buf ( n366425 , n366424 );
xor ( n18649 , n366002 , n366023 );
xor ( n18650 , n18649 , n366234 );
buf ( n366428 , n18650 );
buf ( n366429 , n366428 );
xor ( n18653 , n366425 , n366429 );
buf ( n366431 , n365351 );
not ( n366432 , n366431 );
buf ( n366433 , n366333 );
not ( n18657 , n366433 );
or ( n18658 , n366432 , n18657 );
buf ( n366436 , n586 );
not ( n18660 , n366436 );
buf ( n366438 , n365161 );
not ( n18662 , n366438 );
buf ( n366440 , n18662 );
buf ( n366441 , n366440 );
not ( n18665 , n366441 );
or ( n18666 , n18660 , n18665 );
buf ( n366444 , n360086 );
buf ( n366445 , n365334 );
nand ( n18669 , n366444 , n366445 );
buf ( n366447 , n18669 );
buf ( n366448 , n366447 );
nand ( n18672 , n18666 , n366448 );
buf ( n366450 , n18672 );
buf ( n366451 , n366450 );
buf ( n366452 , n365375 );
nand ( n18676 , n366451 , n366452 );
buf ( n366454 , n18676 );
buf ( n366455 , n366454 );
nand ( n18679 , n18658 , n366455 );
buf ( n366457 , n18679 );
buf ( n366458 , n366457 );
xor ( n18682 , n366095 , n366120 );
xor ( n18683 , n18682 , n366229 );
buf ( n366461 , n18683 );
buf ( n366462 , n366461 );
xor ( n18686 , n366458 , n366462 );
buf ( n366464 , n1121 );
not ( n18688 , n366464 );
buf ( n366466 , n18688 );
buf ( n366467 , n366466 );
not ( n18691 , n366467 );
buf ( n366469 , n18691 );
buf ( n366470 , n366469 );
buf ( n366471 , n576 );
and ( n18695 , n366470 , n366471 );
buf ( n366473 , n18695 );
buf ( n366474 , n366473 );
buf ( n366475 , n364834 );
not ( n18699 , n366475 );
buf ( n366477 , n366155 );
not ( n18701 , n366477 );
or ( n18702 , n18699 , n18701 );
buf ( n366480 , n576 );
not ( n18704 , n366480 );
buf ( n366482 , n366127 );
not ( n18706 , n366482 );
or ( n18707 , n18704 , n18706 );
buf ( n366485 , n366130 );
buf ( n366486 , n354303 );
nand ( n18710 , n366485 , n366486 );
buf ( n366488 , n18710 );
buf ( n366489 , n366488 );
nand ( n18713 , n18707 , n366489 );
buf ( n366491 , n18713 );
buf ( n366492 , n366491 );
buf ( n366493 , n17182 );
nand ( n18717 , n366492 , n366493 );
buf ( n366495 , n18717 );
buf ( n366496 , n366495 );
nand ( n18720 , n18702 , n366496 );
buf ( n366498 , n18720 );
buf ( n366499 , n366498 );
xor ( n18723 , n366474 , n366499 );
buf ( n366501 , n17037 );
not ( n18725 , n366501 );
buf ( n366503 , n366181 );
not ( n18727 , n366503 );
or ( n18728 , n18725 , n18727 );
buf ( n366506 , n578 );
not ( n18730 , n366506 );
buf ( n366508 , n366043 );
not ( n18732 , n366508 );
or ( n18733 , n18730 , n18732 );
buf ( n366511 , n364727 );
buf ( n366512 , n12481 );
nand ( n18736 , n366511 , n366512 );
buf ( n366514 , n18736 );
buf ( n366515 , n366514 );
nand ( n18739 , n18733 , n366515 );
buf ( n366517 , n18739 );
buf ( n366518 , n366517 );
buf ( n366519 , n17082 );
nand ( n18743 , n366518 , n366519 );
buf ( n366521 , n18743 );
buf ( n366522 , n366521 );
nand ( n18746 , n18728 , n366522 );
buf ( n366524 , n18746 );
buf ( n366525 , n366524 );
and ( n18749 , n18723 , n366525 );
and ( n18750 , n366474 , n366499 );
or ( n18751 , n18749 , n18750 );
buf ( n366529 , n18751 );
buf ( n366530 , n366529 );
xor ( n18754 , n366135 , n366163 );
xor ( n18755 , n18754 , n366189 );
buf ( n366533 , n18755 );
buf ( n366534 , n366533 );
xor ( n18758 , n366530 , n366534 );
buf ( n366536 , n17230 );
not ( n18760 , n366536 );
buf ( n366538 , n366211 );
not ( n18762 , n366538 );
or ( n18763 , n18760 , n18762 );
not ( n18764 , n580 );
not ( n18765 , n365063 );
or ( n18766 , n18764 , n18765 );
buf ( n366544 , n17372 );
buf ( n366545 , n364896 );
nand ( n18769 , n366544 , n366545 );
buf ( n366547 , n18769 );
nand ( n18771 , n18766 , n366547 );
nand ( n18772 , n18771 , n364885 );
buf ( n366550 , n18772 );
nand ( n18774 , n18763 , n366550 );
buf ( n366552 , n18774 );
buf ( n366553 , n366552 );
and ( n18777 , n18758 , n366553 );
and ( n18778 , n366530 , n366534 );
or ( n18779 , n18777 , n18778 );
buf ( n366557 , n18779 );
buf ( n366558 , n366557 );
buf ( n366559 , n364779 );
not ( n18783 , n366559 );
buf ( n366561 , n366367 );
not ( n18785 , n366561 );
or ( n18786 , n18783 , n18785 );
buf ( n366564 , n582 );
not ( n18788 , n366564 );
buf ( n366566 , n17725 );
not ( n18790 , n366566 );
or ( n18791 , n18788 , n18790 );
buf ( n366569 , n17174 );
buf ( n366570 , n364797 );
nand ( n18794 , n366569 , n366570 );
buf ( n366572 , n18794 );
buf ( n366573 , n366572 );
nand ( n18797 , n18791 , n366573 );
buf ( n366575 , n18797 );
buf ( n366576 , n366575 );
buf ( n366577 , n17133 );
nand ( n18801 , n366576 , n366577 );
buf ( n366579 , n18801 );
buf ( n366580 , n366579 );
nand ( n18804 , n18786 , n366580 );
buf ( n366582 , n18804 );
buf ( n366583 , n366582 );
xor ( n18807 , n366558 , n366583 );
xor ( n18808 , n366194 , n366219 );
xor ( n18809 , n18808 , n366224 );
buf ( n366587 , n18809 );
buf ( n366588 , n366587 );
and ( n18812 , n18807 , n366588 );
and ( n18813 , n366558 , n366583 );
or ( n18814 , n18812 , n18813 );
buf ( n366592 , n18814 );
buf ( n366593 , n366592 );
and ( n18817 , n18686 , n366593 );
and ( n18818 , n366458 , n366462 );
or ( n18819 , n18817 , n18818 );
buf ( n366597 , n18819 );
buf ( n366598 , n366597 );
and ( n18822 , n18653 , n366598 );
and ( n18823 , n366425 , n366429 );
or ( n18824 , n18822 , n18823 );
buf ( n366602 , n18824 );
buf ( n366603 , n366602 );
and ( n18827 , n366408 , n366603 );
and ( n18828 , n366403 , n366407 );
or ( n18829 , n18827 , n18828 );
buf ( n366607 , n18829 );
buf ( n366608 , n366607 );
xor ( n18832 , n366324 , n366608 );
xor ( n18833 , n366244 , n366248 );
xor ( n18834 , n18833 , n366294 );
buf ( n366612 , n18834 );
buf ( n366613 , n366612 );
and ( n18837 , n18832 , n366613 );
and ( n18838 , n366324 , n366608 );
or ( n18839 , n18837 , n18838 );
buf ( n366617 , n18839 );
nor ( n18841 , n366320 , n366617 );
xor ( n18842 , n366324 , n366608 );
xor ( n18843 , n18842 , n366613 );
buf ( n366621 , n18843 );
buf ( n366622 , n366621 );
xor ( n18846 , n366267 , n366271 );
xor ( n18847 , n18846 , n366289 );
buf ( n366625 , n18847 );
buf ( n366626 , n366625 );
buf ( n366627 , n365738 );
not ( n18851 , n366627 );
and ( n18852 , n590 , n365748 );
not ( n18853 , n590 );
not ( n18854 , n365748 );
and ( n18855 , n18853 , n18854 );
or ( n18856 , n18852 , n18855 );
buf ( n366634 , n18856 );
not ( n18858 , n366634 );
or ( n18859 , n18851 , n18858 );
buf ( n366637 , n366278 );
buf ( n366638 , n591 );
nand ( n18862 , n366637 , n366638 );
buf ( n366640 , n18862 );
buf ( n366641 , n366640 );
nand ( n18865 , n18859 , n366641 );
buf ( n366643 , n18865 );
buf ( n366644 , n366643 );
xor ( n18868 , n366341 , n366345 );
xor ( n18869 , n18868 , n366398 );
buf ( n366647 , n18869 );
buf ( n366648 , n366647 );
xor ( n18872 , n366644 , n366648 );
buf ( n366650 , n365646 );
not ( n18874 , n366650 );
buf ( n366652 , n14498 );
buf ( n18876 , n366652 );
buf ( n366654 , n18876 );
buf ( n366655 , n366654 );
not ( n18879 , n366655 );
buf ( n366657 , n18879 );
and ( n18881 , n588 , n366657 );
not ( n18882 , n588 );
and ( n18883 , n18882 , n366654 );
or ( n18884 , n18881 , n18883 );
buf ( n366662 , n18884 );
not ( n18886 , n366662 );
or ( n18887 , n18874 , n18886 );
buf ( n366665 , n366417 );
buf ( n366666 , n17867 );
nand ( n18890 , n366665 , n366666 );
buf ( n366668 , n18890 );
buf ( n366669 , n366668 );
nand ( n18893 , n18887 , n366669 );
buf ( n366671 , n18893 );
buf ( n366672 , n366671 );
xor ( n18896 , n366350 , n366375 );
xor ( n18897 , n18896 , n366393 );
buf ( n366675 , n18897 );
buf ( n366676 , n366675 );
xor ( n18900 , n366672 , n366676 );
buf ( n366678 , n364925 );
not ( n18902 , n366678 );
buf ( n366680 , n18605 );
not ( n18904 , n366680 );
or ( n18905 , n18902 , n18904 );
and ( n18906 , n584 , n8304 );
not ( n18907 , n584 );
and ( n18908 , n18907 , n8303 );
or ( n18909 , n18906 , n18908 );
buf ( n366687 , n18909 );
buf ( n366688 , n364973 );
nand ( n18912 , n366687 , n366688 );
buf ( n366690 , n18912 );
buf ( n366691 , n366690 );
nand ( n18915 , n18905 , n366691 );
buf ( n366693 , n18915 );
buf ( n366694 , n366693 );
buf ( n366695 , n365351 );
not ( n18919 , n366695 );
buf ( n366697 , n366450 );
not ( n18921 , n366697 );
or ( n18922 , n18919 , n18921 );
buf ( n366700 , n586 );
not ( n18924 , n366700 );
buf ( n366702 , n365176 );
not ( n18926 , n366702 );
or ( n18927 , n18924 , n18926 );
buf ( n366705 , n357316 );
buf ( n366706 , n365334 );
nand ( n18930 , n366705 , n366706 );
buf ( n366708 , n18930 );
buf ( n366709 , n366708 );
nand ( n18933 , n18927 , n366709 );
buf ( n366711 , n18933 );
buf ( n366712 , n366711 );
buf ( n366713 , n365375 );
nand ( n18937 , n366712 , n366713 );
buf ( n366715 , n18937 );
buf ( n366716 , n366715 );
nand ( n18940 , n18922 , n366716 );
buf ( n366718 , n18940 );
buf ( n366719 , n366718 );
xor ( n18943 , n366694 , n366719 );
buf ( n366721 , n364779 );
not ( n18945 , n366721 );
buf ( n366723 , n366575 );
not ( n18947 , n366723 );
or ( n18948 , n18945 , n18947 );
buf ( n366726 , n582 );
not ( n18950 , n366726 );
buf ( n366728 , n364823 );
not ( n18952 , n366728 );
or ( n18953 , n18950 , n18952 );
buf ( n366731 , n365099 );
buf ( n366732 , n364797 );
nand ( n18956 , n366731 , n366732 );
buf ( n366734 , n18956 );
buf ( n366735 , n366734 );
nand ( n18959 , n18953 , n366735 );
buf ( n366737 , n18959 );
buf ( n366738 , n366737 );
buf ( n366739 , n17133 );
nand ( n18963 , n366738 , n366739 );
buf ( n366741 , n18963 );
buf ( n366742 , n366741 );
nand ( n18966 , n18948 , n366742 );
buf ( n366744 , n18966 );
buf ( n366745 , n366744 );
not ( n18969 , n17197 );
not ( n18970 , n18771 );
or ( n18971 , n18969 , n18970 );
and ( n18972 , n365032 , n580 );
not ( n18973 , n365032 );
and ( n18974 , n18973 , n364896 );
or ( n18975 , n18972 , n18974 );
nand ( n18976 , n18975 , n364885 );
nand ( n18977 , n18971 , n18976 );
buf ( n366755 , n18977 );
buf ( n366756 , n576 );
buf ( n366757 , n12484 );
and ( n18981 , n366756 , n366757 );
buf ( n366759 , n18981 );
buf ( n366760 , n366759 );
buf ( n366761 , n364834 );
not ( n18985 , n366761 );
buf ( n366763 , n366491 );
not ( n18987 , n366763 );
or ( n18988 , n18985 , n18987 );
buf ( n366766 , n576 );
not ( n18990 , n366766 );
buf ( n366768 , n366466 );
not ( n18992 , n366768 );
or ( n18993 , n18990 , n18992 );
buf ( n366771 , n366469 );
buf ( n366772 , n354303 );
nand ( n18996 , n366771 , n366772 );
buf ( n366774 , n18996 );
buf ( n366775 , n366774 );
nand ( n18999 , n18993 , n366775 );
buf ( n366777 , n18999 );
buf ( n366778 , n366777 );
buf ( n366779 , n17182 );
nand ( n19003 , n366778 , n366779 );
buf ( n366781 , n19003 );
buf ( n366782 , n366781 );
nand ( n19006 , n18988 , n366782 );
buf ( n366784 , n19006 );
buf ( n366785 , n366784 );
xor ( n19009 , n366760 , n366785 );
buf ( n366787 , n17037 );
not ( n19011 , n366787 );
buf ( n366789 , n366517 );
not ( n19013 , n366789 );
or ( n19014 , n19011 , n19013 );
buf ( n366792 , n578 );
not ( n19016 , n366792 );
buf ( n366794 , n366145 );
not ( n19018 , n366794 );
or ( n19019 , n19016 , n19018 );
buf ( n366797 , n366028 );
buf ( n366798 , n364727 );
nand ( n19022 , n366797 , n366798 );
buf ( n366800 , n19022 );
buf ( n366801 , n366800 );
nand ( n19025 , n19019 , n366801 );
buf ( n366803 , n19025 );
buf ( n366804 , n366803 );
buf ( n366805 , n17082 );
nand ( n19029 , n366804 , n366805 );
buf ( n366807 , n19029 );
buf ( n366808 , n366807 );
nand ( n19032 , n19014 , n366808 );
buf ( n366810 , n19032 );
buf ( n366811 , n366810 );
and ( n19035 , n19009 , n366811 );
and ( n19036 , n366760 , n366785 );
or ( n19037 , n19035 , n19036 );
buf ( n366815 , n19037 );
buf ( n366816 , n366815 );
xor ( n19040 , n366755 , n366816 );
xor ( n19041 , n366474 , n366499 );
xor ( n19042 , n19041 , n366525 );
buf ( n366820 , n19042 );
buf ( n366821 , n366820 );
and ( n19045 , n19040 , n366821 );
and ( n19046 , n366755 , n366816 );
or ( n19047 , n19045 , n19046 );
buf ( n366825 , n19047 );
buf ( n366826 , n366825 );
xor ( n19050 , n366745 , n366826 );
xor ( n19051 , n366530 , n366534 );
xor ( n19052 , n19051 , n366553 );
buf ( n366830 , n19052 );
buf ( n366831 , n366830 );
and ( n19055 , n19050 , n366831 );
and ( n19056 , n366745 , n366826 );
or ( n19057 , n19055 , n19056 );
buf ( n366835 , n19057 );
buf ( n366836 , n366835 );
and ( n19060 , n18943 , n366836 );
and ( n19061 , n366694 , n366719 );
or ( n19062 , n19060 , n19061 );
buf ( n366840 , n19062 );
buf ( n366841 , n366840 );
and ( n19065 , n18900 , n366841 );
and ( n19066 , n366672 , n366676 );
or ( n19067 , n19065 , n19066 );
buf ( n366845 , n19067 );
buf ( n366846 , n366845 );
and ( n19070 , n18872 , n366846 );
and ( n19071 , n366644 , n366648 );
or ( n19072 , n19070 , n19071 );
buf ( n366850 , n19072 );
buf ( n366851 , n366850 );
xor ( n19075 , n366626 , n366851 );
xor ( n19076 , n366403 , n366407 );
xor ( n19077 , n19076 , n366603 );
buf ( n366855 , n19077 );
buf ( n366856 , n366855 );
and ( n19080 , n19075 , n366856 );
and ( n19081 , n366626 , n366851 );
or ( n19082 , n19080 , n19081 );
buf ( n366860 , n19082 );
buf ( n366861 , n366860 );
nor ( n19085 , n366622 , n366861 );
buf ( n366863 , n19085 );
nor ( n19087 , n18841 , n366863 );
buf ( n366865 , n19087 );
not ( n19089 , n366865 );
xor ( n19090 , n366626 , n366851 );
xor ( n19091 , n19090 , n366856 );
buf ( n366869 , n19091 );
xor ( n19093 , n366425 , n366429 );
xor ( n19094 , n19093 , n366598 );
buf ( n366872 , n19094 );
buf ( n366873 , n366872 );
xor ( n19097 , n366458 , n366462 );
xor ( n19098 , n19097 , n366593 );
buf ( n366876 , n19098 );
buf ( n366877 , n366876 );
buf ( n366878 , n591 );
not ( n19102 , n366878 );
buf ( n366880 , n18856 );
not ( n19104 , n366880 );
or ( n19105 , n19102 , n19104 );
not ( n19106 , n17520 );
and ( n19107 , n590 , n19106 );
not ( n19108 , n590 );
and ( n19109 , n19108 , n17520 );
nor ( n19110 , n19107 , n19109 );
buf ( n366888 , n19110 );
buf ( n366889 , n365738 );
nand ( n19113 , n366888 , n366889 );
buf ( n366891 , n19113 );
buf ( n366892 , n366891 );
nand ( n19116 , n19105 , n366892 );
buf ( n366894 , n19116 );
buf ( n366895 , n366894 );
xor ( n19119 , n366877 , n366895 );
xor ( n19120 , n366558 , n366583 );
xor ( n19121 , n19120 , n366588 );
buf ( n366899 , n19121 );
buf ( n366900 , n366899 );
buf ( n366901 , n17867 );
not ( n19125 , n366901 );
buf ( n366903 , n18884 );
not ( n19127 , n366903 );
or ( n19128 , n19125 , n19127 );
xor ( n19129 , n588 , n365403 );
buf ( n366907 , n19129 );
buf ( n366908 , n365646 );
nand ( n19132 , n366907 , n366908 );
buf ( n366910 , n19132 );
buf ( n366911 , n366910 );
nand ( n19135 , n19128 , n366911 );
buf ( n366913 , n19135 );
buf ( n366914 , n366913 );
xor ( n19138 , n366900 , n366914 );
buf ( n366916 , n364925 );
not ( n19140 , n366916 );
buf ( n366918 , n18909 );
not ( n19142 , n366918 );
or ( n19143 , n19140 , n19142 );
buf ( n366921 , n584 );
not ( n19145 , n366921 );
not ( n19146 , n17161 );
buf ( n366924 , n19146 );
not ( n19148 , n366924 );
or ( n19149 , n19145 , n19148 );
buf ( n366927 , n17547 );
buf ( n366928 , n364771 );
nand ( n19152 , n366927 , n366928 );
buf ( n366930 , n19152 );
buf ( n366931 , n366930 );
nand ( n19155 , n19149 , n366931 );
buf ( n366933 , n19155 );
buf ( n366934 , n366933 );
buf ( n366935 , n364973 );
nand ( n19159 , n366934 , n366935 );
buf ( n366937 , n19159 );
buf ( n366938 , n366937 );
nand ( n19162 , n19143 , n366938 );
buf ( n366940 , n19162 );
buf ( n366941 , n366940 );
buf ( n366942 , n576 );
buf ( n19166 , n1093 );
buf ( n366944 , n19166 );
not ( n19168 , n366944 );
buf ( n366946 , n19168 );
buf ( n366947 , n366946 );
not ( n19171 , n366947 );
buf ( n366949 , n19171 );
buf ( n366950 , n366949 );
and ( n19174 , n366942 , n366950 );
buf ( n366952 , n19174 );
buf ( n366953 , n366952 );
buf ( n366954 , n364834 );
not ( n19178 , n366954 );
buf ( n366956 , n366777 );
not ( n19180 , n366956 );
or ( n19181 , n19178 , n19180 );
xor ( n19182 , n366756 , n366757 );
buf ( n366960 , n19182 );
buf ( n366961 , n366960 );
buf ( n366962 , n17182 );
nand ( n19186 , n366961 , n366962 );
buf ( n366964 , n19186 );
buf ( n366965 , n366964 );
nand ( n19189 , n19181 , n366965 );
buf ( n366967 , n19189 );
buf ( n366968 , n366967 );
xor ( n19192 , n366953 , n366968 );
buf ( n366970 , n17037 );
not ( n19194 , n366970 );
buf ( n366972 , n366803 );
not ( n19196 , n366972 );
or ( n19197 , n19194 , n19196 );
buf ( n366975 , n12482 );
not ( n19199 , n366975 );
buf ( n366977 , n19199 );
nand ( n19201 , n366977 , n578 );
not ( n19202 , n19201 );
buf ( n366980 , n12482 );
buf ( n19204 , n366980 );
buf ( n366982 , n19204 );
buf ( n366983 , n366982 );
buf ( n366984 , n364727 );
nand ( n19208 , n366983 , n366984 );
buf ( n366986 , n19208 );
not ( n19210 , n366986 );
or ( n19211 , n19202 , n19210 );
nand ( n19212 , n19211 , n17082 );
buf ( n366990 , n19212 );
nand ( n19214 , n19197 , n366990 );
buf ( n366992 , n19214 );
buf ( n366993 , n366992 );
and ( n19217 , n19192 , n366993 );
and ( n19218 , n366953 , n366968 );
or ( n19219 , n19217 , n19218 );
buf ( n366997 , n19219 );
buf ( n366998 , n366997 );
buf ( n366999 , n17230 );
not ( n19223 , n366999 );
buf ( n367001 , n18975 );
not ( n19225 , n367001 );
or ( n19226 , n19223 , n19225 );
buf ( n367004 , n580 );
not ( n19228 , n367004 );
buf ( n367006 , n365494 );
not ( n19230 , n367006 );
or ( n19231 , n19228 , n19230 );
buf ( n367009 , n365497 );
buf ( n367010 , n364896 );
nand ( n19234 , n367009 , n367010 );
buf ( n367012 , n19234 );
buf ( n367013 , n367012 );
nand ( n19237 , n19231 , n367013 );
buf ( n367015 , n19237 );
buf ( n367016 , n367015 );
buf ( n367017 , n364885 );
nand ( n19241 , n367016 , n367017 );
buf ( n367019 , n19241 );
buf ( n367020 , n367019 );
nand ( n19244 , n19226 , n367020 );
buf ( n367022 , n19244 );
buf ( n367023 , n367022 );
xor ( n19247 , n366998 , n367023 );
xor ( n19248 , n366760 , n366785 );
xor ( n19249 , n19248 , n366811 );
buf ( n367027 , n19249 );
buf ( n367028 , n367027 );
and ( n19252 , n19247 , n367028 );
and ( n19253 , n366998 , n367023 );
or ( n19254 , n19252 , n19253 );
buf ( n367032 , n19254 );
buf ( n367033 , n367032 );
buf ( n367034 , n364779 );
not ( n19258 , n367034 );
buf ( n367036 , n366737 );
not ( n19260 , n367036 );
or ( n19261 , n19258 , n19260 );
buf ( n367039 , n582 );
not ( n19263 , n367039 );
buf ( n367041 , n365516 );
not ( n19265 , n367041 );
or ( n19266 , n19263 , n19265 );
buf ( n367044 , n17301 );
buf ( n367045 , n364797 );
nand ( n19269 , n367044 , n367045 );
buf ( n367047 , n19269 );
buf ( n367048 , n367047 );
nand ( n19272 , n19266 , n367048 );
buf ( n367050 , n19272 );
buf ( n367051 , n367050 );
buf ( n367052 , n17133 );
nand ( n19276 , n367051 , n367052 );
buf ( n367054 , n19276 );
buf ( n367055 , n367054 );
nand ( n19279 , n19261 , n367055 );
buf ( n367057 , n19279 );
buf ( n367058 , n367057 );
xor ( n19282 , n367033 , n367058 );
xor ( n19283 , n366755 , n366816 );
xor ( n19284 , n19283 , n366821 );
buf ( n367062 , n19284 );
buf ( n367063 , n367062 );
and ( n19287 , n19282 , n367063 );
and ( n19288 , n367033 , n367058 );
or ( n19289 , n19287 , n19288 );
buf ( n367067 , n19289 );
buf ( n367068 , n367067 );
xor ( n19292 , n366941 , n367068 );
buf ( n367070 , n365351 );
not ( n19294 , n367070 );
buf ( n367072 , n366711 );
not ( n19296 , n367072 );
or ( n19297 , n19294 , n19296 );
and ( n19298 , n364720 , n586 );
not ( n19299 , n364720 );
and ( n19300 , n19299 , n348260 );
or ( n19301 , n19298 , n19300 );
nand ( n19302 , n19301 , n365375 );
buf ( n367080 , n19302 );
nand ( n19304 , n19297 , n367080 );
buf ( n367082 , n19304 );
buf ( n367083 , n367082 );
and ( n19307 , n19292 , n367083 );
and ( n19308 , n366941 , n367068 );
or ( n19309 , n19307 , n19308 );
buf ( n367087 , n19309 );
buf ( n367088 , n367087 );
and ( n19312 , n19138 , n367088 );
and ( n19313 , n366900 , n366914 );
or ( n19314 , n19312 , n19313 );
buf ( n367092 , n19314 );
buf ( n367093 , n367092 );
and ( n19317 , n19119 , n367093 );
and ( n19318 , n366877 , n366895 );
or ( n19319 , n19317 , n19318 );
buf ( n367097 , n19319 );
buf ( n367098 , n367097 );
xor ( n19322 , n366873 , n367098 );
xor ( n19323 , n366644 , n366648 );
xor ( n19324 , n19323 , n366846 );
buf ( n367102 , n19324 );
buf ( n367103 , n367102 );
and ( n19327 , n19322 , n367103 );
and ( n19328 , n366873 , n367098 );
or ( n19329 , n19327 , n19328 );
buf ( n367107 , n19329 );
nor ( n19331 , n366869 , n367107 );
buf ( n367109 , n591 );
not ( n19333 , n367109 );
buf ( n367111 , n19110 );
not ( n19335 , n367111 );
or ( n19336 , n19333 , n19335 );
buf ( n367114 , n365738 );
not ( n19338 , n367114 );
buf ( n367116 , n19338 );
buf ( n367117 , n367116 );
not ( n19341 , n367117 );
and ( n19342 , n590 , n364936 );
not ( n19343 , n590 );
buf ( n367121 , n365362 );
not ( n19345 , n367121 );
buf ( n367123 , n19345 );
and ( n19347 , n19343 , n367123 );
or ( n19348 , n19342 , n19347 );
buf ( n367126 , n19348 );
nand ( n19350 , n19341 , n367126 );
buf ( n367128 , n19350 );
buf ( n367129 , n367128 );
nand ( n19353 , n19336 , n367129 );
buf ( n367131 , n19353 );
buf ( n367132 , n367131 );
xor ( n19356 , n366694 , n366719 );
xor ( n19357 , n19356 , n366836 );
buf ( n367135 , n19357 );
buf ( n367136 , n367135 );
xor ( n19360 , n367132 , n367136 );
xor ( n19361 , n366745 , n366826 );
xor ( n19362 , n19361 , n366831 );
buf ( n367140 , n19362 );
buf ( n367141 , n367140 );
buf ( n367142 , n17867 );
not ( n19366 , n367142 );
buf ( n367144 , n19129 );
not ( n19368 , n367144 );
or ( n19369 , n19366 , n19368 );
and ( n19370 , n588 , n366440 );
not ( n19371 , n588 );
and ( n19372 , n19371 , n360086 );
or ( n19373 , n19370 , n19372 );
buf ( n367151 , n19373 );
buf ( n367152 , n365646 );
nand ( n19376 , n367151 , n367152 );
buf ( n367154 , n19376 );
buf ( n367155 , n367154 );
nand ( n19379 , n19369 , n367155 );
buf ( n367157 , n19379 );
buf ( n367158 , n367157 );
xor ( n19382 , n367141 , n367158 );
buf ( n367160 , n365738 );
not ( n19384 , n367160 );
and ( n19385 , n590 , n366657 );
not ( n19386 , n590 );
and ( n19387 , n19386 , n366654 );
or ( n19388 , n19385 , n19387 );
buf ( n367166 , n19388 );
not ( n19390 , n367166 );
or ( n19391 , n19384 , n19390 );
buf ( n367169 , n19348 );
buf ( n367170 , n591 );
nand ( n19394 , n367169 , n367170 );
buf ( n367172 , n19394 );
buf ( n367173 , n367172 );
nand ( n19397 , n19391 , n367173 );
buf ( n367175 , n19397 );
buf ( n367176 , n367175 );
and ( n19400 , n19382 , n367176 );
and ( n19401 , n367141 , n367158 );
or ( n19402 , n19400 , n19401 );
buf ( n367180 , n19402 );
buf ( n367181 , n367180 );
and ( n19405 , n19360 , n367181 );
and ( n19406 , n367132 , n367136 );
or ( n19407 , n19405 , n19406 );
buf ( n367185 , n19407 );
buf ( n367186 , n367185 );
xor ( n19410 , n366672 , n366676 );
xor ( n19411 , n19410 , n366841 );
buf ( n367189 , n19411 );
buf ( n367190 , n367189 );
xor ( n19414 , n367186 , n367190 );
xor ( n19415 , n366877 , n366895 );
xor ( n19416 , n19415 , n367093 );
buf ( n367194 , n19416 );
buf ( n367195 , n367194 );
xor ( n19419 , n19414 , n367195 );
buf ( n367197 , n19419 );
xor ( n19421 , n366900 , n366914 );
xor ( n19422 , n19421 , n367088 );
buf ( n367200 , n19422 );
buf ( n367201 , n367200 );
xor ( n19425 , n367132 , n367136 );
xor ( n19426 , n19425 , n367181 );
buf ( n367204 , n19426 );
buf ( n367205 , n367204 );
xor ( n19429 , n367201 , n367205 );
buf ( n367207 , n364925 );
not ( n19431 , n367207 );
buf ( n367209 , n366933 );
not ( n19433 , n367209 );
or ( n19434 , n19431 , n19433 );
buf ( n367212 , n584 );
not ( n19436 , n367212 );
buf ( n367214 , n17725 );
not ( n19438 , n367214 );
or ( n19439 , n19436 , n19438 );
buf ( n367217 , n17174 );
buf ( n367218 , n364771 );
nand ( n19442 , n367217 , n367218 );
buf ( n367220 , n19442 );
buf ( n367221 , n367220 );
nand ( n19445 , n19439 , n367221 );
buf ( n367223 , n19445 );
buf ( n367224 , n367223 );
buf ( n367225 , n364973 );
nand ( n19449 , n367224 , n367225 );
buf ( n367227 , n19449 );
buf ( n367228 , n367227 );
nand ( n19452 , n19434 , n367228 );
buf ( n367230 , n19452 );
buf ( n367231 , n367230 );
buf ( n367232 , C0 );
buf ( n367233 , n367232 );
buf ( n367234 , n364834 );
not ( n19461 , n367234 );
buf ( n367236 , n366960 );
not ( n19463 , n367236 );
or ( n19464 , n19461 , n19463 );
xor ( n19465 , n366942 , n366950 );
buf ( n367240 , n19465 );
buf ( n367241 , n367240 );
buf ( n367242 , n17182 );
nand ( n19469 , n367241 , n367242 );
buf ( n367244 , n19469 );
buf ( n367245 , n367244 );
nand ( n19472 , n19464 , n367245 );
buf ( n367247 , n19472 );
buf ( n367248 , n367247 );
xor ( n19475 , n367233 , n367248 );
buf ( n367250 , C0 );
buf ( n367251 , n367250 );
buf ( n367252 , C0 );
buf ( n367253 , n367252 );
buf ( n367254 , n576 );
not ( n19487 , n367254 );
buf ( n367256 , C1 );
or ( n19493 , n19487 , C0 );
buf ( n367258 , C1 );
buf ( n367259 , n367258 );
nand ( n19499 , n19493 , n367259 );
buf ( n367261 , n19499 );
not ( n19501 , n367261 );
not ( n19502 , n364834 );
or ( n19503 , n19501 , n19502 );
buf ( n367265 , n576 );
not ( n19505 , n367265 );
buf ( n367267 , C1 );
or ( n19511 , n19505 , C0 );
buf ( n367269 , C1 );
buf ( n367270 , n367269 );
nand ( n19520 , n19511 , n367270 );
buf ( n367272 , n19520 );
buf ( n367273 , n367272 );
buf ( n367274 , n17182 );
nand ( n19524 , n367273 , n367274 );
buf ( n367276 , n19524 );
nand ( n19526 , n19503 , n367276 );
buf ( n367278 , n19526 );
xor ( n19528 , n367253 , n367278 );
buf ( n367280 , C1 );
buf ( n367281 , n367280 );
buf ( n367282 , n577 );
buf ( n367283 , n578 );
and ( n19533 , n367282 , n367283 );
buf ( n367285 , n354303 );
nor ( n19535 , n19533 , n367285 );
buf ( n367287 , n19535 );
buf ( n367288 , n367287 );
and ( n19538 , n367281 , n367288 );
buf ( n367290 , n19538 );
buf ( n367291 , n367290 );
not ( n19541 , n367272 );
not ( n19542 , n364834 );
or ( n19543 , n19541 , n19542 );
buf ( n367295 , n576 );
buf ( n367296 , C0 );
xor ( n19546 , n367295 , n367296 );
buf ( n367298 , n19546 );
buf ( n367299 , n367298 );
buf ( n367300 , n17182 );
nand ( n19550 , n367299 , n367300 );
buf ( n367302 , n19550 );
nand ( n19552 , n19543 , n367302 );
buf ( n367304 , n19552 );
and ( n19554 , n367291 , n367304 );
buf ( n367306 , n19554 );
buf ( n367307 , n367306 );
and ( n19557 , n19528 , n367307 );
or ( n19558 , n19557 , C0 );
buf ( n367310 , n19558 );
buf ( n367311 , n367310 );
xor ( n19561 , n367251 , n367311 );
buf ( n367313 , n364834 );
not ( n19563 , n367313 );
buf ( n367315 , n367240 );
not ( n19565 , n367315 );
or ( n19566 , n19563 , n19565 );
buf ( n367318 , n367261 );
buf ( n367319 , n17182 );
nand ( n19569 , n367318 , n367319 );
buf ( n367321 , n19569 );
buf ( n367322 , n367321 );
nand ( n19572 , n19566 , n367322 );
buf ( n367324 , n19572 );
buf ( n367325 , n367324 );
and ( n19575 , n19561 , n367325 );
or ( n19577 , n19575 , C0 );
buf ( n367328 , n19577 );
buf ( n367329 , n367328 );
and ( n19580 , n19475 , n367329 );
or ( n19582 , n19580 , C0 );
buf ( n367332 , n19582 );
buf ( n367333 , n367332 );
xor ( n19585 , n366953 , n366968 );
xor ( n19586 , n19585 , n366993 );
buf ( n367336 , n19586 );
buf ( n367337 , n367336 );
xor ( n19589 , n367333 , n367337 );
buf ( n367339 , n17230 );
not ( n19591 , n367339 );
buf ( n367341 , n367015 );
not ( n19593 , n367341 );
or ( n19594 , n19591 , n19593 );
not ( n19595 , n580 );
not ( n19596 , n365475 );
or ( n19597 , n19595 , n19596 );
buf ( n367347 , n366049 );
buf ( n367348 , n364896 );
nand ( n19600 , n367347 , n367348 );
buf ( n367350 , n19600 );
nand ( n19602 , n19597 , n367350 );
nand ( n19603 , n19602 , n364885 );
buf ( n367353 , n19603 );
nand ( n19605 , n19594 , n367353 );
buf ( n367355 , n19605 );
buf ( n367356 , n367355 );
and ( n19608 , n19589 , n367356 );
and ( n19609 , n367333 , n367337 );
or ( n19610 , n19608 , n19609 );
buf ( n367360 , n19610 );
buf ( n367361 , n367360 );
buf ( n367362 , n364779 );
not ( n19614 , n367362 );
buf ( n367364 , n367050 );
not ( n19616 , n367364 );
or ( n19617 , n19614 , n19616 );
buf ( n367367 , n582 );
not ( n19619 , n367367 );
buf ( n367369 , n365063 );
not ( n19621 , n367369 );
or ( n19622 , n19619 , n19621 );
buf ( n367372 , n17372 );
buf ( n367373 , n364797 );
nand ( n19625 , n367372 , n367373 );
buf ( n367375 , n19625 );
buf ( n367376 , n367375 );
nand ( n19628 , n19622 , n367376 );
buf ( n367378 , n19628 );
buf ( n367379 , n367378 );
buf ( n367380 , n17133 );
nand ( n19632 , n367379 , n367380 );
buf ( n367382 , n19632 );
buf ( n367383 , n367382 );
nand ( n19635 , n19617 , n367383 );
buf ( n367385 , n19635 );
buf ( n367386 , n367385 );
xor ( n19638 , n367361 , n367386 );
xor ( n19639 , n366998 , n367023 );
xor ( n19640 , n19639 , n367028 );
buf ( n367390 , n19640 );
buf ( n367391 , n367390 );
and ( n19643 , n19638 , n367391 );
and ( n19644 , n367361 , n367386 );
or ( n19645 , n19643 , n19644 );
buf ( n367395 , n19645 );
buf ( n367396 , n367395 );
xor ( n19648 , n367231 , n367396 );
xor ( n19649 , n367033 , n367058 );
xor ( n19650 , n19649 , n367063 );
buf ( n367400 , n19650 );
buf ( n367401 , n367400 );
and ( n19653 , n19648 , n367401 );
and ( n19654 , n367231 , n367396 );
or ( n19655 , n19653 , n19654 );
buf ( n367405 , n19655 );
buf ( n367406 , n367405 );
xor ( n19658 , n366941 , n367068 );
xor ( n19659 , n19658 , n367083 );
buf ( n367409 , n19659 );
buf ( n367410 , n367409 );
xor ( n19662 , n367406 , n367410 );
buf ( n367412 , n365351 );
not ( n19664 , n367412 );
buf ( n367414 , n19301 );
not ( n19666 , n367414 );
or ( n19667 , n19664 , n19666 );
buf ( n367417 , n586 );
not ( n19669 , n367417 );
buf ( n367419 , n8304 );
not ( n19671 , n367419 );
or ( n19672 , n19669 , n19671 );
buf ( n367422 , n8303 );
buf ( n367423 , n365334 );
nand ( n19675 , n367422 , n367423 );
buf ( n367425 , n19675 );
buf ( n367426 , n367425 );
nand ( n19678 , n19672 , n367426 );
buf ( n367428 , n19678 );
buf ( n367429 , n367428 );
buf ( n367430 , n365375 );
nand ( n19682 , n367429 , n367430 );
buf ( n367432 , n19682 );
buf ( n367433 , n367432 );
nand ( n19685 , n19667 , n367433 );
buf ( n367435 , n19685 );
buf ( n367436 , n367435 );
buf ( n367437 , n365646 );
not ( n19689 , n367437 );
xnor ( n19690 , n588 , n365176 );
buf ( n367440 , n19690 );
not ( n19692 , n367440 );
or ( n19693 , n19689 , n19692 );
buf ( n367443 , n19373 );
buf ( n367444 , n17867 );
nand ( n19696 , n367443 , n367444 );
buf ( n367446 , n19696 );
buf ( n367447 , n367446 );
nand ( n19699 , n19693 , n367447 );
buf ( n367449 , n19699 );
buf ( n367450 , n367449 );
xor ( n19702 , n367436 , n367450 );
buf ( n367452 , n364925 );
not ( n19704 , n367452 );
buf ( n367454 , n367223 );
not ( n19706 , n367454 );
or ( n19707 , n19704 , n19706 );
buf ( n367457 , n584 );
not ( n19709 , n367457 );
buf ( n367459 , n364823 );
not ( n19711 , n367459 );
or ( n19712 , n19709 , n19711 );
buf ( n367462 , n365093 );
not ( n19714 , n367462 );
buf ( n367464 , n364771 );
nand ( n19716 , n19714 , n367464 );
buf ( n367466 , n19716 );
buf ( n367467 , n367466 );
nand ( n19719 , n19712 , n367467 );
buf ( n367469 , n19719 );
buf ( n367470 , n367469 );
buf ( n367471 , n364973 );
nand ( n19723 , n367470 , n367471 );
buf ( n367473 , n19723 );
buf ( n367474 , n367473 );
nand ( n19726 , n19707 , n367474 );
buf ( n367476 , n19726 );
buf ( n367477 , n367476 );
buf ( n367478 , n17037 );
not ( n19730 , n367478 );
nand ( n19731 , n366986 , n19201 );
buf ( n367481 , n19731 );
not ( n19733 , n367481 );
or ( n19734 , n19730 , n19733 );
buf ( n367484 , n578 );
not ( n19736 , n367484 );
buf ( n367486 , n366466 );
not ( n19738 , n367486 );
or ( n19739 , n19736 , n19738 );
buf ( n367489 , n364727 );
buf ( n367490 , n1121 );
buf ( n19742 , n367490 );
buf ( n367492 , n19742 );
buf ( n367493 , n367492 );
nand ( n19745 , n367489 , n367493 );
buf ( n367495 , n19745 );
buf ( n367496 , n367495 );
nand ( n19748 , n19739 , n367496 );
buf ( n367498 , n19748 );
buf ( n367499 , n367498 );
buf ( n367500 , n17082 );
nand ( n19752 , n367499 , n367500 );
buf ( n367502 , n19752 );
buf ( n367503 , n367502 );
nand ( n19755 , n19734 , n367503 );
buf ( n367505 , n19755 );
buf ( n367506 , n367505 );
xor ( n19758 , n367233 , n367248 );
xor ( n19759 , n19758 , n367329 );
buf ( n367509 , n19759 );
buf ( n367510 , n367509 );
xor ( n19762 , n367506 , n367510 );
not ( n19763 , n17230 );
not ( n19764 , n19602 );
or ( n19765 , n19763 , n19764 );
buf ( n367515 , n580 );
not ( n19767 , n367515 );
buf ( n367517 , n366145 );
not ( n19769 , n367517 );
or ( n19770 , n19767 , n19769 );
buf ( n367520 , n366028 );
buf ( n367521 , n364896 );
nand ( n19773 , n367520 , n367521 );
buf ( n367523 , n19773 );
buf ( n367524 , n367523 );
nand ( n19776 , n19770 , n367524 );
buf ( n367526 , n19776 );
buf ( n367527 , n367526 );
buf ( n367528 , n364885 );
nand ( n19780 , n367527 , n367528 );
buf ( n367530 , n19780 );
nand ( n19782 , n19765 , n367530 );
buf ( n367532 , n19782 );
and ( n19784 , n19762 , n367532 );
and ( n19785 , n367506 , n367510 );
or ( n19786 , n19784 , n19785 );
buf ( n367536 , n19786 );
buf ( n367537 , n367536 );
buf ( n367538 , n364779 );
not ( n19790 , n367538 );
buf ( n367540 , n367378 );
not ( n19792 , n367540 );
or ( n19793 , n19790 , n19792 );
buf ( n367543 , n582 );
not ( n19795 , n367543 );
buf ( n367545 , n365032 );
not ( n19797 , n367545 );
or ( n19798 , n19795 , n19797 );
buf ( n367548 , n365035 );
buf ( n367549 , n364797 );
nand ( n19801 , n367548 , n367549 );
buf ( n367551 , n19801 );
buf ( n367552 , n367551 );
nand ( n19804 , n19798 , n367552 );
buf ( n367554 , n19804 );
buf ( n367555 , n367554 );
buf ( n367556 , n17133 );
nand ( n19808 , n367555 , n367556 );
buf ( n367558 , n19808 );
buf ( n367559 , n367558 );
nand ( n19811 , n19793 , n367559 );
buf ( n367561 , n19811 );
buf ( n367562 , n367561 );
xor ( n19814 , n367537 , n367562 );
xor ( n19815 , n367333 , n367337 );
xor ( n19816 , n19815 , n367356 );
buf ( n367566 , n19816 );
buf ( n367567 , n367566 );
and ( n19819 , n19814 , n367567 );
and ( n19820 , n367537 , n367562 );
or ( n19821 , n19819 , n19820 );
buf ( n367571 , n19821 );
buf ( n367572 , n367571 );
xor ( n19824 , n367477 , n367572 );
xor ( n19825 , n367361 , n367386 );
xor ( n19826 , n19825 , n367391 );
buf ( n367576 , n19826 );
buf ( n367577 , n367576 );
and ( n19829 , n19824 , n367577 );
and ( n19830 , n367477 , n367572 );
or ( n19831 , n19829 , n19830 );
buf ( n367581 , n19831 );
buf ( n367582 , n367581 );
and ( n19834 , n19702 , n367582 );
and ( n19835 , n367436 , n367450 );
or ( n19836 , n19834 , n19835 );
buf ( n367586 , n19836 );
buf ( n367587 , n367586 );
and ( n19839 , n19662 , n367587 );
and ( n19840 , n367406 , n367410 );
or ( n19841 , n19839 , n19840 );
buf ( n367591 , n19841 );
buf ( n367592 , n367591 );
and ( n19844 , n19429 , n367592 );
and ( n19845 , n367201 , n367205 );
or ( n19846 , n19844 , n19845 );
buf ( n367596 , n19846 );
nor ( n19848 , n367197 , n367596 );
xor ( n19849 , n366873 , n367098 );
xor ( n19850 , n19849 , n367103 );
buf ( n367600 , n19850 );
xor ( n19852 , n367186 , n367190 );
and ( n19853 , n19852 , n367195 );
and ( n19854 , n367186 , n367190 );
or ( n19855 , n19853 , n19854 );
buf ( n367605 , n19855 );
nor ( n19857 , n367600 , n367605 );
nor ( n19858 , n19331 , n19848 , n19857 );
not ( n19859 , n19858 );
xor ( n19860 , n367201 , n367205 );
xor ( n19861 , n19860 , n367592 );
buf ( n367611 , n19861 );
buf ( n367612 , n367611 );
not ( n19864 , n367612 );
buf ( n367614 , n19864 );
buf ( n367615 , n367614 );
xor ( n19867 , n367141 , n367158 );
xor ( n19868 , n19867 , n367176 );
buf ( n367618 , n19868 );
buf ( n367619 , n367618 );
buf ( n367620 , n591 );
not ( n19872 , n367620 );
buf ( n367622 , n19388 );
not ( n19874 , n367622 );
or ( n19875 , n19872 , n19874 );
buf ( n367625 , n590 );
not ( n19877 , n367625 );
buf ( n367627 , n365776 );
not ( n19879 , n367627 );
or ( n19880 , n19877 , n19879 );
buf ( n367630 , n590 );
not ( n19882 , n367630 );
buf ( n367632 , n365403 );
nand ( n19884 , n19882 , n367632 );
buf ( n367634 , n19884 );
buf ( n367635 , n367634 );
nand ( n19887 , n19880 , n367635 );
buf ( n367637 , n19887 );
buf ( n367638 , n367637 );
buf ( n19890 , n367638 );
buf ( n367640 , n19890 );
buf ( n367641 , n367640 );
buf ( n367642 , n365738 );
nand ( n19894 , n367641 , n367642 );
buf ( n367644 , n19894 );
buf ( n367645 , n367644 );
nand ( n19897 , n19875 , n367645 );
buf ( n367647 , n19897 );
buf ( n367648 , n367647 );
buf ( n367649 , n365351 );
not ( n19901 , n367649 );
buf ( n367651 , n367428 );
not ( n19903 , n367651 );
or ( n19904 , n19901 , n19903 );
buf ( n367654 , n586 );
not ( n19906 , n367654 );
buf ( n367656 , n19146 );
not ( n19908 , n367656 );
or ( n19909 , n19906 , n19908 );
buf ( n367659 , n17161 );
buf ( n367660 , n365334 );
nand ( n19912 , n367659 , n367660 );
buf ( n367662 , n19912 );
buf ( n367663 , n367662 );
nand ( n19915 , n19909 , n367663 );
buf ( n367665 , n19915 );
buf ( n367666 , n367665 );
buf ( n367667 , n365375 );
nand ( n19919 , n367666 , n367667 );
buf ( n367669 , n19919 );
buf ( n367670 , n367669 );
nand ( n19922 , n19904 , n367670 );
buf ( n367672 , n19922 );
buf ( n367673 , n367672 );
buf ( n367674 , n364925 );
not ( n19926 , n367674 );
buf ( n367676 , n367469 );
not ( n19928 , n367676 );
or ( n19929 , n19926 , n19928 );
buf ( n367679 , n584 );
not ( n19931 , n367679 );
buf ( n367681 , n365516 );
not ( n19933 , n367681 );
or ( n19934 , n19931 , n19933 );
buf ( n367684 , n17301 );
buf ( n367685 , n364771 );
nand ( n19937 , n367684 , n367685 );
buf ( n367687 , n19937 );
buf ( n367688 , n367687 );
nand ( n19940 , n19934 , n367688 );
buf ( n367690 , n19940 );
buf ( n367691 , n367690 );
buf ( n367692 , n364973 );
nand ( n19944 , n367691 , n367692 );
buf ( n367694 , n19944 );
buf ( n367695 , n367694 );
nand ( n19947 , n19929 , n367695 );
buf ( n367697 , n19947 );
buf ( n367698 , n367697 );
buf ( n367699 , n17037 );
not ( n19951 , n367699 );
buf ( n367701 , n367498 );
not ( n19953 , n367701 );
or ( n19954 , n19951 , n19953 );
buf ( n367704 , n578 );
not ( n19956 , n367704 );
buf ( n367706 , n12484 );
not ( n19958 , n367706 );
buf ( n367708 , n19958 );
buf ( n367709 , n367708 );
not ( n19961 , n367709 );
or ( n19962 , n19956 , n19961 );
buf ( n367712 , n12484 );
not ( n19964 , n367712 );
buf ( n367714 , n19964 );
buf ( n367715 , n367714 );
not ( n19967 , n367715 );
buf ( n367717 , n19967 );
buf ( n367718 , n367717 );
buf ( n367719 , n364727 );
nand ( n19971 , n367718 , n367719 );
buf ( n367721 , n19971 );
buf ( n367722 , n367721 );
nand ( n19974 , n19962 , n367722 );
buf ( n367724 , n19974 );
buf ( n367725 , n367724 );
buf ( n367726 , n17082 );
nand ( n19978 , n367725 , n367726 );
buf ( n367728 , n19978 );
buf ( n367729 , n367728 );
nand ( n19981 , n19954 , n367729 );
buf ( n367731 , n19981 );
buf ( n367732 , n367731 );
buf ( n367733 , C0 );
buf ( n367734 , n367733 );
xor ( n19988 , n367732 , n367734 );
buf ( n367736 , n17230 );
not ( n19990 , n367736 );
buf ( n367738 , n367526 );
not ( n19992 , n367738 );
or ( n19993 , n19990 , n19992 );
buf ( n367741 , n580 );
not ( n19995 , n367741 );
buf ( n367743 , n366127 );
not ( n19997 , n367743 );
or ( n19998 , n19995 , n19997 );
buf ( n367746 , n366982 );
buf ( n367747 , n364896 );
nand ( n20001 , n367746 , n367747 );
buf ( n367749 , n20001 );
buf ( n367750 , n367749 );
nand ( n20004 , n19998 , n367750 );
buf ( n367752 , n20004 );
buf ( n367753 , n367752 );
buf ( n367754 , n364885 );
nand ( n20008 , n367753 , n367754 );
buf ( n367756 , n20008 );
buf ( n367757 , n367756 );
nand ( n20011 , n19993 , n367757 );
buf ( n367759 , n20011 );
buf ( n367760 , n367759 );
and ( n20014 , n19988 , n367760 );
or ( n20016 , n20014 , C0 );
buf ( n367763 , n20016 );
buf ( n367764 , n367763 );
buf ( n367765 , n364779 );
not ( n20020 , n367765 );
buf ( n367767 , n367554 );
not ( n20022 , n367767 );
or ( n20023 , n20020 , n20022 );
buf ( n367770 , n582 );
not ( n20025 , n367770 );
buf ( n367772 , n365494 );
not ( n20027 , n367772 );
or ( n20028 , n20025 , n20027 );
buf ( n367775 , n365491 );
buf ( n367776 , n364797 );
nand ( n20031 , n367775 , n367776 );
buf ( n367778 , n20031 );
buf ( n367779 , n367778 );
nand ( n20034 , n20028 , n367779 );
buf ( n367781 , n20034 );
buf ( n367782 , n367781 );
buf ( n367783 , n17133 );
nand ( n20038 , n367782 , n367783 );
buf ( n367785 , n20038 );
buf ( n367786 , n367785 );
nand ( n20041 , n20023 , n367786 );
buf ( n367788 , n20041 );
buf ( n367789 , n367788 );
xor ( n20044 , n367764 , n367789 );
xor ( n20045 , n367506 , n367510 );
xor ( n20046 , n20045 , n367532 );
buf ( n367793 , n20046 );
buf ( n367794 , n367793 );
and ( n20049 , n20044 , n367794 );
and ( n20050 , n367764 , n367789 );
or ( n20051 , n20049 , n20050 );
buf ( n367798 , n20051 );
buf ( n367799 , n367798 );
xor ( n20054 , n367698 , n367799 );
xor ( n20055 , n367537 , n367562 );
xor ( n20056 , n20055 , n367567 );
buf ( n367803 , n20056 );
buf ( n367804 , n367803 );
and ( n20059 , n20054 , n367804 );
and ( n20060 , n367698 , n367799 );
or ( n20061 , n20059 , n20060 );
buf ( n367808 , n20061 );
buf ( n367809 , n367808 );
xor ( n20064 , n367673 , n367809 );
not ( n20065 , n17867 );
not ( n20066 , n19690 );
or ( n20067 , n20065 , n20066 );
buf ( n367814 , n588 );
not ( n20069 , n367814 );
buf ( n367816 , n365388 );
not ( n20071 , n367816 );
or ( n20072 , n20069 , n20071 );
buf ( n367819 , n365388 );
buf ( n367820 , n588 );
or ( n20075 , n367819 , n367820 );
buf ( n367822 , n20075 );
buf ( n367823 , n367822 );
nand ( n20078 , n20072 , n367823 );
buf ( n367825 , n20078 );
nand ( n20080 , n365646 , n367825 );
nand ( n20081 , n20067 , n20080 );
buf ( n367828 , n20081 );
and ( n20083 , n20064 , n367828 );
and ( n20084 , n367673 , n367809 );
or ( n20085 , n20083 , n20084 );
buf ( n367832 , n20085 );
buf ( n367833 , n367832 );
xor ( n20088 , n367648 , n367833 );
xor ( n20089 , n367231 , n367396 );
xor ( n20090 , n20089 , n367401 );
buf ( n367837 , n20090 );
buf ( n367838 , n367837 );
and ( n20093 , n20088 , n367838 );
and ( n20094 , n367648 , n367833 );
or ( n20095 , n20093 , n20094 );
buf ( n367842 , n20095 );
buf ( n367843 , n367842 );
xor ( n20098 , n367619 , n367843 );
xor ( n20099 , n367406 , n367410 );
xor ( n20100 , n20099 , n367587 );
buf ( n367847 , n20100 );
buf ( n367848 , n367847 );
and ( n20103 , n20098 , n367848 );
and ( n20104 , n367619 , n367843 );
or ( n20105 , n20103 , n20104 );
buf ( n367852 , n20105 );
buf ( n367853 , n367852 );
not ( n20108 , n367853 );
buf ( n367855 , n20108 );
buf ( n367856 , n367855 );
nand ( n20111 , n367615 , n367856 );
buf ( n367858 , n20111 );
not ( n20113 , n367858 );
xor ( n20114 , n367619 , n367843 );
xor ( n20115 , n20114 , n367848 );
buf ( n367862 , n20115 );
buf ( n367863 , n367862 );
xor ( n20118 , n367436 , n367450 );
xor ( n20119 , n20118 , n367582 );
buf ( n367866 , n20119 );
buf ( n367867 , n367866 );
buf ( n367868 , n591 );
not ( n20123 , n367868 );
buf ( n367870 , n367637 );
not ( n20125 , n367870 );
or ( n20126 , n20123 , n20125 );
and ( n20127 , n590 , n12418 );
not ( n20128 , n590 );
and ( n20129 , n20128 , n360086 );
or ( n20130 , n20127 , n20129 );
buf ( n367877 , n20130 );
buf ( n367878 , n365738 );
nand ( n20133 , n367877 , n367878 );
buf ( n367880 , n20133 );
buf ( n367881 , n367880 );
nand ( n20136 , n20126 , n367881 );
buf ( n367883 , n20136 );
buf ( n367884 , n367883 );
xor ( n20139 , n367477 , n367572 );
xor ( n20140 , n20139 , n367577 );
buf ( n367887 , n20140 );
buf ( n367888 , n367887 );
xor ( n20143 , n367884 , n367888 );
buf ( n367890 , C0 );
buf ( n367891 , n367890 );
buf ( n367892 , n17037 );
not ( n20149 , n367892 );
buf ( n367894 , n367724 );
not ( n20151 , n367894 );
or ( n20152 , n20149 , n20151 );
not ( n20153 , n578 );
buf ( n367898 , n19166 );
not ( n20155 , n367898 );
buf ( n367900 , n20155 );
not ( n20157 , n367900 );
or ( n20158 , n20153 , n20157 );
buf ( n367903 , n364727 );
buf ( n367904 , n19166 );
nand ( n20161 , n367903 , n367904 );
buf ( n367906 , n20161 );
nand ( n20163 , n20158 , n367906 );
buf ( n367908 , n20163 );
buf ( n367909 , n17082 );
nand ( n20166 , n367908 , n367909 );
buf ( n367911 , n20166 );
buf ( n367912 , n367911 );
nand ( n20169 , n20152 , n367912 );
buf ( n367914 , n20169 );
buf ( n367915 , n367914 );
xor ( n20172 , n367891 , n367915 );
buf ( n367917 , C0 );
buf ( n367918 , n367917 );
not ( n20176 , n17037 );
not ( n20177 , n20163 );
or ( n20178 , n20176 , n20177 );
buf ( n367922 , n578 );
not ( n20180 , n367922 );
or ( n20183 , n20180 , C0 );
buf ( n367925 , C1 );
buf ( n367926 , n367925 );
nand ( n20189 , n20183 , n367926 );
buf ( n367928 , n20189 );
nand ( n20191 , n367928 , n17082 );
nand ( n20192 , n20178 , n20191 );
buf ( n367931 , n20192 );
xor ( n20194 , n367918 , n367931 );
buf ( n367933 , C0 );
buf ( n367934 , n367933 );
buf ( n367935 , n17037 );
not ( n20198 , n367935 );
buf ( n367937 , n367928 );
not ( n20200 , n367937 );
or ( n20201 , n20198 , n20200 );
buf ( n367940 , n578 );
not ( n20203 , n367940 );
or ( n20206 , n20203 , C0 );
buf ( n367943 , C1 );
buf ( n367944 , n367943 );
nand ( n20212 , n20206 , n367944 );
buf ( n367946 , n20212 );
buf ( n367947 , n367946 );
buf ( n367948 , n17082 );
nand ( n20216 , n367947 , n367948 );
buf ( n367950 , n20216 );
buf ( n367951 , n367950 );
nand ( n20219 , n20201 , n367951 );
buf ( n367953 , n20219 );
buf ( n367954 , n367953 );
xor ( n20222 , n367934 , n367954 );
buf ( n367956 , C1 );
buf ( n367957 , n367956 );
buf ( n367958 , n579 );
buf ( n367959 , n580 );
and ( n20227 , n367958 , n367959 );
buf ( n367961 , n364727 );
nor ( n20229 , n20227 , n367961 );
buf ( n367963 , n20229 );
buf ( n367964 , n367963 );
and ( n20232 , n367957 , n367964 );
buf ( n367966 , n20232 );
buf ( n367967 , n367966 );
buf ( n367968 , n17037 );
not ( n20236 , n367968 );
buf ( n367970 , n367946 );
not ( n20238 , n367970 );
or ( n20239 , n20236 , n20238 );
buf ( n367973 , C0 );
buf ( n367974 , n364727 );
or ( n20242 , n367973 , n367974 );
nand ( n20243 , n20242 , C1 );
buf ( n367977 , n20243 );
buf ( n367978 , n367977 );
buf ( n367979 , n17082 );
nand ( n20247 , n367978 , n367979 );
buf ( n367981 , n20247 );
buf ( n367982 , n367981 );
nand ( n20250 , n20239 , n367982 );
buf ( n367984 , n20250 );
buf ( n367985 , n367984 );
and ( n20253 , n367967 , n367985 );
buf ( n367987 , n20253 );
buf ( n367988 , n367987 );
and ( n20256 , n20222 , n367988 );
or ( n20257 , n20256 , C0 );
buf ( n367991 , n20257 );
buf ( n367992 , n367991 );
and ( n20260 , n20194 , n367992 );
or ( n20262 , n20260 , C0 );
buf ( n367995 , n20262 );
buf ( n367996 , n367995 );
and ( n20265 , n20172 , n367996 );
or ( n20267 , n20265 , C0 );
buf ( n367999 , n20267 );
buf ( n368000 , n367999 );
xor ( n20270 , n367732 , n367734 );
xor ( n20271 , n20270 , n367760 );
buf ( n368003 , n20271 );
buf ( n368004 , n368003 );
xor ( n20274 , n368000 , n368004 );
buf ( n368006 , n364779 );
not ( n20276 , n368006 );
buf ( n368008 , n367781 );
not ( n20278 , n368008 );
or ( n20279 , n20276 , n20278 );
and ( n20280 , n12481 , n364797 );
not ( n20281 , n12481 );
and ( n20282 , n20281 , n582 );
or ( n20283 , n20280 , n20282 );
buf ( n368015 , n20283 );
buf ( n368016 , n17133 );
nand ( n20286 , n368015 , n368016 );
buf ( n368018 , n20286 );
buf ( n368019 , n368018 );
nand ( n20289 , n20279 , n368019 );
buf ( n368021 , n20289 );
buf ( n368022 , n368021 );
and ( n20292 , n20274 , n368022 );
and ( n20293 , n368000 , n368004 );
or ( n20294 , n20292 , n20293 );
buf ( n368026 , n20294 );
buf ( n368027 , n368026 );
buf ( n368028 , n364925 );
not ( n20298 , n368028 );
buf ( n368030 , n367690 );
not ( n20300 , n368030 );
or ( n20301 , n20298 , n20300 );
buf ( n368033 , n584 );
not ( n20303 , n368033 );
buf ( n368035 , n365063 );
not ( n20305 , n368035 );
or ( n20306 , n20303 , n20305 );
buf ( n368038 , n17372 );
buf ( n368039 , n364771 );
nand ( n20309 , n368038 , n368039 );
buf ( n368041 , n20309 );
buf ( n368042 , n368041 );
nand ( n20312 , n20306 , n368042 );
buf ( n368044 , n20312 );
buf ( n368045 , n368044 );
buf ( n368046 , n364973 );
nand ( n20316 , n368045 , n368046 );
buf ( n368048 , n20316 );
buf ( n368049 , n368048 );
nand ( n20319 , n20301 , n368049 );
buf ( n368051 , n20319 );
buf ( n368052 , n368051 );
xor ( n20322 , n368027 , n368052 );
xor ( n20323 , n367764 , n367789 );
xor ( n20324 , n20323 , n367794 );
buf ( n368056 , n20324 );
buf ( n368057 , n368056 );
and ( n20327 , n20322 , n368057 );
and ( n20328 , n368027 , n368052 );
or ( n20329 , n20327 , n20328 );
buf ( n368061 , n20329 );
buf ( n368062 , n368061 );
buf ( n368063 , n365351 );
not ( n20333 , n368063 );
buf ( n368065 , n367665 );
not ( n20335 , n368065 );
or ( n20336 , n20333 , n20335 );
and ( n20337 , n586 , n17725 );
not ( n20338 , n586 );
and ( n20339 , n20338 , n17174 );
or ( n20340 , n20337 , n20339 );
buf ( n368072 , n20340 );
buf ( n368073 , n365375 );
nand ( n20343 , n368072 , n368073 );
buf ( n368075 , n20343 );
buf ( n368076 , n368075 );
nand ( n20346 , n20336 , n368076 );
buf ( n368078 , n20346 );
buf ( n368079 , n368078 );
xor ( n20349 , n368062 , n368079 );
buf ( n368081 , n17867 );
not ( n20351 , n368081 );
buf ( n368083 , n367825 );
not ( n20353 , n368083 );
or ( n20354 , n20351 , n20353 );
buf ( n368086 , n365129 );
buf ( n368087 , n588 );
nand ( n20357 , n368086 , n368087 );
buf ( n368089 , n20357 );
buf ( n368090 , n368089 );
not ( n20360 , n368090 );
buf ( n368092 , n588 );
not ( n20362 , n368092 );
buf ( n368094 , n8303 );
nand ( n20364 , n20362 , n368094 );
buf ( n368096 , n20364 );
buf ( n368097 , n368096 );
not ( n20367 , n368097 );
or ( n20368 , n20360 , n20367 );
buf ( n368100 , n365646 );
nand ( n20370 , n20368 , n368100 );
buf ( n368102 , n20370 );
buf ( n368103 , n368102 );
nand ( n20373 , n20354 , n368103 );
buf ( n368105 , n20373 );
buf ( n368106 , n368105 );
and ( n20376 , n20349 , n368106 );
and ( n20377 , n368062 , n368079 );
or ( n20378 , n20376 , n20377 );
buf ( n368110 , n20378 );
buf ( n368111 , n368110 );
and ( n20381 , n20143 , n368111 );
and ( n20382 , n367884 , n367888 );
or ( n20383 , n20381 , n20382 );
buf ( n368115 , n20383 );
buf ( n368116 , n368115 );
xor ( n20386 , n367867 , n368116 );
xor ( n20387 , n367648 , n367833 );
xor ( n20388 , n20387 , n367838 );
buf ( n368120 , n20388 );
buf ( n368121 , n368120 );
and ( n20391 , n20386 , n368121 );
and ( n20392 , n367867 , n368116 );
or ( n20393 , n20391 , n20392 );
buf ( n368125 , n20393 );
buf ( n368126 , n368125 );
nor ( n20396 , n367863 , n368126 );
buf ( n368128 , n20396 );
buf ( n368129 , n368128 );
xor ( n20399 , n367867 , n368116 );
xor ( n20400 , n20399 , n368121 );
buf ( n368132 , n20400 );
xor ( n20402 , n367673 , n367809 );
xor ( n20403 , n20402 , n367828 );
buf ( n368135 , n20403 );
buf ( n368136 , n368135 );
xor ( n20406 , n367698 , n367799 );
xor ( n20407 , n20406 , n367804 );
buf ( n368139 , n20407 );
buf ( n368140 , n368139 );
buf ( n368141 , n365738 );
not ( n20411 , n368141 );
xor ( n20412 , n590 , n357316 );
buf ( n368144 , n20412 );
not ( n20414 , n368144 );
or ( n20415 , n20411 , n20414 );
buf ( n368147 , n20130 );
buf ( n368148 , n591 );
nand ( n20418 , n368147 , n368148 );
buf ( n368150 , n20418 );
buf ( n368151 , n368150 );
nand ( n20421 , n20415 , n368151 );
buf ( n368153 , n20421 );
buf ( n368154 , n368153 );
xor ( n20424 , n368140 , n368154 );
buf ( n368156 , n365351 );
not ( n20426 , n368156 );
buf ( n368158 , n20340 );
not ( n20428 , n368158 );
or ( n20429 , n20426 , n20428 );
buf ( n368161 , n586 );
not ( n20431 , n368161 );
buf ( n368163 , n364823 );
not ( n20433 , n368163 );
or ( n20434 , n20431 , n20433 );
buf ( n368166 , n365099 );
buf ( n368167 , n365334 );
nand ( n20437 , n368166 , n368167 );
buf ( n368169 , n20437 );
buf ( n368170 , n368169 );
nand ( n20440 , n20434 , n368170 );
buf ( n368172 , n20440 );
buf ( n368173 , n368172 );
buf ( n368174 , n365375 );
nand ( n20444 , n368173 , n368174 );
buf ( n368176 , n20444 );
buf ( n368177 , n368176 );
nand ( n20447 , n20429 , n368177 );
buf ( n368179 , n20447 );
buf ( n368180 , n368179 );
buf ( n368181 , n17230 );
not ( n20451 , n368181 );
buf ( n368183 , n367752 );
not ( n20453 , n368183 );
or ( n20454 , n20451 , n20453 );
buf ( n368186 , n580 );
not ( n20456 , n368186 );
buf ( n368188 , n366466 );
not ( n20458 , n368188 );
or ( n20459 , n20456 , n20458 );
buf ( n368191 , n364896 );
buf ( n368192 , n367492 );
nand ( n20462 , n368191 , n368192 );
buf ( n368194 , n20462 );
buf ( n368195 , n368194 );
nand ( n20465 , n20459 , n368195 );
buf ( n368197 , n20465 );
buf ( n368198 , n368197 );
buf ( n368199 , n364885 );
nand ( n20469 , n368198 , n368199 );
buf ( n368201 , n20469 );
buf ( n368202 , n368201 );
nand ( n20472 , n20454 , n368202 );
buf ( n368204 , n20472 );
buf ( n368205 , n368204 );
xor ( n20475 , n367891 , n367915 );
xor ( n20476 , n20475 , n367996 );
buf ( n368208 , n20476 );
buf ( n368209 , n368208 );
xor ( n20479 , n368205 , n368209 );
buf ( n368211 , n364779 );
not ( n20481 , n368211 );
buf ( n368213 , n20283 );
not ( n20483 , n368213 );
or ( n20484 , n20481 , n20483 );
buf ( n368216 , n582 );
not ( n20486 , n368216 );
buf ( n368218 , n18248 );
not ( n20488 , n368218 );
buf ( n368220 , n20488 );
buf ( n368221 , n368220 );
not ( n20491 , n368221 );
or ( n20492 , n20486 , n20491 );
nand ( n20493 , n364797 , n3564 );
buf ( n368225 , n20493 );
nand ( n20495 , n20492 , n368225 );
buf ( n368227 , n20495 );
buf ( n368228 , n368227 );
buf ( n368229 , n17133 );
nand ( n20499 , n368228 , n368229 );
buf ( n368231 , n20499 );
buf ( n368232 , n368231 );
nand ( n20502 , n20484 , n368232 );
buf ( n368234 , n20502 );
buf ( n368235 , n368234 );
and ( n20505 , n20479 , n368235 );
and ( n20506 , n368205 , n368209 );
or ( n20507 , n20505 , n20506 );
buf ( n368239 , n20507 );
buf ( n368240 , n368239 );
buf ( n368241 , n364925 );
not ( n20511 , n368241 );
buf ( n368243 , n368044 );
not ( n20513 , n368243 );
or ( n20514 , n20511 , n20513 );
and ( n20515 , n12483 , n364771 );
not ( n20516 , n12483 );
and ( n20517 , n20516 , n584 );
or ( n20518 , n20515 , n20517 );
buf ( n368250 , n20518 );
buf ( n368251 , n364973 );
nand ( n20521 , n368250 , n368251 );
buf ( n368253 , n20521 );
buf ( n368254 , n368253 );
nand ( n20524 , n20514 , n368254 );
buf ( n368256 , n20524 );
buf ( n368257 , n368256 );
xor ( n20527 , n368240 , n368257 );
xor ( n20528 , n368000 , n368004 );
xor ( n20529 , n20528 , n368022 );
buf ( n368261 , n20529 );
buf ( n368262 , n368261 );
and ( n20532 , n20527 , n368262 );
and ( n20533 , n368240 , n368257 );
or ( n20534 , n20532 , n20533 );
buf ( n368266 , n20534 );
buf ( n368267 , n368266 );
xor ( n20537 , n368180 , n368267 );
xor ( n20538 , n368027 , n368052 );
xor ( n20539 , n20538 , n368057 );
buf ( n368271 , n20539 );
buf ( n368272 , n368271 );
and ( n20542 , n20537 , n368272 );
and ( n20543 , n368180 , n368267 );
or ( n20544 , n20542 , n20543 );
buf ( n368276 , n20544 );
buf ( n368277 , n368276 );
and ( n20547 , n20424 , n368277 );
and ( n20548 , n368140 , n368154 );
or ( n20549 , n20547 , n20548 );
buf ( n368281 , n20549 );
buf ( n368282 , n368281 );
xor ( n20552 , n368136 , n368282 );
xor ( n20553 , n367884 , n367888 );
xor ( n20554 , n20553 , n368111 );
buf ( n368286 , n20554 );
buf ( n368287 , n368286 );
and ( n20557 , n20552 , n368287 );
and ( n20558 , n368136 , n368282 );
or ( n20559 , n20557 , n20558 );
buf ( n368291 , n20559 );
nor ( n20561 , n368132 , n368291 );
buf ( n368293 , n20561 );
nor ( n20563 , n368129 , n368293 );
buf ( n368295 , n20563 );
not ( n20565 , n368295 );
xor ( n20566 , n368136 , n368282 );
xor ( n20567 , n20566 , n368287 );
buf ( n368299 , n20567 );
buf ( n368300 , n368299 );
not ( n20570 , n368300 );
buf ( n368302 , n365129 );
buf ( n368303 , n588 );
not ( n20573 , n368303 );
buf ( n368305 , n17867 );
not ( n20575 , n368305 );
buf ( n368307 , n20575 );
buf ( n368308 , n368307 );
nor ( n20578 , n20573 , n368308 );
buf ( n368310 , n20578 );
buf ( n368311 , n368310 );
nand ( n20581 , n368302 , n368311 );
buf ( n368313 , n20581 );
buf ( n368314 , n368313 );
buf ( n368315 , n365129 );
not ( n20585 , n368315 );
buf ( n368317 , n368307 );
buf ( n368318 , n588 );
nor ( n20588 , n368317 , n368318 );
buf ( n368320 , n20588 );
buf ( n368321 , n368320 );
nand ( n20591 , n20585 , n368321 );
buf ( n368323 , n20591 );
buf ( n368324 , n368323 );
and ( n20594 , n588 , n19146 );
not ( n20595 , n588 );
and ( n20596 , n20595 , n17547 );
or ( n20597 , n20594 , n20596 );
buf ( n368329 , n20597 );
buf ( n368330 , n365646 );
nand ( n20600 , n368329 , n368330 );
buf ( n368332 , n20600 );
buf ( n368333 , n368332 );
nand ( n20603 , n368314 , n368324 , n368333 );
buf ( n368335 , n20603 );
buf ( n368336 , n368335 );
buf ( n368337 , n365351 );
not ( n20607 , n368337 );
buf ( n368339 , n368172 );
not ( n20609 , n368339 );
or ( n20610 , n20607 , n20609 );
buf ( n368342 , n586 );
not ( n20612 , n368342 );
buf ( n368344 , n365516 );
not ( n20614 , n368344 );
or ( n20615 , n20612 , n20614 );
buf ( n368347 , n17301 );
buf ( n368348 , n365334 );
nand ( n20618 , n368347 , n368348 );
buf ( n368350 , n20618 );
buf ( n368351 , n368350 );
nand ( n20621 , n20615 , n368351 );
buf ( n368353 , n20621 );
buf ( n368354 , n368353 );
buf ( n368355 , n365375 );
nand ( n20625 , n368354 , n368355 );
buf ( n368357 , n20625 );
buf ( n368358 , n368357 );
nand ( n20628 , n20610 , n368358 );
buf ( n368360 , n20628 );
buf ( n368361 , n368360 );
buf ( n368362 , n17230 );
not ( n20632 , n368362 );
buf ( n368364 , n368197 );
not ( n20634 , n368364 );
or ( n20635 , n20632 , n20634 );
buf ( n368367 , n580 );
not ( n20637 , n368367 );
buf ( n368369 , n367714 );
not ( n20639 , n368369 );
or ( n20640 , n20637 , n20639 );
buf ( n368372 , n364896 );
buf ( n368373 , n12484 );
nand ( n20643 , n368372 , n368373 );
buf ( n368375 , n20643 );
buf ( n368376 , n368375 );
nand ( n20646 , n20640 , n368376 );
buf ( n368378 , n20646 );
buf ( n368379 , n368378 );
buf ( n368380 , n364885 );
nand ( n20650 , n368379 , n368380 );
buf ( n368382 , n20650 );
buf ( n368383 , n368382 );
nand ( n20653 , n20635 , n368383 );
buf ( n368385 , n20653 );
buf ( n368386 , n368385 );
xor ( n20656 , n367918 , n367931 );
xor ( n20657 , n20656 , n367992 );
buf ( n368389 , n20657 );
buf ( n368390 , n368389 );
xor ( n20660 , n368386 , n368390 );
buf ( n368392 , n364779 );
not ( n20662 , n368392 );
buf ( n368394 , n368227 );
not ( n20664 , n368394 );
or ( n20665 , n20662 , n20664 );
buf ( n368397 , n582 );
not ( n20667 , n368397 );
buf ( n368399 , n12482 );
not ( n20669 , n368399 );
buf ( n368401 , n20669 );
buf ( n368402 , n368401 );
not ( n20672 , n368402 );
or ( n20673 , n20667 , n20672 );
buf ( n368405 , n12482 );
buf ( n368406 , n364797 );
nand ( n20676 , n368405 , n368406 );
buf ( n368408 , n20676 );
buf ( n368409 , n368408 );
nand ( n20679 , n20673 , n368409 );
buf ( n368411 , n20679 );
buf ( n368412 , n368411 );
buf ( n368413 , n17133 );
nand ( n20683 , n368412 , n368413 );
buf ( n368415 , n20683 );
buf ( n368416 , n368415 );
nand ( n20686 , n20665 , n368416 );
buf ( n368418 , n20686 );
buf ( n368419 , n368418 );
and ( n20689 , n20660 , n368419 );
and ( n20690 , n368386 , n368390 );
or ( n20691 , n20689 , n20690 );
buf ( n368423 , n20691 );
buf ( n368424 , n368423 );
nand ( n20694 , n364925 , n20518 );
and ( n20695 , n365491 , n364771 );
not ( n20696 , n365491 );
and ( n20697 , n20696 , n584 );
or ( n20698 , n20695 , n20697 );
buf ( n368430 , n20698 );
buf ( n368431 , n364973 );
nand ( n20701 , n368430 , n368431 );
buf ( n368433 , n20701 );
nand ( n20703 , n20694 , n368433 );
buf ( n368435 , n20703 );
xor ( n20705 , n368424 , n368435 );
xor ( n20706 , n368205 , n368209 );
xor ( n20707 , n20706 , n368235 );
buf ( n368439 , n20707 );
buf ( n368440 , n368439 );
and ( n20710 , n20705 , n368440 );
and ( n20711 , n368424 , n368435 );
or ( n20712 , n20710 , n20711 );
buf ( n368444 , n20712 );
buf ( n368445 , n368444 );
xor ( n20715 , n368361 , n368445 );
xor ( n20716 , n368240 , n368257 );
xor ( n20717 , n20716 , n368262 );
buf ( n368449 , n20717 );
buf ( n368450 , n368449 );
and ( n20720 , n20715 , n368450 );
and ( n20721 , n368361 , n368445 );
or ( n20722 , n20720 , n20721 );
buf ( n368454 , n20722 );
buf ( n368455 , n368454 );
xor ( n20725 , n368336 , n368455 );
buf ( n368457 , n365738 );
not ( n20727 , n368457 );
and ( n20728 , n590 , n365388 );
not ( n20729 , n590 );
and ( n20730 , n20729 , n357348 );
or ( n20731 , n20728 , n20730 );
buf ( n368463 , n20731 );
not ( n20733 , n368463 );
or ( n20734 , n20727 , n20733 );
buf ( n368466 , n20412 );
buf ( n368467 , n591 );
nand ( n20737 , n368466 , n368467 );
buf ( n368469 , n20737 );
buf ( n368470 , n368469 );
nand ( n20740 , n20734 , n368470 );
buf ( n368472 , n20740 );
buf ( n368473 , n368472 );
and ( n20743 , n20725 , n368473 );
and ( n20744 , n368336 , n368455 );
or ( n20745 , n20743 , n20744 );
buf ( n368477 , n20745 );
buf ( n368478 , n368477 );
xor ( n20748 , n368062 , n368079 );
xor ( n20749 , n20748 , n368106 );
buf ( n368481 , n20749 );
buf ( n368482 , n368481 );
xor ( n20752 , n368478 , n368482 );
xor ( n20753 , n368140 , n368154 );
xor ( n20754 , n20753 , n368277 );
buf ( n368486 , n20754 );
buf ( n368487 , n368486 );
and ( n20757 , n20752 , n368487 );
and ( n20758 , n368478 , n368482 );
or ( n20759 , n20757 , n20758 );
buf ( n368491 , n20759 );
buf ( n368492 , n368491 );
not ( n20762 , n368492 );
buf ( n368494 , n20762 );
buf ( n368495 , n368494 );
nand ( n20765 , n20570 , n368495 );
buf ( n368497 , n20765 );
xor ( n20767 , n368180 , n368267 );
xor ( n20768 , n20767 , n368272 );
buf ( n368500 , n20768 );
buf ( n368501 , n368500 );
buf ( n368502 , C0 );
buf ( n368503 , n368502 );
buf ( n368504 , n17230 );
not ( n20776 , n368504 );
buf ( n368506 , n368378 );
not ( n20778 , n368506 );
or ( n20779 , n20776 , n20778 );
and ( n20780 , n19166 , n364896 );
not ( n20781 , n19166 );
and ( n20782 , n20781 , n580 );
or ( n20783 , n20780 , n20782 );
buf ( n368513 , n20783 );
buf ( n368514 , n364885 );
nand ( n20786 , n368513 , n368514 );
buf ( n368516 , n20786 );
buf ( n368517 , n368516 );
nand ( n20789 , n20779 , n368517 );
buf ( n368519 , n20789 );
buf ( n368520 , n368519 );
xor ( n20792 , n368503 , n368520 );
buf ( n368522 , C0 );
buf ( n368523 , n368522 );
buf ( n368524 , n17197 );
not ( n20797 , n368524 );
buf ( n368526 , n20783 );
not ( n20799 , n368526 );
or ( n20800 , n20797 , n20799 );
buf ( n368529 , n580 );
not ( n20802 , n368529 );
or ( n20805 , n20802 , C0 );
buf ( n368532 , C1 );
buf ( n368533 , n368532 );
nand ( n20811 , n20805 , n368533 );
buf ( n368535 , n20811 );
buf ( n368536 , n368535 );
buf ( n368537 , n364885 );
nand ( n20815 , n368536 , n368537 );
buf ( n368539 , n20815 );
buf ( n368540 , n368539 );
nand ( n20818 , n20800 , n368540 );
buf ( n368542 , n20818 );
buf ( n368543 , n368542 );
xor ( n20821 , n368523 , n368543 );
buf ( n368545 , C0 );
buf ( n368546 , n368545 );
buf ( n368547 , n17197 );
not ( n20825 , n368547 );
buf ( n368549 , n368535 );
not ( n20827 , n368549 );
or ( n20828 , n20825 , n20827 );
buf ( n368552 , n580 );
not ( n20830 , n368552 );
or ( n20833 , n20830 , C0 );
buf ( n368555 , C1 );
buf ( n368556 , n368555 );
nand ( n20839 , n20833 , n368556 );
buf ( n368558 , n20839 );
buf ( n368559 , n368558 );
buf ( n368560 , n364885 );
nand ( n20843 , n368559 , n368560 );
buf ( n368562 , n20843 );
buf ( n368563 , n368562 );
nand ( n20846 , n20828 , n368563 );
buf ( n368565 , n20846 );
buf ( n368566 , n368565 );
xor ( n20849 , n368546 , n368566 );
buf ( n368568 , n17197 );
not ( n20851 , n368568 );
buf ( n368570 , n368558 );
not ( n20853 , n368570 );
or ( n20854 , n20851 , n20853 );
buf ( n368573 , C0 );
buf ( n368574 , n364896 );
or ( n20857 , n368573 , n368574 );
nand ( n20858 , n20857 , C1 );
buf ( n368577 , n20858 );
buf ( n368578 , n368577 );
buf ( n368579 , n364882 );
nand ( n20862 , n368578 , n368579 );
buf ( n368581 , n20862 );
buf ( n368582 , n368581 );
nand ( n20865 , n20854 , n368582 );
buf ( n368584 , n20865 );
buf ( n368585 , n368584 );
not ( n20868 , n368585 );
buf ( n368587 , C1 );
buf ( n368588 , n368587 );
buf ( n368589 , n581 );
buf ( n368590 , n582 );
nand ( n20873 , n368589 , n368590 );
buf ( n368592 , n20873 );
buf ( n368593 , n368592 );
buf ( n368594 , n580 );
nand ( n20877 , n368588 , n368593 , n368594 );
buf ( n368596 , n20877 );
buf ( n368597 , n368596 );
nor ( n20880 , n20868 , n368597 );
buf ( n368599 , n20880 );
buf ( n368600 , n368599 );
and ( n20883 , n20849 , n368600 );
or ( n20884 , n20883 , C0 );
buf ( n368603 , n20884 );
buf ( n368604 , n368603 );
and ( n20887 , n20821 , n368604 );
or ( n20889 , n20887 , C0 );
buf ( n368607 , n20889 );
buf ( n368608 , n368607 );
and ( n20892 , n20792 , n368608 );
or ( n20894 , n20892 , C0 );
buf ( n368611 , n20894 );
buf ( n368612 , n368611 );
xor ( n20897 , n368386 , n368390 );
xor ( n20898 , n20897 , n368419 );
buf ( n368615 , n20898 );
buf ( n368616 , n368615 );
xor ( n20901 , n368612 , n368616 );
buf ( n368618 , n364925 );
not ( n20903 , n368618 );
buf ( n368620 , n20698 );
not ( n20905 , n368620 );
or ( n20906 , n20903 , n20905 );
buf ( n368623 , n584 );
not ( n20908 , n368623 );
buf ( n368625 , n365475 );
not ( n20910 , n368625 );
or ( n20911 , n20908 , n20910 );
buf ( n368628 , n364771 );
buf ( n368629 , n12481 );
nand ( n20914 , n368628 , n368629 );
buf ( n368631 , n20914 );
buf ( n368632 , n368631 );
nand ( n20917 , n20911 , n368632 );
buf ( n368634 , n20917 );
buf ( n368635 , n368634 );
buf ( n368636 , n364973 );
nand ( n20921 , n368635 , n368636 );
buf ( n368638 , n20921 );
buf ( n368639 , n368638 );
nand ( n20924 , n20906 , n368639 );
buf ( n368641 , n20924 );
buf ( n368642 , n368641 );
and ( n20927 , n20901 , n368642 );
and ( n20928 , n368612 , n368616 );
or ( n20929 , n20927 , n20928 );
buf ( n368646 , n20929 );
buf ( n368647 , n368646 );
xor ( n20932 , n368424 , n368435 );
xor ( n20933 , n20932 , n368440 );
buf ( n368650 , n20933 );
buf ( n368651 , n368650 );
xor ( n20936 , n368647 , n368651 );
buf ( n368653 , n365351 );
not ( n20938 , n368653 );
buf ( n368655 , n368353 );
not ( n20940 , n368655 );
or ( n20941 , n20938 , n20940 );
buf ( n368658 , n586 );
buf ( n368659 , n17372 );
and ( n20944 , n368658 , n368659 );
not ( n20945 , n368658 );
buf ( n368662 , n365063 );
and ( n20947 , n20945 , n368662 );
nor ( n20948 , n20944 , n20947 );
buf ( n368665 , n20948 );
buf ( n368666 , n368665 );
buf ( n368667 , n365375 );
nand ( n20952 , n368666 , n368667 );
buf ( n368669 , n20952 );
buf ( n368670 , n368669 );
nand ( n20955 , n20941 , n368670 );
buf ( n368672 , n20955 );
buf ( n368673 , n368672 );
and ( n20958 , n20936 , n368673 );
and ( n20959 , n368647 , n368651 );
or ( n20960 , n20958 , n20959 );
buf ( n368677 , n20960 );
buf ( n368678 , n368677 );
buf ( n368679 , n17867 );
not ( n20964 , n368679 );
buf ( n368681 , n20597 );
not ( n20966 , n368681 );
or ( n20967 , n20964 , n20966 );
xnor ( n20968 , n588 , n17725 );
buf ( n368685 , n20968 );
buf ( n368686 , n365646 );
nand ( n20971 , n368685 , n368686 );
buf ( n368688 , n20971 );
buf ( n368689 , n368688 );
nand ( n20974 , n20967 , n368689 );
buf ( n368691 , n20974 );
buf ( n368692 , n368691 );
xor ( n20977 , n368678 , n368692 );
buf ( n368694 , n365738 );
not ( n20979 , n368694 );
and ( n20980 , n590 , n365129 );
not ( n20981 , n590 );
and ( n20982 , n20981 , n8303 );
or ( n20983 , n20980 , n20982 );
buf ( n368700 , n20983 );
not ( n20985 , n368700 );
or ( n20986 , n20979 , n20985 );
buf ( n368703 , n20731 );
buf ( n368704 , n591 );
nand ( n20989 , n368703 , n368704 );
buf ( n368706 , n20989 );
buf ( n368707 , n368706 );
nand ( n20992 , n20986 , n368707 );
buf ( n368709 , n20992 );
buf ( n368710 , n368709 );
and ( n20995 , n20977 , n368710 );
and ( n20996 , n368678 , n368692 );
or ( n20997 , n20995 , n20996 );
buf ( n368714 , n20997 );
buf ( n368715 , n368714 );
xor ( n21000 , n368501 , n368715 );
xor ( n21001 , n368336 , n368455 );
xor ( n21002 , n21001 , n368473 );
buf ( n368719 , n21002 );
buf ( n368720 , n368719 );
xor ( n21005 , n21000 , n368720 );
buf ( n368722 , n21005 );
not ( n21007 , n368722 );
xor ( n21008 , n368361 , n368445 );
xor ( n21009 , n21008 , n368450 );
buf ( n368726 , n21009 );
buf ( n368727 , n368726 );
buf ( n368728 , n17867 );
not ( n21013 , n368728 );
buf ( n368730 , n20968 );
not ( n21015 , n368730 );
or ( n21016 , n21013 , n21015 );
and ( n21017 , n588 , n365093 );
not ( n21018 , n588 );
and ( n21019 , n21018 , n17143 );
or ( n21020 , n21017 , n21019 );
buf ( n368737 , n21020 );
buf ( n368738 , n365646 );
nand ( n21023 , n368737 , n368738 );
buf ( n368740 , n21023 );
buf ( n368741 , n368740 );
nand ( n21026 , n21016 , n368741 );
buf ( n368743 , n21026 );
buf ( n368744 , n368743 );
buf ( n368745 , n364779 );
not ( n21030 , n368745 );
buf ( n368747 , n368411 );
not ( n21032 , n368747 );
or ( n21033 , n21030 , n21032 );
buf ( n368750 , n582 );
not ( n21035 , n368750 );
buf ( n368752 , n367492 );
not ( n21037 , n368752 );
buf ( n368754 , n21037 );
buf ( n368755 , n368754 );
not ( n21040 , n368755 );
or ( n21041 , n21035 , n21040 );
buf ( n368758 , n366469 );
buf ( n368759 , n364797 );
nand ( n21044 , n368758 , n368759 );
buf ( n368761 , n21044 );
buf ( n368762 , n368761 );
nand ( n21047 , n21041 , n368762 );
buf ( n368764 , n21047 );
buf ( n368765 , n368764 );
buf ( n368766 , n17133 );
nand ( n21051 , n368765 , n368766 );
buf ( n368768 , n21051 );
buf ( n368769 , n368768 );
nand ( n21054 , n21033 , n368769 );
buf ( n368771 , n21054 );
buf ( n368772 , n368771 );
xor ( n21057 , n368503 , n368520 );
xor ( n21058 , n21057 , n368608 );
buf ( n368775 , n21058 );
buf ( n368776 , n368775 );
xor ( n21061 , n368772 , n368776 );
buf ( n368778 , n364925 );
not ( n21063 , n368778 );
buf ( n368780 , n368634 );
not ( n21065 , n368780 );
or ( n21066 , n21063 , n21065 );
buf ( n368783 , n584 );
not ( n21068 , n368783 );
buf ( n368785 , n366145 );
not ( n21070 , n368785 );
or ( n21071 , n21068 , n21070 );
buf ( n368788 , n366028 );
buf ( n368789 , n364771 );
nand ( n21074 , n368788 , n368789 );
buf ( n368791 , n21074 );
buf ( n368792 , n368791 );
nand ( n21077 , n21071 , n368792 );
buf ( n368794 , n21077 );
buf ( n368795 , n368794 );
buf ( n368796 , n364973 );
nand ( n21081 , n368795 , n368796 );
buf ( n368798 , n21081 );
buf ( n368799 , n368798 );
nand ( n21084 , n21066 , n368799 );
buf ( n368801 , n21084 );
buf ( n368802 , n368801 );
and ( n21087 , n21061 , n368802 );
and ( n21088 , n368772 , n368776 );
or ( n21089 , n21087 , n21088 );
buf ( n368806 , n21089 );
buf ( n368807 , n368806 );
buf ( n368808 , n365351 );
not ( n21093 , n368808 );
buf ( n368810 , n368665 );
not ( n21095 , n368810 );
or ( n21096 , n21093 , n21095 );
and ( n21097 , n12483 , n365334 );
not ( n21098 , n12483 );
and ( n21099 , n21098 , n586 );
or ( n21100 , n21097 , n21099 );
buf ( n368817 , n21100 );
buf ( n368818 , n365375 );
nand ( n21103 , n368817 , n368818 );
buf ( n368820 , n21103 );
buf ( n368821 , n368820 );
nand ( n21106 , n21096 , n368821 );
buf ( n368823 , n21106 );
buf ( n368824 , n368823 );
xor ( n21109 , n368807 , n368824 );
xor ( n21110 , n368612 , n368616 );
xor ( n21111 , n21110 , n368642 );
buf ( n368828 , n21111 );
buf ( n368829 , n368828 );
and ( n21114 , n21109 , n368829 );
and ( n21115 , n368807 , n368824 );
or ( n21116 , n21114 , n21115 );
buf ( n368833 , n21116 );
buf ( n368834 , n368833 );
xor ( n21119 , n368744 , n368834 );
xor ( n21120 , n368647 , n368651 );
xor ( n21121 , n21120 , n368673 );
buf ( n368838 , n21121 );
buf ( n368839 , n368838 );
and ( n21124 , n21119 , n368839 );
and ( n21125 , n368744 , n368834 );
or ( n21126 , n21124 , n21125 );
buf ( n368843 , n21126 );
buf ( n368844 , n368843 );
xor ( n21129 , n368727 , n368844 );
xor ( n21130 , n368678 , n368692 );
xor ( n21131 , n21130 , n368710 );
buf ( n368848 , n21131 );
buf ( n368849 , n368848 );
and ( n21134 , n21129 , n368849 );
and ( n21135 , n368727 , n368844 );
or ( n21136 , n21134 , n21135 );
buf ( n368853 , n21136 );
not ( n21138 , n368853 );
and ( n21139 , n21007 , n21138 );
xor ( n21140 , n368478 , n368482 );
xor ( n21141 , n21140 , n368487 );
buf ( n368858 , n21141 );
buf ( n368859 , n368858 );
xor ( n21144 , n368501 , n368715 );
and ( n21145 , n21144 , n368720 );
and ( n21146 , n368501 , n368715 );
or ( n21147 , n21145 , n21146 );
buf ( n368864 , n21147 );
buf ( n368865 , n368864 );
nor ( n21150 , n368859 , n368865 );
buf ( n368867 , n21150 );
nor ( n21152 , n21139 , n368867 );
xor ( n21153 , n368727 , n368844 );
xor ( n21154 , n21153 , n368849 );
buf ( n368871 , n21154 );
buf ( n368872 , n368871 );
not ( n21157 , n368872 );
buf ( n368874 , n591 );
not ( n21159 , n368874 );
buf ( n368876 , n20983 );
not ( n21161 , n368876 );
or ( n21162 , n21159 , n21161 );
and ( n21163 , n590 , n19146 );
not ( n21164 , n590 );
and ( n21165 , n21164 , n17161 );
or ( n21166 , n21163 , n21165 );
buf ( n368883 , n21166 );
buf ( n368884 , n365738 );
nand ( n21169 , n368883 , n368884 );
buf ( n368886 , n21169 );
buf ( n368887 , n368886 );
nand ( n21172 , n21162 , n368887 );
buf ( n368889 , n21172 );
buf ( n368890 , n368889 );
buf ( n368891 , n17867 );
not ( n21176 , n368891 );
buf ( n368893 , n21020 );
not ( n21178 , n368893 );
or ( n21179 , n21176 , n21178 );
and ( n21180 , n588 , n364986 );
not ( n21181 , n588 );
and ( n21182 , n21181 , n17301 );
or ( n21183 , n21180 , n21182 );
buf ( n368900 , n21183 );
buf ( n368901 , n365646 );
nand ( n21186 , n368900 , n368901 );
buf ( n368903 , n21186 );
buf ( n368904 , n368903 );
nand ( n21189 , n21179 , n368904 );
buf ( n368906 , n21189 );
buf ( n368907 , n368906 );
buf ( n368908 , n364779 );
not ( n21193 , n368908 );
buf ( n368910 , n368764 );
not ( n21195 , n368910 );
or ( n21196 , n21193 , n21195 );
buf ( n368913 , n582 );
not ( n21198 , n368913 );
buf ( n368915 , n367708 );
not ( n21200 , n368915 );
or ( n21201 , n21198 , n21200 );
buf ( n368918 , n12484 );
buf ( n368919 , n364797 );
nand ( n21204 , n368918 , n368919 );
buf ( n368921 , n21204 );
buf ( n368922 , n368921 );
nand ( n21207 , n21201 , n368922 );
buf ( n368924 , n21207 );
buf ( n368925 , n368924 );
buf ( n368926 , n17133 );
nand ( n21211 , n368925 , n368926 );
buf ( n368928 , n21211 );
buf ( n368929 , n368928 );
nand ( n21214 , n21196 , n368929 );
buf ( n368931 , n21214 );
buf ( n368932 , n368931 );
xor ( n21217 , n368523 , n368543 );
xor ( n21218 , n21217 , n368604 );
buf ( n368935 , n21218 );
buf ( n368936 , n368935 );
xor ( n21221 , n368932 , n368936 );
buf ( n368938 , C0 );
buf ( n368939 , n368938 );
buf ( n368940 , n364779 );
not ( n21227 , n368940 );
buf ( n368942 , n368924 );
not ( n21229 , n368942 );
or ( n21230 , n21227 , n21229 );
and ( n21231 , n19166 , n364797 );
not ( n21232 , n19166 );
and ( n21233 , n21232 , n582 );
or ( n21234 , n21231 , n21233 );
buf ( n368949 , n21234 );
buf ( n368950 , n17133 );
nand ( n21237 , n368949 , n368950 );
buf ( n368952 , n21237 );
buf ( n368953 , n368952 );
nand ( n21240 , n21230 , n368953 );
buf ( n368955 , n21240 );
buf ( n368956 , n368955 );
xor ( n21243 , n368939 , n368956 );
buf ( n368958 , C0 );
buf ( n368959 , n368958 );
buf ( n368960 , n364779 );
not ( n21256 , n368960 );
buf ( n368962 , n21234 );
not ( n21258 , n368962 );
or ( n21259 , n21256 , n21258 );
buf ( n368965 , n582 );
not ( n21261 , n368965 );
or ( n21264 , n21261 , C0 );
buf ( n368968 , C1 );
buf ( n368969 , n368968 );
nand ( n21270 , n21264 , n368969 );
buf ( n368971 , n21270 );
buf ( n368972 , n368971 );
buf ( n368973 , n17133 );
nand ( n21274 , n368972 , n368973 );
buf ( n368975 , n21274 );
buf ( n368976 , n368975 );
nand ( n21277 , n21259 , n368976 );
buf ( n368978 , n21277 );
buf ( n368979 , n368978 );
xor ( n21280 , n368959 , n368979 );
buf ( n368981 , C0 );
buf ( n368982 , n368981 );
buf ( n368983 , n364779 );
not ( n21284 , n368983 );
buf ( n368985 , n368971 );
not ( n21286 , n368985 );
or ( n21287 , n21284 , n21286 );
buf ( n368988 , n582 );
not ( n21289 , n368988 );
or ( n21295 , n21289 , C0 );
buf ( n368991 , C1 );
buf ( n368992 , n368991 );
nand ( n21301 , n21295 , n368992 );
buf ( n368994 , n21301 );
buf ( n368995 , n368994 );
buf ( n368996 , n17133 );
nand ( n21305 , n368995 , n368996 );
buf ( n368998 , n21305 );
buf ( n368999 , n368998 );
nand ( n21308 , n21287 , n368999 );
buf ( n369001 , n21308 );
buf ( n369002 , n369001 );
xor ( n21311 , n368982 , n369002 );
buf ( n369004 , n364779 );
not ( n21313 , n369004 );
buf ( n369006 , n368994 );
not ( n21315 , n369006 );
or ( n21316 , n21313 , n21315 );
buf ( n369009 , C0 );
buf ( n369010 , n364797 );
or ( n21319 , n369009 , n369010 );
nand ( n21320 , n21319 , C1 );
buf ( n369013 , n21320 );
buf ( n369014 , n369013 );
buf ( n369015 , n17133 );
nand ( n21324 , n369014 , n369015 );
buf ( n369017 , n21324 );
buf ( n369018 , n369017 );
nand ( n21327 , n21316 , n369018 );
buf ( n369020 , n21327 );
buf ( n369021 , n369020 );
not ( n21330 , n369021 );
buf ( n369023 , C1 );
buf ( n369024 , n369023 );
buf ( n369025 , n583 );
buf ( n369026 , n584 );
and ( n21335 , n369025 , n369026 );
buf ( n369028 , n364797 );
nor ( n21337 , n21335 , n369028 );
buf ( n369030 , n21337 );
buf ( n369031 , n369030 );
and ( n21340 , n369024 , n369031 );
buf ( n369033 , n21340 );
buf ( n369034 , n369033 );
not ( n21343 , n369034 );
buf ( n369036 , n21343 );
buf ( n369037 , n369036 );
nor ( n21346 , n21330 , n369037 );
buf ( n369039 , n21346 );
buf ( n369040 , n369039 );
and ( n21349 , n21311 , n369040 );
or ( n21350 , n21349 , C0 );
buf ( n369043 , n21350 );
buf ( n369044 , n369043 );
and ( n21353 , n21280 , n369044 );
or ( n21355 , n21353 , C0 );
buf ( n369047 , n21355 );
buf ( n369048 , n369047 );
and ( n21358 , n21243 , n369048 );
or ( n21360 , n21358 , C0 );
buf ( n369051 , n21360 );
buf ( n369052 , n369051 );
and ( n21363 , n21221 , n369052 );
or ( n21365 , n21363 , C0 );
buf ( n369055 , n21365 );
buf ( n369056 , n369055 );
buf ( n369057 , n365351 );
not ( n21369 , n369057 );
buf ( n369059 , n21100 );
not ( n21371 , n369059 );
or ( n21372 , n21369 , n21371 );
buf ( n369062 , n586 );
not ( n21374 , n369062 );
buf ( n369064 , n365494 );
not ( n21376 , n369064 );
or ( n21377 , n21374 , n21376 );
buf ( n369067 , n365491 );
buf ( n369068 , n365334 );
nand ( n21380 , n369067 , n369068 );
buf ( n369070 , n21380 );
buf ( n369071 , n369070 );
nand ( n21383 , n21377 , n369071 );
buf ( n369073 , n21383 );
buf ( n369074 , n369073 );
buf ( n369075 , n365375 );
nand ( n21387 , n369074 , n369075 );
buf ( n369077 , n21387 );
buf ( n369078 , n369077 );
nand ( n21390 , n21372 , n369078 );
buf ( n369080 , n21390 );
buf ( n369081 , n369080 );
xor ( n21393 , n369056 , n369081 );
xor ( n21394 , n368772 , n368776 );
xor ( n21395 , n21394 , n368802 );
buf ( n369085 , n21395 );
buf ( n369086 , n369085 );
and ( n21398 , n21393 , n369086 );
and ( n21399 , n369056 , n369081 );
or ( n21400 , n21398 , n21399 );
buf ( n369090 , n21400 );
buf ( n369091 , n369090 );
xor ( n21403 , n368907 , n369091 );
xor ( n21404 , n368807 , n368824 );
xor ( n21405 , n21404 , n368829 );
buf ( n369095 , n21405 );
buf ( n369096 , n369095 );
and ( n21408 , n21403 , n369096 );
and ( n21409 , n368907 , n369091 );
or ( n21410 , n21408 , n21409 );
buf ( n369100 , n21410 );
buf ( n369101 , n369100 );
xor ( n21413 , n368890 , n369101 );
xor ( n21414 , n368744 , n368834 );
xor ( n21415 , n21414 , n368839 );
buf ( n369105 , n21415 );
buf ( n369106 , n369105 );
and ( n21418 , n21413 , n369106 );
and ( n21419 , n368890 , n369101 );
or ( n21420 , n21418 , n21419 );
buf ( n369110 , n21420 );
buf ( n369111 , n369110 );
not ( n21423 , n369111 );
buf ( n369113 , n21423 );
buf ( n369114 , n369113 );
nand ( n21426 , n21157 , n369114 );
buf ( n369116 , n21426 );
buf ( n369117 , n369116 );
not ( n21429 , n369117 );
buf ( n369119 , n591 );
not ( n21431 , n369119 );
and ( n21432 , n590 , n17725 );
not ( n21433 , n590 );
and ( n21434 , n21433 , n17174 );
or ( n21435 , n21432 , n21434 );
buf ( n369125 , n21435 );
not ( n21437 , n369125 );
or ( n21438 , n21431 , n21437 );
and ( n21439 , n590 , n364823 );
not ( n21440 , n590 );
and ( n21441 , n21440 , n364826 );
or ( n21442 , n21439 , n21441 );
buf ( n369132 , n21442 );
buf ( n369133 , n365738 );
nand ( n21445 , n369132 , n369133 );
buf ( n369135 , n21445 );
buf ( n369136 , n369135 );
nand ( n21448 , n21438 , n369136 );
buf ( n369138 , n21448 );
buf ( n369139 , n369138 );
buf ( n369140 , n364925 );
not ( n21452 , n369140 );
and ( n21453 , n366977 , n584 );
not ( n21454 , n366977 );
and ( n21455 , n21454 , n364771 );
or ( n21456 , n21453 , n21455 );
buf ( n369146 , n21456 );
not ( n21458 , n369146 );
or ( n21459 , n21452 , n21458 );
buf ( n369149 , n584 );
not ( n21461 , n369149 );
buf ( n369151 , n366466 );
not ( n21463 , n369151 );
or ( n21464 , n21461 , n21463 );
buf ( n369154 , n364771 );
buf ( n369155 , n367492 );
nand ( n21467 , n369154 , n369155 );
buf ( n369157 , n21467 );
buf ( n369158 , n369157 );
nand ( n21470 , n21464 , n369158 );
buf ( n369160 , n21470 );
buf ( n369161 , n369160 );
buf ( n369162 , n364973 );
nand ( n21474 , n369161 , n369162 );
buf ( n369164 , n21474 );
buf ( n369165 , n369164 );
nand ( n21477 , n21459 , n369165 );
buf ( n369167 , n21477 );
buf ( n369168 , n369167 );
xor ( n21480 , n368939 , n368956 );
xor ( n21481 , n21480 , n369048 );
buf ( n369171 , n21481 );
buf ( n369172 , n369171 );
xor ( n21484 , n369168 , n369172 );
buf ( n369174 , n365351 );
not ( n21486 , n369174 );
buf ( n369176 , n586 );
not ( n21488 , n369176 );
buf ( n369178 , n366043 );
not ( n21490 , n369178 );
or ( n21491 , n21488 , n21490 );
buf ( n369181 , n365334 );
buf ( n369182 , n12481 );
nand ( n21494 , n369181 , n369182 );
buf ( n369184 , n21494 );
buf ( n369185 , n369184 );
nand ( n21497 , n21491 , n369185 );
buf ( n369187 , n21497 );
buf ( n369188 , n369187 );
not ( n21500 , n369188 );
or ( n21501 , n21486 , n21500 );
buf ( n369191 , n586 );
not ( n21503 , n369191 );
buf ( n369193 , n368220 );
not ( n21505 , n369193 );
or ( n21506 , n21503 , n21505 );
buf ( n369196 , n368220 );
not ( n21508 , n369196 );
buf ( n369198 , n21508 );
buf ( n369199 , n369198 );
buf ( n369200 , n365334 );
nand ( n21512 , n369199 , n369200 );
buf ( n369202 , n21512 );
buf ( n369203 , n369202 );
nand ( n21515 , n21506 , n369203 );
buf ( n369205 , n21515 );
buf ( n369206 , n369205 );
buf ( n369207 , n365375 );
nand ( n21519 , n369206 , n369207 );
buf ( n369209 , n21519 );
buf ( n369210 , n369209 );
nand ( n21522 , n21501 , n369210 );
buf ( n369212 , n21522 );
buf ( n369213 , n369212 );
and ( n21525 , n21484 , n369213 );
and ( n21526 , n369168 , n369172 );
or ( n21527 , n21525 , n21526 );
buf ( n369217 , n21527 );
buf ( n369218 , n369217 );
buf ( n369219 , n17867 );
not ( n21531 , n369219 );
buf ( n369221 , n588 );
not ( n21533 , n369221 );
buf ( n369223 , n365063 );
not ( n21535 , n369223 );
or ( n21536 , n21533 , n21535 );
buf ( n369226 , n588 );
not ( n21538 , n369226 );
buf ( n369228 , n17372 );
nand ( n21540 , n21538 , n369228 );
buf ( n369230 , n21540 );
buf ( n369231 , n369230 );
nand ( n21543 , n21536 , n369231 );
buf ( n369233 , n21543 );
buf ( n369234 , n369233 );
not ( n21546 , n369234 );
or ( n21547 , n21531 , n21546 );
not ( n21548 , n365032 );
not ( n21549 , n588 );
or ( n21550 , n21548 , n21549 );
not ( n21551 , n588 );
nand ( n21552 , n21551 , n12483 );
nand ( n21553 , n21550 , n21552 );
nand ( n21554 , n21553 , n365646 );
buf ( n369244 , n21554 );
nand ( n21556 , n21547 , n369244 );
buf ( n369246 , n21556 );
buf ( n369247 , n369246 );
xor ( n21559 , n369218 , n369247 );
buf ( n369249 , n364925 );
not ( n21561 , n369249 );
buf ( n369251 , n368794 );
not ( n21563 , n369251 );
or ( n21564 , n21561 , n21563 );
buf ( n369254 , n21456 );
buf ( n369255 , n364973 );
nand ( n21567 , n369254 , n369255 );
buf ( n369257 , n21567 );
buf ( n369258 , n369257 );
nand ( n21570 , n21564 , n369258 );
buf ( n369260 , n21570 );
buf ( n369261 , n369260 );
xor ( n21573 , n368932 , n368936 );
xor ( n21574 , n21573 , n369052 );
buf ( n369264 , n21574 );
buf ( n369265 , n369264 );
xor ( n21577 , n369261 , n369265 );
buf ( n369267 , n365351 );
not ( n21579 , n369267 );
buf ( n369269 , n369073 );
not ( n21581 , n369269 );
or ( n21582 , n21579 , n21581 );
buf ( n369272 , n369187 );
buf ( n369273 , n365375 );
nand ( n21585 , n369272 , n369273 );
buf ( n369275 , n21585 );
buf ( n369276 , n369275 );
nand ( n21588 , n21582 , n369276 );
buf ( n369278 , n21588 );
buf ( n369279 , n369278 );
xor ( n21591 , n21577 , n369279 );
buf ( n369281 , n21591 );
buf ( n369282 , n369281 );
and ( n21594 , n21559 , n369282 );
and ( n21595 , n369218 , n369247 );
or ( n21596 , n21594 , n21595 );
buf ( n369286 , n21596 );
buf ( n369287 , n369286 );
xor ( n21599 , n369139 , n369287 );
xor ( n21600 , n369261 , n369265 );
and ( n21601 , n21600 , n369279 );
and ( n21602 , n369261 , n369265 );
or ( n21603 , n21601 , n21602 );
buf ( n369293 , n21603 );
buf ( n369294 , n369293 );
xor ( n21606 , n369056 , n369081 );
xor ( n21607 , n21606 , n369086 );
buf ( n369297 , n21607 );
buf ( n369298 , n369297 );
xor ( n21610 , n369294 , n369298 );
buf ( n369300 , n17867 );
not ( n21612 , n369300 );
buf ( n369302 , n21183 );
not ( n21614 , n369302 );
or ( n21615 , n21612 , n21614 );
buf ( n369305 , n369233 );
buf ( n369306 , n365646 );
nand ( n21618 , n369305 , n369306 );
buf ( n369308 , n21618 );
buf ( n369309 , n369308 );
nand ( n21621 , n21615 , n369309 );
buf ( n369311 , n21621 );
buf ( n369312 , n369311 );
xor ( n21624 , n21610 , n369312 );
buf ( n369314 , n21624 );
buf ( n369315 , n369314 );
and ( n21627 , n21599 , n369315 );
and ( n21628 , n369139 , n369287 );
or ( n21629 , n21627 , n21628 );
buf ( n369319 , n21629 );
not ( n21631 , n369319 );
xor ( n21632 , n369294 , n369298 );
and ( n21633 , n21632 , n369312 );
and ( n21634 , n369294 , n369298 );
or ( n21635 , n21633 , n21634 );
buf ( n369325 , n21635 );
buf ( n369326 , n369325 );
buf ( n369327 , n591 );
not ( n21639 , n369327 );
buf ( n369329 , n21166 );
not ( n21641 , n369329 );
or ( n21642 , n21639 , n21641 );
buf ( n369332 , n21435 );
buf ( n369333 , n365738 );
nand ( n21645 , n369332 , n369333 );
buf ( n369335 , n21645 );
buf ( n369336 , n369335 );
nand ( n21648 , n21642 , n369336 );
buf ( n369338 , n21648 );
buf ( n369339 , n369338 );
xor ( n21651 , n369326 , n369339 );
xor ( n21652 , n368907 , n369091 );
xor ( n21653 , n21652 , n369096 );
buf ( n369343 , n21653 );
buf ( n369344 , n369343 );
xor ( n21656 , n21651 , n369344 );
buf ( n369346 , n21656 );
not ( n21658 , n369346 );
and ( n21659 , n21631 , n21658 );
xor ( n21660 , n369139 , n369287 );
xor ( n21661 , n21660 , n369315 );
buf ( n369351 , n21661 );
buf ( n369352 , n369351 );
buf ( n369353 , n591 );
not ( n21665 , n369353 );
buf ( n369355 , n21442 );
not ( n21667 , n369355 );
or ( n21668 , n21665 , n21667 );
buf ( n369358 , n590 );
not ( n21670 , n369358 );
buf ( n369360 , n365516 );
not ( n21672 , n369360 );
or ( n21673 , n21670 , n21672 );
buf ( n369363 , n17301 );
buf ( n369364 , n590 );
not ( n21676 , n369364 );
buf ( n369366 , n21676 );
buf ( n369367 , n369366 );
nand ( n21679 , n369363 , n369367 );
buf ( n369369 , n21679 );
buf ( n369370 , n369369 );
nand ( n21682 , n21673 , n369370 );
buf ( n369372 , n21682 );
buf ( n369373 , n369372 );
buf ( n369374 , n365738 );
nand ( n21686 , n369373 , n369374 );
buf ( n369376 , n21686 );
buf ( n369377 , n369376 );
nand ( n21689 , n21668 , n369377 );
buf ( n369379 , n21689 );
buf ( n369380 , n369379 );
buf ( n369381 , n364925 );
not ( n21693 , n369381 );
buf ( n369383 , n369160 );
not ( n21695 , n369383 );
or ( n21696 , n21693 , n21695 );
buf ( n369386 , n584 );
not ( n21698 , n369386 );
buf ( n369388 , n367714 );
not ( n21700 , n369388 );
or ( n21701 , n21698 , n21700 );
buf ( n369391 , n367717 );
buf ( n369392 , n364771 );
nand ( n21704 , n369391 , n369392 );
buf ( n369394 , n21704 );
buf ( n369395 , n369394 );
nand ( n21707 , n21701 , n369395 );
buf ( n369397 , n21707 );
buf ( n369398 , n369397 );
buf ( n369399 , n364973 );
nand ( n21711 , n369398 , n369399 );
buf ( n369401 , n21711 );
buf ( n369402 , n369401 );
nand ( n21714 , n21696 , n369402 );
buf ( n369404 , n21714 );
buf ( n369405 , n369404 );
buf ( n369406 , C0 );
buf ( n369407 , n369406 );
xor ( n21721 , n369405 , n369407 );
buf ( n369409 , n365351 );
not ( n21723 , n369409 );
buf ( n369411 , n369205 );
not ( n21725 , n369411 );
or ( n21726 , n21723 , n21725 );
buf ( n369414 , n586 );
not ( n21728 , n369414 );
buf ( n369416 , n368401 );
not ( n21730 , n369416 );
or ( n21731 , n21728 , n21730 );
buf ( n369419 , n12482 );
buf ( n369420 , n365334 );
nand ( n21734 , n369419 , n369420 );
buf ( n369422 , n21734 );
buf ( n369423 , n369422 );
nand ( n21737 , n21731 , n369423 );
buf ( n369425 , n21737 );
buf ( n369426 , n369425 );
buf ( n369427 , n365375 );
nand ( n21741 , n369426 , n369427 );
buf ( n369429 , n21741 );
buf ( n369430 , n369429 );
nand ( n21744 , n21726 , n369430 );
buf ( n369432 , n21744 );
buf ( n369433 , n369432 );
and ( n21747 , n21721 , n369433 );
or ( n21749 , n21747 , C0 );
buf ( n369436 , n21749 );
buf ( n369437 , n369436 );
not ( n21752 , n365646 );
and ( n21753 , n588 , n365494 );
not ( n21754 , n588 );
and ( n21755 , n21754 , n365491 );
or ( n21756 , n21753 , n21755 );
not ( n21757 , n21756 );
or ( n21758 , n21752 , n21757 );
nand ( n21759 , n21553 , n17867 );
nand ( n21760 , n21758 , n21759 );
buf ( n369447 , n21760 );
xor ( n21762 , n369437 , n369447 );
xor ( n21763 , n369168 , n369172 );
xor ( n21764 , n21763 , n369213 );
buf ( n369451 , n21764 );
buf ( n369452 , n369451 );
and ( n21767 , n21762 , n369452 );
and ( n21768 , n369437 , n369447 );
or ( n21769 , n21767 , n21768 );
buf ( n369456 , n21769 );
buf ( n369457 , n369456 );
xor ( n21772 , n369380 , n369457 );
xor ( n21773 , n369218 , n369247 );
xor ( n21774 , n21773 , n369282 );
buf ( n369461 , n21774 );
buf ( n369462 , n369461 );
and ( n21777 , n21772 , n369462 );
and ( n21778 , n369380 , n369457 );
or ( n21779 , n21777 , n21778 );
buf ( n369466 , n21779 );
buf ( n369467 , n369466 );
nor ( n21782 , n369352 , n369467 );
buf ( n369469 , n21782 );
nor ( n21784 , n21659 , n369469 );
xor ( n21785 , n369380 , n369457 );
xor ( n21786 , n21785 , n369462 );
buf ( n369473 , n21786 );
buf ( n369474 , n369473 );
not ( n21789 , n369474 );
buf ( n369476 , C0 );
buf ( n369477 , n369476 );
buf ( n369478 , n364925 );
not ( n21795 , n369478 );
buf ( n369480 , n369397 );
not ( n21797 , n369480 );
or ( n21798 , n21795 , n21797 );
buf ( n369483 , n584 );
not ( n21800 , n369483 );
buf ( n369485 , n366946 );
not ( n21802 , n369485 );
or ( n21803 , n21800 , n21802 );
buf ( n369488 , n366949 );
buf ( n369489 , n364771 );
nand ( n21806 , n369488 , n369489 );
buf ( n369491 , n21806 );
buf ( n369492 , n369491 );
nand ( n21809 , n21803 , n369492 );
buf ( n369494 , n21809 );
buf ( n369495 , n369494 );
buf ( n369496 , n364973 );
nand ( n21813 , n369495 , n369496 );
buf ( n369498 , n21813 );
buf ( n369499 , n369498 );
nand ( n21816 , n21798 , n369499 );
buf ( n369501 , n21816 );
buf ( n369502 , n369501 );
xor ( n21819 , n369477 , n369502 );
buf ( n369504 , C0 );
buf ( n369505 , n369504 );
buf ( n369506 , C0 );
buf ( n369507 , n369506 );
buf ( n369508 , n584 );
not ( n21832 , n369508 );
or ( n21835 , n21832 , C0 );
buf ( n369511 , C1 );
buf ( n369512 , n369511 );
nand ( n21841 , n21835 , n369512 );
buf ( n369514 , n21841 );
not ( n21843 , n369514 );
not ( n21844 , n364925 );
or ( n21845 , n21843 , n21844 );
buf ( n369518 , n584 );
buf ( n369519 , n367267 );
and ( n21848 , n369518 , n369519 );
nor ( n21852 , n21848 , C0 );
buf ( n369522 , n21852 );
buf ( n369523 , n369522 );
not ( n21855 , n369523 );
buf ( n369525 , n364973 );
nand ( n21857 , n21855 , n369525 );
buf ( n369527 , n21857 );
nand ( n21859 , n21845 , n369527 );
buf ( n369529 , n21859 );
xor ( n21861 , n369507 , n369529 );
buf ( n369531 , C1 );
buf ( n369532 , n369531 );
buf ( n369533 , n585 );
buf ( n369534 , n586 );
and ( n21866 , n369533 , n369534 );
buf ( n369536 , n364771 );
nor ( n21868 , n21866 , n369536 );
buf ( n369538 , n21868 );
buf ( n369539 , n369538 );
and ( n21871 , n369532 , n369539 );
buf ( n369541 , n21871 );
buf ( n369542 , n369541 );
buf ( n369543 , n369522 );
buf ( n369544 , n365406 );
or ( n21876 , n369543 , n369544 );
buf ( n369546 , C1 );
buf ( n369547 , n369546 );
buf ( n369548 , n364973 );
not ( n21880 , n369548 );
buf ( n369550 , n21880 );
buf ( n369551 , n369550 );
buf ( n369552 , n364771 );
nor ( n21884 , n369551 , n369552 );
buf ( n369554 , n21884 );
buf ( n369555 , n369554 );
and ( n21887 , n369547 , n369555 );
nor ( n21888 , C0 , n21887 );
buf ( n369558 , n21888 );
buf ( n369559 , n369558 );
nand ( n21891 , n21876 , n369559 );
buf ( n369561 , n21891 );
buf ( n369562 , n369561 );
and ( n21894 , n369542 , n369562 );
buf ( n369564 , n21894 );
buf ( n369565 , n369564 );
and ( n21897 , n21861 , n369565 );
or ( n21898 , n21897 , C0 );
buf ( n369568 , n21898 );
buf ( n369569 , n369568 );
xor ( n21901 , n369505 , n369569 );
buf ( n369571 , n364925 );
not ( n21903 , n369571 );
buf ( n369573 , n369494 );
not ( n21905 , n369573 );
or ( n21906 , n21903 , n21905 );
buf ( n369576 , n369514 );
buf ( n369577 , n364973 );
nand ( n21909 , n369576 , n369577 );
buf ( n369579 , n21909 );
buf ( n369580 , n369579 );
nand ( n21912 , n21906 , n369580 );
buf ( n369582 , n21912 );
buf ( n369583 , n369582 );
and ( n21915 , n21901 , n369583 );
or ( n21917 , n21915 , C0 );
buf ( n369586 , n21917 );
buf ( n369587 , n369586 );
and ( n21920 , n21819 , n369587 );
or ( n21922 , n21920 , C0 );
buf ( n369590 , n21922 );
buf ( n369591 , n369590 );
xor ( n21925 , n369405 , n369407 );
xor ( n21926 , n21925 , n369433 );
buf ( n369594 , n21926 );
buf ( n369595 , n369594 );
xor ( n21929 , n369591 , n369595 );
buf ( n369597 , n17867 );
not ( n21931 , n369597 );
buf ( n369599 , n21756 );
not ( n21933 , n369599 );
or ( n21934 , n21931 , n21933 );
and ( n21935 , n588 , n366043 );
not ( n21936 , n588 );
and ( n21937 , n21936 , n12481 );
or ( n21938 , n21935 , n21937 );
buf ( n369606 , n21938 );
buf ( n369607 , n365646 );
nand ( n21941 , n369606 , n369607 );
buf ( n369609 , n21941 );
buf ( n369610 , n369609 );
nand ( n21944 , n21934 , n369610 );
buf ( n369612 , n21944 );
buf ( n369613 , n369612 );
and ( n21947 , n21929 , n369613 );
and ( n21948 , n369591 , n369595 );
or ( n21949 , n21947 , n21948 );
buf ( n369617 , n21949 );
buf ( n369618 , n369617 );
xor ( n21952 , n369437 , n369447 );
xor ( n21953 , n21952 , n369452 );
buf ( n369621 , n21953 );
buf ( n369622 , n369621 );
xor ( n21956 , n369618 , n369622 );
buf ( n369624 , n591 );
not ( n21958 , n369624 );
buf ( n369626 , n369372 );
not ( n21960 , n369626 );
or ( n21961 , n21958 , n21960 );
buf ( n369629 , n590 );
not ( n21963 , n369629 );
buf ( n369631 , n365063 );
not ( n21965 , n369631 );
or ( n21966 , n21963 , n21965 );
buf ( n369634 , n590 );
not ( n21968 , n369634 );
buf ( n369636 , n17372 );
nand ( n21970 , n21968 , n369636 );
buf ( n369638 , n21970 );
buf ( n369639 , n369638 );
nand ( n21973 , n21966 , n369639 );
buf ( n369641 , n21973 );
buf ( n369642 , n369641 );
buf ( n369643 , n365738 );
nand ( n21977 , n369642 , n369643 );
buf ( n369645 , n21977 );
buf ( n369646 , n369645 );
nand ( n21980 , n21961 , n369646 );
buf ( n369648 , n21980 );
buf ( n369649 , n369648 );
and ( n21983 , n21956 , n369649 );
and ( n21984 , n369618 , n369622 );
or ( n21985 , n21983 , n21984 );
buf ( n369653 , n21985 );
buf ( n369654 , n369653 );
not ( n21988 , n369654 );
buf ( n369656 , n21988 );
buf ( n369657 , n369656 );
nand ( n21991 , n21789 , n369657 );
buf ( n369659 , n21991 );
not ( n21993 , n369659 );
buf ( n369661 , C0 );
buf ( n369662 , n369661 );
buf ( n369663 , n365347 );
not ( n21999 , n369663 );
buf ( n369665 , n586 );
not ( n22001 , n369665 );
buf ( n369667 , n367708 );
not ( n22003 , n369667 );
or ( n22004 , n22001 , n22003 );
buf ( n369670 , n12484 );
buf ( n369671 , n365334 );
nand ( n22007 , n369670 , n369671 );
buf ( n369673 , n22007 );
buf ( n369674 , n369673 );
nand ( n22010 , n22004 , n369674 );
buf ( n369676 , n22010 );
buf ( n369677 , n369676 );
not ( n22013 , n369677 );
or ( n22014 , n21999 , n22013 );
buf ( n369680 , n586 );
not ( n22016 , n369680 );
buf ( n369682 , n367900 );
not ( n22018 , n369682 );
or ( n22019 , n22016 , n22018 );
buf ( n369685 , n366949 );
buf ( n369686 , n365334 );
nand ( n22022 , n369685 , n369686 );
buf ( n369688 , n22022 );
buf ( n369689 , n369688 );
nand ( n22025 , n22019 , n369689 );
buf ( n369691 , n22025 );
buf ( n369692 , n369691 );
buf ( n369693 , n365375 );
nand ( n22029 , n369692 , n369693 );
buf ( n369695 , n22029 );
buf ( n369696 , n369695 );
nand ( n22032 , n22014 , n369696 );
buf ( n369698 , n22032 );
buf ( n369699 , n369698 );
xor ( n22035 , n369662 , n369699 );
buf ( n369701 , C0 );
buf ( n369702 , n369701 );
buf ( n369703 , C0 );
buf ( n369704 , n369703 );
not ( n22043 , n365347 );
nor ( n22044 , n22043 , n365334 );
nand ( n22045 , C1 , n22044 );
buf ( n369708 , n586 );
not ( n22048 , n369708 );
or ( n22051 , n22048 , C0 );
buf ( n369711 , C1 );
buf ( n369712 , n369711 );
nand ( n22057 , n22051 , n369712 );
buf ( n369714 , n22057 );
nand ( n22059 , n369714 , n365375 );
nand ( n22060 , n22045 , C1 , n22059 );
buf ( n369717 , n22060 );
xor ( n22062 , n369704 , n369717 );
buf ( n369719 , C1 );
buf ( n369720 , n369719 );
buf ( n369721 , n587 );
buf ( n369722 , n588 );
and ( n22067 , n369721 , n369722 );
buf ( n369724 , n365334 );
nor ( n22069 , n22067 , n369724 );
buf ( n369726 , n22069 );
buf ( n369727 , n369726 );
and ( n22072 , n369720 , n369727 );
buf ( n369729 , n22072 );
buf ( n369730 , n369729 );
not ( n22075 , n369730 );
buf ( n369732 , n369714 );
buf ( n369733 , n365347 );
and ( n22078 , n369732 , n369733 );
buf ( n369735 , n369546 );
buf ( n369736 , n586 );
and ( n22081 , n369735 , n369736 );
nor ( n22082 , n22081 , C0 );
buf ( n369739 , n22082 );
buf ( n369740 , n369739 );
buf ( n369741 , n365375 );
not ( n22086 , n369741 );
buf ( n369743 , n22086 );
buf ( n369744 , n369743 );
nor ( n22089 , n369740 , n369744 );
buf ( n369746 , n22089 );
buf ( n369747 , n369746 );
nor ( n22092 , n22078 , n369747 );
buf ( n369749 , n22092 );
buf ( n369750 , n369749 );
nor ( n22095 , n22075 , n369750 );
buf ( n369752 , n22095 );
buf ( n369753 , n369752 );
and ( n22098 , n22062 , n369753 );
or ( n22099 , n22098 , C0 );
buf ( n369756 , n22099 );
buf ( n369757 , n369756 );
xor ( n22102 , n369702 , n369757 );
buf ( n369759 , n365347 );
not ( n22104 , n369759 );
buf ( n369761 , n369691 );
not ( n22106 , n369761 );
or ( n22107 , n22104 , n22106 );
and ( n22108 , n365334 , C1 );
nor ( n22111 , n22108 , C0 );
nand ( n22112 , n22111 , n365375 );
buf ( n369767 , n22112 );
nand ( n22114 , n22107 , n369767 );
buf ( n369769 , n22114 );
buf ( n369770 , n369769 );
and ( n22117 , n22102 , n369770 );
or ( n22119 , n22117 , C0 );
buf ( n369773 , n22119 );
buf ( n369774 , n369773 );
and ( n22122 , n22035 , n369774 );
or ( n22124 , n22122 , C0 );
buf ( n369777 , n22124 );
buf ( n369778 , n369777 );
buf ( n369779 , n365351 );
not ( n22128 , n369779 );
buf ( n369781 , n586 );
not ( n22130 , n369781 );
buf ( n369783 , n368754 );
not ( n22132 , n369783 );
or ( n22133 , n22130 , n22132 );
buf ( n369786 , n366469 );
buf ( n369787 , n365334 );
nand ( n22136 , n369786 , n369787 );
buf ( n369789 , n22136 );
buf ( n369790 , n369789 );
nand ( n22139 , n22133 , n369790 );
buf ( n369792 , n22139 );
buf ( n369793 , n369792 );
not ( n22142 , n369793 );
or ( n22143 , n22128 , n22142 );
buf ( n369796 , n369676 );
buf ( n369797 , n365375 );
nand ( n22146 , n369796 , n369797 );
buf ( n369799 , n22146 );
buf ( n369800 , n369799 );
nand ( n22149 , n22143 , n369800 );
buf ( n369802 , n22149 );
buf ( n369803 , n369802 );
buf ( n369804 , C0 );
buf ( n369805 , n369804 );
xor ( n22156 , n369803 , n369805 );
buf ( n369807 , n17867 );
not ( n22158 , n369807 );
xor ( n22159 , n588 , n18248 );
buf ( n369810 , n22159 );
not ( n22161 , n369810 );
or ( n22162 , n22158 , n22161 );
buf ( n369813 , n588 );
not ( n22164 , n369813 );
buf ( n369815 , n366124 );
not ( n22166 , n369815 );
or ( n22167 , n22164 , n22166 );
buf ( n369818 , n588 );
not ( n22169 , n369818 );
buf ( n369820 , n12482 );
nand ( n22171 , n22169 , n369820 );
buf ( n369822 , n22171 );
buf ( n369823 , n369822 );
nand ( n22174 , n22167 , n369823 );
buf ( n369825 , n22174 );
buf ( n369826 , n369825 );
buf ( n369827 , n365646 );
nand ( n22178 , n369826 , n369827 );
buf ( n369829 , n22178 );
buf ( n369830 , n369829 );
nand ( n22181 , n22162 , n369830 );
buf ( n369832 , n22181 );
buf ( n369833 , n369832 );
xor ( n22184 , n22156 , n369833 );
buf ( n369835 , n22184 );
buf ( n369836 , n369835 );
xor ( n22187 , n369778 , n369836 );
buf ( n369838 , n591 );
not ( n22189 , n369838 );
and ( n22190 , n590 , n365494 );
not ( n22191 , n590 );
and ( n22192 , n22191 , n365491 );
or ( n22193 , n22190 , n22192 );
buf ( n369844 , n22193 );
not ( n22195 , n369844 );
or ( n22196 , n22189 , n22195 );
buf ( n369847 , n590 );
not ( n22198 , n369847 );
buf ( n369849 , n365475 );
not ( n22200 , n369849 );
or ( n22201 , n22198 , n22200 );
buf ( n369852 , n590 );
not ( n22203 , n369852 );
buf ( n369854 , n12481 );
nand ( n22205 , n22203 , n369854 );
buf ( n369856 , n22205 );
buf ( n369857 , n369856 );
nand ( n22208 , n22201 , n369857 );
buf ( n369859 , n22208 );
buf ( n369860 , n369859 );
buf ( n369861 , n365735 );
nand ( n22212 , n369860 , n369861 );
buf ( n369863 , n22212 );
buf ( n369864 , n369863 );
nand ( n22215 , n22196 , n369864 );
buf ( n369866 , n22215 );
buf ( n369867 , n369866 );
xor ( n22218 , n22187 , n369867 );
buf ( n369869 , n22218 );
not ( n22220 , n369869 );
buf ( n369871 , n17867 );
not ( n22222 , n369871 );
buf ( n369873 , n369825 );
not ( n22224 , n369873 );
or ( n22225 , n22222 , n22224 );
and ( n22226 , n588 , n366466 );
not ( n22227 , n588 );
and ( n22228 , n22227 , n367492 );
or ( n22229 , n22226 , n22228 );
buf ( n369880 , n22229 );
buf ( n369881 , n365646 );
nand ( n22232 , n369880 , n369881 );
buf ( n369883 , n22232 );
buf ( n369884 , n369883 );
nand ( n22235 , n22225 , n369884 );
buf ( n369886 , n22235 );
buf ( n369887 , n369886 );
xor ( n22238 , n369662 , n369699 );
xor ( n22239 , n22238 , n369774 );
buf ( n369890 , n22239 );
buf ( n369891 , n369890 );
xor ( n22242 , n369887 , n369891 );
buf ( n369893 , n591 );
not ( n22244 , n369893 );
buf ( n369895 , n369859 );
not ( n22246 , n369895 );
or ( n22247 , n22244 , n22246 );
and ( n22248 , n18248 , n590 );
not ( n22249 , n18248 );
and ( n22250 , n22249 , n347484 );
nor ( n22251 , n22248 , n22250 );
buf ( n369902 , n22251 );
buf ( n369903 , n365735 );
nand ( n22254 , n369902 , n369903 );
buf ( n369905 , n22254 );
buf ( n369906 , n369905 );
nand ( n22257 , n22247 , n369906 );
buf ( n369908 , n22257 );
buf ( n369909 , n369908 );
and ( n22260 , n22242 , n369909 );
and ( n22261 , n369887 , n369891 );
or ( n22262 , n22260 , n22261 );
buf ( n369913 , n22262 );
not ( n22264 , n369913 );
nand ( n22265 , n22220 , n22264 );
buf ( n369916 , n22265 );
not ( n22267 , n369916 );
buf ( n369918 , C0 );
buf ( n369919 , n17867 );
not ( n22271 , n369919 );
buf ( n369921 , n588 );
not ( n22275 , n369921 );
buf ( n369923 , n367900 );
and ( n22277 , n22275 , n369923 );
nor ( n22278 , C0 , n22277 );
buf ( n369926 , n22278 );
buf ( n369927 , n369926 );
not ( n22281 , n369927 );
or ( n22282 , n22271 , n22281 );
and ( n22283 , n588 , n367256 );
or ( n22286 , n22283 , C0 );
buf ( n369932 , n22286 );
buf ( n369933 , n365646 );
nand ( n22289 , n369932 , n369933 );
buf ( n369935 , n22289 );
buf ( n369936 , n369935 );
nand ( n22292 , n22282 , n369936 );
buf ( n369938 , n22292 );
buf ( n369939 , n369938 );
buf ( n369940 , C0 );
buf ( n369941 , n369940 );
not ( n22298 , n365646 );
buf ( n369943 , n588 );
not ( n22300 , n369943 );
buf ( n369945 , n369546 );
and ( n22302 , n22300 , n369945 );
nor ( n22303 , C0 , n22302 );
buf ( n369948 , n22303 );
not ( n22305 , n369948 );
or ( n22306 , n22298 , n22305 );
and ( n22309 , C1 , n17631 );
nor ( n22310 , C0 , n22309 );
nand ( n22311 , n22310 , n17867 );
nand ( n22312 , n22306 , n22311 );
buf ( n369955 , n22312 );
not ( n22314 , n369955 );
buf ( n369957 , C1 );
buf ( n369958 , n369957 );
buf ( n369959 , n589 );
buf ( n369960 , n590 );
nand ( n22319 , n369959 , n369960 );
buf ( n369962 , n22319 );
buf ( n369963 , n369962 );
buf ( n369964 , n588 );
nand ( n22323 , n369958 , n369963 , n369964 );
buf ( n369966 , n22323 );
buf ( n369967 , n369966 );
nor ( n22326 , n22314 , n369967 );
buf ( n369969 , n22326 );
buf ( n369970 , n369969 );
xor ( n22329 , n369941 , n369970 );
buf ( n369972 , n17867 );
not ( n22331 , n369972 );
buf ( n369974 , n22286 );
not ( n22333 , n369974 );
or ( n22334 , n22331 , n22333 );
buf ( n369977 , n22310 );
buf ( n369978 , n365646 );
nand ( n22337 , n369977 , n369978 );
buf ( n369980 , n22337 );
buf ( n369981 , n369980 );
nand ( n22340 , n22334 , n369981 );
buf ( n369983 , n22340 );
buf ( n369984 , n369983 );
and ( n22343 , n22329 , n369984 );
or ( n22344 , n22343 , C0 );
buf ( n369987 , n22344 );
buf ( n369988 , n369987 );
buf ( n369989 , C0 );
buf ( n369990 , n591 );
not ( n22351 , n369990 );
buf ( n369992 , n590 );
not ( n22353 , n369992 );
buf ( n369994 , n366466 );
not ( n22355 , n369994 );
or ( n22356 , n22353 , n22355 );
buf ( n369997 , n590 );
not ( n22358 , n369997 );
buf ( n369999 , n367492 );
nand ( n22360 , n22358 , n369999 );
buf ( n370001 , n22360 );
buf ( n370002 , n370001 );
nand ( n22363 , n22356 , n370002 );
buf ( n370004 , n22363 );
buf ( n370005 , n370004 );
not ( n22366 , n370005 );
or ( n22367 , n22351 , n22366 );
buf ( n370008 , n365732 );
buf ( n370009 , n590 );
not ( n22370 , n370009 );
buf ( n370011 , n12484 );
not ( n22372 , n370011 );
buf ( n370013 , n22372 );
buf ( n370014 , n370013 );
not ( n22375 , n370014 );
or ( n22376 , n22370 , n22375 );
buf ( n370017 , n590 );
not ( n22378 , n370017 );
buf ( n370019 , n12484 );
nand ( n22380 , n22378 , n370019 );
buf ( n370021 , n22380 );
buf ( n370022 , n370021 );
nand ( n22383 , n22376 , n370022 );
buf ( n370024 , n22383 );
buf ( n370025 , n370024 );
nand ( n22386 , n370008 , n370025 );
buf ( n370027 , n22386 );
buf ( n370028 , n370027 );
nand ( n22389 , n22367 , n370028 );
buf ( n370030 , n22389 );
buf ( n370031 , C1 );
buf ( n370032 , n370030 );
buf ( n370033 , n369989 );
nor ( n22396 , n370032 , n370033 );
buf ( n370035 , n22396 );
not ( n22398 , n370035 );
buf ( n370037 , n370024 );
buf ( n370038 , n591 );
and ( n22401 , n370037 , n370038 );
buf ( n370040 , n365732 );
not ( n22403 , n370040 );
buf ( n370042 , n19166 );
not ( n22405 , n370042 );
buf ( n370044 , n369366 );
not ( n22407 , n370044 );
and ( n22408 , n22405 , n22407 );
nor ( n22412 , n22408 , C0 );
buf ( n370048 , n22412 );
buf ( n370049 , n370048 );
nor ( n22415 , n22403 , n370049 );
buf ( n370051 , n22415 );
buf ( n370052 , n370051 );
nor ( n22418 , n22401 , n370052 );
buf ( n370054 , n22418 );
buf ( n370055 , C1 );
buf ( n370056 , n370054 );
buf ( n370057 , n370055 );
nand ( n22434 , n370056 , n370057 );
buf ( n370059 , n22434 );
buf ( n370060 , n591 );
not ( n22437 , n370060 );
buf ( n370062 , n22437 );
or ( n22439 , n370048 , n370062 );
buf ( n370064 , C0 );
buf ( n370065 , n590 );
xnor ( n22442 , n370064 , n370065 );
buf ( n370067 , n22442 );
buf ( n370068 , n370067 );
not ( n22445 , n370068 );
buf ( n370070 , n365732 );
nand ( n22447 , n22445 , n370070 );
buf ( n370072 , n22447 );
nand ( n22449 , n22439 , n370072 );
not ( n22450 , n22449 );
buf ( n370075 , C0 );
buf ( n370076 , n370075 );
xor ( n22453 , n590 , C0 );
buf ( n370078 , n22453 );
buf ( n370079 , n591 );
and ( n22456 , n370078 , n370079 );
buf ( n370081 , n365729 );
not ( n22458 , n370081 );
buf ( n370083 , C0 );
nor ( n22460 , n22458 , n370083 );
buf ( n370085 , n22460 );
buf ( n370086 , n370085 );
nor ( n22463 , n22456 , n370086 );
buf ( n370088 , n22463 );
buf ( n370089 , n370088 );
nand ( n22466 , C1 , n590 );
buf ( n370091 , n22466 );
nor ( n22468 , n370089 , n370091 );
buf ( n370093 , n22468 );
buf ( n370094 , n370093 );
xor ( n22471 , n370076 , n370094 );
not ( n22472 , n22453 );
not ( n22473 , n365732 );
or ( n22474 , n22472 , n22473 );
or ( n22475 , n370067 , n370062 );
nand ( n22476 , n22474 , n22475 );
buf ( n370101 , n22476 );
and ( n22478 , n22471 , n370101 );
or ( n22479 , n22478 , C0 );
buf ( n370104 , n22479 );
not ( n22481 , n370104 );
nand ( n22493 , n22481 , C1 );
not ( n22494 , n22493 );
or ( n22495 , n22450 , n22494 );
nand ( n22497 , n22495 , C1 );
nand ( n22498 , n370059 , n22497 );
buf ( n370111 , n22498 );
nand ( n22500 , C1 , n370111 );
buf ( n370113 , n22500 );
nand ( n22502 , n22398 , n370113 );
nand ( n22503 , n370031 , n22502 );
not ( n22504 , n22503 );
buf ( n370117 , C0 );
buf ( n370118 , n370117 );
buf ( n370119 , n17867 );
not ( n22510 , n370119 );
buf ( n370121 , n588 );
buf ( n370122 , n12484 );
and ( n22513 , n370121 , n370122 );
not ( n22514 , n370121 );
buf ( n370125 , n367708 );
and ( n22516 , n22514 , n370125 );
nor ( n22517 , n22513 , n22516 );
buf ( n370128 , n22517 );
buf ( n370129 , n370128 );
not ( n22520 , n370129 );
or ( n22521 , n22510 , n22520 );
buf ( n370132 , n365646 );
buf ( n370133 , n369926 );
nand ( n22524 , n370132 , n370133 );
buf ( n370135 , n22524 );
buf ( n370136 , n370135 );
nand ( n22527 , n22521 , n370136 );
buf ( n370138 , n22527 );
buf ( n370139 , n370138 );
xor ( n22530 , n370118 , n370139 );
xor ( n22531 , n369918 , n369939 );
and ( n22532 , n22531 , n369988 );
or ( n22534 , n22532 , C0 );
buf ( n370144 , n22534 );
buf ( n370145 , n370144 );
xor ( n22537 , n22530 , n370145 );
buf ( n370147 , n22537 );
buf ( n370148 , n591 );
not ( n22540 , n370148 );
xor ( n22541 , n12482 , n590 );
buf ( n370151 , n22541 );
not ( n22543 , n370151 );
or ( n22544 , n22540 , n22543 );
buf ( n370154 , n365735 );
buf ( n370155 , n370004 );
nand ( n22547 , n370154 , n370155 );
buf ( n370157 , n22547 );
buf ( n370158 , n370157 );
nand ( n22550 , n22544 , n370158 );
buf ( n370160 , n22550 );
nor ( n22552 , n370147 , n370160 );
not ( n22553 , n22552 );
not ( n22554 , n22553 );
or ( n22555 , n22504 , n22554 );
nand ( n22556 , n370147 , n370160 );
nand ( n22557 , n22555 , n22556 );
buf ( n370167 , n22557 );
not ( n22559 , n370167 );
buf ( n370169 , n22559 );
buf ( n370170 , n370169 );
buf ( n370171 , n17867 );
not ( n22563 , n370171 );
buf ( n370173 , n22229 );
not ( n22565 , n370173 );
or ( n22566 , n22563 , n22565 );
buf ( n370176 , n370128 );
buf ( n370177 , n365646 );
nand ( n22569 , n370176 , n370177 );
buf ( n370179 , n22569 );
buf ( n370180 , n370179 );
nand ( n22572 , n22566 , n370180 );
buf ( n370182 , n22572 );
buf ( n370183 , n370182 );
buf ( n370184 , C0 );
buf ( n370185 , n370184 );
xor ( n22579 , n370183 , n370185 );
buf ( n370187 , n591 );
not ( n22581 , n370187 );
buf ( n370189 , n22251 );
not ( n22583 , n370189 );
or ( n22584 , n22581 , n22583 );
buf ( n370192 , n22541 );
buf ( n370193 , n365732 );
nand ( n22587 , n370192 , n370193 );
buf ( n370195 , n22587 );
buf ( n370196 , n370195 );
nand ( n22590 , n22584 , n370196 );
buf ( n370198 , n22590 );
buf ( n370199 , n370198 );
xor ( n22593 , n22579 , n370199 );
buf ( n370201 , n22593 );
buf ( n370202 , n370201 );
buf ( n22596 , n370202 );
buf ( n370204 , n22596 );
buf ( n370205 , n370204 );
xor ( n22599 , n370118 , n370139 );
and ( n22600 , n22599 , n370145 );
or ( n22602 , n22600 , C0 );
buf ( n370209 , n22602 );
buf ( n370210 , n370209 );
nor ( n22605 , n370205 , n370210 );
buf ( n370212 , n22605 );
buf ( n370213 , n370212 );
or ( n22608 , n370170 , n370213 );
buf ( n370215 , n370204 );
buf ( n370216 , n370209 );
nand ( n22611 , n370215 , n370216 );
buf ( n370218 , n22611 );
buf ( n370219 , n370218 );
nand ( n22614 , n22608 , n370219 );
buf ( n370221 , n22614 );
buf ( n370222 , n370221 );
not ( n22617 , n370222 );
xor ( n22618 , n369887 , n369891 );
xor ( n22619 , n22618 , n369909 );
buf ( n370226 , n22619 );
not ( n22621 , n370226 );
xor ( n22622 , n370183 , n370185 );
and ( n22623 , n22622 , n370199 );
or ( n22625 , n22623 , C0 );
buf ( n370231 , n22625 );
buf ( n370232 , n370231 );
not ( n22628 , n370232 );
buf ( n370234 , n22628 );
nand ( n22630 , n22621 , n370234 );
buf ( n370236 , n22630 );
not ( n22632 , n370236 );
or ( n22633 , n22617 , n22632 );
buf ( n370239 , n370226 );
buf ( n370240 , n370231 );
nand ( n22636 , n370239 , n370240 );
buf ( n370242 , n22636 );
buf ( n370243 , n370242 );
nand ( n22639 , n22633 , n370243 );
buf ( n370245 , n22639 );
buf ( n370246 , n370245 );
not ( n22642 , n370246 );
or ( n22643 , n22267 , n22642 );
buf ( n370249 , n369869 );
buf ( n370250 , n369913 );
nand ( n22646 , n370249 , n370250 );
buf ( n370252 , n22646 );
buf ( n370253 , n370252 );
nand ( n22649 , n22643 , n370253 );
buf ( n370255 , n22649 );
buf ( n370256 , n370255 );
not ( n22652 , n370256 );
xor ( n22653 , n369803 , n369805 );
and ( n22654 , n22653 , n369833 );
or ( n22656 , n22654 , C0 );
buf ( n370261 , n22656 );
buf ( n370262 , n370261 );
buf ( n370263 , n591 );
not ( n22660 , n370263 );
and ( n22661 , n590 , n365032 );
not ( n22662 , n590 );
and ( n22663 , n22662 , n12483 );
or ( n22664 , n22661 , n22663 );
buf ( n370269 , n22664 );
not ( n22666 , n370269 );
or ( n22667 , n22660 , n22666 );
buf ( n370272 , n22193 );
buf ( n370273 , n365735 );
nand ( n22670 , n370272 , n370273 );
buf ( n370275 , n22670 );
buf ( n370276 , n370275 );
nand ( n22673 , n22667 , n370276 );
buf ( n370278 , n22673 );
buf ( n370279 , n370278 );
xor ( n22676 , n370262 , n370279 );
buf ( n370281 , n365351 );
not ( n22678 , n370281 );
buf ( n370283 , n369425 );
not ( n22680 , n370283 );
or ( n22681 , n22678 , n22680 );
buf ( n370286 , n369792 );
buf ( n370287 , n365375 );
nand ( n22684 , n370286 , n370287 );
buf ( n370289 , n22684 );
buf ( n370290 , n370289 );
nand ( n22687 , n22681 , n370290 );
buf ( n370292 , n22687 );
buf ( n370293 , n370292 );
xor ( n22690 , n369477 , n369502 );
xor ( n22691 , n22690 , n369587 );
buf ( n370296 , n22691 );
buf ( n370297 , n370296 );
xor ( n22694 , n370293 , n370297 );
buf ( n370299 , n17867 );
not ( n22696 , n370299 );
buf ( n370301 , n21938 );
not ( n22698 , n370301 );
or ( n22699 , n22696 , n22698 );
buf ( n370304 , n22159 );
buf ( n370305 , n365646 );
nand ( n22702 , n370304 , n370305 );
buf ( n370307 , n22702 );
buf ( n370308 , n370307 );
nand ( n22705 , n22699 , n370308 );
buf ( n370310 , n22705 );
buf ( n370311 , n370310 );
xor ( n22708 , n22694 , n370311 );
buf ( n370313 , n22708 );
buf ( n370314 , n370313 );
xor ( n22711 , n22676 , n370314 );
buf ( n370316 , n22711 );
xor ( n22713 , n369778 , n369836 );
and ( n22714 , n22713 , n369867 );
and ( n22715 , n369778 , n369836 );
or ( n22716 , n22714 , n22715 );
buf ( n370321 , n22716 );
or ( n22718 , n370316 , n370321 );
buf ( n370323 , n22718 );
not ( n22720 , n370323 );
or ( n22721 , n22652 , n22720 );
buf ( n370326 , n370316 );
buf ( n370327 , n370321 );
nand ( n22724 , n370326 , n370327 );
buf ( n370329 , n22724 );
buf ( n370330 , n370329 );
nand ( n22727 , n22721 , n370330 );
buf ( n370332 , n22727 );
not ( n22729 , n370332 );
buf ( n370334 , n591 );
not ( n22731 , n370334 );
buf ( n370336 , n369641 );
not ( n22733 , n370336 );
or ( n22734 , n22731 , n22733 );
buf ( n370339 , n22664 );
buf ( n370340 , n365738 );
nand ( n22737 , n370339 , n370340 );
buf ( n370342 , n22737 );
buf ( n370343 , n370342 );
nand ( n22740 , n22734 , n370343 );
buf ( n370345 , n22740 );
buf ( n370346 , n370345 );
xor ( n22743 , n370293 , n370297 );
and ( n22744 , n22743 , n370311 );
and ( n22745 , n370293 , n370297 );
or ( n22746 , n22744 , n22745 );
buf ( n370351 , n22746 );
buf ( n370352 , n370351 );
xor ( n22749 , n370346 , n370352 );
xor ( n22750 , n369591 , n369595 );
xor ( n22751 , n22750 , n369613 );
buf ( n370356 , n22751 );
buf ( n370357 , n370356 );
xor ( n22754 , n22749 , n370357 );
buf ( n370359 , n22754 );
buf ( n370360 , n370359 );
xor ( n22757 , n370262 , n370279 );
and ( n22758 , n22757 , n370314 );
and ( n22759 , n370262 , n370279 );
or ( n22760 , n22758 , n22759 );
buf ( n370365 , n22760 );
buf ( n370366 , n370365 );
or ( n22763 , n370360 , n370366 );
buf ( n370368 , n22763 );
not ( n22765 , n370368 );
or ( n22766 , n22729 , n22765 );
buf ( n370371 , n370359 );
buf ( n370372 , n370365 );
nand ( n22769 , n370371 , n370372 );
buf ( n370374 , n22769 );
nand ( n22771 , n22766 , n370374 );
buf ( n370376 , n22771 );
not ( n22773 , n370376 );
xor ( n22774 , n369618 , n369622 );
xor ( n22775 , n22774 , n369649 );
buf ( n370380 , n22775 );
not ( n22777 , n370380 );
buf ( n370382 , n22777 );
xor ( n22779 , n370346 , n370352 );
and ( n22780 , n22779 , n370357 );
and ( n22781 , n370346 , n370352 );
or ( n22782 , n22780 , n22781 );
buf ( n370387 , n22782 );
buf ( n370388 , n370387 );
not ( n22785 , n370388 );
buf ( n370390 , n22785 );
buf ( n370391 , n370390 );
nand ( n22788 , n370382 , n370391 );
buf ( n370393 , n22788 );
buf ( n370394 , n370393 );
not ( n22791 , n370394 );
or ( n22792 , n22773 , n22791 );
buf ( n370397 , n370380 );
buf ( n370398 , n370387 );
nand ( n22795 , n370397 , n370398 );
buf ( n370400 , n22795 );
buf ( n370401 , n370400 );
nand ( n22798 , n22792 , n370401 );
buf ( n370403 , n22798 );
not ( n22800 , n370403 );
or ( n22801 , n21993 , n22800 );
buf ( n370406 , n369473 );
buf ( n22803 , n370406 );
buf ( n370408 , n22803 );
buf ( n370409 , n370408 );
buf ( n370410 , n369653 );
nand ( n22807 , n370409 , n370410 );
buf ( n370412 , n22807 );
nand ( n22809 , n22801 , n370412 );
buf ( n22810 , n22809 );
and ( n22811 , n21784 , n22810 );
buf ( n370416 , n369351 );
not ( n22813 , n370416 );
buf ( n370418 , n369466 );
not ( n22815 , n370418 );
buf ( n370420 , n22815 );
buf ( n370421 , n370420 );
nor ( n22818 , n22813 , n370421 );
buf ( n370423 , n22818 );
not ( n22820 , n370423 );
buf ( n370425 , n369346 );
not ( n22822 , n370425 );
buf ( n370427 , n22822 );
buf ( n370428 , n370427 );
buf ( n370429 , n369319 );
not ( n22826 , n370429 );
buf ( n370431 , n22826 );
buf ( n370432 , n370431 );
nand ( n22829 , n370428 , n370432 );
buf ( n370434 , n22829 );
not ( n22831 , n370434 );
or ( n22832 , n22820 , n22831 );
buf ( n370437 , n369346 );
buf ( n370438 , n369319 );
nand ( n22835 , n370437 , n370438 );
buf ( n370440 , n22835 );
nand ( n22837 , n22832 , n370440 );
nor ( n22838 , n22811 , n22837 );
buf ( n370443 , n22838 );
xor ( n22840 , n368890 , n369101 );
xor ( n22841 , n22840 , n369106 );
buf ( n370446 , n22841 );
buf ( n370447 , n370446 );
xor ( n22844 , n369326 , n369339 );
and ( n22845 , n22844 , n369344 );
and ( n22846 , n369326 , n369339 );
or ( n22847 , n22845 , n22846 );
buf ( n370452 , n22847 );
buf ( n370453 , n370452 );
nor ( n22850 , n370447 , n370453 );
buf ( n370455 , n22850 );
buf ( n370456 , n370455 );
nor ( n22853 , n370443 , n370456 );
buf ( n370458 , n22853 );
buf ( n370459 , n370458 );
not ( n22856 , n370459 );
or ( n22857 , n21429 , n22856 );
buf ( n370462 , n369116 );
buf ( n370463 , n370446 );
buf ( n370464 , n370452 );
nand ( n22861 , n370463 , n370464 );
buf ( n370466 , n22861 );
buf ( n370467 , n370466 );
not ( n22864 , n370467 );
buf ( n370469 , n22864 );
buf ( n370470 , n370469 );
and ( n22867 , n370462 , n370470 );
buf ( n370472 , n368871 );
buf ( n370473 , n369110 );
nand ( n22870 , n370472 , n370473 );
buf ( n370475 , n22870 );
buf ( n370476 , n370475 );
not ( n22873 , n370476 );
buf ( n370478 , n22873 );
buf ( n370479 , n370478 );
nor ( n22876 , n22867 , n370479 );
buf ( n370481 , n22876 );
buf ( n370482 , n370481 );
nand ( n22879 , n22857 , n370482 );
buf ( n370484 , n22879 );
nand ( n22881 , n368497 , n21152 , n370484 );
buf ( n370486 , n368299 );
not ( n22883 , n370486 );
buf ( n370488 , n368494 );
nand ( n22885 , n22883 , n370488 );
buf ( n370490 , n22885 );
or ( n22887 , n368858 , n368864 );
buf ( n370492 , n368858 );
buf ( n370493 , n368864 );
nand ( n22890 , n370492 , n370493 );
buf ( n370495 , n22890 );
buf ( n370496 , n370495 );
buf ( n370497 , n368722 );
buf ( n370498 , n368853 );
nand ( n22895 , n370497 , n370498 );
buf ( n370500 , n22895 );
buf ( n370501 , n370500 );
nand ( n22898 , n370496 , n370501 );
buf ( n370503 , n22898 );
nand ( n22900 , n370490 , n22887 , n370503 );
buf ( n370505 , n368299 );
buf ( n22902 , n370505 );
buf ( n370507 , n22902 );
nand ( n22904 , n370507 , n368491 );
nand ( n22905 , n22881 , n22900 , n22904 );
not ( n22906 , n22905 );
or ( n22907 , n20565 , n22906 );
buf ( n370512 , n367862 );
not ( n22909 , n370512 );
buf ( n370514 , n22909 );
buf ( n370515 , n370514 );
buf ( n370516 , n368125 );
not ( n22913 , n370516 );
buf ( n370518 , n22913 );
buf ( n370519 , n370518 );
nand ( n22916 , n370515 , n370519 );
buf ( n370521 , n22916 );
buf ( n370522 , n370521 );
buf ( n370523 , n368132 );
not ( n22920 , n370523 );
buf ( n370525 , n368291 );
not ( n22922 , n370525 );
buf ( n370527 , n22922 );
buf ( n370528 , n370527 );
nor ( n22925 , n22920 , n370528 );
buf ( n370530 , n22925 );
buf ( n370531 , n370530 );
and ( n22928 , n370522 , n370531 );
buf ( n370533 , n367862 );
buf ( n370534 , n368125 );
and ( n22931 , n370533 , n370534 );
buf ( n370536 , n22931 );
buf ( n370537 , n370536 );
nor ( n22934 , n22928 , n370537 );
buf ( n370539 , n22934 );
nand ( n22936 , n22907 , n370539 );
not ( n22937 , n22936 );
or ( n22938 , n20113 , n22937 );
buf ( n370543 , n367611 );
buf ( n370544 , n367852 );
nand ( n22941 , n370543 , n370544 );
buf ( n370546 , n22941 );
buf ( n22943 , n370546 );
nand ( n22944 , n22938 , n22943 );
not ( n22945 , n22944 );
or ( n22946 , n19859 , n22945 );
not ( n22947 , n367600 );
not ( n22948 , n367605 );
and ( n22949 , n22947 , n22948 );
nor ( n22950 , n366869 , n367107 );
nor ( n22951 , n22949 , n22950 );
nand ( n22952 , n367596 , n367197 );
not ( n22953 , n22952 );
and ( n22954 , n22951 , n22953 );
nand ( n22955 , n367600 , n367605 );
or ( n22956 , n19331 , n22955 );
nand ( n22957 , n366869 , n367107 );
nand ( n22958 , n22956 , n22957 );
nor ( n22959 , n22954 , n22958 );
nand ( n22960 , n22946 , n22959 );
buf ( n370565 , n22960 );
not ( n22962 , n370565 );
or ( n22963 , n19089 , n22962 );
not ( n22964 , n366320 );
not ( n22965 , n366617 );
or ( n22966 , n22964 , n22965 );
nor ( n22967 , n366617 , n366320 );
nand ( n22968 , n366860 , n366621 );
or ( n22969 , n22967 , n22968 );
nand ( n22970 , n22966 , n22969 );
buf ( n370575 , n22970 );
not ( n22972 , n370575 );
buf ( n370577 , n22972 );
buf ( n370578 , n370577 );
nand ( n22975 , n22963 , n370578 );
buf ( n370580 , n22975 );
not ( n22977 , n370580 );
not ( n22978 , n22977 );
or ( n22979 , n366317 , n22978 );
nand ( n22980 , n370580 , n18538 );
nand ( n22981 , n22979 , n22980 );
buf ( n22982 , n22981 );
buf ( n370587 , n22982 );
xor ( n22984 , n364708 , n364709 );
xor ( n22985 , n22984 , n370587 );
buf ( n370590 , n22985 );
xor ( n22987 , n364708 , n364709 );
and ( n22988 , n22987 , n370587 );
and ( n22989 , n364708 , n364709 );
or ( n22990 , n22988 , n22989 );
buf ( n370595 , n22990 );
buf ( n370596 , n364127 );
buf ( n370597 , n364097 );
buf ( n370598 , n17230 );
not ( n22995 , n370598 );
xor ( n22996 , n580 , n14498 );
buf ( n370601 , n22996 );
not ( n22998 , n370601 );
or ( n22999 , n22995 , n22998 );
not ( n23000 , n580 );
not ( n23001 , n364790 );
or ( n23002 , n23000 , n23001 );
nand ( n23003 , n365403 , n364896 );
nand ( n23004 , n23002 , n23003 );
buf ( n370609 , n23004 );
buf ( n370610 , n17209 );
nand ( n23007 , n370609 , n370610 );
buf ( n370612 , n23007 );
buf ( n370613 , n370612 );
nand ( n23010 , n22999 , n370613 );
buf ( n370615 , n23010 );
buf ( n370616 , n370615 );
buf ( n370617 , n17519 );
not ( n23014 , n370617 );
buf ( n370619 , n364779 );
not ( n23016 , n370619 );
buf ( n370621 , n23016 );
buf ( n370622 , n370621 );
buf ( n370623 , n364797 );
nor ( n23020 , n370622 , n370623 );
buf ( n370625 , n23020 );
buf ( n370626 , n370625 );
nand ( n23023 , n23014 , n370626 );
buf ( n370628 , n23023 );
not ( n23025 , n17519 );
buf ( n370630 , n23025 );
not ( n23027 , n370630 );
buf ( n370632 , n365151 );
not ( n23029 , n370632 );
buf ( n370634 , n582 );
nor ( n23031 , n23029 , n370634 );
buf ( n370636 , n23031 );
buf ( n370637 , n370636 );
nand ( n23034 , n23027 , n370637 );
buf ( n370639 , n23034 );
buf ( n370640 , n582 );
not ( n23037 , n370640 );
buf ( n370642 , n365362 );
not ( n23039 , n370642 );
or ( n23040 , n23037 , n23039 );
buf ( n370645 , n364797 );
buf ( n370646 , n17251 );
nand ( n23043 , n370645 , n370646 );
buf ( n370648 , n23043 );
buf ( n370649 , n370648 );
nand ( n23046 , n23040 , n370649 );
buf ( n370651 , n23046 );
buf ( n370652 , n370651 );
buf ( n370653 , n17133 );
nand ( n23050 , n370652 , n370653 );
buf ( n370655 , n23050 );
nand ( n23052 , n370628 , n370639 , n370655 );
buf ( n370657 , n23052 );
xor ( n23054 , n370616 , n370657 );
and ( n23055 , n364845 , n364852 );
buf ( n370660 , n23055 );
buf ( n370661 , n370660 );
buf ( n370662 , n17082 );
not ( n23059 , n370662 );
buf ( n370664 , n364733 );
not ( n23061 , n370664 );
or ( n23062 , n23059 , n23061 );
and ( n23063 , n9625 , n364727 );
not ( n23064 , n9625 );
and ( n23065 , n23064 , n578 );
or ( n23066 , n23063 , n23065 );
buf ( n370671 , n23066 );
buf ( n370672 , n17037 );
nand ( n23069 , n370671 , n370672 );
buf ( n370674 , n23069 );
buf ( n370675 , n370674 );
nand ( n23072 , n23062 , n370675 );
buf ( n370677 , n23072 );
buf ( n370678 , n370677 );
xor ( n23075 , n370661 , n370678 );
buf ( n370680 , n364834 );
not ( n23077 , n370680 );
buf ( n370682 , n576 );
buf ( n370683 , n8303 );
xor ( n23080 , n370682 , n370683 );
buf ( n370685 , n23080 );
buf ( n370686 , n370685 );
not ( n23083 , n370686 );
or ( n23084 , n23077 , n23083 );
buf ( n370689 , n364841 );
buf ( n370690 , n17182 );
nand ( n23087 , n370689 , n370690 );
buf ( n370692 , n23087 );
buf ( n370693 , n370692 );
nand ( n23090 , n23084 , n370693 );
buf ( n370695 , n23090 );
buf ( n370696 , n370695 );
and ( n23093 , n23075 , n370696 );
and ( n23094 , n370661 , n370678 );
or ( n23095 , n23093 , n23094 );
buf ( n370700 , n23095 );
buf ( n370701 , n370700 );
xor ( n23098 , n23054 , n370701 );
buf ( n370703 , n23098 );
buf ( n370704 , n370703 );
xor ( n23101 , n370661 , n370678 );
xor ( n23102 , n23101 , n370696 );
buf ( n370707 , n23102 );
buf ( n370708 , n370707 );
buf ( n370709 , n364925 );
not ( n23106 , n370709 );
buf ( n370711 , n364771 );
not ( n23108 , n16900 );
buf ( n370713 , n23108 );
and ( n23110 , n370711 , n370713 );
not ( n23111 , n370711 );
buf ( n370716 , n16900 );
and ( n23113 , n23111 , n370716 );
nor ( n23114 , n23110 , n23113 );
buf ( n370719 , n23114 );
buf ( n370720 , n370719 );
not ( n23117 , n370720 );
or ( n23118 , n23106 , n23117 );
buf ( n370723 , n365230 );
buf ( n370724 , n364973 );
nand ( n23121 , n370723 , n370724 );
buf ( n370726 , n23121 );
buf ( n370727 , n370726 );
nand ( n23124 , n23118 , n370727 );
buf ( n370729 , n23124 );
buf ( n370730 , n370729 );
xor ( n23127 , n370708 , n370730 );
buf ( n370732 , n365351 );
not ( n23129 , n370732 );
buf ( n370734 , n365712 );
buf ( n370735 , n586 );
and ( n23132 , n370734 , n370735 );
not ( n23133 , n370734 );
buf ( n370738 , n365334 );
and ( n23135 , n23133 , n370738 );
or ( n23136 , n23132 , n23135 );
buf ( n370741 , n23136 );
buf ( n370742 , n370741 );
not ( n23139 , n370742 );
or ( n23140 , n23129 , n23139 );
buf ( n370745 , n365375 );
buf ( n370746 , n365867 );
nand ( n23143 , n370745 , n370746 );
buf ( n370748 , n23143 );
buf ( n370749 , n370748 );
nand ( n23146 , n23140 , n370749 );
buf ( n370751 , n23146 );
buf ( n370752 , n370751 );
and ( n23149 , n23127 , n370752 );
and ( n23150 , n370708 , n370730 );
or ( n23151 , n23149 , n23150 );
buf ( n370756 , n23151 );
buf ( n370757 , n370756 );
xor ( n23154 , n370704 , n370757 );
and ( n23155 , n364837 , n364839 );
buf ( n370760 , n23155 );
buf ( n370761 , n370760 );
buf ( n370762 , n17082 );
not ( n23159 , n370762 );
buf ( n370764 , n23066 );
not ( n23161 , n370764 );
or ( n23162 , n23159 , n23161 );
nand ( n23163 , n364903 , n578 );
not ( n23164 , n23163 );
buf ( n370769 , n360086 );
buf ( n370770 , n364727 );
nand ( n23167 , n370769 , n370770 );
buf ( n370772 , n23167 );
not ( n23169 , n370772 );
or ( n23170 , n23164 , n23169 );
nand ( n23171 , n23170 , n17037 );
buf ( n370776 , n23171 );
nand ( n23173 , n23162 , n370776 );
buf ( n370778 , n23173 );
buf ( n370779 , n370778 );
xor ( n23176 , n370761 , n370779 );
not ( n23177 , n364834 );
not ( n23178 , n576 );
not ( n23179 , n365388 );
or ( n23180 , n23178 , n23179 );
buf ( n370785 , n8990 );
buf ( n370786 , n354303 );
nand ( n23183 , n370785 , n370786 );
buf ( n370788 , n23183 );
nand ( n23185 , n23180 , n370788 );
not ( n23186 , n23185 );
or ( n23187 , n23177 , n23186 );
buf ( n370792 , n370685 );
buf ( n370793 , n17182 );
nand ( n23190 , n370792 , n370793 );
buf ( n370795 , n23190 );
nand ( n23192 , n23187 , n370795 );
buf ( n370797 , n23192 );
xor ( n23194 , n23176 , n370797 );
buf ( n370799 , n23194 );
buf ( n370800 , n370799 );
buf ( n370801 , n365748 );
not ( n23198 , n370801 );
buf ( n370803 , n369550 );
buf ( n370804 , n584 );
nor ( n23201 , n370803 , n370804 );
buf ( n370806 , n23201 );
buf ( n370807 , n370806 );
nand ( n23204 , n23198 , n370807 );
buf ( n370809 , n23204 );
buf ( n370810 , n370809 );
buf ( n370811 , n365661 );
not ( n23208 , n370811 );
buf ( n370813 , n17687 );
not ( n23210 , n370813 );
and ( n23211 , n23208 , n23210 );
buf ( n370816 , n16955 );
not ( n23213 , n370816 );
buf ( n370818 , n23213 );
buf ( n370819 , n370818 );
not ( n23216 , n370819 );
buf ( n370821 , n23216 );
buf ( n370822 , n370821 );
buf ( n370823 , n365430 );
and ( n23220 , n370822 , n370823 );
nor ( n23221 , n23211 , n23220 );
buf ( n370826 , n23221 );
buf ( n370827 , n370826 );
nand ( n23224 , n23108 , n369554 );
buf ( n370829 , n23224 );
nand ( n23226 , n370810 , n370827 , n370829 );
buf ( n370831 , n23226 );
buf ( n370832 , n370831 );
xor ( n23229 , n370800 , n370832 );
not ( n23230 , n370741 );
not ( n23231 , n365375 );
or ( n23232 , n23230 , n23231 );
not ( n23233 , n365350 );
buf ( n370838 , n586 );
not ( n23235 , n370838 );
not ( n23236 , n17933 );
buf ( n370841 , n23236 );
not ( n23238 , n370841 );
or ( n23239 , n23235 , n23238 );
buf ( n370844 , n365881 );
buf ( n370845 , n365334 );
nand ( n23242 , n370844 , n370845 );
buf ( n370847 , n23242 );
buf ( n370848 , n370847 );
nand ( n23245 , n23239 , n370848 );
buf ( n370850 , n23245 );
nand ( n23247 , n23233 , n370850 );
nand ( n23248 , n23232 , n23247 );
buf ( n370853 , n23248 );
xor ( n23250 , n23229 , n370853 );
buf ( n370855 , n23250 );
buf ( n370856 , n370855 );
xor ( n23253 , n23154 , n370856 );
buf ( n370858 , n23253 );
buf ( n370859 , n370858 );
xor ( n23256 , n365875 , n365888 );
and ( n23257 , n23256 , n365909 );
and ( n23258 , n365875 , n365888 );
or ( n23259 , n23257 , n23258 );
buf ( n370864 , n23259 );
buf ( n370865 , n370864 );
not ( n23262 , n365646 );
not ( n23263 , n365883 );
or ( n23264 , n23262 , n23263 );
and ( n23265 , n365897 , n368320 );
not ( n23266 , n365897 );
and ( n23267 , n23266 , n368310 );
nor ( n23268 , n23265 , n23267 );
nand ( n23269 , n23264 , n23268 );
buf ( n370874 , n23269 );
xor ( n23271 , n364765 , n364817 );
and ( n23272 , n23271 , n364918 );
and ( n23273 , n364765 , n364817 );
or ( n23274 , n23272 , n23273 );
buf ( n370879 , n23274 );
buf ( n370880 , n370879 );
xor ( n23277 , n370874 , n370880 );
not ( n23278 , n17230 );
not ( n23279 , n23004 );
or ( n23280 , n23278 , n23279 );
not ( n23281 , n364909 );
not ( n23282 , n364904 );
or ( n23283 , n23281 , n23282 );
nand ( n23284 , n23283 , n17209 );
nand ( n23285 , n23280 , n23284 );
buf ( n370890 , n23285 );
buf ( n370891 , n17133 );
not ( n23288 , n370891 );
buf ( n370893 , n17106 );
not ( n23290 , n370893 );
or ( n23291 , n23288 , n23290 );
buf ( n370896 , n370651 );
buf ( n370897 , n365151 );
nand ( n23294 , n370896 , n370897 );
buf ( n370899 , n23294 );
buf ( n370900 , n370899 );
nand ( n23297 , n23291 , n370900 );
buf ( n370902 , n23297 );
buf ( n370903 , n370902 );
xor ( n23300 , n370890 , n370903 );
xor ( n23301 , n364830 , n364866 );
and ( n23302 , n23301 , n364915 );
and ( n23303 , n364830 , n364866 );
or ( n23304 , n23302 , n23303 );
buf ( n370909 , n23304 );
buf ( n370910 , n370909 );
xor ( n23307 , n23300 , n370910 );
buf ( n370912 , n23307 );
buf ( n370913 , n370912 );
xor ( n23310 , n23277 , n370913 );
buf ( n370915 , n23310 );
buf ( n370916 , n370915 );
xor ( n23313 , n370865 , n370916 );
xor ( n23314 , n364921 , n365201 );
and ( n23315 , n23314 , n365327 );
and ( n23316 , n364921 , n365201 );
or ( n23317 , n23315 , n23316 );
buf ( n370922 , n23317 );
buf ( n370923 , n370922 );
and ( n23320 , n23313 , n370923 );
and ( n23321 , n370865 , n370916 );
or ( n23322 , n23320 , n23321 );
buf ( n370927 , n23322 );
buf ( n370928 , n370927 );
xor ( n23325 , n370859 , n370928 );
xor ( n23326 , n370874 , n370880 );
and ( n23327 , n23326 , n370913 );
and ( n23328 , n370874 , n370880 );
or ( n23329 , n23327 , n23328 );
buf ( n370934 , n23329 );
buf ( n370935 , n370934 );
buf ( n370936 , n365646 );
not ( n23333 , n370936 );
buf ( n370938 , n588 );
buf ( n370939 , n365897 );
and ( n23336 , n370938 , n370939 );
not ( n23337 , n370938 );
buf ( n370942 , n365897 );
not ( n23339 , n370942 );
buf ( n370944 , n23339 );
buf ( n370945 , n370944 );
and ( n23342 , n23337 , n370945 );
nor ( n23343 , n23336 , n23342 );
buf ( n370948 , n23343 );
buf ( n370949 , n370948 );
not ( n23346 , n370949 );
or ( n23347 , n23333 , n23346 );
buf ( n370952 , n588 );
not ( n23349 , n370952 );
buf ( n370954 , n365892 );
not ( n23351 , n370954 );
buf ( n370956 , n23351 );
buf ( n370957 , n370956 );
not ( n23354 , n370957 );
or ( n23355 , n23349 , n23354 );
buf ( n370960 , n588 );
not ( n23357 , n370960 );
buf ( n370962 , n365892 );
nand ( n23359 , n23357 , n370962 );
buf ( n370964 , n23359 );
buf ( n370965 , n370964 );
nand ( n23362 , n23355 , n370965 );
buf ( n370967 , n23362 );
buf ( n370968 , n370967 );
buf ( n370969 , n17867 );
nand ( n23366 , n370968 , n370969 );
buf ( n370971 , n23366 );
buf ( n370972 , n370971 );
nand ( n23369 , n23347 , n370972 );
buf ( n370974 , n23369 );
buf ( n370975 , n370974 );
xor ( n23372 , n370890 , n370903 );
and ( n23373 , n23372 , n370910 );
and ( n23374 , n370890 , n370903 );
or ( n23375 , n23373 , n23374 );
buf ( n370980 , n23375 );
buf ( n370981 , n370980 );
xor ( n23378 , n370975 , n370981 );
buf ( n370983 , n590 );
not ( n23380 , n370983 );
buf ( n23381 , n16613 );
nand ( n23382 , n16793 , n16792 );
not ( n23383 , n23382 );
and ( n23384 , n23381 , n23383 );
not ( n23385 , n23381 );
and ( n23386 , n23385 , n23382 );
nor ( n23387 , n23384 , n23386 );
not ( n23388 , n23387 );
buf ( n370993 , n23388 );
not ( n23390 , n370993 );
or ( n23391 , n23380 , n23390 );
not ( n23392 , n590 );
nand ( n23393 , n23392 , n23387 );
buf ( n370998 , n23393 );
nand ( n23395 , n23391 , n370998 );
buf ( n371000 , n23395 );
not ( n23397 , n371000 );
not ( n23398 , n591 );
or ( n23399 , n23397 , n23398 );
buf ( n371004 , n16815 );
not ( n23401 , n371004 );
buf ( n371006 , n23401 );
and ( n23403 , n590 , n371006 );
not ( n23404 , n590 );
and ( n23405 , n23404 , n16815 );
or ( n23406 , n23403 , n23405 );
buf ( n371011 , n23406 );
buf ( n371012 , n365738 );
nand ( n23409 , n371011 , n371012 );
buf ( n371014 , n23409 );
nand ( n23411 , n23399 , n371014 );
buf ( n371016 , n23411 );
xor ( n23413 , n23378 , n371016 );
buf ( n371018 , n23413 );
buf ( n371019 , n371018 );
xor ( n23416 , n370935 , n371019 );
buf ( n371021 , n591 );
not ( n23418 , n371021 );
buf ( n371023 , n23406 );
not ( n23420 , n371023 );
or ( n23421 , n23418 , n23420 );
buf ( n371026 , n365893 );
buf ( n371027 , n365738 );
nand ( n23424 , n371026 , n371027 );
buf ( n371029 , n23424 );
buf ( n371030 , n371029 );
nand ( n23427 , n23421 , n371030 );
buf ( n371032 , n23427 );
buf ( n371033 , n371032 );
xor ( n23430 , n365208 , n365241 );
and ( n23431 , n23430 , n365324 );
and ( n23432 , n365208 , n365241 );
or ( n23433 , n23431 , n23432 );
buf ( n371038 , n23433 );
buf ( n371039 , n371038 );
xor ( n23436 , n371033 , n371039 );
xor ( n23437 , n370708 , n370730 );
xor ( n23438 , n23437 , n370752 );
buf ( n371043 , n23438 );
buf ( n371044 , n371043 );
and ( n23441 , n23436 , n371044 );
and ( n23442 , n371033 , n371039 );
or ( n23443 , n23441 , n23442 );
buf ( n371048 , n23443 );
buf ( n371049 , n371048 );
xor ( n23446 , n23416 , n371049 );
buf ( n371051 , n23446 );
buf ( n371052 , n371051 );
xor ( n23449 , n23325 , n371052 );
buf ( n371054 , n23449 );
buf ( n371055 , n371054 );
xor ( n23452 , n371033 , n371039 );
xor ( n23453 , n23452 , n371044 );
buf ( n371058 , n23453 );
buf ( n371059 , n371058 );
xor ( n23456 , n365846 , n365912 );
and ( n23457 , n23456 , n365938 );
and ( n23458 , n365846 , n365912 );
or ( n23459 , n23457 , n23458 );
buf ( n371064 , n23459 );
buf ( n371065 , n371064 );
xor ( n23462 , n371059 , n371065 );
xor ( n23463 , n370865 , n370916 );
xor ( n23464 , n23463 , n370923 );
buf ( n371069 , n23464 );
buf ( n371070 , n371069 );
and ( n23467 , n23462 , n371070 );
and ( n23468 , n371059 , n371065 );
or ( n23469 , n23467 , n23468 );
buf ( n371074 , n23469 );
buf ( n371075 , n371074 );
or ( n23472 , n371055 , n371075 );
buf ( n371077 , n23472 );
buf ( n371078 , n371054 );
buf ( n371079 , n371074 );
nand ( n23476 , n371078 , n371079 );
buf ( n371081 , n23476 );
and ( n23478 , n371077 , n371081 );
buf ( n371083 , n22960 );
not ( n23480 , n371083 );
xor ( n23481 , n371059 , n371065 );
xor ( n23482 , n23481 , n371070 );
buf ( n371087 , n23482 );
not ( n23484 , n371087 );
xor ( n23485 , n365330 , n365839 );
and ( n23486 , n23485 , n365941 );
and ( n23487 , n365330 , n365839 );
or ( n23488 , n23486 , n23487 );
buf ( n371093 , n23488 );
not ( n23490 , n371093 );
and ( n23491 , n23484 , n23490 );
buf ( n371096 , n365943 );
buf ( n371097 , n366308 );
nor ( n23494 , n371096 , n371097 );
buf ( n371099 , n23494 );
nor ( n23496 , n23491 , n371099 );
and ( n23497 , n19087 , n23496 );
buf ( n371102 , n23497 );
not ( n23499 , n371102 );
or ( n23500 , n23480 , n23499 );
not ( n23501 , n22970 );
not ( n23502 , n23496 );
or ( n23503 , n23501 , n23502 );
buf ( n371108 , n371093 );
buf ( n371109 , n371087 );
nor ( n23506 , n371108 , n371109 );
buf ( n371111 , n23506 );
buf ( n371112 , n365943 );
buf ( n371113 , n366308 );
nand ( n23510 , n371112 , n371113 );
buf ( n371115 , n23510 );
nor ( n23512 , n371111 , n371115 );
buf ( n371117 , n371087 );
buf ( n371118 , n371093 );
and ( n23515 , n371117 , n371118 );
buf ( n371120 , n23515 );
nor ( n23517 , n23512 , n371120 );
nand ( n23518 , n23503 , n23517 );
buf ( n371123 , n23518 );
not ( n23520 , n371123 );
buf ( n371125 , n23520 );
buf ( n371126 , n371125 );
nand ( n23523 , n23500 , n371126 );
buf ( n371128 , n23523 );
buf ( n371129 , n371128 );
buf ( n23526 , n371129 );
buf ( n371131 , n23526 );
xor ( n23528 , n23478 , n371131 );
buf ( n371133 , n23528 );
xor ( n23530 , n370596 , n370597 );
xor ( n23531 , n23530 , n371133 );
buf ( n371136 , n23531 );
xor ( n23533 , n370596 , n370597 );
and ( n23534 , n23533 , n371133 );
and ( n23535 , n370596 , n370597 );
or ( n23536 , n23534 , n23535 );
buf ( n371141 , n23536 );
buf ( n371142 , n347471 );
buf ( n371143 , n347729 );
not ( n23540 , n370113 );
not ( n23541 , n23540 );
buf ( n371146 , n370035 );
not ( n23543 , n371146 );
buf ( n371148 , n370031 );
nand ( n23545 , n23543 , n371148 );
buf ( n371150 , n23545 );
not ( n23547 , n371150 );
not ( n23548 , n23547 );
or ( n23549 , n23541 , n23548 );
nand ( n23550 , n370113 , n371150 );
nand ( n23551 , n23549 , n23550 );
buf ( n371156 , n23551 );
xor ( n23553 , n371142 , n371143 );
xor ( n23554 , n23553 , n371156 );
buf ( n371159 , n23554 );
xor ( n23556 , n371142 , n371143 );
and ( n23557 , n23556 , n371156 );
and ( n23558 , n371142 , n371143 );
or ( n23559 , n23557 , n23558 );
buf ( n371164 , n23559 );
buf ( n371165 , n347637 );
buf ( n371166 , n12496 );
buf ( n371167 , n22552 );
not ( n23564 , n371167 );
buf ( n371169 , n22556 );
nand ( n23566 , n23564 , n371169 );
buf ( n371171 , n23566 );
buf ( n371172 , n371171 );
not ( n23569 , n22503 );
buf ( n371174 , n23569 );
and ( n23571 , n371172 , n371174 );
not ( n23572 , n371172 );
buf ( n371177 , n23569 );
not ( n23574 , n371177 );
buf ( n371179 , n23574 );
buf ( n371180 , n371179 );
and ( n23577 , n23572 , n371180 );
nor ( n23578 , n23571 , n23577 );
buf ( n371183 , n23578 );
buf ( n371184 , n371183 );
xor ( n23581 , n371165 , n371166 );
xor ( n23582 , n23581 , n371184 );
buf ( n371187 , n23582 );
xor ( n23584 , n371165 , n371166 );
and ( n23585 , n23584 , n371184 );
and ( n23586 , n371165 , n371166 );
or ( n23587 , n23585 , n23586 );
buf ( n371192 , n23587 );
buf ( n371193 , n348551 );
buf ( n371194 , n12495 );
not ( n23591 , n22557 );
and ( n23592 , n370201 , n370209 );
not ( n23593 , n370201 );
buf ( n371198 , n370209 );
not ( n23595 , n371198 );
buf ( n371200 , n23595 );
and ( n23597 , n23593 , n371200 );
or ( n23598 , n23592 , n23597 );
not ( n23599 , n23598 );
not ( n23600 , n23599 );
or ( n23601 , n23591 , n23600 );
nand ( n23602 , n370169 , n23598 );
nand ( n23603 , n23601 , n23602 );
not ( n23604 , n23603 );
buf ( n371209 , n23604 );
xor ( n23606 , n371193 , n371194 );
xor ( n23607 , n23606 , n371209 );
buf ( n371212 , n23607 );
xor ( n23609 , n371193 , n371194 );
and ( n23610 , n23609 , n371209 );
and ( n23611 , n371193 , n371194 );
or ( n23612 , n23610 , n23611 );
buf ( n371217 , n23612 );
buf ( n371218 , n350028 );
buf ( n371219 , n12494 );
buf ( n371220 , n370221 );
not ( n23617 , n371220 );
buf ( n371222 , n370226 );
not ( n23619 , n371222 );
buf ( n371224 , n370234 );
nand ( n23621 , n23619 , n371224 );
buf ( n371226 , n23621 );
buf ( n371227 , n371226 );
buf ( n371228 , n370242 );
nand ( n23625 , n371227 , n371228 );
buf ( n371230 , n23625 );
buf ( n371231 , n371230 );
not ( n23628 , n371231 );
or ( n23629 , n23617 , n23628 );
buf ( n371234 , n370221 );
not ( n23631 , n371234 );
buf ( n371236 , n371230 );
not ( n23633 , n371236 );
buf ( n371238 , n23633 );
buf ( n371239 , n371238 );
nand ( n23636 , n23631 , n371239 );
buf ( n371241 , n23636 );
buf ( n371242 , n371241 );
nand ( n23639 , n23629 , n371242 );
buf ( n371244 , n23639 );
buf ( n371245 , n371244 );
xor ( n23642 , n371218 , n371219 );
xor ( n23643 , n23642 , n371245 );
buf ( n371248 , n23643 );
xor ( n23645 , n371218 , n371219 );
and ( n23646 , n23645 , n371245 );
and ( n23647 , n371218 , n371219 );
or ( n23648 , n23646 , n23647 );
buf ( n371253 , n23648 );
buf ( n23650 , n350645 );
buf ( n371255 , n23650 );
buf ( n371256 , n350632 );
buf ( n371257 , n370255 );
not ( n23654 , n371257 );
buf ( n371259 , n22718 );
buf ( n371260 , n370329 );
nand ( n23657 , n371259 , n371260 );
buf ( n371262 , n23657 );
buf ( n371263 , n371262 );
not ( n23660 , n371263 );
or ( n23661 , n23654 , n23660 );
buf ( n371266 , n371262 );
not ( n23663 , n371266 );
buf ( n371268 , n23663 );
buf ( n371269 , n371268 );
buf ( n371270 , n370255 );
not ( n23667 , n371270 );
buf ( n371272 , n23667 );
buf ( n371273 , n371272 );
nand ( n23670 , n371269 , n371273 );
buf ( n371275 , n23670 );
buf ( n371276 , n371275 );
nand ( n23673 , n23661 , n371276 );
buf ( n371278 , n23673 );
buf ( n371279 , n371278 );
xor ( n23676 , n371255 , n371256 );
xor ( n23677 , n23676 , n371279 );
buf ( n371282 , n23677 );
xor ( n23679 , n371255 , n371256 );
and ( n23680 , n23679 , n371279 );
and ( n23681 , n371255 , n371256 );
or ( n23682 , n23680 , n23681 );
buf ( n371287 , n23682 );
buf ( n371288 , n12502 );
buf ( n371289 , n350958 );
not ( n23686 , n370332 );
buf ( n371291 , n370368 );
buf ( n371292 , n370374 );
nand ( n23689 , n371291 , n371292 );
buf ( n371294 , n23689 );
not ( n23691 , n371294 );
or ( n23692 , n23686 , n23691 );
buf ( n371297 , n370332 );
not ( n23694 , n371297 );
buf ( n371299 , n371294 );
not ( n23696 , n371299 );
buf ( n371301 , n23696 );
buf ( n371302 , n371301 );
nand ( n23699 , n23694 , n371302 );
buf ( n371304 , n23699 );
nand ( n23701 , n23692 , n371304 );
buf ( n371306 , n23701 );
xor ( n23703 , n371288 , n371289 );
xor ( n23704 , n23703 , n371306 );
buf ( n371309 , n23704 );
xor ( n23706 , n371288 , n371289 );
and ( n23707 , n23706 , n371306 );
and ( n23708 , n371288 , n371289 );
or ( n23709 , n23707 , n23708 );
buf ( n371314 , n23709 );
buf ( n371315 , n351500 );
buf ( n371316 , n351487 );
buf ( n371317 , n370380 );
buf ( n371318 , n370387 );
nand ( n23715 , n371317 , n371318 );
buf ( n371320 , n23715 );
nand ( n23717 , n370393 , n371320 );
buf ( n23718 , n22771 );
not ( n23719 , n23718 );
and ( n23720 , n23717 , n23719 );
not ( n23721 , n23717 );
and ( n23722 , n23721 , n23718 );
nor ( n23723 , n23720 , n23722 );
not ( n23724 , n23723 );
not ( n23725 , n23724 );
buf ( n371330 , n23725 );
xor ( n23727 , n371315 , n371316 );
xor ( n23728 , n23727 , n371330 );
buf ( n371333 , n23728 );
xor ( n23730 , n371315 , n371316 );
and ( n23731 , n23730 , n371330 );
and ( n23732 , n371315 , n371316 );
or ( n23733 , n23731 , n23732 );
buf ( n371338 , n23733 );
buf ( n371339 , n361565 );
buf ( n371340 , n13728 );
buf ( n371341 , n22936 );
buf ( n23738 , n371341 );
buf ( n371343 , n23738 );
buf ( n371344 , n371343 );
buf ( n371345 , n370546 );
buf ( n371346 , n367858 );
nand ( n23743 , n371345 , n371346 );
buf ( n371348 , n23743 );
not ( n23745 , n371348 );
buf ( n371350 , n23745 );
and ( n23747 , n371344 , n371350 );
not ( n23748 , n371344 );
buf ( n371353 , n371348 );
and ( n23750 , n23748 , n371353 );
nor ( n23751 , n23747 , n23750 );
buf ( n371356 , n23751 );
buf ( n371357 , n371356 );
xor ( n23754 , n371339 , n371340 );
xor ( n23755 , n23754 , n371357 );
buf ( n371360 , n23755 );
xor ( n23757 , n371339 , n371340 );
and ( n23758 , n23757 , n371357 );
and ( n23759 , n371339 , n371340 );
or ( n23760 , n23758 , n23759 );
buf ( n371365 , n23760 );
buf ( n371366 , n354602 );
buf ( n371367 , n12491 );
buf ( n371368 , n370446 );
buf ( n371369 , n370452 );
or ( n23766 , n371368 , n371369 );
buf ( n371371 , n23766 );
buf ( n371372 , n371371 );
buf ( n371373 , n370466 );
nand ( n23770 , n371372 , n371373 );
buf ( n371375 , n23770 );
buf ( n23772 , n22838 );
xor ( n23773 , n371375 , n23772 );
not ( n23774 , n23773 );
not ( n23775 , n23774 );
buf ( n371380 , n23775 );
xor ( n23777 , n371366 , n371367 );
xor ( n23778 , n23777 , n371380 );
buf ( n371383 , n23778 );
xor ( n23780 , n371366 , n371367 );
and ( n23781 , n23780 , n371380 );
and ( n23782 , n371366 , n371367 );
or ( n23783 , n23781 , n23782 );
buf ( n371388 , n23783 );
buf ( n371389 , n359724 );
buf ( n371390 , n359711 );
not ( n23787 , n370507 );
not ( n23788 , n368491 );
or ( n23789 , n23787 , n23788 );
buf ( n371394 , n368497 );
buf ( n23791 , n371394 );
buf ( n371396 , n23791 );
nand ( n23793 , n23789 , n371396 );
not ( n23794 , n22887 );
buf ( n371399 , n370484 );
buf ( n371400 , n368722 );
buf ( n371401 , n368853 );
or ( n23798 , n371400 , n371401 );
buf ( n371403 , n23798 );
buf ( n371404 , n371403 );
nand ( n23801 , n371399 , n371404 );
buf ( n371406 , n23801 );
buf ( n371407 , n371406 );
not ( n23804 , n371407 );
buf ( n371409 , n23804 );
not ( n23806 , n371409 );
or ( n23807 , n23794 , n23806 );
buf ( n371412 , n22887 );
buf ( n371413 , n370503 );
nand ( n23810 , n371412 , n371413 );
buf ( n371415 , n23810 );
nand ( n23812 , n23807 , n371415 );
xor ( n23813 , n23793 , n23812 );
buf ( n371418 , n23813 );
not ( n23815 , n371418 );
buf ( n371420 , n23815 );
buf ( n371421 , n371420 );
xor ( n23818 , n371389 , n371390 );
xor ( n23819 , n23818 , n371421 );
buf ( n371424 , n23819 );
xor ( n23821 , n371389 , n371390 );
and ( n23822 , n23821 , n371421 );
and ( n23823 , n371389 , n371390 );
or ( n23824 , n23822 , n23823 );
buf ( n371429 , n23824 );
buf ( n371430 , n360515 );
buf ( n371431 , n360502 );
buf ( n23828 , n22905 );
not ( n23829 , n368132 );
not ( n23830 , n23829 );
not ( n23831 , n370527 );
and ( n23832 , n23830 , n23831 );
and ( n23833 , n23829 , n370527 );
nor ( n23834 , n23832 , n23833 );
and ( n23835 , n23828 , n23834 );
not ( n23836 , n23828 );
not ( n23837 , n23834 );
and ( n23838 , n23836 , n23837 );
nor ( n23839 , n23835 , n23838 );
not ( n23840 , n23839 );
not ( n23841 , n23840 );
buf ( n371446 , n23841 );
xor ( n23843 , n371430 , n371431 );
xor ( n23844 , n23843 , n371446 );
buf ( n371449 , n23844 );
xor ( n23846 , n371430 , n371431 );
and ( n23847 , n23846 , n371446 );
and ( n23848 , n371430 , n371431 );
or ( n23849 , n23847 , n23848 );
buf ( n371454 , n23849 );
buf ( n371455 , n12500 );
buf ( n371456 , n12492 );
buf ( n371457 , n369351 );
not ( n23854 , n371457 );
buf ( n371459 , n23854 );
buf ( n371460 , n371459 );
buf ( n371461 , n370420 );
nand ( n23858 , n371460 , n371461 );
buf ( n371463 , n23858 );
buf ( n371464 , n371463 );
buf ( n371465 , n369351 );
buf ( n371466 , n369466 );
nand ( n23863 , n371465 , n371466 );
buf ( n371468 , n23863 );
buf ( n371469 , n371468 );
nand ( n23866 , n371464 , n371469 );
buf ( n371471 , n23866 );
xnor ( n23868 , n22809 , n371471 );
buf ( n371473 , n23868 );
xor ( n23870 , n371455 , n371456 );
xor ( n23871 , n23870 , n371473 );
buf ( n371476 , n23871 );
xor ( n23873 , n371455 , n371456 );
and ( n23874 , n23873 , n371473 );
and ( n23875 , n371455 , n371456 );
or ( n23876 , n23874 , n23875 );
buf ( n371481 , n23876 );
buf ( n371482 , n361039 );
buf ( n371483 , n361195 );
buf ( n371484 , n370536 );
buf ( n371485 , n368128 );
nor ( n23882 , n371484 , n371485 );
buf ( n371487 , n23882 );
buf ( n23884 , n371487 );
not ( n23885 , n23884 );
nor ( n23886 , n23829 , n370527 );
not ( n23887 , n23886 );
nor ( n23888 , n368132 , n368291 );
not ( n23889 , n23888 );
nand ( n23890 , n23889 , n23828 );
nand ( n23891 , n23887 , n23890 );
buf ( n371496 , n23891 );
not ( n23893 , n371496 );
buf ( n371498 , n23893 );
not ( n23895 , n371498 );
or ( n23896 , n23885 , n23895 );
not ( n23897 , n371487 );
nand ( n23898 , n23897 , n23891 );
nand ( n23899 , n23896 , n23898 );
buf ( n23900 , n23899 );
buf ( n371505 , n23900 );
xor ( n23902 , n371482 , n371483 );
xor ( n23903 , n23902 , n371505 );
buf ( n371508 , n23903 );
xor ( n23905 , n371482 , n371483 );
and ( n23906 , n23905 , n371505 );
and ( n23907 , n371482 , n371483 );
or ( n23908 , n23906 , n23907 );
buf ( n371513 , n23908 );
buf ( n371514 , n361981 );
buf ( n371515 , n14441 );
buf ( n23912 , n22944 );
buf ( n371517 , n23912 );
or ( n23914 , n367596 , n367197 );
nand ( n23915 , n23914 , n22952 );
buf ( n371520 , n23915 );
xnor ( n23917 , n371517 , n371520 );
buf ( n371522 , n23917 );
buf ( n371523 , n371522 );
xor ( n23920 , n371514 , n371515 );
xor ( n23921 , n23920 , n371523 );
buf ( n371526 , n23921 );
xor ( n23923 , n371514 , n371515 );
and ( n23924 , n23923 , n371523 );
and ( n23925 , n371514 , n371515 );
or ( n23926 , n23924 , n23925 );
buf ( n371531 , n23926 );
buf ( n371532 , n362696 );
buf ( n371533 , n362909 );
buf ( n371534 , n22950 );
not ( n23931 , n371534 );
buf ( n371536 , n366869 );
buf ( n371537 , n367107 );
nand ( n23934 , n371536 , n371537 );
buf ( n371539 , n23934 );
buf ( n371540 , n371539 );
nand ( n23937 , n23931 , n371540 );
buf ( n371542 , n23937 );
not ( n23939 , n371542 );
not ( n23940 , n23939 );
nand ( n23941 , n22947 , n22948 );
buf ( n371546 , n23941 );
not ( n23943 , n371546 );
not ( n23944 , n19848 );
not ( n23945 , n23944 );
not ( n23946 , n22944 );
or ( n23947 , n23945 , n23946 );
buf ( n23948 , n22952 );
nand ( n23949 , n23947 , n23948 );
buf ( n371554 , n23949 );
not ( n23951 , n371554 );
or ( n23952 , n23943 , n23951 );
buf ( n371557 , n22955 );
nand ( n23954 , n23952 , n371557 );
buf ( n371559 , n23954 );
not ( n23956 , n371559 );
not ( n23957 , n23956 );
or ( n23958 , n23940 , n23957 );
nand ( n23959 , n371542 , n371559 );
nand ( n23960 , n23958 , n23959 );
buf ( n371565 , n23960 );
xor ( n23962 , n371532 , n371533 );
xor ( n23963 , n23962 , n371565 );
buf ( n371568 , n23963 );
xor ( n23965 , n371532 , n371533 );
and ( n23966 , n23965 , n371565 );
and ( n23967 , n371532 , n371533 );
or ( n23968 , n23966 , n23967 );
buf ( n371573 , n23968 );
buf ( n371574 , n363482 );
buf ( n371575 , n363411 );
or ( n23972 , n366860 , n366621 );
buf ( n371577 , n23972 );
not ( n23974 , n371577 );
buf ( n371579 , n22960 );
not ( n23976 , n371579 );
or ( n23977 , n23974 , n23976 );
buf ( n371582 , n22968 );
nand ( n23979 , n23977 , n371582 );
buf ( n371584 , n23979 );
not ( n23981 , n366617 );
xor ( n23982 , n366320 , n23981 );
and ( n23983 , n371584 , n23982 );
not ( n23984 , n371584 );
not ( n23985 , n23982 );
and ( n23986 , n23984 , n23985 );
nor ( n23987 , n23983 , n23986 );
not ( n23988 , n23987 );
buf ( n371593 , n23988 );
xor ( n23990 , n371574 , n371575 );
xor ( n23991 , n23990 , n371593 );
buf ( n371596 , n23991 );
xor ( n23993 , n371574 , n371575 );
and ( n23994 , n23993 , n371593 );
and ( n23995 , n371574 , n371575 );
or ( n23996 , n23994 , n23995 );
buf ( n371601 , n23996 );
buf ( n371602 , n347747 );
buf ( n371603 , n347830 );
buf ( n371604 , n347830 );
buf ( n371605 , n347747 );
or ( n24002 , n371604 , n371605 );
buf ( n371607 , n24002 );
buf ( n371608 , n371607 );
not ( n24005 , n371602 );
not ( n24006 , n371603 );
or ( n24007 , n24005 , n24006 );
nand ( n24008 , n24007 , n371608 );
buf ( n371613 , n24008 );
buf ( n371614 , n364445 );
buf ( n371615 , n364422 );
xor ( n24012 , n371614 , n371615 );
buf ( n371617 , n24012 );
xor ( n24014 , n363959 , n363918 );
buf ( n24015 , n371111 );
buf ( n371620 , n24015 );
buf ( n371621 , n371120 );
or ( n24018 , n371620 , n371621 );
buf ( n371623 , n24018 );
not ( n24020 , n371623 );
not ( n24021 , n18533 );
not ( n24022 , n370580 );
or ( n24023 , n24021 , n24022 );
nand ( n24024 , n24023 , n366314 );
not ( n24025 , n24024 );
not ( n24026 , n24025 );
or ( n24027 , n24020 , n24026 );
or ( n24028 , n371623 , n24025 );
nand ( n24029 , n24027 , n24028 );
not ( n24030 , n24029 );
xor ( n24031 , n24014 , n24030 );
buf ( n371636 , n24031 );
buf ( n371637 , n370595 );
xor ( n24034 , n371636 , n371637 );
buf ( n371639 , n371601 );
buf ( n371640 , n370590 );
xor ( n24037 , n371639 , n371640 );
buf ( n371642 , n371596 );
xor ( n24039 , n363037 , n363126 );
xor ( n24040 , n366860 , n366621 );
not ( n24041 , n24040 );
not ( n24042 , n24041 );
not ( n24043 , n22960 );
not ( n24044 , n24043 );
not ( n24045 , n24044 );
or ( n24046 , n24042 , n24045 );
nand ( n24047 , n24043 , n24040 );
nand ( n24048 , n24046 , n24047 );
buf ( n24049 , n24048 );
buf ( n24050 , n24049 );
and ( n24051 , n24039 , n24050 );
and ( n24052 , n363037 , n363126 );
or ( n24053 , n24051 , n24052 );
buf ( n371658 , n24053 );
xor ( n24055 , n371642 , n371658 );
buf ( n371660 , n371573 );
xor ( n24057 , n363037 , n363126 );
xor ( n24058 , n24057 , n24050 );
buf ( n371663 , n24058 );
xor ( n24060 , n371660 , n371663 );
buf ( n371665 , n362576 );
buf ( n371666 , n362309 );
xor ( n24063 , n371665 , n371666 );
and ( n24064 , n23941 , n22955 );
and ( n24065 , n23949 , n24064 );
not ( n24066 , n23949 );
not ( n24067 , n24064 );
and ( n24068 , n24066 , n24067 );
nor ( n24069 , n24065 , n24068 );
buf ( n24070 , n24069 );
not ( n24071 , n24070 );
not ( n24072 , n24071 );
not ( n24073 , n24072 );
not ( n24074 , n24073 );
buf ( n371679 , n24074 );
and ( n24076 , n24063 , n371679 );
and ( n24077 , n371665 , n371666 );
or ( n24078 , n24076 , n24077 );
buf ( n371683 , n24078 );
buf ( n371684 , n371683 );
buf ( n371685 , n371568 );
xor ( n24082 , n371684 , n371685 );
buf ( n371687 , n371531 );
xor ( n24084 , n371665 , n371666 );
xor ( n24085 , n24084 , n371679 );
buf ( n371690 , n24085 );
buf ( n371691 , n371690 );
xor ( n24088 , n371687 , n371691 );
buf ( n371693 , n371365 );
buf ( n371694 , n371526 );
xor ( n24091 , n371693 , n371694 );
buf ( n371696 , n371513 );
buf ( n371697 , n371360 );
xor ( n24094 , n371696 , n371697 );
buf ( n371699 , n371508 );
buf ( n371700 , n371454 );
xor ( n24097 , n371699 , n371700 );
buf ( n371702 , n371429 );
buf ( n371703 , n371449 );
xor ( n24100 , n371702 , n371703 );
buf ( n371705 , n9377 );
buf ( n371706 , n357048 );
xor ( n24103 , n371705 , n371706 );
buf ( n371708 , n371406 );
buf ( n371709 , n370500 );
nand ( n24106 , n371708 , n371709 );
buf ( n371711 , n24106 );
buf ( n371712 , n371711 );
buf ( n371713 , n22887 );
buf ( n371714 , n370495 );
and ( n24111 , n371713 , n371714 );
buf ( n371716 , n24111 );
buf ( n371717 , n371716 );
xor ( n24114 , n371712 , n371717 );
buf ( n371719 , n24114 );
buf ( n24116 , n371719 );
not ( n24117 , n24116 );
not ( n24118 , n24117 );
buf ( n371723 , n24118 );
and ( n24120 , n24103 , n371723 );
and ( n24121 , n371705 , n371706 );
or ( n24122 , n24120 , n24121 );
buf ( n371727 , n24122 );
buf ( n371728 , n371727 );
buf ( n371729 , n371424 );
xor ( n24126 , n371728 , n371729 );
buf ( n371731 , n356419 );
buf ( n371732 , n8700 );
xor ( n24129 , n371731 , n371732 );
buf ( n371734 , n370484 );
buf ( n24131 , n371734 );
buf ( n371736 , n24131 );
buf ( n371737 , n371736 );
buf ( n371738 , n371403 );
buf ( n371739 , n370500 );
nand ( n24136 , n371738 , n371739 );
buf ( n371741 , n24136 );
buf ( n371742 , n371741 );
not ( n24139 , n371742 );
buf ( n371744 , n24139 );
buf ( n371745 , n371744 );
and ( n24142 , n371737 , n371745 );
not ( n24143 , n371737 );
buf ( n371748 , n371741 );
and ( n24145 , n24143 , n371748 );
nor ( n24146 , n24142 , n24145 );
buf ( n371751 , n24146 );
buf ( n371752 , n371751 );
and ( n24149 , n24129 , n371752 );
and ( n24150 , n371731 , n371732 );
or ( n24151 , n24149 , n24150 );
buf ( n371756 , n24151 );
buf ( n371757 , n371756 );
xor ( n24154 , n371705 , n371706 );
xor ( n24155 , n24154 , n371723 );
buf ( n371760 , n24155 );
buf ( n371761 , n371760 );
xor ( n24158 , n371757 , n371761 );
xor ( n24159 , n371731 , n371732 );
xor ( n24160 , n24159 , n371752 );
buf ( n371765 , n24160 );
not ( n24162 , n7814 );
not ( n24163 , n355536 );
or ( n24164 , n24162 , n24163 );
buf ( n371769 , n370458 );
not ( n24166 , n371769 );
buf ( n371771 , n370466 );
nand ( n24168 , n24166 , n371771 );
buf ( n371773 , n24168 );
buf ( n371774 , n371773 );
buf ( n371775 , n369116 );
buf ( n371776 , n370475 );
and ( n24173 , n371775 , n371776 );
buf ( n371778 , n24173 );
buf ( n371779 , n371778 );
xor ( n24176 , n371774 , n371779 );
buf ( n371781 , n24176 );
buf ( n371782 , n371781 );
buf ( n24179 , n371782 );
buf ( n371784 , n24179 );
buf ( n371785 , n371784 );
not ( n24182 , n371785 );
buf ( n371787 , n24182 );
nor ( n24184 , n7814 , n355536 );
or ( n24185 , n371787 , n24184 );
nand ( n24186 , n24164 , n24185 );
or ( n24187 , n371765 , n24186 );
buf ( n371792 , n24187 );
not ( n24189 , n371792 );
xor ( n24190 , n7814 , n355536 );
buf ( n371795 , n371781 );
not ( n24192 , n371795 );
buf ( n371797 , n24192 );
buf ( n371798 , n371797 );
not ( n24195 , n371798 );
buf ( n371800 , n24195 );
and ( n24197 , n24190 , n371800 );
not ( n24198 , n24190 );
and ( n24199 , n24198 , n371787 );
nor ( n24200 , n24197 , n24199 );
buf ( n371805 , n24200 );
not ( n24202 , n371805 );
buf ( n371807 , n371388 );
not ( n24204 , n371807 );
buf ( n371809 , n24204 );
buf ( n371810 , n371809 );
nand ( n24207 , n24202 , n371810 );
buf ( n371812 , n24207 );
buf ( n371813 , n371812 );
not ( n24210 , n371813 );
buf ( n371815 , n371383 );
not ( n24212 , n371815 );
buf ( n24213 , n5486 );
xor ( n24214 , n5471 , n24213 );
not ( n24215 , n371463 );
not ( n24216 , n22809 );
or ( n24217 , n24215 , n24216 );
nand ( n24218 , n24217 , n371468 );
not ( n24219 , n24218 );
not ( n24220 , n24219 );
xnor ( n24221 , n369346 , n369319 );
not ( n24222 , n24221 );
not ( n24223 , n24222 );
or ( n24224 , n24220 , n24223 );
nand ( n24225 , n24221 , n24218 );
nand ( n24226 , n24224 , n24225 );
and ( n24227 , n24214 , n24226 );
and ( n24228 , n5471 , n24213 );
or ( n24229 , n24227 , n24228 );
buf ( n371834 , n24229 );
not ( n24231 , n371834 );
buf ( n371836 , n24231 );
buf ( n371837 , n371836 );
nand ( n24234 , n24212 , n371837 );
buf ( n371839 , n24234 );
buf ( n371840 , n371839 );
not ( n24237 , n371840 );
xor ( n24238 , n5471 , n24213 );
xor ( n24239 , n24238 , n24226 );
buf ( n371844 , n24239 );
buf ( n371845 , n371481 );
or ( n24242 , n371844 , n371845 );
buf ( n371847 , n24242 );
buf ( n371848 , n371847 );
not ( n24245 , n371848 );
buf ( n371850 , n371476 );
buf ( n371851 , n12501 );
buf ( n371852 , n5220 );
xor ( n24249 , n371851 , n371852 );
buf ( n371854 , n370408 );
not ( n24251 , n371854 );
buf ( n371856 , n24251 );
buf ( n371857 , n371856 );
buf ( n371858 , n369656 );
nand ( n24255 , n371857 , n371858 );
buf ( n371860 , n24255 );
nand ( n24257 , n371860 , n370412 );
not ( n24258 , n24257 );
not ( n24259 , n24258 );
buf ( n371864 , n370403 );
buf ( n24261 , n371864 );
buf ( n371866 , n24261 );
buf ( n371867 , n371866 );
not ( n24264 , n371867 );
buf ( n371869 , n24264 );
not ( n24266 , n371869 );
or ( n24267 , n24259 , n24266 );
nand ( n24268 , n24257 , n371866 );
nand ( n24269 , n24267 , n24268 );
buf ( n371874 , n24269 );
not ( n24271 , n371874 );
buf ( n371876 , n24271 );
buf ( n371877 , n371876 );
not ( n24274 , n371877 );
buf ( n371879 , n24274 );
buf ( n371880 , n371879 );
and ( n24277 , n24249 , n371880 );
and ( n24278 , n371851 , n371852 );
or ( n24279 , n24277 , n24278 );
buf ( n371884 , n24279 );
buf ( n371885 , n371884 );
or ( n24282 , n371850 , n371885 );
buf ( n371887 , n24282 );
buf ( n371888 , n371887 );
not ( n24285 , n371888 );
xor ( n24286 , n371851 , n371852 );
xor ( n24287 , n24286 , n371880 );
buf ( n371892 , n24287 );
not ( n24289 , n371892 );
not ( n24290 , n371338 );
nand ( n24291 , n24289 , n24290 );
not ( n24292 , n24291 );
not ( n24293 , n371314 );
not ( n24294 , n24293 );
not ( n24295 , n371333 );
not ( n24296 , n24295 );
or ( n24297 , n24294 , n24296 );
buf ( n371902 , n371309 );
buf ( n371903 , n371287 );
nor ( n24300 , n371902 , n371903 );
buf ( n371905 , n24300 );
buf ( n371906 , n371905 );
buf ( n371907 , n371282 );
buf ( n371908 , n2672 );
buf ( n371909 , n350336 );
xor ( n24306 , n371908 , n371909 );
buf ( n371911 , n22265 );
buf ( n371912 , n370252 );
nand ( n24309 , n371911 , n371912 );
buf ( n371914 , n24309 );
buf ( n371915 , n371914 );
buf ( n371916 , n370245 );
not ( n24313 , n371916 );
buf ( n371918 , n24313 );
buf ( n371919 , n371918 );
and ( n24316 , n371915 , n371919 );
not ( n24317 , n371915 );
buf ( n371922 , n370245 );
and ( n24319 , n24317 , n371922 );
nor ( n24320 , n24316 , n24319 );
buf ( n371925 , n24320 );
buf ( n371926 , n371925 );
and ( n24323 , n24306 , n371926 );
and ( n24324 , n371908 , n371909 );
or ( n24325 , n24323 , n24324 );
buf ( n371930 , n24325 );
buf ( n371931 , n371930 );
or ( n24328 , n371907 , n371931 );
buf ( n371933 , n24328 );
not ( n24330 , n371933 );
buf ( n371935 , n371253 );
xor ( n24332 , n371908 , n371909 );
xor ( n24333 , n24332 , n371926 );
buf ( n371938 , n24333 );
buf ( n371939 , n371938 );
xor ( n24336 , n371935 , n371939 );
xor ( n24337 , n371212 , n371192 );
xor ( n24338 , n371187 , n371164 );
buf ( n371943 , n371159 );
not ( n24340 , n371943 );
buf ( n371945 , n24340 );
buf ( n371946 , n371945 );
buf ( n371947 , n371607 );
not ( n24344 , n371947 );
buf ( n371949 , n24344 );
buf ( n371950 , n371949 );
nand ( n24347 , n371946 , n371950 );
buf ( n371952 , n24347 );
not ( n24349 , n347973 );
buf ( n371954 , n24349 );
buf ( n371955 , n348052 );
and ( n24352 , n371954 , n371955 );
buf ( n371957 , n24352 );
buf ( n371958 , n371957 );
buf ( n371959 , n347976 );
or ( n24356 , n371958 , n371959 );
xor ( n24357 , n347818 , n347901 );
buf ( n371962 , n24357 );
nand ( n24359 , n24356 , n371962 );
buf ( n371964 , n24359 );
buf ( n371965 , n371964 );
not ( n24362 , n371965 );
buf ( n371967 , n24362 );
buf ( n371968 , n371967 );
and ( n24365 , n347818 , n347901 );
buf ( n371970 , n24365 );
xor ( n24367 , n371968 , n371970 );
buf ( n371972 , n371613 );
and ( n24369 , n24367 , n371972 );
or ( n24370 , n24369 , C0 );
buf ( n371975 , n24370 );
and ( n24372 , n371952 , n371975 );
buf ( n371977 , n371945 );
buf ( n371978 , n371949 );
nor ( n24375 , n371977 , n371978 );
buf ( n371980 , n24375 );
nor ( n24377 , n24372 , n371980 );
not ( n24378 , n24377 );
and ( n24379 , n24338 , n24378 );
and ( n24380 , n371187 , n371164 );
or ( n24381 , n24379 , n24380 );
and ( n24382 , n24337 , n24381 );
and ( n24383 , n371212 , n371192 );
nor ( n24384 , n24382 , n24383 );
buf ( n371989 , n24384 );
buf ( n371990 , n371248 );
buf ( n371991 , n371217 );
nor ( n24388 , n371990 , n371991 );
buf ( n371993 , n24388 );
buf ( n371994 , n371993 );
or ( n24391 , n371989 , n371994 );
buf ( n371996 , n371248 );
buf ( n371997 , n371217 );
nand ( n24394 , n371996 , n371997 );
buf ( n371999 , n24394 );
buf ( n372000 , n371999 );
nand ( n24397 , n24391 , n372000 );
buf ( n372002 , n24397 );
buf ( n372003 , n372002 );
and ( n24400 , n24336 , n372003 );
and ( n24401 , n371935 , n371939 );
or ( n24402 , n24400 , n24401 );
buf ( n372007 , n24402 );
not ( n24404 , n372007 );
or ( n24405 , n24330 , n24404 );
nand ( n24406 , n371282 , n371930 );
nand ( n24407 , n24405 , n24406 );
not ( n24408 , n24407 );
buf ( n372013 , n24408 );
or ( n24410 , n371906 , n372013 );
buf ( n372015 , n371309 );
buf ( n372016 , n371287 );
nand ( n24413 , n372015 , n372016 );
buf ( n372018 , n24413 );
buf ( n372019 , n372018 );
nand ( n24416 , n24410 , n372019 );
buf ( n372021 , n24416 );
nand ( n24418 , n24297 , n372021 );
nand ( n24419 , n371333 , n371314 );
nand ( n24420 , n24418 , n24419 );
not ( n24421 , n24420 );
or ( n24422 , n24292 , n24421 );
nand ( n24423 , n371892 , n371338 );
nand ( n24424 , n24422 , n24423 );
buf ( n372029 , n24424 );
not ( n24426 , n372029 );
or ( n24427 , n24285 , n24426 );
buf ( n372032 , n371476 );
buf ( n372033 , n371884 );
nand ( n24430 , n372032 , n372033 );
buf ( n372035 , n24430 );
buf ( n372036 , n372035 );
nand ( n24433 , n24427 , n372036 );
buf ( n372038 , n24433 );
buf ( n372039 , n372038 );
not ( n24436 , n372039 );
or ( n24437 , n24245 , n24436 );
buf ( n372042 , n24239 );
buf ( n372043 , n371481 );
nand ( n24440 , n372042 , n372043 );
buf ( n372045 , n24440 );
buf ( n372046 , n372045 );
nand ( n24443 , n24437 , n372046 );
buf ( n372048 , n24443 );
buf ( n372049 , n372048 );
not ( n24446 , n372049 );
or ( n24447 , n24237 , n24446 );
buf ( n372052 , n371383 );
buf ( n372053 , n24229 );
nand ( n24450 , n372052 , n372053 );
buf ( n372055 , n24450 );
buf ( n372056 , n372055 );
nand ( n24453 , n24447 , n372056 );
buf ( n372058 , n24453 );
buf ( n372059 , n372058 );
not ( n24456 , n372059 );
or ( n24457 , n24210 , n24456 );
buf ( n372062 , n24200 );
buf ( n372063 , n371388 );
nand ( n24460 , n372062 , n372063 );
buf ( n372065 , n24460 );
buf ( n372066 , n372065 );
nand ( n24463 , n24457 , n372066 );
buf ( n372068 , n24463 );
buf ( n372069 , n372068 );
not ( n24466 , n372069 );
or ( n24467 , n24189 , n24466 );
buf ( n372072 , n371765 );
buf ( n372073 , n24186 );
nand ( n24470 , n372072 , n372073 );
buf ( n372075 , n24470 );
buf ( n372076 , n372075 );
nand ( n24473 , n24467 , n372076 );
buf ( n372078 , n24473 );
buf ( n372079 , n372078 );
and ( n24476 , n24158 , n372079 );
and ( n24477 , n371757 , n371761 );
or ( n24478 , n24476 , n24477 );
buf ( n372083 , n24478 );
buf ( n372084 , n372083 );
and ( n24481 , n24126 , n372084 );
and ( n24482 , n371728 , n371729 );
or ( n24483 , n24481 , n24482 );
buf ( n372088 , n24483 );
buf ( n372089 , n372088 );
and ( n24486 , n24100 , n372089 );
and ( n24487 , n371702 , n371703 );
or ( n24488 , n24486 , n24487 );
buf ( n372093 , n24488 );
buf ( n372094 , n372093 );
and ( n24491 , n24097 , n372094 );
and ( n24492 , n371699 , n371700 );
or ( n24493 , n24491 , n24492 );
buf ( n372098 , n24493 );
buf ( n372099 , n372098 );
and ( n24496 , n24094 , n372099 );
and ( n24497 , n371696 , n371697 );
or ( n24498 , n24496 , n24497 );
buf ( n372103 , n24498 );
buf ( n372104 , n372103 );
and ( n24501 , n24091 , n372104 );
and ( n24502 , n371693 , n371694 );
or ( n24503 , n24501 , n24502 );
buf ( n372108 , n24503 );
buf ( n372109 , n372108 );
and ( n24506 , n24088 , n372109 );
and ( n24507 , n371687 , n371691 );
or ( n24508 , n24506 , n24507 );
buf ( n372113 , n24508 );
buf ( n372114 , n372113 );
and ( n24511 , n24082 , n372114 );
and ( n24512 , n371684 , n371685 );
or ( n24513 , n24511 , n24512 );
buf ( n372118 , n24513 );
buf ( n372119 , n372118 );
and ( n24516 , n24060 , n372119 );
and ( n24517 , n371660 , n371663 );
or ( n24518 , n24516 , n24517 );
buf ( n372123 , n24518 );
buf ( n372124 , n372123 );
and ( n24521 , n24055 , n372124 );
and ( n24522 , n371642 , n371658 );
or ( n24523 , n24521 , n24522 );
buf ( n372128 , n24523 );
buf ( n372129 , n372128 );
and ( n24526 , n24037 , n372129 );
and ( n24527 , n371639 , n371640 );
or ( n24528 , n24526 , n24527 );
buf ( n372133 , n24528 );
buf ( n372134 , n372133 );
and ( n24531 , n24034 , n372134 );
and ( n24532 , n371636 , n371637 );
or ( n24533 , n24531 , n24532 );
buf ( n372138 , n24533 );
buf ( n372139 , n372138 );
buf ( n372140 , n371136 );
not ( n24537 , n372140 );
buf ( n372142 , n24537 );
buf ( n372143 , n372142 );
xor ( n24540 , n363959 , n363918 );
and ( n24541 , n24540 , n24030 );
and ( n24542 , n363959 , n363918 );
or ( n24543 , n24541 , n24542 );
buf ( n372148 , n24543 );
not ( n24545 , n372148 );
buf ( n372150 , n24545 );
buf ( n372151 , n372150 );
nand ( n24548 , n372143 , n372151 );
buf ( n372153 , n24548 );
buf ( n372154 , n372153 );
and ( n24551 , n372139 , n372154 );
buf ( n372156 , n372142 );
buf ( n372157 , n372150 );
nor ( n24554 , n372156 , n372157 );
buf ( n372159 , n24554 );
buf ( n372160 , n372159 );
nor ( n24557 , n24551 , n372160 );
buf ( n372162 , n24557 );
buf ( n372163 , n372162 );
buf ( n372164 , n372138 );
not ( n24561 , n372164 );
buf ( n372166 , n372159 );
not ( n24563 , n372166 );
and ( n24564 , n24561 , n24563 );
buf ( n372169 , n372153 );
not ( n24566 , n372169 );
buf ( n372171 , n24566 );
buf ( n372172 , n372171 );
nor ( n24569 , n24564 , n372172 );
buf ( n372174 , n24569 );
buf ( n372175 , n372174 );
buf ( n372176 , n371141 );
buf ( n372177 , n371617 );
xor ( n24574 , n372176 , n372177 );
buf ( n372179 , n24574 );
buf ( n372180 , n372179 );
and ( n24577 , n372180 , n372175 );
not ( n24578 , n372180 );
and ( n24579 , n24578 , n372163 );
nor ( n24580 , n24577 , n24579 );
buf ( n372185 , n24580 );
buf ( n372186 , n372150 );
buf ( n372187 , n371136 );
and ( n24584 , n372186 , n372187 );
not ( n24585 , n372186 );
buf ( n372190 , n372142 );
and ( n24587 , n24585 , n372190 );
nor ( n24588 , n24584 , n24587 );
buf ( n372193 , n24588 );
buf ( n372194 , n372193 );
buf ( n372195 , n372138 );
buf ( n372196 , n372193 );
buf ( n372197 , n372138 );
not ( n24594 , n372194 );
not ( n24595 , n372195 );
or ( n24596 , n24594 , n24595 );
or ( n24597 , n372196 , n372197 );
nand ( n24598 , n24596 , n24597 );
buf ( n372203 , n24598 );
xor ( n24600 , n371636 , n371637 );
xor ( n24601 , n24600 , n372134 );
buf ( n372206 , n24601 );
xor ( n24603 , n371639 , n371640 );
xor ( n24604 , n24603 , n372129 );
buf ( n372209 , n24604 );
xor ( n24606 , n371642 , n371658 );
xor ( n24607 , n24606 , n372124 );
buf ( n372212 , n24607 );
xor ( n24609 , n371660 , n371663 );
xor ( n24610 , n24609 , n372119 );
buf ( n372215 , n24610 );
xor ( n24612 , n371684 , n371685 );
xor ( n24613 , n24612 , n372114 );
buf ( n372218 , n24613 );
xor ( n24615 , n371687 , n371691 );
xor ( n24616 , n24615 , n372109 );
buf ( n372221 , n24616 );
xor ( n24618 , n371693 , n371694 );
xor ( n24619 , n24618 , n372104 );
buf ( n372224 , n24619 );
xor ( n24621 , n371696 , n371697 );
xor ( n24622 , n24621 , n372099 );
buf ( n372227 , n24622 );
xor ( n24624 , n371699 , n371700 );
xor ( n24625 , n24624 , n372094 );
buf ( n372230 , n24625 );
xor ( n24627 , n371702 , n371703 );
xor ( n24628 , n24627 , n372089 );
buf ( n372233 , n24628 );
xor ( n24630 , n371728 , n371729 );
xor ( n24631 , n24630 , n372084 );
buf ( n372236 , n24631 );
xor ( n24633 , n371757 , n371761 );
xor ( n24634 , n24633 , n372079 );
buf ( n372239 , n24634 );
buf ( n372240 , n372068 );
buf ( n372241 , n371765 );
buf ( n372242 , n24186 );
xnor ( n24639 , n372241 , n372242 );
buf ( n372244 , n24639 );
buf ( n372245 , n372244 );
buf ( n372246 , n372244 );
buf ( n372247 , n372068 );
not ( n24644 , n372240 );
not ( n24645 , n372245 );
or ( n24646 , n24644 , n24645 );
or ( n24647 , n372246 , n372247 );
nand ( n24648 , n24646 , n24647 );
buf ( n372253 , n24648 );
buf ( n372254 , n372058 );
and ( n24651 , n24200 , n371809 );
not ( n24652 , n24200 );
and ( n24653 , n24652 , n371388 );
nor ( n24654 , n24651 , n24653 );
buf ( n372259 , n24654 );
buf ( n372260 , n24654 );
buf ( n372261 , n372058 );
not ( n24658 , n372254 );
not ( n24659 , n372259 );
or ( n24660 , n24658 , n24659 );
or ( n24661 , n372260 , n372261 );
nand ( n24662 , n24660 , n24661 );
buf ( n372267 , n24662 );
buf ( n372268 , n372048 );
buf ( n372269 , n371383 );
buf ( n372270 , n24229 );
xnor ( n24667 , n372269 , n372270 );
buf ( n372272 , n24667 );
buf ( n372273 , n372272 );
buf ( n372274 , n372272 );
buf ( n372275 , n372048 );
not ( n24672 , n372268 );
not ( n24673 , n372273 );
or ( n24674 , n24672 , n24673 );
or ( n24675 , n372274 , n372275 );
nand ( n24676 , n24674 , n24675 );
buf ( n372281 , n24676 );
buf ( n372282 , n372038 );
buf ( n372283 , n24239 );
buf ( n372284 , n371481 );
xor ( n24681 , n372283 , n372284 );
buf ( n372286 , n24681 );
buf ( n372287 , n372286 );
xor ( n24684 , n372282 , n372287 );
buf ( n372289 , n24684 );
buf ( n372290 , n24424 );
buf ( n372291 , n371476 );
buf ( n372292 , n371884 );
xor ( n24689 , n372291 , n372292 );
buf ( n372294 , n24689 );
buf ( n372295 , n372294 );
xor ( n24692 , n372290 , n372295 );
buf ( n372297 , n24692 );
buf ( n372298 , n24408 );
buf ( n372299 , n24407 );
buf ( n372300 , n371309 );
buf ( n372301 , n371287 );
xor ( n24698 , n372300 , n372301 );
buf ( n372303 , n24698 );
buf ( n372304 , n372303 );
and ( n24701 , n372304 , n372299 );
not ( n24702 , n372304 );
and ( n24703 , n24702 , n372298 );
nor ( n24704 , n24701 , n24703 );
buf ( n372309 , n24704 );
buf ( n372310 , n372007 );
buf ( n372311 , n371282 );
buf ( n372312 , n371930 );
xor ( n24709 , n372311 , n372312 );
buf ( n372314 , n24709 );
buf ( n372315 , n372314 );
xor ( n24712 , n372310 , n372315 );
buf ( n372317 , n24712 );
xor ( n24714 , n371935 , n371939 );
xor ( n24715 , n24714 , n372003 );
buf ( n372320 , n24715 );
buf ( n372321 , n371159 );
buf ( n372322 , n371607 );
xor ( n24719 , n372321 , n372322 );
buf ( n372324 , n24719 );
buf ( n372325 , n372324 );
buf ( n372326 , n371975 );
xor ( n24723 , n372325 , n372326 );
buf ( n372328 , n24723 );
xor ( n24725 , n371968 , n371970 );
xor ( n24726 , n24725 , n371972 );
buf ( n372331 , n24726 );
buf ( n372332 , n371957 );
not ( n24729 , n347901 );
and ( n24730 , n347818 , n347976 );
not ( n24731 , n347818 );
and ( n24732 , n24731 , n24349 );
nor ( n24733 , n24730 , n24732 );
not ( n24734 , n24733 );
or ( n24735 , n24729 , n24734 );
or ( n24736 , n347901 , n24733 );
nand ( n24737 , n24735 , n24736 );
buf ( n372342 , n24737 );
buf ( n372343 , n371957 );
buf ( n372344 , n24737 );
not ( n24741 , n372332 );
not ( n24742 , n372342 );
or ( n24743 , n24741 , n24742 );
or ( n24744 , n372343 , n372344 );
nand ( n24745 , n24743 , n24744 );
buf ( n372350 , n24745 );
xor ( n24747 , n371954 , n371955 );
buf ( n372352 , n24747 );
buf ( n372353 , n371333 );
buf ( n372354 , n371314 );
xor ( n24751 , n372353 , n372354 );
buf ( n372356 , n24751 );
buf ( n372357 , n371892 );
buf ( n372358 , n371338 );
xor ( n24755 , n372357 , n372358 );
buf ( n372360 , n24755 );
buf ( n372361 , n371248 );
buf ( n372362 , n371217 );
xor ( n24759 , n372361 , n372362 );
buf ( n372364 , n24759 );
buf ( n372365 , n24384 );
buf ( n372366 , n372364 );
xnor ( n24763 , n372365 , n372366 );
buf ( n372368 , n24763 );
buf ( n372369 , n347515 );
buf ( n372370 , n12493 );
xor ( n24767 , n358917 , n358921 );
xor ( n24768 , n24767 , n359044 );
buf ( n372373 , n24768 );
buf ( n372374 , n372373 );
xor ( n24771 , n372369 , n372370 );
xor ( n24772 , n24771 , n372374 );
buf ( n372377 , n24772 );
xor ( n24774 , n372369 , n372370 );
and ( n24775 , n24774 , n372374 );
and ( n24776 , n372369 , n372370 );
or ( n24777 , n24775 , n24776 );
buf ( n372382 , n24777 );
buf ( n372383 , n347591 );
buf ( n372384 , n12498 );
nor ( n24781 , n11225 , n358872 );
not ( n24782 , n359048 );
nand ( n24783 , n24781 , n24782 );
not ( n24784 , n11226 );
nand ( n24785 , n24784 , n359048 );
not ( n24786 , n358872 );
nor ( n24787 , n24786 , n358901 );
nand ( n24788 , n24782 , n24787 );
nand ( n24789 , n11374 , n359048 );
nand ( n24790 , n24783 , n24785 , n24788 , n24789 );
buf ( n372395 , n24790 );
xor ( n24792 , n372383 , n372384 );
xor ( n24793 , n24792 , n372395 );
buf ( n372398 , n24793 );
xor ( n24795 , n372383 , n372384 );
and ( n24796 , n24795 , n372395 );
and ( n24797 , n372383 , n372384 );
or ( n24798 , n24796 , n24797 );
buf ( n372403 , n24798 );
buf ( n372404 , n348556 );
buf ( n372405 , n12485 );
buf ( n372406 , n359067 );
not ( n24803 , n372406 );
buf ( n372408 , n359073 );
nand ( n24805 , n24803 , n372408 );
buf ( n372410 , n24805 );
buf ( n372411 , n372410 );
buf ( n372412 , n11375 );
and ( n24809 , n372411 , n372412 );
not ( n24810 , n372411 );
not ( n24811 , n11375 );
buf ( n372416 , n24811 );
and ( n24813 , n24810 , n372416 );
nor ( n24814 , n24809 , n24813 );
buf ( n372419 , n24814 );
buf ( n372420 , n372419 );
xor ( n24817 , n372404 , n372405 );
xor ( n24818 , n24817 , n372420 );
buf ( n372423 , n24818 );
xor ( n24820 , n372404 , n372405 );
and ( n24821 , n24820 , n372420 );
and ( n24822 , n372404 , n372405 );
or ( n24823 , n24821 , n24822 );
buf ( n372428 , n24823 );
buf ( n372429 , n350044 );
buf ( n372430 , n12499 );
xor ( n24827 , n358865 , n358868 );
xor ( n24828 , n24827 , n359076 );
buf ( n372433 , n24828 );
xor ( n24830 , n372429 , n372430 );
xor ( n24831 , n24830 , n372433 );
buf ( n372436 , n24831 );
xor ( n24833 , n372429 , n372430 );
and ( n24834 , n24833 , n372433 );
and ( n24835 , n372429 , n372430 );
or ( n24836 , n24834 , n24835 );
buf ( n372441 , n24836 );
buf ( n372442 , n350365 );
buf ( n372443 , n12490 );
xor ( n24840 , n358685 , n358688 );
xor ( n24841 , n24840 , n11403 );
buf ( n372446 , n24841 );
xor ( n24843 , n372442 , n372443 );
xor ( n24844 , n24843 , n372446 );
buf ( n372449 , n24844 );
xor ( n24846 , n372442 , n372443 );
and ( n24847 , n24846 , n372446 );
and ( n24848 , n372442 , n372443 );
or ( n24849 , n24847 , n24848 );
buf ( n372454 , n24849 );
buf ( n372455 , n350651 );
buf ( n372456 , n12503 );
buf ( n372457 , n358640 );
buf ( n372458 , n359088 );
nand ( n24855 , n372457 , n372458 );
buf ( n372460 , n24855 );
buf ( n372461 , n372460 );
not ( n24858 , n372461 );
buf ( n372463 , n11406 );
not ( n24860 , n372463 );
or ( n24861 , n24858 , n24860 );
not ( n24862 , n372460 );
not ( n24863 , n11406 );
nand ( n24864 , n24862 , n24863 );
buf ( n372469 , n24864 );
nand ( n24866 , n24861 , n372469 );
buf ( n372471 , n24866 );
buf ( n372472 , n372471 );
xor ( n24869 , n372455 , n372456 );
xor ( n24870 , n24869 , n372472 );
buf ( n372475 , n24870 );
xor ( n24872 , n372455 , n372456 );
and ( n24873 , n24872 , n372472 );
and ( n24874 , n372455 , n372456 );
or ( n24875 , n24873 , n24874 );
buf ( n372480 , n24875 );
buf ( n372481 , n350977 );
buf ( n372482 , n12489 );
not ( n24879 , n359160 );
not ( n24880 , n359096 );
or ( n24881 , n24879 , n24880 );
nand ( n24882 , n24881 , n11488 );
not ( n24883 , n24882 );
not ( n24884 , n11413 );
or ( n24885 , n24883 , n24884 );
or ( n24886 , n11413 , n24882 );
nand ( n24887 , n24885 , n24886 );
buf ( n372492 , n24887 );
xor ( n24889 , n372481 , n372482 );
xor ( n24890 , n24889 , n372492 );
buf ( n372495 , n24890 );
xor ( n24892 , n372481 , n372482 );
and ( n24893 , n24892 , n372492 );
and ( n24894 , n372481 , n372482 );
or ( n24895 , n24893 , n24894 );
buf ( n372500 , n24895 );
buf ( n372501 , n351506 );
buf ( n372502 , n12488 );
buf ( n372503 , n359175 );
not ( n24900 , n372503 );
buf ( n372505 , n359203 );
buf ( n372506 , n359209 );
nor ( n24903 , n372505 , n372506 );
buf ( n372508 , n24903 );
buf ( n372509 , n372508 );
not ( n24906 , n372509 );
buf ( n372511 , n359222 );
nand ( n24908 , n24906 , n372511 );
buf ( n372513 , n24908 );
buf ( n372514 , n372513 );
not ( n24911 , n372514 );
or ( n24912 , n24900 , n24911 );
buf ( n372517 , n359175 );
not ( n24914 , n372517 );
buf ( n372519 , n372513 );
not ( n24916 , n372519 );
buf ( n372521 , n24916 );
buf ( n372522 , n372521 );
nand ( n24919 , n24914 , n372522 );
buf ( n372524 , n24919 );
buf ( n372525 , n372524 );
nand ( n24922 , n24912 , n372525 );
buf ( n372527 , n24922 );
buf ( n372528 , n372527 );
xor ( n24925 , n372501 , n372502 );
xor ( n24926 , n24925 , n372528 );
buf ( n372531 , n24926 );
xor ( n24928 , n372501 , n372502 );
and ( n24929 , n24928 , n372528 );
and ( n24930 , n372501 , n372502 );
or ( n24931 , n24929 , n24930 );
buf ( n372536 , n24931 );
buf ( n372537 , n15521 );
buf ( n372538 , n363204 );
buf ( n372539 , n357376 );
not ( n24936 , n372539 );
buf ( n372541 , n606 );
not ( n24938 , n372541 );
or ( n24939 , n17012 , n23108 );
not ( n24940 , n17011 );
nand ( n24941 , n24940 , n23108 );
nand ( n24942 , n24939 , n24941 );
buf ( n24943 , n24942 );
buf ( n372548 , n24943 );
not ( n24945 , n372548 );
buf ( n372550 , n24945 );
buf ( n372551 , n372550 );
not ( n24948 , n372551 );
or ( n24949 , n24938 , n24948 );
buf ( n372554 , n24943 );
not ( n24951 , n372554 );
buf ( n372556 , n24951 );
buf ( n372557 , n372556 );
not ( n24954 , n372557 );
buf ( n372559 , n24954 );
buf ( n372560 , n372559 );
buf ( n372561 , n9642 );
nand ( n24958 , n372560 , n372561 );
buf ( n372563 , n24958 );
buf ( n372564 , n372563 );
nand ( n24961 , n24949 , n372564 );
buf ( n372566 , n24961 );
buf ( n372567 , n372566 );
not ( n24964 , n372567 );
or ( n24965 , n24936 , n24964 );
buf ( n372570 , n606 );
not ( n24967 , n372570 );
not ( n24968 , n370821 );
nand ( n24969 , n14500 , n8323 , n16900 );
not ( n24970 , n24969 );
or ( n24971 , n24968 , n24970 );
not ( n24972 , n8323 );
nor ( n24973 , n16955 , n24972 );
nand ( n24974 , n14500 , n24973 , n16900 );
nand ( n24975 , n24971 , n24974 );
buf ( n372580 , n24975 );
not ( n24977 , n372580 );
buf ( n372582 , n24977 );
buf ( n372583 , n372582 );
not ( n24980 , n372583 );
or ( n24981 , n24967 , n24980 );
buf ( n372586 , n372582 );
not ( n24983 , n372586 );
buf ( n372588 , n24983 );
buf ( n372589 , n372588 );
buf ( n372590 , n9642 );
nand ( n24987 , n372589 , n372590 );
buf ( n372592 , n24987 );
buf ( n372593 , n372592 );
nand ( n24990 , n24981 , n372593 );
buf ( n372595 , n24990 );
buf ( n372596 , n372595 );
buf ( n372597 , n607 );
nand ( n24994 , n372596 , n372597 );
buf ( n372599 , n24994 );
buf ( n372600 , n372599 );
nand ( n24997 , n24965 , n372600 );
buf ( n372602 , n24997 );
buf ( n372603 , n372602 );
buf ( n372604 , n348855 );
buf ( n372605 , n592 );
and ( n25002 , n372604 , n372605 );
buf ( n372607 , n25002 );
buf ( n372608 , n372607 );
buf ( n372609 , n348946 );
not ( n25006 , n372609 );
buf ( n372611 , n592 );
not ( n25008 , n372611 );
buf ( n372613 , n354248 );
not ( n25010 , n372613 );
or ( n25011 , n25008 , n25010 );
buf ( n372616 , n348910 );
buf ( n372617 , n6561 );
nand ( n25014 , n372616 , n372617 );
buf ( n372619 , n25014 );
buf ( n372620 , n372619 );
nand ( n25017 , n25011 , n372620 );
buf ( n372622 , n25017 );
buf ( n372623 , n372622 );
not ( n25020 , n372623 );
or ( n25021 , n25006 , n25020 );
buf ( n372626 , n592 );
not ( n25023 , n372626 );
buf ( n372628 , n351952 );
not ( n25025 , n372628 );
or ( n25026 , n25023 , n25025 );
buf ( n372631 , n348910 );
buf ( n372632 , n351958 );
nand ( n25029 , n372631 , n372632 );
buf ( n372634 , n25029 );
buf ( n372635 , n372634 );
nand ( n25032 , n25026 , n372635 );
buf ( n372637 , n25032 );
buf ( n372638 , n372637 );
buf ( n372639 , n1250 );
nand ( n25036 , n372638 , n372639 );
buf ( n372641 , n25036 );
buf ( n372642 , n372641 );
nand ( n25039 , n25021 , n372642 );
buf ( n372644 , n25039 );
buf ( n372645 , n372644 );
xor ( n25042 , n372608 , n372645 );
buf ( n372647 , n349035 );
not ( n25044 , n372647 );
buf ( n372649 , n594 );
not ( n25046 , n372649 );
buf ( n372651 , n351901 );
not ( n25048 , n372651 );
or ( n25049 , n25046 , n25048 );
buf ( n372654 , n4221 );
buf ( n372655 , n348975 );
nand ( n25052 , n372654 , n372655 );
buf ( n372657 , n25052 );
buf ( n372658 , n372657 );
nand ( n25055 , n25049 , n372658 );
buf ( n372660 , n25055 );
buf ( n372661 , n372660 );
not ( n25058 , n372661 );
or ( n25059 , n25044 , n25058 );
buf ( n372664 , n594 );
not ( n25061 , n372664 );
buf ( n372666 , n7445 );
not ( n25063 , n372666 );
or ( n25064 , n25061 , n25063 );
not ( n25065 , n352066 );
buf ( n372670 , n25065 );
buf ( n372671 , n348975 );
nand ( n25068 , n372670 , n372671 );
buf ( n372673 , n25068 );
buf ( n372674 , n372673 );
nand ( n25071 , n25064 , n372674 );
buf ( n372676 , n25071 );
buf ( n372677 , n372676 );
buf ( n372678 , n1397 );
nand ( n25075 , n372677 , n372678 );
buf ( n372680 , n25075 );
buf ( n372681 , n372680 );
nand ( n25078 , n25059 , n372681 );
buf ( n372683 , n25078 );
buf ( n372684 , n372683 );
and ( n25081 , n25042 , n372684 );
and ( n25082 , n372608 , n372645 );
or ( n25083 , n25081 , n25082 );
buf ( n372688 , n25083 );
buf ( n372689 , n372688 );
buf ( n372690 , n592 );
not ( n25087 , n372690 );
buf ( n372692 , n355089 );
nor ( n25089 , n25087 , n372692 );
buf ( n372694 , n25089 );
buf ( n372695 , n372694 );
buf ( n372696 , n348946 );
not ( n25093 , n372696 );
buf ( n372698 , n592 );
not ( n25095 , n372698 );
buf ( n372700 , n7445 );
not ( n25097 , n372700 );
or ( n25098 , n25095 , n25097 );
buf ( n372703 , n25065 );
buf ( n372704 , n348910 );
nand ( n25101 , n372703 , n372704 );
buf ( n372706 , n25101 );
buf ( n372707 , n372706 );
nand ( n25104 , n25098 , n372707 );
buf ( n372709 , n25104 );
buf ( n372710 , n372709 );
not ( n25107 , n372710 );
or ( n25108 , n25093 , n25107 );
buf ( n372713 , n372622 );
buf ( n372714 , n1250 );
nand ( n25111 , n372713 , n372714 );
buf ( n372716 , n25111 );
buf ( n372717 , n372716 );
nand ( n25114 , n25108 , n372717 );
buf ( n372719 , n25114 );
buf ( n372720 , n372719 );
xor ( n25117 , n372695 , n372720 );
buf ( n372722 , n349035 );
not ( n25119 , n372722 );
and ( n25120 , n594 , n351870 );
not ( n25121 , n594 );
and ( n25122 , n25121 , n4183 );
or ( n25123 , n25120 , n25122 );
buf ( n372728 , n25123 );
not ( n25125 , n372728 );
or ( n25126 , n25119 , n25125 );
buf ( n372731 , n372660 );
buf ( n372732 , n1397 );
nand ( n25129 , n372731 , n372732 );
buf ( n372734 , n25129 );
buf ( n372735 , n372734 );
nand ( n25132 , n25126 , n372735 );
buf ( n372737 , n25132 );
buf ( n372738 , n372737 );
xor ( n25135 , n25117 , n372738 );
buf ( n372740 , n25135 );
buf ( n372741 , n372740 );
xor ( n25138 , n372689 , n372741 );
buf ( n372743 , n347319 );
not ( n25140 , n372743 );
buf ( n372745 , n596 );
not ( n25142 , n372745 );
buf ( n372747 , n354087 );
not ( n25144 , n372747 );
or ( n25145 , n25142 , n25144 );
nand ( n25146 , n9814 , n348865 );
buf ( n372751 , n25146 );
nand ( n25148 , n25145 , n372751 );
buf ( n372753 , n25148 );
buf ( n372754 , n372753 );
not ( n25151 , n372754 );
or ( n25152 , n25140 , n25151 );
buf ( n372757 , n596 );
not ( n25154 , n372757 );
buf ( n372759 , n355178 );
not ( n25156 , n372759 );
or ( n25157 , n25154 , n25156 );
buf ( n372762 , n6458 );
buf ( n372763 , n348865 );
nand ( n25160 , n372762 , n372763 );
buf ( n372765 , n25160 );
buf ( n372766 , n372765 );
nand ( n25163 , n25157 , n372766 );
buf ( n372768 , n25163 );
buf ( n372769 , n372768 );
buf ( n372770 , n348898 );
buf ( n25167 , n372770 );
buf ( n372772 , n25167 );
buf ( n372773 , n372772 );
nand ( n25170 , n372769 , n372773 );
buf ( n372775 , n25170 );
buf ( n372776 , n372775 );
nand ( n25173 , n25152 , n372776 );
buf ( n372778 , n25173 );
buf ( n372779 , n372778 );
and ( n25176 , n25138 , n372779 );
and ( n25177 , n372689 , n372741 );
or ( n25178 , n25176 , n25177 );
buf ( n372783 , n25178 );
buf ( n372784 , n372783 );
not ( n25181 , n4362 );
not ( n25182 , n347312 );
not ( n25183 , n8333 );
or ( n25184 , n25182 , n25183 );
nand ( n25185 , n598 , n8330 );
nand ( n25186 , n25184 , n25185 );
not ( n25187 , n25186 );
or ( n25188 , n25181 , n25187 );
buf ( n372793 , n598 );
not ( n25190 , n372793 );
not ( n25191 , n7359 );
buf ( n372796 , n25191 );
not ( n25193 , n372796 );
or ( n25194 , n25190 , n25193 );
buf ( n372799 , n7359 );
buf ( n372800 , n347312 );
nand ( n25197 , n372799 , n372800 );
buf ( n372802 , n25197 );
buf ( n372803 , n372802 );
nand ( n25200 , n25194 , n372803 );
buf ( n372805 , n25200 );
buf ( n372806 , n372805 );
buf ( n372807 , n4443 );
nand ( n25204 , n372806 , n372807 );
buf ( n372809 , n25204 );
nand ( n25206 , n25188 , n372809 );
buf ( n372811 , n25206 );
xor ( n25208 , n372784 , n372811 );
xor ( n25209 , n372695 , n372720 );
and ( n25210 , n25209 , n372738 );
and ( n25211 , n372695 , n372720 );
or ( n25212 , n25210 , n25211 );
buf ( n372817 , n25212 );
buf ( n372818 , n372817 );
not ( n25215 , n372753 );
not ( n25216 , n372772 );
or ( n25217 , n25215 , n25216 );
buf ( n372822 , n357712 );
buf ( n372823 , n596 );
nor ( n25220 , n372822 , n372823 );
buf ( n372825 , n25220 );
and ( n25222 , n354053 , n372825 );
not ( n25223 , n354053 );
buf ( n372828 , n357712 );
buf ( n372829 , n348865 );
nor ( n25226 , n372828 , n372829 );
buf ( n372831 , n25226 );
and ( n25228 , n25223 , n372831 );
nor ( n25229 , n25222 , n25228 );
nand ( n25230 , n25217 , n25229 );
buf ( n372835 , n25230 );
xor ( n25232 , n372818 , n372835 );
buf ( n372837 , n352101 );
buf ( n372838 , n592 );
and ( n25235 , n372837 , n372838 );
buf ( n372840 , n25235 );
buf ( n372841 , n372840 );
buf ( n372842 , n348946 );
not ( n25239 , n372842 );
buf ( n372844 , n592 );
not ( n25241 , n372844 );
buf ( n372846 , n351901 );
not ( n25243 , n372846 );
or ( n25244 , n25241 , n25243 );
buf ( n372849 , n4221 );
buf ( n372850 , n348910 );
nand ( n25247 , n372849 , n372850 );
buf ( n372852 , n25247 );
buf ( n372853 , n372852 );
nand ( n25250 , n25244 , n372853 );
buf ( n372855 , n25250 );
buf ( n372856 , n372855 );
not ( n25253 , n372856 );
or ( n25254 , n25239 , n25253 );
buf ( n372859 , n372709 );
buf ( n372860 , n1250 );
nand ( n25257 , n372859 , n372860 );
buf ( n372862 , n25257 );
buf ( n372863 , n372862 );
nand ( n25260 , n25254 , n372863 );
buf ( n372865 , n25260 );
buf ( n372866 , n372865 );
xor ( n25263 , n372841 , n372866 );
buf ( n372868 , n1335 );
buf ( n372869 , n594 );
nor ( n25266 , n372868 , n372869 );
buf ( n372871 , n25266 );
nand ( n25268 , n372871 , n6458 );
buf ( n372873 , n25123 );
buf ( n372874 , n1397 );
nand ( n25271 , n372873 , n372874 );
buf ( n372876 , n25271 );
buf ( n372877 , n1335 );
buf ( n372878 , n348975 );
nor ( n25275 , n372877 , n372878 );
buf ( n372880 , n25275 );
nand ( n25277 , n10617 , n372880 );
nand ( n25278 , n25268 , n372876 , n25277 );
buf ( n372883 , n25278 );
xor ( n25280 , n25263 , n372883 );
buf ( n372885 , n25280 );
buf ( n372886 , n372885 );
xor ( n25283 , n25232 , n372886 );
buf ( n372888 , n25283 );
buf ( n372889 , n372888 );
and ( n25286 , n25208 , n372889 );
and ( n25287 , n372784 , n372811 );
or ( n25288 , n25286 , n25287 );
buf ( n372893 , n25288 );
buf ( n372894 , n372893 );
xor ( n25291 , n372603 , n372894 );
xor ( n25292 , n372818 , n372835 );
and ( n25293 , n25292 , n372886 );
and ( n25294 , n372818 , n372835 );
or ( n25295 , n25293 , n25294 );
buf ( n372900 , n25295 );
buf ( n372901 , n372900 );
not ( n25298 , n4443 );
not ( n25299 , n25186 );
or ( n25300 , n25298 , n25299 );
nand ( n25301 , n4362 , n598 );
buf ( n372906 , n25301 );
not ( n25303 , n372906 );
buf ( n372908 , n25303 );
or ( n25305 , n372908 , n9664 );
not ( n25306 , n9661 );
not ( n25307 , n9662 );
or ( n25308 , n25306 , n25307 );
nor ( n25309 , n352112 , n598 );
not ( n25310 , n25309 );
nand ( n25311 , n25308 , n25310 );
nand ( n25312 , n25305 , n25311 );
nand ( n25313 , n25300 , n25312 );
buf ( n372918 , n25313 );
xor ( n25315 , n372901 , n372918 );
and ( n25316 , n7359 , n372825 );
not ( n25317 , n7359 );
and ( n25318 , n25317 , n372831 );
nor ( n25319 , n25316 , n25318 );
buf ( n372924 , n596 );
not ( n25321 , n372924 );
buf ( n372926 , n354056 );
not ( n25323 , n372926 );
or ( n25324 , n25321 , n25323 );
buf ( n372929 , n354053 );
buf ( n372930 , n348865 );
nand ( n25327 , n372929 , n372930 );
buf ( n372932 , n25327 );
buf ( n372933 , n372932 );
nand ( n25330 , n25324 , n372933 );
buf ( n372935 , n25330 );
buf ( n372936 , n372935 );
buf ( n372937 , n372772 );
nand ( n25334 , n372936 , n372937 );
buf ( n372939 , n25334 );
nand ( n25336 , n25319 , n372939 );
buf ( n372941 , n25336 );
xor ( n25338 , n372841 , n372866 );
and ( n25339 , n25338 , n372883 );
and ( n25340 , n372841 , n372866 );
or ( n25341 , n25339 , n25340 );
buf ( n372946 , n25341 );
buf ( n372947 , n372946 );
xor ( n25344 , n372941 , n372947 );
buf ( n372949 , n25065 );
buf ( n372950 , n592 );
and ( n25347 , n372949 , n372950 );
buf ( n372952 , n25347 );
buf ( n372953 , n372952 );
buf ( n372954 , n348946 );
not ( n25351 , n372954 );
not ( n25352 , n4179 );
xor ( n25353 , n592 , n25352 );
buf ( n372958 , n25353 );
not ( n25355 , n372958 );
or ( n25356 , n25351 , n25355 );
buf ( n372961 , n372855 );
buf ( n372962 , n1250 );
nand ( n25359 , n372961 , n372962 );
buf ( n372964 , n25359 );
buf ( n372965 , n372964 );
nand ( n25362 , n25356 , n372965 );
buf ( n372967 , n25362 );
buf ( n372968 , n372967 );
xor ( n25365 , n372953 , n372968 );
buf ( n372970 , n349035 );
not ( n25367 , n372970 );
buf ( n372972 , n594 );
not ( n25369 , n372972 );
buf ( n372974 , n354087 );
not ( n25371 , n372974 );
or ( n25372 , n25369 , n25371 );
buf ( n372977 , n9814 );
buf ( n372978 , n348975 );
nand ( n25375 , n372977 , n372978 );
buf ( n372980 , n25375 );
buf ( n372981 , n372980 );
nand ( n25378 , n25372 , n372981 );
buf ( n372983 , n25378 );
buf ( n372984 , n372983 );
not ( n25381 , n372984 );
or ( n25382 , n25367 , n25381 );
buf ( n372987 , n6458 );
buf ( n372988 , n349153 );
and ( n25385 , n372987 , n372988 );
buf ( n372990 , n355178 );
buf ( n372991 , n349163 );
and ( n25388 , n372990 , n372991 );
nor ( n25389 , n25385 , n25388 );
buf ( n372994 , n25389 );
buf ( n372995 , n372994 );
nand ( n25392 , n25382 , n372995 );
buf ( n372997 , n25392 );
buf ( n372998 , n372997 );
xor ( n25395 , n25365 , n372998 );
buf ( n373000 , n25395 );
buf ( n373001 , n373000 );
xor ( n25398 , n25344 , n373001 );
buf ( n373003 , n25398 );
buf ( n373004 , n373003 );
xor ( n25401 , n25315 , n373004 );
buf ( n373006 , n25401 );
buf ( n373007 , n373006 );
and ( n25404 , n25291 , n373007 );
and ( n25405 , n372603 , n372894 );
or ( n25406 , n25404 , n25405 );
buf ( n373011 , n25406 );
buf ( n373012 , n373011 );
buf ( n373013 , n351924 );
not ( n25410 , n373013 );
and ( n25411 , n600 , n357355 );
not ( n25412 , n600 );
and ( n25413 , n25412 , n9664 );
or ( n25414 , n25411 , n25413 );
buf ( n373019 , n25414 );
not ( n25416 , n373019 );
or ( n25417 , n25410 , n25416 );
buf ( n373022 , n600 );
not ( n25419 , n373022 );
not ( n25420 , n9635 );
buf ( n373025 , n25420 );
not ( n25422 , n373025 );
or ( n25423 , n25419 , n25422 );
buf ( n373028 , n9635 );
buf ( n373029 , n6460 );
nand ( n25426 , n373028 , n373029 );
buf ( n373031 , n25426 );
buf ( n373032 , n373031 );
nand ( n25429 , n25423 , n373032 );
buf ( n373034 , n25429 );
buf ( n373035 , n373034 );
buf ( n373036 , n1722 );
nand ( n25433 , n373035 , n373036 );
buf ( n373038 , n25433 );
buf ( n373039 , n373038 );
nand ( n25436 , n25417 , n373039 );
buf ( n373041 , n25436 );
buf ( n373042 , n373041 );
and ( n25439 , n359430 , n359432 );
buf ( n373044 , n25439 );
buf ( n373045 , n373044 );
buf ( n373046 , n348946 );
not ( n25443 , n373046 );
buf ( n373048 , n372637 );
not ( n25445 , n373048 );
or ( n25446 , n25443 , n25445 );
buf ( n373051 , n592 );
not ( n25448 , n373051 );
buf ( n373053 , n348858 );
not ( n25450 , n373053 );
or ( n25451 , n25448 , n25450 );
buf ( n373056 , n348855 );
buf ( n373057 , n348910 );
nand ( n25454 , n373056 , n373057 );
buf ( n373059 , n25454 );
buf ( n373060 , n373059 );
nand ( n25457 , n25451 , n373060 );
buf ( n373062 , n25457 );
buf ( n373063 , n373062 );
buf ( n373064 , n1250 );
nand ( n25461 , n373063 , n373064 );
buf ( n373066 , n25461 );
buf ( n373067 , n373066 );
nand ( n25464 , n25446 , n373067 );
buf ( n373069 , n25464 );
buf ( n373070 , n373069 );
xor ( n25467 , n373045 , n373070 );
buf ( n373072 , n349035 );
not ( n25469 , n373072 );
buf ( n373074 , n372676 );
not ( n25471 , n373074 );
or ( n25472 , n25469 , n25471 );
buf ( n373077 , n594 );
not ( n25474 , n373077 );
buf ( n373079 , n354248 );
not ( n25476 , n373079 );
or ( n25477 , n25474 , n25476 );
buf ( n373082 , n348975 );
buf ( n373083 , n6561 );
nand ( n25480 , n373082 , n373083 );
buf ( n373085 , n25480 );
buf ( n373086 , n373085 );
nand ( n25483 , n25477 , n373086 );
buf ( n373088 , n25483 );
buf ( n373089 , n373088 );
buf ( n373090 , n1397 );
nand ( n25487 , n373089 , n373090 );
buf ( n373092 , n25487 );
buf ( n373093 , n373092 );
nand ( n25490 , n25472 , n373093 );
buf ( n373095 , n25490 );
buf ( n373096 , n373095 );
and ( n25493 , n25467 , n373096 );
and ( n25494 , n373045 , n373070 );
or ( n25495 , n25493 , n25494 );
buf ( n373100 , n25495 );
buf ( n373101 , n373100 );
xor ( n25498 , n372608 , n372645 );
xor ( n25499 , n25498 , n372684 );
buf ( n373104 , n25499 );
buf ( n373105 , n373104 );
xor ( n25502 , n373101 , n373105 );
buf ( n373107 , n347319 );
not ( n25504 , n373107 );
buf ( n373109 , n372768 );
not ( n25506 , n373109 );
or ( n25507 , n25504 , n25506 );
and ( n25508 , n4183 , n348865 );
not ( n25509 , n4183 );
and ( n25510 , n25509 , n596 );
or ( n25511 , n25508 , n25510 );
buf ( n373116 , n25511 );
buf ( n373117 , n372772 );
nand ( n25514 , n373116 , n373117 );
buf ( n373119 , n25514 );
buf ( n373120 , n373119 );
nand ( n25517 , n25507 , n373120 );
buf ( n373122 , n25517 );
buf ( n373123 , n373122 );
and ( n25520 , n25502 , n373123 );
and ( n25521 , n373101 , n373105 );
or ( n25522 , n25520 , n25521 );
buf ( n373127 , n25522 );
buf ( n373128 , n373127 );
buf ( n373129 , n4362 );
not ( n25526 , n373129 );
buf ( n373131 , n372805 );
not ( n25528 , n373131 );
or ( n25529 , n25526 , n25528 );
buf ( n373134 , n598 );
not ( n25531 , n373134 );
buf ( n373136 , n354056 );
not ( n25533 , n373136 );
or ( n25534 , n25531 , n25533 );
buf ( n373139 , n354053 );
buf ( n373140 , n347312 );
nand ( n25537 , n373139 , n373140 );
buf ( n373142 , n25537 );
buf ( n373143 , n373142 );
nand ( n25540 , n25534 , n373143 );
buf ( n373145 , n25540 );
buf ( n373146 , n373145 );
buf ( n373147 , n4443 );
nand ( n25544 , n373146 , n373147 );
buf ( n373149 , n25544 );
buf ( n373150 , n373149 );
nand ( n25547 , n25529 , n373150 );
buf ( n373152 , n25547 );
buf ( n373153 , n373152 );
xor ( n25550 , n373128 , n373153 );
xor ( n25551 , n372689 , n372741 );
xor ( n25552 , n25551 , n372779 );
buf ( n373157 , n25552 );
buf ( n373158 , n373157 );
and ( n25555 , n25550 , n373158 );
and ( n25556 , n373128 , n373153 );
or ( n25557 , n25555 , n25556 );
buf ( n373162 , n25557 );
buf ( n373163 , n373162 );
xor ( n25560 , n373042 , n373163 );
not ( n25561 , n17020 );
not ( n25562 , n17022 );
and ( n25563 , n25561 , n25562 );
and ( n25564 , n17022 , n17020 );
nor ( n25565 , n25563 , n25564 );
not ( n25566 , n25565 );
buf ( n373171 , n25566 );
not ( n25568 , n373171 );
buf ( n373173 , n4464 );
buf ( n373174 , n349406 );
nor ( n25571 , n373173 , n373174 );
buf ( n373176 , n25571 );
buf ( n373177 , n373176 );
not ( n25574 , n373177 );
buf ( n373179 , n25574 );
buf ( n373180 , n373179 );
not ( n25577 , n373180 );
and ( n25578 , n25568 , n25577 );
buf ( n373183 , n25566 );
buf ( n373184 , n352149 );
buf ( n373185 , n349406 );
and ( n25582 , n373184 , n373185 );
buf ( n373187 , n25582 );
buf ( n373188 , n373187 );
and ( n25585 , n373183 , n373188 );
nor ( n25586 , n25578 , n25585 );
buf ( n373191 , n25586 );
buf ( n373192 , n373191 );
buf ( n373193 , n602 );
not ( n25590 , n373193 );
buf ( n373195 , n360099 );
not ( n25592 , n373195 );
or ( n25593 , n25590 , n25592 );
buf ( n373198 , n12420 );
buf ( n373199 , n349406 );
nand ( n25596 , n373198 , n373199 );
buf ( n373201 , n25596 );
buf ( n373202 , n373201 );
nand ( n25599 , n25593 , n373202 );
buf ( n373204 , n25599 );
buf ( n373205 , n373204 );
buf ( n373206 , n354113 );
nand ( n25603 , n373205 , n373206 );
buf ( n373208 , n25603 );
buf ( n373209 , n373208 );
nand ( n25606 , n373192 , n373209 );
buf ( n373211 , n25606 );
buf ( n373212 , n373211 );
and ( n25609 , n25560 , n373212 );
and ( n25610 , n373042 , n373163 );
or ( n25611 , n25609 , n25610 );
buf ( n373216 , n25611 );
buf ( n373217 , n373216 );
buf ( n373218 , n25566 );
not ( n25615 , n373218 );
buf ( n373220 , n358424 );
nand ( n25617 , n25615 , n373220 );
buf ( n373222 , n25617 );
buf ( n373223 , n25566 );
buf ( n373224 , n358417 );
nand ( n25621 , n373223 , n373224 );
buf ( n373226 , n25621 );
and ( n25623 , n17023 , n366657 );
not ( n25624 , n17023 );
and ( n25625 , n25624 , n366654 );
nor ( n25626 , n25623 , n25625 );
buf ( n25627 , n25626 );
buf ( n373232 , n25627 );
not ( n25629 , n373232 );
buf ( n373234 , n25629 );
buf ( n373235 , n373234 );
buf ( n373236 , n373176 );
nand ( n25633 , n373235 , n373236 );
buf ( n373238 , n25633 );
buf ( n373239 , n25627 );
buf ( n373240 , n373187 );
nand ( n25637 , n373239 , n373240 );
buf ( n373242 , n25637 );
nand ( n25639 , n373222 , n373226 , n373238 , n373242 );
buf ( n373244 , n25639 );
not ( n25641 , n373034 );
not ( n25642 , n351924 );
or ( n25643 , n25641 , n25642 );
buf ( n373248 , n358041 );
buf ( n373249 , n600 );
nor ( n25646 , n373248 , n373249 );
buf ( n373251 , n25646 );
and ( n25648 , n360105 , n373251 );
not ( n25649 , n360105 );
buf ( n373254 , n358041 );
buf ( n373255 , n6460 );
nor ( n25652 , n373254 , n373255 );
buf ( n373257 , n25652 );
and ( n25654 , n25649 , n373257 );
nor ( n25655 , n25648 , n25654 );
nand ( n25656 , n25643 , n25655 );
buf ( n373261 , n25656 );
xor ( n25658 , n373244 , n373261 );
not ( n25659 , n355075 );
not ( n25660 , n604 );
buf ( n373265 , n25660 );
not ( n25662 , n373265 );
not ( n25663 , n13074 );
nand ( n25664 , n25663 , n17017 );
not ( n25665 , n25664 );
nor ( n25666 , n8326 , n17031 );
nand ( n25667 , n25665 , n25666 );
and ( n25668 , n25667 , n17025 );
not ( n25669 , n25667 );
and ( n25670 , n25669 , n17026 );
nor ( n25671 , n25668 , n25670 );
buf ( n25672 , n25671 );
buf ( n373277 , n25672 );
not ( n25674 , n373277 );
or ( n25675 , n25662 , n25674 );
not ( n25676 , n25671 );
buf ( n373281 , n25676 );
not ( n25678 , n373281 );
buf ( n373283 , n25678 );
buf ( n373284 , n373283 );
not ( n25681 , n373284 );
buf ( n373286 , n604 );
nand ( n25683 , n25681 , n373286 );
buf ( n373288 , n25683 );
buf ( n373289 , n373288 );
nand ( n25686 , n25675 , n373289 );
buf ( n373291 , n25686 );
not ( n25688 , n373291 );
or ( n25689 , n25659 , n25688 );
not ( n25690 , n11145 );
not ( n25691 , n17018 );
not ( n25692 , n17028 );
nand ( n25693 , n25691 , n25692 , n17026 , n8327 );
not ( n25694 , n17024 );
and ( n25695 , n25693 , n25694 );
not ( n25696 , n25693 );
buf ( n25697 , n17519 );
and ( n25698 , n25696 , n25697 );
nor ( n25699 , n25695 , n25698 );
buf ( n25700 , n25699 );
not ( n25701 , n25700 );
or ( n25702 , n25690 , n25701 );
not ( n25703 , n25700 );
not ( n25704 , n25703 );
or ( n25705 , n25704 , n11145 );
nand ( n25706 , n25702 , n25705 );
nand ( n25707 , n25706 , n6599 );
nand ( n25708 , n25689 , n25707 );
buf ( n373313 , n25708 );
xor ( n25710 , n25658 , n373313 );
buf ( n373315 , n25710 );
buf ( n373316 , n373315 );
xor ( n25713 , n373217 , n373316 );
buf ( n373318 , n355075 );
not ( n25715 , n373318 );
buf ( n373320 , n25627 );
not ( n25717 , n373320 );
buf ( n373322 , n25717 );
and ( n25719 , n604 , n373322 );
not ( n25720 , n604 );
and ( n25721 , n25720 , n25627 );
or ( n25722 , n25719 , n25721 );
buf ( n373327 , n25722 );
not ( n25724 , n373327 );
or ( n25725 , n25715 , n25724 );
buf ( n373330 , n373291 );
buf ( n373331 , n6600 );
nand ( n25728 , n373330 , n373331 );
buf ( n373333 , n25728 );
buf ( n373334 , n373333 );
nand ( n25731 , n25725 , n373334 );
buf ( n373336 , n25731 );
buf ( n373337 , n373336 );
buf ( n373338 , n607 );
not ( n25735 , n373338 );
buf ( n373340 , n372566 );
not ( n25737 , n373340 );
or ( n25738 , n25735 , n25737 );
buf ( n373343 , n606 );
not ( n25740 , n373343 );
not ( n25741 , n25700 );
buf ( n373346 , n25741 );
not ( n25743 , n373346 );
or ( n25744 , n25740 , n25743 );
buf ( n373349 , n25700 );
buf ( n373350 , n9642 );
nand ( n25747 , n373349 , n373350 );
buf ( n373352 , n25747 );
buf ( n373353 , n373352 );
nand ( n25750 , n25744 , n373353 );
buf ( n373355 , n25750 );
buf ( n373356 , n373355 );
buf ( n373357 , n357376 );
nand ( n25754 , n373356 , n373357 );
buf ( n373359 , n25754 );
buf ( n373360 , n373359 );
nand ( n25757 , n25738 , n373360 );
buf ( n373362 , n25757 );
buf ( n373363 , n373362 );
xor ( n25760 , n373337 , n373363 );
xor ( n25761 , n372784 , n372811 );
xor ( n25762 , n25761 , n372889 );
buf ( n373367 , n25762 );
buf ( n373368 , n373367 );
and ( n25765 , n25760 , n373368 );
and ( n25766 , n373337 , n373363 );
or ( n25767 , n25765 , n25766 );
buf ( n373372 , n25767 );
buf ( n373373 , n373372 );
and ( n25770 , n25713 , n373373 );
and ( n25771 , n373217 , n373316 );
or ( n25772 , n25770 , n25771 );
buf ( n373377 , n25772 );
buf ( n373378 , n373377 );
xor ( n25775 , n373012 , n373378 );
xor ( n25776 , n372941 , n372947 );
and ( n25777 , n25776 , n373001 );
and ( n25778 , n372941 , n372947 );
or ( n25779 , n25777 , n25778 );
buf ( n373384 , n25779 );
buf ( n373385 , n373384 );
not ( n25782 , n4362 );
not ( n25783 , n598 );
not ( n25784 , n9635 );
not ( n25785 , n25784 );
or ( n25786 , n25783 , n25785 );
buf ( n373391 , n9635 );
buf ( n373392 , n347312 );
nand ( n25789 , n373391 , n373392 );
buf ( n373394 , n25789 );
nand ( n25791 , n25786 , n373394 );
not ( n25792 , n25791 );
or ( n25793 , n25782 , n25792 );
buf ( n373398 , n9664 );
not ( n25795 , n373398 );
buf ( n373400 , n357731 );
not ( n25797 , n373400 );
and ( n25798 , n25795 , n25797 );
buf ( n373403 , n9664 );
buf ( n373404 , n357742 );
and ( n25801 , n373403 , n373404 );
nor ( n25802 , n25798 , n25801 );
buf ( n373407 , n25802 );
nand ( n25804 , n25793 , n373407 );
buf ( n373409 , n25804 );
xor ( n25806 , n373385 , n373409 );
buf ( n373411 , n9751 );
not ( n25808 , n373411 );
buf ( n373413 , n600 );
not ( n25810 , n373413 );
buf ( n25811 , n25565 );
buf ( n373416 , n25811 );
not ( n25813 , n373416 );
or ( n25814 , n25810 , n25813 );
buf ( n373419 , n25566 );
buf ( n373420 , n6460 );
nand ( n25817 , n373419 , n373420 );
buf ( n373422 , n25817 );
buf ( n373423 , n373422 );
nand ( n25820 , n25814 , n373423 );
buf ( n373425 , n25820 );
buf ( n373426 , n373425 );
not ( n25823 , n373426 );
or ( n25824 , n25808 , n25823 );
buf ( n373429 , n360105 );
not ( n25826 , n373429 );
buf ( n373431 , n358062 );
not ( n25828 , n373431 );
and ( n25829 , n25826 , n25828 );
buf ( n373434 , n360105 );
buf ( n373435 , n358055 );
and ( n25832 , n373434 , n373435 );
nor ( n25833 , n25829 , n25832 );
buf ( n373438 , n25833 );
buf ( n373439 , n373438 );
nand ( n25836 , n25824 , n373439 );
buf ( n373441 , n25836 );
buf ( n373442 , n373441 );
xor ( n25839 , n25806 , n373442 );
buf ( n373444 , n25839 );
buf ( n373445 , n373444 );
buf ( n373446 , n352149 );
not ( n25843 , n373446 );
buf ( n373448 , n602 );
not ( n25845 , n373448 );
buf ( n373450 , n25676 );
not ( n25847 , n373450 );
or ( n25848 , n25845 , n25847 );
buf ( n373453 , n25672 );
buf ( n373454 , n349406 );
nand ( n25851 , n373453 , n373454 );
buf ( n373456 , n25851 );
buf ( n373457 , n373456 );
nand ( n25854 , n25848 , n373457 );
buf ( n373459 , n25854 );
buf ( n373460 , n373459 );
not ( n25857 , n373460 );
or ( n25858 , n25843 , n25857 );
buf ( n373463 , n358424 );
not ( n25860 , n373463 );
buf ( n373465 , n25860 );
not ( n25862 , n373465 );
not ( n25863 , n25627 );
not ( n25864 , n25863 );
or ( n25865 , n25862 , n25864 );
not ( n25866 , n25627 );
or ( n25867 , n25866 , n358417 );
nand ( n25868 , n25865 , n25867 );
buf ( n373473 , n25868 );
nand ( n25870 , n25858 , n373473 );
buf ( n373475 , n25870 );
buf ( n373476 , n373475 );
not ( n25873 , n6598 );
not ( n25874 , n604 );
not ( n25875 , n372556 );
or ( n25876 , n25874 , n25875 );
nand ( n25877 , n24943 , n25660 );
nand ( n25878 , n25876 , n25877 );
not ( n25879 , n25878 );
or ( n25880 , n25873 , n25879 );
nand ( n25881 , n25706 , n355075 );
nand ( n25882 , n25880 , n25881 );
buf ( n373487 , n25882 );
xor ( n25884 , n373476 , n373487 );
not ( n25885 , n607 );
buf ( n373490 , n606 );
not ( n25887 , n373490 );
buf ( n373492 , n17009 );
not ( n25889 , n373492 );
buf ( n373494 , n25889 );
buf ( n373495 , n373494 );
not ( n25892 , n373495 );
or ( n25893 , n25887 , n25892 );
buf ( n373498 , n17009 );
buf ( n373499 , n9642 );
nand ( n25896 , n373498 , n373499 );
buf ( n373501 , n25896 );
buf ( n373502 , n373501 );
nand ( n25899 , n25893 , n373502 );
buf ( n373504 , n25899 );
not ( n25901 , n373504 );
or ( n25902 , n25885 , n25901 );
nand ( n25903 , n372595 , n357376 );
nand ( n25904 , n25902 , n25903 );
buf ( n373509 , n25904 );
xor ( n25906 , n25884 , n373509 );
buf ( n373511 , n25906 );
buf ( n373512 , n373511 );
xor ( n25909 , n373445 , n373512 );
xor ( n25910 , n372953 , n372968 );
and ( n25911 , n25910 , n372998 );
and ( n25912 , n372953 , n372968 );
or ( n25913 , n25911 , n25912 );
buf ( n373518 , n25913 );
buf ( n373519 , n373518 );
buf ( n373520 , n4221 );
buf ( n373521 , n592 );
and ( n25918 , n373520 , n373521 );
buf ( n373523 , n25918 );
buf ( n373524 , n373523 );
buf ( n373525 , n348946 );
not ( n25922 , n373525 );
buf ( n373527 , n592 );
not ( n25924 , n373527 );
buf ( n373529 , n355178 );
not ( n25926 , n373529 );
or ( n25927 , n25924 , n25926 );
buf ( n373532 , n6458 );
buf ( n373533 , n348910 );
nand ( n25930 , n373532 , n373533 );
buf ( n373535 , n25930 );
buf ( n373536 , n373535 );
nand ( n25933 , n25927 , n373536 );
buf ( n373538 , n25933 );
buf ( n373539 , n373538 );
not ( n25936 , n373539 );
or ( n25937 , n25922 , n25936 );
buf ( n373542 , n25353 );
buf ( n373543 , n1250 );
nand ( n25940 , n373542 , n373543 );
buf ( n373545 , n25940 );
buf ( n373546 , n373545 );
nand ( n25943 , n25937 , n373546 );
buf ( n373548 , n25943 );
buf ( n373549 , n373548 );
xor ( n25946 , n373524 , n373549 );
buf ( n373551 , n349035 );
not ( n25948 , n373551 );
and ( n25949 , n594 , n354056 );
not ( n25950 , n594 );
and ( n25951 , n25950 , n354053 );
or ( n25952 , n25949 , n25951 );
buf ( n373557 , n25952 );
not ( n25954 , n373557 );
or ( n25955 , n25948 , n25954 );
buf ( n373560 , n372983 );
buf ( n373561 , n1397 );
nand ( n25958 , n373560 , n373561 );
buf ( n373563 , n25958 );
buf ( n373564 , n373563 );
nand ( n25961 , n25955 , n373564 );
buf ( n373566 , n25961 );
buf ( n373567 , n373566 );
xor ( n25964 , n25946 , n373567 );
buf ( n373569 , n25964 );
buf ( n373570 , n373569 );
xor ( n25967 , n373519 , n373570 );
not ( n25968 , n347319 );
not ( n25969 , n596 );
not ( n25970 , n9708 );
or ( n25971 , n25969 , n25970 );
buf ( n373576 , n8333 );
buf ( n373577 , n348865 );
nand ( n25974 , n373576 , n373577 );
buf ( n373579 , n25974 );
nand ( n25976 , n25971 , n373579 );
not ( n25977 , n25976 );
or ( n25978 , n25968 , n25977 );
and ( n25979 , n7359 , n1651 );
not ( n25980 , n7359 );
and ( n25981 , n25980 , n1649 );
nor ( n25982 , n25979 , n25981 );
nand ( n25983 , n25978 , n25982 );
buf ( n373588 , n25983 );
xor ( n25985 , n25967 , n373588 );
buf ( n373590 , n25985 );
buf ( n373591 , n373590 );
xor ( n25988 , n372901 , n372918 );
and ( n25989 , n25988 , n373004 );
and ( n25990 , n372901 , n372918 );
or ( n25991 , n25989 , n25990 );
buf ( n373596 , n25991 );
buf ( n373597 , n373596 );
xor ( n25994 , n373591 , n373597 );
xor ( n25995 , n373244 , n373261 );
and ( n25996 , n25995 , n373313 );
and ( n25997 , n373244 , n373261 );
or ( n25998 , n25996 , n25997 );
buf ( n373603 , n25998 );
buf ( n373604 , n373603 );
xor ( n26001 , n25994 , n373604 );
buf ( n373606 , n26001 );
buf ( n373607 , n373606 );
xor ( n26004 , n25909 , n373607 );
buf ( n373609 , n26004 );
buf ( n373610 , n373609 );
xor ( n26007 , n25775 , n373610 );
buf ( n373612 , n26007 );
buf ( n373613 , n373612 );
not ( n26010 , n373613 );
buf ( n373615 , n26010 );
buf ( n373616 , n373615 );
buf ( n373617 , n347319 );
not ( n26014 , n373617 );
and ( n26015 , n4183 , n348865 );
not ( n26016 , n4183 );
and ( n26017 , n26016 , n596 );
or ( n26018 , n26015 , n26017 );
buf ( n373623 , n26018 );
not ( n26020 , n373623 );
or ( n26021 , n26014 , n26020 );
buf ( n373626 , n596 );
not ( n26023 , n373626 );
buf ( n373628 , n351901 );
not ( n26025 , n373628 );
or ( n26026 , n26023 , n26025 );
buf ( n373631 , n4221 );
buf ( n373632 , n348865 );
nand ( n26029 , n373631 , n373632 );
buf ( n373634 , n26029 );
buf ( n373635 , n373634 );
nand ( n26032 , n26026 , n373635 );
buf ( n373637 , n26032 );
buf ( n373638 , n373637 );
buf ( n373639 , n348898 );
nand ( n26036 , n373638 , n373639 );
buf ( n373641 , n26036 );
buf ( n373642 , n373641 );
nand ( n26039 , n26021 , n373642 );
buf ( n373644 , n26039 );
buf ( n373645 , n373644 );
buf ( n373646 , n354213 );
not ( n26043 , n373646 );
buf ( n373648 , n348910 );
nor ( n26045 , n26043 , n373648 );
buf ( n373650 , n26045 );
buf ( n373651 , n373650 );
buf ( n373652 , n348946 );
not ( n26049 , n373652 );
buf ( n373654 , n373062 );
not ( n26051 , n373654 );
or ( n26052 , n26049 , n26051 );
buf ( n373657 , n359434 );
buf ( n373658 , n1250 );
nand ( n26055 , n373657 , n373658 );
buf ( n373660 , n26055 );
buf ( n373661 , n373660 );
nand ( n26058 , n26052 , n373661 );
buf ( n373663 , n26058 );
buf ( n373664 , n373663 );
xor ( n26061 , n373651 , n373664 );
not ( n26062 , n349035 );
not ( n26063 , n373088 );
or ( n26064 , n26062 , n26063 );
not ( n26065 , n1396 );
nand ( n26066 , n26065 , n11738 );
nand ( n26067 , n26064 , n26066 );
buf ( n373672 , n26067 );
and ( n26069 , n26061 , n373672 );
and ( n26070 , n373651 , n373664 );
or ( n26071 , n26069 , n26070 );
buf ( n373676 , n26071 );
buf ( n373677 , n373676 );
xor ( n26074 , n373645 , n373677 );
xor ( n26075 , n373045 , n373070 );
xor ( n26076 , n26075 , n373096 );
buf ( n373681 , n26076 );
buf ( n373682 , n373681 );
and ( n26079 , n26074 , n373682 );
and ( n26080 , n373645 , n373677 );
or ( n26081 , n26079 , n26080 );
buf ( n373686 , n26081 );
buf ( n373687 , n373686 );
buf ( n373688 , n4362 );
not ( n26085 , n373688 );
buf ( n373690 , n373145 );
not ( n26087 , n373690 );
or ( n26088 , n26085 , n26087 );
and ( n26089 , n598 , n354087 );
not ( n26090 , n598 );
and ( n26091 , n26090 , n9814 );
or ( n26092 , n26089 , n26091 );
buf ( n373697 , n26092 );
buf ( n373698 , n4443 );
nand ( n26095 , n373697 , n373698 );
buf ( n373700 , n26095 );
buf ( n373701 , n373700 );
nand ( n26098 , n26088 , n373701 );
buf ( n373703 , n26098 );
buf ( n373704 , n373703 );
xor ( n26101 , n373687 , n373704 );
xor ( n26102 , n373101 , n373105 );
xor ( n26103 , n26102 , n373123 );
buf ( n373708 , n26103 );
buf ( n373709 , n373708 );
and ( n26106 , n26101 , n373709 );
and ( n26107 , n373687 , n373704 );
or ( n26108 , n26106 , n26107 );
buf ( n373713 , n26108 );
buf ( n373714 , n373713 );
buf ( n373715 , n9751 );
not ( n26112 , n373715 );
buf ( n373717 , n25414 );
not ( n26114 , n373717 );
or ( n26115 , n26112 , n26114 );
not ( n26116 , n8333 );
not ( n26117 , n600 );
not ( n26118 , n26117 );
or ( n26119 , n26116 , n26118 );
nand ( n26120 , n8330 , n600 );
nand ( n26121 , n26119 , n26120 );
buf ( n373726 , n26121 );
buf ( n373727 , n351924 );
nand ( n26124 , n373726 , n373727 );
buf ( n373729 , n26124 );
buf ( n373730 , n373729 );
nand ( n26127 , n26115 , n373730 );
buf ( n373732 , n26127 );
buf ( n373733 , n373732 );
xor ( n26130 , n373714 , n373733 );
xor ( n26131 , n373128 , n373153 );
xor ( n26132 , n26131 , n373158 );
buf ( n373737 , n26132 );
buf ( n373738 , n373737 );
and ( n26135 , n26130 , n373738 );
and ( n26136 , n373714 , n373733 );
or ( n26137 , n26135 , n26136 );
buf ( n373742 , n26137 );
buf ( n373743 , n373742 );
xor ( n26140 , n373042 , n373163 );
xor ( n26141 , n26140 , n373212 );
buf ( n373746 , n26141 );
buf ( n373747 , n373746 );
xor ( n26144 , n373743 , n373747 );
buf ( n373749 , n354113 );
not ( n26146 , n373749 );
buf ( n373751 , n602 );
not ( n26148 , n373751 );
buf ( n373753 , n25784 );
not ( n26150 , n373753 );
or ( n26151 , n26148 , n26150 );
buf ( n373756 , n9635 );
buf ( n373757 , n349406 );
nand ( n26154 , n373756 , n373757 );
buf ( n373759 , n26154 );
buf ( n373760 , n373759 );
nand ( n26157 , n26151 , n373760 );
buf ( n373762 , n26157 );
buf ( n373763 , n373762 );
not ( n26160 , n373763 );
or ( n26161 , n26146 , n26160 );
buf ( n373766 , n373204 );
buf ( n373767 , n352149 );
nand ( n26164 , n373766 , n373767 );
buf ( n373769 , n26164 );
buf ( n373770 , n373769 );
nand ( n26167 , n26161 , n373770 );
buf ( n373772 , n26167 );
buf ( n373773 , n373772 );
buf ( n373774 , n357376 );
not ( n26171 , n373774 );
buf ( n373776 , n9642 );
not ( n26173 , n373776 );
buf ( n373778 , n25672 );
not ( n26175 , n373778 );
or ( n26176 , n26173 , n26175 );
buf ( n373781 , n25676 );
buf ( n373782 , n606 );
nand ( n26179 , n373781 , n373782 );
buf ( n373784 , n26179 );
buf ( n373785 , n373784 );
nand ( n26182 , n26176 , n373785 );
buf ( n373787 , n26182 );
buf ( n373788 , n373787 );
not ( n26185 , n373788 );
or ( n26186 , n26171 , n26185 );
buf ( n373791 , n373355 );
buf ( n373792 , n607 );
nand ( n26189 , n373791 , n373792 );
buf ( n373794 , n26189 );
buf ( n373795 , n373794 );
nand ( n26192 , n26186 , n373795 );
buf ( n373797 , n26192 );
buf ( n373798 , n373797 );
xor ( n26195 , n373773 , n373798 );
buf ( n373800 , n355075 );
not ( n26197 , n373800 );
and ( n26198 , n604 , n25811 );
not ( n26199 , n604 );
buf ( n373804 , n25811 );
not ( n26201 , n373804 );
buf ( n373806 , n26201 );
and ( n26203 , n26199 , n373806 );
or ( n26204 , n26198 , n26203 );
buf ( n373809 , n26204 );
not ( n26206 , n373809 );
or ( n26207 , n26197 , n26206 );
buf ( n373812 , n25722 );
buf ( n373813 , n6600 );
nand ( n26210 , n373812 , n373813 );
buf ( n373815 , n26210 );
buf ( n373816 , n373815 );
nand ( n26213 , n26207 , n373816 );
buf ( n373818 , n26213 );
buf ( n373819 , n373818 );
and ( n26216 , n26195 , n373819 );
and ( n26217 , n373773 , n373798 );
or ( n26218 , n26216 , n26217 );
buf ( n373823 , n26218 );
buf ( n373824 , n373823 );
and ( n26221 , n26144 , n373824 );
and ( n26222 , n373743 , n373747 );
or ( n26223 , n26221 , n26222 );
buf ( n373828 , n26223 );
buf ( n373829 , n373828 );
xor ( n26226 , n372603 , n372894 );
xor ( n26227 , n26226 , n373007 );
buf ( n373832 , n26227 );
buf ( n373833 , n373832 );
xor ( n26230 , n373829 , n373833 );
xor ( n26231 , n373217 , n373316 );
xor ( n26232 , n26231 , n373373 );
buf ( n373837 , n26232 );
buf ( n373838 , n373837 );
and ( n26235 , n26230 , n373838 );
and ( n26236 , n373829 , n373833 );
or ( n26237 , n26235 , n26236 );
buf ( n373842 , n26237 );
buf ( n373843 , n373842 );
not ( n26240 , n373843 );
buf ( n373845 , n26240 );
buf ( n373846 , n373845 );
nand ( n26243 , n373616 , n373846 );
buf ( n373848 , n26243 );
xor ( n26245 , n373829 , n373833 );
xor ( n26246 , n26245 , n373838 );
buf ( n373851 , n26246 );
not ( n26248 , n373851 );
xor ( n26249 , n373337 , n373363 );
xor ( n26250 , n26249 , n373368 );
buf ( n373855 , n26250 );
buf ( n373856 , n373855 );
xor ( n26253 , n359427 , n359445 );
and ( n26254 , n26253 , n359452 );
and ( n26255 , n359427 , n359445 );
or ( n26256 , n26254 , n26255 );
buf ( n373861 , n26256 );
buf ( n373862 , n373861 );
buf ( n373863 , n347319 );
not ( n26260 , n373863 );
buf ( n373865 , n373637 );
not ( n26262 , n373865 );
or ( n26263 , n26260 , n26262 );
buf ( n373868 , n359470 );
buf ( n373869 , n348898 );
nand ( n26266 , n373868 , n373869 );
buf ( n373871 , n26266 );
buf ( n373872 , n373871 );
nand ( n26269 , n26263 , n373872 );
buf ( n373874 , n26269 );
buf ( n373875 , n373874 );
xor ( n26272 , n373862 , n373875 );
xor ( n26273 , n373651 , n373664 );
xor ( n26274 , n26273 , n373672 );
buf ( n373879 , n26274 );
buf ( n373880 , n373879 );
and ( n26277 , n26272 , n373880 );
and ( n26278 , n373862 , n373875 );
or ( n26279 , n26277 , n26278 );
buf ( n373884 , n26279 );
buf ( n373885 , n373884 );
buf ( n373886 , n4362 );
not ( n26283 , n373886 );
buf ( n373888 , n26092 );
not ( n26285 , n373888 );
or ( n26286 , n26283 , n26285 );
buf ( n373891 , n598 );
not ( n26288 , n373891 );
buf ( n373893 , n355178 );
not ( n26290 , n373893 );
or ( n26291 , n26288 , n26290 );
buf ( n373896 , n6458 );
buf ( n373897 , n347312 );
nand ( n26294 , n373896 , n373897 );
buf ( n373899 , n26294 );
buf ( n373900 , n373899 );
nand ( n26297 , n26291 , n373900 );
buf ( n373902 , n26297 );
buf ( n373903 , n373902 );
buf ( n373904 , n4443 );
nand ( n26301 , n373903 , n373904 );
buf ( n373906 , n26301 );
buf ( n373907 , n373906 );
nand ( n26304 , n26286 , n373907 );
buf ( n373909 , n26304 );
buf ( n373910 , n373909 );
xor ( n26307 , n373885 , n373910 );
xor ( n26308 , n373645 , n373677 );
xor ( n26309 , n26308 , n373682 );
buf ( n373914 , n26309 );
buf ( n373915 , n373914 );
and ( n26312 , n26307 , n373915 );
and ( n26313 , n373885 , n373910 );
or ( n26314 , n26312 , n26313 );
buf ( n373919 , n26314 );
buf ( n373920 , n373919 );
not ( n26317 , n9751 );
not ( n26318 , n26121 );
or ( n26319 , n26317 , n26318 );
buf ( n373924 , n600 );
not ( n26321 , n373924 );
buf ( n373926 , n25191 );
not ( n26323 , n373926 );
or ( n26324 , n26321 , n26323 );
buf ( n373929 , n7359 );
buf ( n373930 , n4193 );
nand ( n26327 , n373929 , n373930 );
buf ( n373932 , n26327 );
buf ( n373933 , n373932 );
nand ( n26330 , n26324 , n373933 );
buf ( n373935 , n26330 );
nand ( n26332 , n373935 , n351924 );
nand ( n26333 , n26319 , n26332 );
buf ( n373938 , n26333 );
xor ( n26335 , n373920 , n373938 );
xor ( n26336 , n373687 , n373704 );
xor ( n26337 , n26336 , n373709 );
buf ( n373942 , n26337 );
buf ( n373943 , n373942 );
and ( n26340 , n26335 , n373943 );
and ( n26341 , n373920 , n373938 );
or ( n26342 , n26340 , n26341 );
buf ( n373947 , n26342 );
buf ( n373948 , n373947 );
xor ( n26345 , n373714 , n373733 );
xor ( n26346 , n26345 , n373738 );
buf ( n373951 , n26346 );
buf ( n373952 , n373951 );
xor ( n26349 , n373948 , n373952 );
buf ( n373954 , n354113 );
not ( n26351 , n373954 );
buf ( n373956 , n602 );
not ( n26353 , n373956 );
buf ( n373958 , n357355 );
not ( n26355 , n373958 );
or ( n26356 , n26353 , n26355 );
buf ( n373961 , n9664 );
buf ( n373962 , n349406 );
nand ( n26359 , n373961 , n373962 );
buf ( n373964 , n26359 );
buf ( n373965 , n373964 );
nand ( n26362 , n26356 , n373965 );
buf ( n373967 , n26362 );
buf ( n373968 , n373967 );
not ( n26365 , n373968 );
or ( n26366 , n26351 , n26365 );
buf ( n373971 , n373762 );
buf ( n373972 , n352149 );
nand ( n26369 , n373971 , n373972 );
buf ( n373974 , n26369 );
buf ( n373975 , n373974 );
nand ( n26372 , n26366 , n373975 );
buf ( n373977 , n26372 );
buf ( n373978 , n373977 );
buf ( n373979 , n1722 );
not ( n26376 , n373979 );
buf ( n373981 , n373935 );
not ( n26378 , n373981 );
or ( n26379 , n26376 , n26378 );
buf ( n373984 , n354053 );
buf ( n373985 , n600 );
and ( n26382 , n373984 , n373985 );
not ( n26383 , n373984 );
buf ( n373988 , n6460 );
and ( n26385 , n26383 , n373988 );
nor ( n26386 , n26382 , n26385 );
buf ( n373991 , n26386 );
buf ( n373992 , n373991 );
buf ( n373993 , n351924 );
nand ( n26390 , n373992 , n373993 );
buf ( n373995 , n26390 );
buf ( n373996 , n373995 );
nand ( n26393 , n26379 , n373996 );
buf ( n373998 , n26393 );
buf ( n373999 , n373998 );
xor ( n26396 , n359422 , n359455 );
and ( n26397 , n26396 , n359481 );
and ( n26398 , n359422 , n359455 );
or ( n26399 , n26397 , n26398 );
buf ( n374004 , n26399 );
buf ( n374005 , n374004 );
buf ( n374006 , n4362 );
not ( n26403 , n374006 );
buf ( n374008 , n373902 );
not ( n26405 , n374008 );
or ( n26406 , n26403 , n26405 );
buf ( n374011 , n11726 );
buf ( n374012 , n4443 );
nand ( n26409 , n374011 , n374012 );
buf ( n374014 , n26409 );
buf ( n374015 , n374014 );
nand ( n26412 , n26406 , n374015 );
buf ( n374017 , n26412 );
buf ( n374018 , n374017 );
xor ( n26415 , n374005 , n374018 );
xor ( n26416 , n373862 , n373875 );
xor ( n26417 , n26416 , n373880 );
buf ( n374022 , n26417 );
buf ( n374023 , n374022 );
and ( n26420 , n26415 , n374023 );
and ( n26421 , n374005 , n374018 );
or ( n26422 , n26420 , n26421 );
buf ( n374027 , n26422 );
buf ( n374028 , n374027 );
xor ( n26425 , n373999 , n374028 );
xor ( n26426 , n373885 , n373910 );
xor ( n26427 , n26426 , n373915 );
buf ( n374032 , n26427 );
buf ( n374033 , n374032 );
and ( n26430 , n26425 , n374033 );
and ( n26431 , n373999 , n374028 );
or ( n26432 , n26430 , n26431 );
buf ( n374037 , n26432 );
buf ( n374038 , n374037 );
xor ( n26435 , n373978 , n374038 );
buf ( n374040 , n25627 );
not ( n26437 , n374040 );
buf ( n374042 , n26437 );
and ( n26439 , n9642 , n374042 );
not ( n26440 , n9642 );
buf ( n374045 , n25627 );
buf ( n26442 , n374045 );
buf ( n374047 , n26442 );
and ( n26444 , n26440 , n374047 );
nor ( n26445 , n26439 , n26444 );
not ( n26446 , n26445 );
not ( n26447 , n357376 );
or ( n26448 , n26446 , n26447 );
buf ( n374053 , n373787 );
buf ( n374054 , n607 );
nand ( n26451 , n374053 , n374054 );
buf ( n374056 , n26451 );
nand ( n26453 , n26448 , n374056 );
buf ( n374058 , n26453 );
and ( n26455 , n26435 , n374058 );
and ( n26456 , n373978 , n374038 );
or ( n26457 , n26455 , n26456 );
buf ( n374062 , n26457 );
buf ( n374063 , n374062 );
and ( n26460 , n26349 , n374063 );
and ( n26461 , n373948 , n373952 );
or ( n26462 , n26460 , n26461 );
buf ( n374067 , n26462 );
buf ( n374068 , n374067 );
xor ( n26465 , n373856 , n374068 );
xor ( n26466 , n373743 , n373747 );
xor ( n26467 , n26466 , n373824 );
buf ( n374072 , n26467 );
buf ( n374073 , n374072 );
and ( n26470 , n26465 , n374073 );
and ( n26471 , n373856 , n374068 );
or ( n26472 , n26470 , n26471 );
buf ( n374077 , n26472 );
not ( n26474 , n374077 );
nand ( n26475 , n26248 , n26474 );
nand ( n26476 , n373848 , n26475 );
not ( n26477 , n26476 );
not ( n26478 , n26477 );
xor ( n26479 , n359364 , n359386 );
and ( n26480 , n26479 , n359487 );
and ( n26481 , n359364 , n359386 );
or ( n26482 , n26480 , n26481 );
buf ( n374087 , n26482 );
buf ( n374088 , n374087 );
buf ( n374089 , n352149 );
not ( n26486 , n374089 );
buf ( n374091 , n602 );
not ( n26488 , n374091 );
buf ( n374093 , n9708 );
not ( n26490 , n374093 );
or ( n26491 , n26488 , n26490 );
buf ( n374096 , n8333 );
buf ( n374097 , n349406 );
nand ( n26494 , n374096 , n374097 );
buf ( n374099 , n26494 );
buf ( n374100 , n374099 );
nand ( n26497 , n26491 , n374100 );
buf ( n374102 , n26497 );
buf ( n374103 , n374102 );
not ( n26500 , n374103 );
or ( n26501 , n26486 , n26500 );
buf ( n374106 , n354113 );
buf ( n374107 , n359346 );
nand ( n26504 , n374106 , n374107 );
buf ( n374109 , n26504 );
buf ( n374110 , n374109 );
nand ( n26507 , n26501 , n374110 );
buf ( n374112 , n26507 );
buf ( n374113 , n374112 );
xor ( n26510 , n374088 , n374113 );
xor ( n26511 , n359393 , n359407 );
and ( n26512 , n26511 , n359484 );
and ( n26513 , n359393 , n359407 );
or ( n26514 , n26512 , n26513 );
buf ( n374119 , n26514 );
buf ( n374120 , n374119 );
buf ( n374121 , n1722 );
not ( n26518 , n374121 );
buf ( n374123 , n373991 );
not ( n26520 , n374123 );
or ( n26521 , n26518 , n26520 );
buf ( n374126 , n359378 );
buf ( n374127 , n351924 );
nand ( n26524 , n374126 , n374127 );
buf ( n374129 , n26524 );
buf ( n374130 , n374129 );
nand ( n26527 , n26521 , n374130 );
buf ( n374132 , n26527 );
buf ( n374133 , n374132 );
xor ( n26530 , n374120 , n374133 );
xor ( n26531 , n374005 , n374018 );
xor ( n26532 , n26531 , n374023 );
buf ( n374137 , n26532 );
buf ( n374138 , n374137 );
xor ( n26535 , n26530 , n374138 );
buf ( n374140 , n26535 );
buf ( n374141 , n374140 );
xor ( n26538 , n26510 , n374141 );
buf ( n374143 , n26538 );
buf ( n374144 , n374143 );
xor ( n26541 , n359506 , n359523 );
and ( n26542 , n26541 , n360123 );
and ( n26543 , n359506 , n359523 );
or ( n26544 , n26542 , n26543 );
buf ( n374149 , n26544 );
buf ( n374150 , n374149 );
xor ( n26547 , n374144 , n374150 );
buf ( n374152 , n6600 );
not ( n26549 , n374152 );
buf ( n374154 , n604 );
not ( n26551 , n374154 );
buf ( n374156 , n9637 );
not ( n26553 , n374156 );
or ( n26554 , n26551 , n26553 );
buf ( n374159 , n604 );
not ( n26556 , n374159 );
buf ( n374161 , n9636 );
nand ( n26558 , n26556 , n374161 );
buf ( n374163 , n26558 );
buf ( n374164 , n374163 );
nand ( n26561 , n26554 , n374164 );
buf ( n374166 , n26561 );
buf ( n374167 , n374166 );
not ( n26564 , n374167 );
or ( n26565 , n26549 , n26564 );
buf ( n374170 , n11836 );
buf ( n374171 , n355075 );
nand ( n26568 , n374170 , n374171 );
buf ( n374173 , n26568 );
buf ( n374174 , n374173 );
nand ( n26571 , n26565 , n374174 );
buf ( n374176 , n26571 );
buf ( n374177 , n374176 );
xor ( n26574 , n359332 , n359357 );
and ( n26575 , n26574 , n359490 );
and ( n26576 , n359332 , n359357 );
or ( n26577 , n26575 , n26576 );
buf ( n374182 , n26577 );
buf ( n374183 , n374182 );
xor ( n26580 , n374177 , n374183 );
buf ( n374185 , n607 );
not ( n26582 , n374185 );
buf ( n374187 , n606 );
not ( n26584 , n374187 );
buf ( n374189 , n25811 );
not ( n26586 , n374189 );
or ( n26587 , n26584 , n26586 );
buf ( n374192 , n373806 );
buf ( n374193 , n9642 );
nand ( n26590 , n374192 , n374193 );
buf ( n374195 , n26590 );
buf ( n374196 , n374195 );
nand ( n26593 , n26587 , n374196 );
buf ( n374198 , n26593 );
buf ( n374199 , n374198 );
not ( n26596 , n374199 );
or ( n26597 , n26582 , n26596 );
buf ( n374202 , n360112 );
buf ( n374203 , n357376 );
nand ( n26600 , n374202 , n374203 );
buf ( n374205 , n26600 );
buf ( n374206 , n374205 );
nand ( n26603 , n26597 , n374206 );
buf ( n374208 , n26603 );
buf ( n374209 , n374208 );
xor ( n26606 , n26580 , n374209 );
buf ( n374211 , n26606 );
buf ( n374212 , n374211 );
xor ( n26609 , n26547 , n374212 );
buf ( n374214 , n26609 );
buf ( n374215 , n374214 );
xor ( n26612 , n359493 , n359499 );
and ( n26613 , n26612 , n360126 );
and ( n26614 , n359493 , n359499 );
or ( n26615 , n26613 , n26614 );
buf ( n374220 , n26615 );
buf ( n374221 , n374220 );
nor ( n26618 , n374215 , n374221 );
buf ( n374223 , n26618 );
buf ( n374224 , n374223 );
not ( n26621 , n374224 );
buf ( n374226 , n12458 );
buf ( n374227 , n357542 );
nand ( n26624 , n26621 , n374226 , n374227 );
buf ( n374229 , n26624 );
not ( n26626 , n11645 );
or ( n26627 , n374229 , n26626 );
buf ( n374232 , n374214 );
not ( n26629 , n374232 );
buf ( n374234 , n26629 );
buf ( n374235 , n374234 );
buf ( n374236 , n374220 );
not ( n26633 , n374236 );
buf ( n374238 , n26633 );
buf ( n374239 , n374238 );
nand ( n26636 , n374235 , n374239 );
buf ( n374241 , n26636 );
buf ( n374242 , n374241 );
buf ( n374243 , n360128 );
buf ( n374244 , n360133 );
nor ( n26641 , n374243 , n374244 );
buf ( n374246 , n26641 );
or ( n26643 , n374246 , n11648 );
nand ( n26644 , n26643 , n360139 );
buf ( n374249 , n26644 );
and ( n26646 , n374242 , n374249 );
buf ( n374251 , n374214 );
buf ( n374252 , n374220 );
nand ( n26649 , n374251 , n374252 );
buf ( n374254 , n26649 );
buf ( n374255 , n374254 );
not ( n26652 , n374255 );
buf ( n374257 , n26652 );
buf ( n374258 , n374257 );
nor ( n26655 , n26646 , n374258 );
buf ( n374260 , n26655 );
nand ( n26657 , n26627 , n374260 );
not ( n26658 , n26657 );
xor ( n26659 , n373856 , n374068 );
xor ( n26660 , n26659 , n374073 );
buf ( n374265 , n26660 );
buf ( n374266 , n374265 );
not ( n26663 , n374266 );
buf ( n374268 , n26663 );
buf ( n374269 , n374268 );
xor ( n26666 , n373773 , n373798 );
xor ( n26667 , n26666 , n373819 );
buf ( n374272 , n26667 );
buf ( n374273 , n374272 );
buf ( n374274 , n6600 );
not ( n26671 , n374274 );
buf ( n374276 , n26204 );
not ( n26673 , n374276 );
or ( n26674 , n26671 , n26673 );
buf ( n374279 , n360105 );
not ( n26676 , n374279 );
buf ( n374281 , n26676 );
and ( n26678 , n604 , n374281 );
not ( n26679 , n604 );
and ( n26680 , n26679 , n360105 );
or ( n26681 , n26678 , n26680 );
buf ( n374286 , n26681 );
buf ( n374287 , n355075 );
nand ( n26684 , n374286 , n374287 );
buf ( n374289 , n26684 );
buf ( n374290 , n374289 );
nand ( n26687 , n26674 , n374290 );
buf ( n374292 , n26687 );
buf ( n374293 , n374292 );
xor ( n26690 , n373920 , n373938 );
xor ( n26691 , n26690 , n373943 );
buf ( n374296 , n26691 );
buf ( n374297 , n374296 );
xor ( n26694 , n374293 , n374297 );
xor ( n26695 , n374120 , n374133 );
and ( n26696 , n26695 , n374138 );
and ( n26697 , n374120 , n374133 );
or ( n26698 , n26696 , n26697 );
buf ( n374303 , n26698 );
buf ( n374304 , n374303 );
buf ( n374305 , n352149 );
not ( n26702 , n374305 );
buf ( n374307 , n373967 );
not ( n26704 , n374307 );
or ( n26705 , n26702 , n26704 );
buf ( n374310 , n374102 );
buf ( n374311 , n354113 );
nand ( n26708 , n374310 , n374311 );
buf ( n374313 , n26708 );
buf ( n374314 , n374313 );
nand ( n26711 , n26705 , n374314 );
buf ( n374316 , n26711 );
buf ( n374317 , n374316 );
xor ( n26714 , n374304 , n374317 );
buf ( n374319 , n6600 );
not ( n26716 , n374319 );
buf ( n374321 , n26681 );
not ( n26718 , n374321 );
or ( n26719 , n26716 , n26718 );
buf ( n374324 , n374166 );
buf ( n374325 , n355075 );
nand ( n26722 , n374324 , n374325 );
buf ( n374327 , n26722 );
buf ( n374328 , n374327 );
nand ( n26725 , n26719 , n374328 );
buf ( n374330 , n26725 );
buf ( n374331 , n374330 );
and ( n26728 , n26714 , n374331 );
and ( n26729 , n374304 , n374317 );
or ( n26730 , n26728 , n26729 );
buf ( n374335 , n26730 );
buf ( n374336 , n374335 );
and ( n26733 , n26694 , n374336 );
and ( n26734 , n374293 , n374297 );
or ( n26735 , n26733 , n26734 );
buf ( n374340 , n26735 );
buf ( n374341 , n374340 );
xor ( n26738 , n374273 , n374341 );
xor ( n26739 , n373948 , n373952 );
xor ( n26740 , n26739 , n374063 );
buf ( n374345 , n26740 );
buf ( n374346 , n374345 );
and ( n26743 , n26738 , n374346 );
and ( n26744 , n374273 , n374341 );
or ( n26745 , n26743 , n26744 );
buf ( n374350 , n26745 );
buf ( n374351 , n374350 );
not ( n26748 , n374351 );
buf ( n374353 , n26748 );
buf ( n374354 , n374353 );
nand ( n26751 , n374269 , n374354 );
buf ( n374356 , n26751 );
buf ( n374357 , n374356 );
xor ( n26754 , n374273 , n374341 );
xor ( n26755 , n26754 , n374346 );
buf ( n374360 , n26755 );
buf ( n374361 , n374360 );
not ( n26758 , n374361 );
xor ( n26759 , n373978 , n374038 );
xor ( n26760 , n26759 , n374058 );
buf ( n374365 , n26760 );
buf ( n374366 , n374365 );
xor ( n26763 , n373999 , n374028 );
xor ( n26764 , n26763 , n374033 );
buf ( n374369 , n26764 );
buf ( n374370 , n374369 );
buf ( n374371 , n357376 );
not ( n26768 , n374371 );
buf ( n374373 , n374198 );
not ( n26770 , n374373 );
or ( n26771 , n26768 , n26770 );
buf ( n374376 , n9642 );
buf ( n374377 , n374042 );
and ( n26774 , n374376 , n374377 );
not ( n26775 , n374376 );
buf ( n374380 , n374047 );
and ( n26777 , n26775 , n374380 );
nor ( n26778 , n26774 , n26777 );
buf ( n374383 , n26778 );
buf ( n374384 , n374383 );
buf ( n374385 , n607 );
nand ( n26782 , n374384 , n374385 );
buf ( n374387 , n26782 );
buf ( n374388 , n374387 );
nand ( n26785 , n26771 , n374388 );
buf ( n374390 , n26785 );
buf ( n374391 , n374390 );
xor ( n26788 , n374370 , n374391 );
xor ( n26789 , n374088 , n374113 );
and ( n26790 , n26789 , n374141 );
and ( n26791 , n374088 , n374113 );
or ( n26792 , n26790 , n26791 );
buf ( n374397 , n26792 );
buf ( n374398 , n374397 );
and ( n26795 , n26788 , n374398 );
and ( n26796 , n374370 , n374391 );
or ( n26797 , n26795 , n26796 );
buf ( n374402 , n26797 );
buf ( n374403 , n374402 );
xor ( n26800 , n374366 , n374403 );
xor ( n26801 , n374293 , n374297 );
xor ( n26802 , n26801 , n374336 );
buf ( n374407 , n26802 );
buf ( n374408 , n374407 );
and ( n26805 , n26800 , n374408 );
and ( n26806 , n374366 , n374403 );
or ( n26807 , n26805 , n26806 );
buf ( n374412 , n26807 );
buf ( n374413 , n374412 );
not ( n26810 , n374413 );
buf ( n374415 , n26810 );
buf ( n374416 , n374415 );
nand ( n26813 , n26758 , n374416 );
buf ( n374418 , n26813 );
buf ( n374419 , n374418 );
nand ( n26816 , n374357 , n374419 );
buf ( n374421 , n26816 );
buf ( n374422 , n374421 );
xor ( n26819 , n374366 , n374403 );
xor ( n26820 , n26819 , n374408 );
buf ( n374425 , n26820 );
xor ( n26822 , n374177 , n374183 );
and ( n26823 , n26822 , n374209 );
and ( n26824 , n374177 , n374183 );
or ( n26825 , n26823 , n26824 );
buf ( n374430 , n26825 );
buf ( n374431 , n374430 );
xor ( n26828 , n374304 , n374317 );
xor ( n26829 , n26828 , n374331 );
buf ( n374434 , n26829 );
buf ( n374435 , n374434 );
xor ( n26832 , n374431 , n374435 );
xor ( n26833 , n374370 , n374391 );
xor ( n26834 , n26833 , n374398 );
buf ( n374439 , n26834 );
buf ( n374440 , n374439 );
and ( n26837 , n26832 , n374440 );
and ( n26838 , n374431 , n374435 );
or ( n26839 , n26837 , n26838 );
buf ( n374444 , n26839 );
or ( n26841 , n374425 , n374444 );
xor ( n26842 , n374431 , n374435 );
xor ( n26843 , n26842 , n374440 );
buf ( n374448 , n26843 );
buf ( n374449 , n374448 );
not ( n26846 , n374449 );
xor ( n26847 , n374144 , n374150 );
and ( n26848 , n26847 , n374212 );
and ( n26849 , n374144 , n374150 );
or ( n26850 , n26848 , n26849 );
buf ( n374455 , n26850 );
buf ( n374456 , n374455 );
not ( n26853 , n374456 );
buf ( n374458 , n26853 );
buf ( n374459 , n374458 );
nand ( n26856 , n26846 , n374459 );
buf ( n374461 , n26856 );
nand ( n26858 , n26841 , n374461 );
buf ( n374463 , n26858 );
nor ( n26860 , n374422 , n374463 );
buf ( n374465 , n26860 );
not ( n26862 , n374465 );
or ( n26863 , n26658 , n26862 );
buf ( n374468 , n374421 );
not ( n26865 , n374468 );
buf ( n374470 , n26865 );
buf ( n374471 , n374470 );
buf ( n374472 , n374425 );
buf ( n374473 , n374444 );
nor ( n26870 , n374472 , n374473 );
buf ( n374475 , n26870 );
buf ( n374476 , n374475 );
buf ( n374477 , n374448 );
buf ( n374478 , n374455 );
nand ( n26875 , n374477 , n374478 );
buf ( n374480 , n26875 );
buf ( n374481 , n374480 );
or ( n26878 , n374476 , n374481 );
buf ( n374483 , n374425 );
buf ( n374484 , n374444 );
nand ( n26881 , n374483 , n374484 );
buf ( n374486 , n26881 );
buf ( n374487 , n374486 );
nand ( n26884 , n26878 , n374487 );
buf ( n374489 , n26884 );
buf ( n374490 , n374489 );
and ( n26887 , n374471 , n374490 );
buf ( n374492 , n374360 );
not ( n26889 , n374492 );
buf ( n374494 , n26889 );
buf ( n374495 , n374494 );
buf ( n374496 , n374415 );
nor ( n26893 , n374495 , n374496 );
buf ( n374498 , n26893 );
buf ( n374499 , n374498 );
not ( n26896 , n374499 );
buf ( n374501 , n374268 );
buf ( n374502 , n374353 );
nand ( n26899 , n374501 , n374502 );
buf ( n374504 , n26899 );
buf ( n374505 , n374504 );
not ( n26902 , n374505 );
or ( n26903 , n26896 , n26902 );
not ( n26904 , n374268 );
nand ( n26905 , n26904 , n374350 );
buf ( n374510 , n26905 );
nand ( n26907 , n26903 , n374510 );
buf ( n374512 , n26907 );
buf ( n374513 , n374512 );
nor ( n26910 , n26887 , n374513 );
buf ( n374515 , n26910 );
nand ( n26912 , n26863 , n374515 );
not ( n26913 , n26912 );
or ( n26914 , n26478 , n26913 );
not ( n26915 , n373612 );
not ( n26916 , n373842 );
or ( n26917 , n26915 , n26916 );
buf ( n374522 , n374077 );
buf ( n374523 , n373851 );
nand ( n26920 , n374522 , n374523 );
buf ( n374525 , n26920 );
nand ( n26922 , n26917 , n374525 );
buf ( n374527 , n26922 );
buf ( n374528 , n373848 );
and ( n26925 , n374527 , n374528 );
buf ( n374530 , n26925 );
buf ( n374531 , n374530 );
not ( n26928 , n374531 );
buf ( n374533 , n26928 );
nand ( n26930 , n26914 , n374533 );
xor ( n26931 , n373524 , n373549 );
and ( n26932 , n26931 , n373567 );
and ( n26933 , n373524 , n373549 );
or ( n26934 , n26932 , n26933 );
buf ( n374539 , n26934 );
buf ( n374540 , n374539 );
and ( n26937 , n592 , n25352 );
buf ( n374542 , n26937 );
buf ( n374543 , n348946 );
not ( n26940 , n374543 );
buf ( n374545 , n592 );
not ( n26942 , n374545 );
buf ( n374547 , n357505 );
not ( n26944 , n374547 );
or ( n26945 , n26942 , n26944 );
buf ( n374550 , n354093 );
buf ( n374551 , n348910 );
nand ( n26948 , n374550 , n374551 );
buf ( n374553 , n26948 );
buf ( n374554 , n374553 );
nand ( n26951 , n26945 , n374554 );
buf ( n374556 , n26951 );
buf ( n374557 , n374556 );
not ( n26954 , n374557 );
or ( n26955 , n26940 , n26954 );
buf ( n374560 , n373538 );
buf ( n374561 , n1250 );
nand ( n26958 , n374560 , n374561 );
buf ( n374563 , n26958 );
buf ( n374564 , n374563 );
nand ( n26961 , n26955 , n374564 );
buf ( n374566 , n26961 );
buf ( n374567 , n374566 );
xor ( n26964 , n374542 , n374567 );
buf ( n374569 , n349035 );
not ( n26966 , n374569 );
xor ( n26967 , n594 , n7359 );
buf ( n374572 , n26967 );
not ( n26969 , n374572 );
or ( n26970 , n26966 , n26969 );
buf ( n374575 , n25952 );
buf ( n374576 , n1397 );
nand ( n26973 , n374575 , n374576 );
buf ( n374578 , n26973 );
buf ( n374579 , n374578 );
nand ( n26976 , n26970 , n374579 );
buf ( n374581 , n26976 );
buf ( n374582 , n374581 );
xor ( n26979 , n26964 , n374582 );
buf ( n374584 , n26979 );
buf ( n374585 , n374584 );
xor ( n26982 , n374540 , n374585 );
buf ( n374587 , n372772 );
not ( n26984 , n374587 );
buf ( n374589 , n25976 );
not ( n26986 , n374589 );
or ( n26987 , n26984 , n26986 );
buf ( n374592 , n596 );
not ( n26989 , n374592 );
buf ( n374594 , n357355 );
not ( n26991 , n374594 );
or ( n26992 , n26989 , n26991 );
buf ( n374597 , n9664 );
buf ( n374598 , n348865 );
nand ( n26995 , n374597 , n374598 );
buf ( n374600 , n26995 );
buf ( n374601 , n374600 );
nand ( n26998 , n26992 , n374601 );
buf ( n374603 , n26998 );
buf ( n374604 , n374603 );
buf ( n374605 , n347319 );
nand ( n27002 , n374604 , n374605 );
buf ( n374607 , n27002 );
buf ( n374608 , n374607 );
nand ( n27005 , n26987 , n374608 );
buf ( n374610 , n27005 );
buf ( n374611 , n374610 );
xor ( n27008 , n26982 , n374611 );
buf ( n374613 , n27008 );
buf ( n374614 , n374613 );
xor ( n27011 , n373385 , n373409 );
and ( n27012 , n27011 , n373442 );
and ( n27013 , n373385 , n373409 );
or ( n27014 , n27012 , n27013 );
buf ( n374619 , n27014 );
buf ( n374620 , n374619 );
xor ( n27017 , n374614 , n374620 );
xor ( n27018 , n373476 , n373487 );
and ( n27019 , n27018 , n373509 );
and ( n27020 , n373476 , n373487 );
or ( n27021 , n27019 , n27020 );
buf ( n374626 , n27021 );
buf ( n374627 , n374626 );
xor ( n27024 , n27017 , n374627 );
buf ( n374629 , n27024 );
buf ( n374630 , n374629 );
buf ( n374631 , n354113 );
not ( n27028 , n374631 );
buf ( n374633 , n373459 );
not ( n27030 , n374633 );
or ( n27031 , n27028 , n27030 );
buf ( n374636 , n25700 );
not ( n27033 , n374636 );
buf ( n374638 , n373179 );
not ( n27035 , n374638 );
and ( n27036 , n27033 , n27035 );
buf ( n374641 , n25700 );
buf ( n374642 , n373187 );
and ( n27039 , n374641 , n374642 );
nor ( n27040 , n27036 , n27039 );
buf ( n374645 , n27040 );
buf ( n374646 , n374645 );
nand ( n27043 , n27031 , n374646 );
buf ( n374648 , n27043 );
buf ( n374649 , n374648 );
not ( n27046 , n4443 );
not ( n27047 , n25791 );
or ( n27048 , n27046 , n27047 );
not ( n27049 , n347312 );
buf ( n374654 , n360099 );
not ( n27051 , n374654 );
buf ( n374656 , n27051 );
not ( n27053 , n374656 );
or ( n27054 , n27049 , n27053 );
buf ( n374659 , n12420 );
not ( n27056 , n374659 );
buf ( n374661 , n598 );
nand ( n27058 , n27056 , n374661 );
buf ( n374663 , n27058 );
nand ( n27060 , n27054 , n374663 );
nand ( n27061 , n27060 , n4362 );
nand ( n27062 , n27048 , n27061 );
buf ( n374667 , n27062 );
xor ( n27064 , n374649 , n374667 );
buf ( n374669 , n9751 );
not ( n27066 , n374669 );
buf ( n374671 , n600 );
buf ( n374672 , n25627 );
buf ( n27069 , n374672 );
buf ( n374674 , n27069 );
buf ( n374675 , n374674 );
and ( n27072 , n374671 , n374675 );
not ( n27073 , n374671 );
buf ( n374678 , n373322 );
and ( n27075 , n27073 , n374678 );
nor ( n27076 , n27072 , n27075 );
buf ( n374681 , n27076 );
buf ( n374682 , n374681 );
not ( n27079 , n374682 );
or ( n27080 , n27066 , n27079 );
buf ( n374685 , n373425 );
buf ( n374686 , n351924 );
nand ( n27083 , n374685 , n374686 );
buf ( n374688 , n27083 );
buf ( n374689 , n374688 );
nand ( n27086 , n27080 , n374689 );
buf ( n374691 , n27086 );
buf ( n374692 , n374691 );
xor ( n27089 , n27064 , n374692 );
buf ( n374694 , n27089 );
buf ( n374695 , n374694 );
buf ( n374696 , n355075 );
not ( n27093 , n374696 );
buf ( n374698 , n25878 );
not ( n27095 , n374698 );
or ( n27096 , n27093 , n27095 );
and ( n27097 , n604 , n372582 );
not ( n27098 , n604 );
buf ( n374703 , n24975 );
buf ( n27100 , n374703 );
buf ( n374705 , n27100 );
and ( n27102 , n27098 , n374705 );
or ( n27103 , n27097 , n27102 );
buf ( n374708 , n27103 );
buf ( n374709 , n6600 );
nand ( n27106 , n374708 , n374709 );
buf ( n374711 , n27106 );
buf ( n374712 , n374711 );
nand ( n27109 , n27096 , n374712 );
buf ( n374714 , n27109 );
buf ( n374715 , n374714 );
xor ( n27112 , n373519 , n373570 );
and ( n27113 , n27112 , n373588 );
and ( n27114 , n373519 , n373570 );
or ( n27115 , n27113 , n27114 );
buf ( n374720 , n27115 );
buf ( n374721 , n374720 );
xor ( n27118 , n374715 , n374721 );
buf ( n374723 , n357376 );
not ( n27120 , n374723 );
buf ( n374725 , n373504 );
not ( n27122 , n374725 );
or ( n27123 , n27120 , n27122 );
not ( n27124 , n606 );
nand ( n27125 , n16929 , n8323 );
not ( n27126 , n27125 );
nand ( n27127 , n27126 , n14500 , n16900 , n16955 );
buf ( n27128 , n365878 );
and ( n27129 , n27127 , n27128 );
not ( n27130 , n27127 );
not ( n27131 , n23236 );
and ( n27132 , n27130 , n27131 );
nor ( n27133 , n27129 , n27132 );
not ( n27134 , n27133 );
not ( n27135 , n27134 );
or ( n27136 , n27124 , n27135 );
buf ( n27137 , n27133 );
nand ( n27138 , n27137 , n9642 );
nand ( n27139 , n27136 , n27138 );
buf ( n374744 , n27139 );
buf ( n374745 , n607 );
nand ( n27142 , n374744 , n374745 );
buf ( n374747 , n27142 );
buf ( n374748 , n374747 );
nand ( n27145 , n27123 , n374748 );
buf ( n374750 , n27145 );
buf ( n374751 , n374750 );
xor ( n27148 , n27118 , n374751 );
buf ( n374753 , n27148 );
buf ( n374754 , n374753 );
xor ( n27151 , n374695 , n374754 );
xor ( n27152 , n373591 , n373597 );
and ( n27153 , n27152 , n373604 );
and ( n27154 , n373591 , n373597 );
or ( n27155 , n27153 , n27154 );
buf ( n374760 , n27155 );
buf ( n374761 , n374760 );
xor ( n27158 , n27151 , n374761 );
buf ( n374763 , n27158 );
buf ( n374764 , n374763 );
xor ( n27161 , n374630 , n374764 );
xor ( n27162 , n373445 , n373512 );
and ( n27163 , n27162 , n373607 );
and ( n27164 , n373445 , n373512 );
or ( n27165 , n27163 , n27164 );
buf ( n374770 , n27165 );
buf ( n374771 , n374770 );
xor ( n27168 , n27161 , n374771 );
buf ( n374773 , n27168 );
buf ( n374774 , n374773 );
not ( n27171 , n374774 );
buf ( n374776 , n27171 );
buf ( n374777 , n374776 );
xor ( n27174 , n373012 , n373378 );
and ( n27175 , n27174 , n373610 );
and ( n27176 , n373012 , n373378 );
or ( n27177 , n27175 , n27176 );
buf ( n374782 , n27177 );
buf ( n374783 , n374782 );
not ( n27180 , n374783 );
buf ( n374785 , n27180 );
buf ( n374786 , n374785 );
nand ( n27183 , n374777 , n374786 );
buf ( n374788 , n27183 );
buf ( n374789 , n374788 );
buf ( n374790 , n374776 );
not ( n27187 , n374790 );
buf ( n374792 , n374782 );
nand ( n27189 , n27187 , n374792 );
buf ( n374794 , n27189 );
buf ( n374795 , n374794 );
nand ( n27192 , n374789 , n374795 );
buf ( n374797 , n27192 );
xnor ( n27194 , n26930 , n374797 );
buf ( n27195 , n27194 );
buf ( n27196 , n27195 );
buf ( n374801 , n27196 );
xor ( n27198 , n372537 , n372538 );
xor ( n27199 , n27198 , n374801 );
buf ( n374804 , n27199 );
xor ( n27201 , n372537 , n372538 );
and ( n27202 , n27201 , n374801 );
and ( n27203 , n372537 , n372538 );
or ( n27204 , n27202 , n27203 );
buf ( n374809 , n27204 );
buf ( n374810 , n355519 );
buf ( n374811 , n355728 );
buf ( n374812 , n12479 );
xor ( n27209 , n374810 , n374811 );
xor ( n27210 , n27209 , n374812 );
buf ( n374815 , n27210 );
xor ( n27212 , n374810 , n374811 );
and ( n27213 , n27212 , n374812 );
and ( n27214 , n374810 , n374811 );
or ( n27215 , n27213 , n27214 );
buf ( n374820 , n27215 );
buf ( n374821 , n356425 );
buf ( n374822 , n356647 );
not ( n27219 , n26626 );
not ( n27220 , n357539 );
not ( n27221 , n357388 );
not ( n27222 , n27221 );
or ( n27223 , n27220 , n27222 );
nand ( n27224 , n27223 , n11648 );
buf ( n374829 , n27224 );
not ( n27226 , n374829 );
buf ( n374831 , n27226 );
not ( n27228 , n374831 );
or ( n27229 , n27219 , n27228 );
buf ( n374834 , n27224 );
buf ( n374835 , n11645 );
nand ( n27232 , n374834 , n374835 );
buf ( n374837 , n27232 );
nand ( n27234 , n27229 , n374837 );
buf ( n374839 , n27234 );
xor ( n27236 , n374821 , n374822 );
xor ( n27237 , n27236 , n374839 );
buf ( n374842 , n27237 );
xor ( n27239 , n374821 , n374822 );
and ( n27240 , n27239 , n374839 );
and ( n27241 , n374821 , n374822 );
or ( n27242 , n27240 , n27241 );
buf ( n374847 , n27242 );
buf ( n374848 , n360673 );
buf ( n374849 , n360521 );
not ( n27246 , n26657 );
buf ( n374851 , n374461 );
buf ( n374852 , n374480 );
nand ( n27249 , n374851 , n374852 );
buf ( n374854 , n27249 );
and ( n27251 , n27246 , n374854 );
not ( n27252 , n27246 );
buf ( n374857 , n374854 );
not ( n27254 , n374857 );
buf ( n374859 , n27254 );
and ( n27256 , n27252 , n374859 );
nor ( n27257 , n27251 , n27256 );
buf ( n27258 , n27257 );
buf ( n374863 , n27258 );
xor ( n27260 , n374848 , n374849 );
xor ( n27261 , n27260 , n374863 );
buf ( n374866 , n27261 );
xor ( n27263 , n374848 , n374849 );
and ( n27264 , n27263 , n374863 );
and ( n27265 , n374848 , n374849 );
or ( n27266 , n27264 , n27265 );
buf ( n374871 , n27266 );
buf ( n374872 , n361414 );
buf ( n374873 , n361559 );
not ( n27270 , n26657 );
buf ( n374875 , n26858 );
not ( n27272 , n374875 );
buf ( n374877 , n27272 );
not ( n27274 , n374877 );
or ( n27275 , n27270 , n27274 );
buf ( n374880 , n374489 );
not ( n27277 , n374880 );
buf ( n374882 , n27277 );
nand ( n27279 , n27275 , n374882 );
not ( n27280 , n27279 );
buf ( n374885 , n374494 );
buf ( n374886 , n374415 );
nand ( n27283 , n374885 , n374886 );
buf ( n374888 , n27283 );
buf ( n374889 , n374888 );
buf ( n374890 , n374494 );
not ( n27287 , n374890 );
buf ( n374892 , n374412 );
nand ( n27289 , n27287 , n374892 );
buf ( n374894 , n27289 );
buf ( n374895 , n374894 );
nand ( n27292 , n374889 , n374895 );
buf ( n374897 , n27292 );
and ( n27294 , n27280 , n374897 );
not ( n27295 , n27280 );
buf ( n374900 , n374897 );
not ( n27297 , n374900 );
buf ( n374902 , n27297 );
and ( n27299 , n27295 , n374902 );
nor ( n27300 , n27294 , n27299 );
buf ( n27301 , n27300 );
buf ( n374906 , n27301 );
xor ( n27303 , n374872 , n374873 );
xor ( n27304 , n27303 , n374906 );
buf ( n374909 , n27304 );
xor ( n27306 , n374872 , n374873 );
and ( n27307 , n27306 , n374906 );
and ( n27308 , n374872 , n374873 );
or ( n27309 , n27307 , n27308 );
buf ( n374914 , n27309 );
buf ( n374915 , n353173 );
buf ( n374916 , n353360 );
and ( n27313 , n358215 , n359259 );
buf ( n27314 , n11577 );
and ( n27315 , n27313 , n27314 );
not ( n27316 , n27313 );
not ( n27317 , n27314 );
and ( n27318 , n27316 , n27317 );
nor ( n27319 , n27315 , n27318 );
buf ( n27320 , n27319 );
buf ( n374925 , n27320 );
xor ( n27322 , n374915 , n374916 );
xor ( n27323 , n27322 , n374925 );
buf ( n374928 , n27323 );
xor ( n27325 , n374915 , n374916 );
and ( n27326 , n27325 , n374925 );
and ( n27327 , n374915 , n374916 );
or ( n27328 , n27326 , n27327 );
buf ( n374933 , n27328 );
buf ( n374934 , n15871 );
buf ( n374935 , n15877 );
not ( n27332 , n374788 );
not ( n27333 , n26930 );
or ( n27334 , n27332 , n27333 );
nand ( n27335 , n27334 , n374794 );
xor ( n27336 , n374630 , n374764 );
and ( n27337 , n27336 , n374771 );
and ( n27338 , n374630 , n374764 );
or ( n27339 , n27337 , n27338 );
buf ( n374944 , n27339 );
buf ( n374945 , n374944 );
not ( n27342 , n374945 );
buf ( n374947 , n27342 );
buf ( n374948 , n374947 );
not ( n27345 , n374948 );
buf ( n374950 , n27345 );
buf ( n374951 , n374950 );
xor ( n27348 , n374649 , n374667 );
and ( n27349 , n27348 , n374692 );
and ( n27350 , n374649 , n374667 );
or ( n27351 , n27349 , n27350 );
buf ( n374956 , n27351 );
buf ( n374957 , n374956 );
xor ( n27354 , n374542 , n374567 );
and ( n27355 , n27354 , n374582 );
and ( n27356 , n374542 , n374567 );
or ( n27357 , n27355 , n27356 );
buf ( n374962 , n27357 );
buf ( n374963 , n374962 );
buf ( n374964 , n372772 );
not ( n27361 , n374964 );
buf ( n374966 , n374603 );
not ( n27363 , n374966 );
or ( n27364 , n27361 , n27363 );
and ( n27365 , n9635 , n348865 );
not ( n27366 , n9635 );
and ( n27367 , n27366 , n596 );
or ( n27368 , n27365 , n27367 );
buf ( n374973 , n27368 );
buf ( n374974 , n347319 );
nand ( n27371 , n374973 , n374974 );
buf ( n374976 , n27371 );
buf ( n374977 , n374976 );
nand ( n27374 , n27364 , n374977 );
buf ( n374979 , n27374 );
buf ( n374980 , n374979 );
xor ( n27377 , n374963 , n374980 );
not ( n27378 , n4443 );
not ( n27379 , n27060 );
or ( n27380 , n27378 , n27379 );
buf ( n374985 , n373806 );
not ( n27382 , n374985 );
buf ( n374987 , n25301 );
not ( n27384 , n374987 );
and ( n27385 , n27382 , n27384 );
buf ( n374990 , n25566 );
buf ( n374991 , n25309 );
and ( n27388 , n374990 , n374991 );
nor ( n27389 , n27385 , n27388 );
buf ( n374994 , n27389 );
nand ( n27391 , n27380 , n374994 );
buf ( n374996 , n27391 );
xor ( n27393 , n27377 , n374996 );
buf ( n374998 , n27393 );
buf ( n374999 , n374998 );
xor ( n27396 , n374957 , n374999 );
not ( n27397 , n9751 );
buf ( n375002 , n600 );
not ( n27399 , n375002 );
buf ( n375004 , n25676 );
not ( n27401 , n375004 );
or ( n27402 , n27399 , n27401 );
buf ( n375007 , n25672 );
buf ( n375008 , n6460 );
nand ( n27405 , n375007 , n375008 );
buf ( n375010 , n27405 );
buf ( n375011 , n375010 );
nand ( n27408 , n27402 , n375011 );
buf ( n375013 , n27408 );
not ( n27410 , n375013 );
or ( n27411 , n27397 , n27410 );
or ( n27412 , n25866 , n358055 );
nand ( n27413 , n25866 , n358062 );
nand ( n27414 , n27412 , n27413 );
nand ( n27415 , n27411 , n27414 );
buf ( n375020 , n27415 );
buf ( n375021 , n6458 );
buf ( n375022 , n592 );
and ( n27419 , n375021 , n375022 );
buf ( n375024 , n27419 );
buf ( n375025 , n375024 );
buf ( n375026 , n348946 );
not ( n27423 , n375026 );
buf ( n375028 , n592 );
buf ( n375029 , n354053 );
xor ( n27426 , n375028 , n375029 );
buf ( n375031 , n27426 );
buf ( n375032 , n375031 );
not ( n27429 , n375032 );
or ( n27430 , n27423 , n27429 );
buf ( n375035 , n374556 );
buf ( n375036 , n1250 );
buf ( n27433 , n375036 );
buf ( n375038 , n27433 );
buf ( n375039 , n375038 );
nand ( n27436 , n375035 , n375039 );
buf ( n375041 , n27436 );
buf ( n375042 , n375041 );
nand ( n27439 , n27430 , n375042 );
buf ( n375044 , n27439 );
buf ( n375045 , n375044 );
xor ( n27442 , n375025 , n375045 );
and ( n27443 , n8333 , n372871 );
not ( n27444 , n8333 );
and ( n27445 , n27444 , n372880 );
nor ( n27446 , n27443 , n27445 );
buf ( n375051 , n26967 );
buf ( n375052 , n1397 );
nand ( n27449 , n375051 , n375052 );
buf ( n375054 , n27449 );
nand ( n27451 , n27446 , n375054 );
buf ( n375056 , n27451 );
xor ( n27453 , n27442 , n375056 );
buf ( n375058 , n27453 );
buf ( n375059 , n375058 );
xor ( n27456 , n375020 , n375059 );
buf ( n375061 , n6600 );
not ( n27458 , n375061 );
not ( n27459 , n604 );
not ( n27460 , n373494 );
or ( n27461 , n27459 , n27460 );
not ( n27462 , n604 );
nand ( n27463 , n27462 , n17009 );
nand ( n27464 , n27461 , n27463 );
buf ( n375069 , n27464 );
not ( n27466 , n375069 );
or ( n27467 , n27458 , n27466 );
buf ( n375072 , n27103 );
buf ( n375073 , n355075 );
nand ( n27470 , n375072 , n375073 );
buf ( n375075 , n27470 );
buf ( n375076 , n375075 );
nand ( n27473 , n27467 , n375076 );
buf ( n375078 , n27473 );
buf ( n375079 , n375078 );
xor ( n27476 , n27456 , n375079 );
buf ( n375081 , n27476 );
buf ( n375082 , n375081 );
xor ( n27479 , n27396 , n375082 );
buf ( n375084 , n27479 );
buf ( n375085 , n375084 );
xor ( n27482 , n374695 , n374754 );
and ( n27483 , n27482 , n374761 );
and ( n27484 , n374695 , n374754 );
or ( n27485 , n27483 , n27484 );
buf ( n375090 , n27485 );
buf ( n375091 , n375090 );
xor ( n27488 , n375085 , n375091 );
xor ( n27489 , n374715 , n374721 );
and ( n27490 , n27489 , n374751 );
and ( n27491 , n374715 , n374721 );
or ( n27492 , n27490 , n27491 );
buf ( n375097 , n27492 );
buf ( n375098 , n375097 );
buf ( n375099 , n352149 );
not ( n27496 , n375099 );
buf ( n375101 , n602 );
not ( n27498 , n375101 );
buf ( n375103 , n24943 );
not ( n27500 , n375103 );
buf ( n375105 , n27500 );
buf ( n375106 , n375105 );
not ( n27503 , n375106 );
or ( n27504 , n27498 , n27503 );
buf ( n375109 , n24943 );
buf ( n375110 , n349406 );
nand ( n27507 , n375109 , n375110 );
buf ( n375112 , n27507 );
buf ( n375113 , n375112 );
nand ( n27510 , n27504 , n375113 );
buf ( n375115 , n27510 );
buf ( n375116 , n375115 );
not ( n27513 , n375116 );
or ( n27514 , n27496 , n27513 );
not ( n27515 , n25700 );
not ( n27516 , n27515 );
buf ( n375121 , n27516 );
buf ( n375122 , n358417 );
and ( n27519 , n375121 , n375122 );
buf ( n375124 , n27515 );
buf ( n375125 , n358424 );
and ( n27522 , n375124 , n375125 );
nor ( n27523 , n27519 , n27522 );
buf ( n375128 , n27523 );
buf ( n375129 , n375128 );
nand ( n27526 , n27514 , n375129 );
buf ( n375131 , n27526 );
buf ( n375132 , n375131 );
xor ( n27529 , n374540 , n374585 );
and ( n27530 , n27529 , n374611 );
and ( n27531 , n374540 , n374585 );
or ( n27532 , n27530 , n27531 );
buf ( n375137 , n27532 );
buf ( n375138 , n375137 );
xor ( n27535 , n375132 , n375138 );
buf ( n375140 , n357376 );
not ( n27537 , n375140 );
buf ( n375142 , n27139 );
not ( n27539 , n375142 );
or ( n27540 , n27537 , n27539 );
buf ( n375145 , n606 );
not ( n27542 , n375145 );
not ( n27543 , n17013 );
and ( n27544 , n16900 , n365877 );
and ( n27545 , n17002 , n17019 , n16958 );
nand ( n27546 , n27544 , n17030 , n27545 );
not ( n27547 , n27546 );
or ( n27548 , n27543 , n27547 );
buf ( n375153 , n17013 );
not ( n27550 , n375153 );
buf ( n375155 , n27550 );
nand ( n27552 , n27544 , n17030 , n27545 , n375155 );
nand ( n27553 , n27548 , n27552 );
buf ( n27554 , n27553 );
buf ( n375159 , n27554 );
not ( n27556 , n375159 );
buf ( n375161 , n27556 );
buf ( n375162 , n375161 );
not ( n27559 , n375162 );
or ( n27560 , n27542 , n27559 );
buf ( n375165 , n27554 );
buf ( n375166 , n9642 );
nand ( n27563 , n375165 , n375166 );
buf ( n375168 , n27563 );
buf ( n375169 , n375168 );
nand ( n27566 , n27560 , n375169 );
buf ( n375171 , n27566 );
buf ( n375172 , n375171 );
buf ( n375173 , n607 );
nand ( n27570 , n375172 , n375173 );
buf ( n375175 , n27570 );
buf ( n375176 , n375175 );
nand ( n27573 , n27540 , n375176 );
buf ( n375178 , n27573 );
buf ( n375179 , n375178 );
xor ( n27576 , n27535 , n375179 );
buf ( n375181 , n27576 );
buf ( n375182 , n375181 );
xor ( n27579 , n375098 , n375182 );
xor ( n27580 , n374614 , n374620 );
and ( n27581 , n27580 , n374627 );
and ( n27582 , n374614 , n374620 );
or ( n27583 , n27581 , n27582 );
buf ( n375188 , n27583 );
buf ( n375189 , n375188 );
xor ( n27586 , n27579 , n375189 );
buf ( n375191 , n27586 );
buf ( n375192 , n375191 );
xor ( n27589 , n27488 , n375192 );
buf ( n375194 , n27589 );
buf ( n375195 , n375194 );
not ( n27592 , n375195 );
buf ( n375197 , n27592 );
buf ( n375198 , n375197 );
not ( n27595 , n375198 );
buf ( n375200 , n27595 );
buf ( n375201 , n375200 );
nand ( n27598 , n374951 , n375201 );
buf ( n375203 , n27598 );
buf ( n375204 , n375197 );
buf ( n375205 , n374947 );
nand ( n27602 , n375204 , n375205 );
buf ( n375207 , n27602 );
buf ( n27604 , n375207 );
nand ( n27605 , n375203 , n27604 );
not ( n27606 , n27605 );
and ( n27607 , n27335 , n27606 );
not ( n27608 , n27335 );
and ( n27609 , n27608 , n27605 );
nor ( n27610 , n27607 , n27609 );
buf ( n27611 , n27610 );
not ( n27612 , n27611 );
not ( n27613 , n27612 );
buf ( n375218 , n27613 );
xor ( n27615 , n374934 , n374935 );
xor ( n27616 , n27615 , n375218 );
buf ( n375221 , n27616 );
xor ( n27618 , n374934 , n374935 );
and ( n27619 , n27618 , n375218 );
and ( n27620 , n374934 , n374935 );
or ( n27621 , n27619 , n27620 );
buf ( n375226 , n27621 );
buf ( n375227 , n347768 );
buf ( n375228 , n347771 );
xor ( n27625 , n375227 , n375228 );
buf ( n375230 , n27625 );
and ( n27627 , n375227 , n375228 );
buf ( n375232 , n27627 );
buf ( n375233 , n364397 );
buf ( n375234 , n364390 );
xor ( n27631 , n375233 , n375234 );
buf ( n375236 , n27631 );
buf ( n375237 , n364002 );
buf ( n375238 , n364009 );
xor ( n27635 , n375237 , n375238 );
and ( n27636 , n9635 , n348865 );
not ( n27637 , n9635 );
and ( n27638 , n27637 , n596 );
or ( n27639 , n27636 , n27638 );
not ( n27640 , n27639 );
not ( n27641 , n372772 );
or ( n27642 , n27640 , n27641 );
and ( n27643 , n12420 , n372825 );
not ( n27644 , n12420 );
and ( n27645 , n27644 , n372831 );
nor ( n27646 , n27643 , n27645 );
nand ( n27647 , n27642 , n27646 );
buf ( n375252 , n27647 );
buf ( n375253 , n25566 );
buf ( n375254 , n357731 );
or ( n27651 , n375253 , n375254 );
buf ( n375256 , n27651 );
buf ( n375257 , n375256 );
buf ( n375258 , n25627 );
not ( n27655 , n375258 );
buf ( n375260 , n372908 );
nand ( n27657 , n27655 , n375260 );
buf ( n375262 , n27657 );
buf ( n375263 , n375262 );
buf ( n375264 , n25627 );
buf ( n375265 , n25309 );
nand ( n27662 , n375264 , n375265 );
buf ( n375267 , n27662 );
buf ( n375268 , n375267 );
buf ( n375269 , n25566 );
buf ( n375270 , n357742 );
nand ( n27667 , n375269 , n375270 );
buf ( n375272 , n27667 );
buf ( n375273 , n375272 );
nand ( n27670 , n375257 , n375263 , n375268 , n375273 );
buf ( n375275 , n27670 );
buf ( n375276 , n375275 );
xor ( n27673 , n375252 , n375276 );
not ( n27674 , n1722 );
and ( n27675 , n25700 , n6460 );
not ( n27676 , n25700 );
and ( n27677 , n27676 , n600 );
or ( n27678 , n27675 , n27677 );
not ( n27679 , n27678 );
or ( n27680 , n27674 , n27679 );
nand ( n27681 , n375013 , n351924 );
nand ( n27682 , n27680 , n27681 );
buf ( n375287 , n27682 );
xor ( n27684 , n27673 , n375287 );
buf ( n375289 , n27684 );
buf ( n375290 , n375289 );
xor ( n27687 , n375020 , n375059 );
and ( n27688 , n27687 , n375079 );
and ( n27689 , n375020 , n375059 );
or ( n27690 , n27688 , n27689 );
buf ( n375295 , n27690 );
buf ( n375296 , n375295 );
xor ( n27693 , n375290 , n375296 );
buf ( n375298 , n374705 );
not ( n27695 , n375298 );
buf ( n375300 , n373179 );
not ( n27697 , n375300 );
and ( n27698 , n27695 , n27697 );
buf ( n375303 , n372588 );
buf ( n375304 , n373187 );
and ( n27701 , n375303 , n375304 );
nor ( n27702 , n27698 , n27701 );
buf ( n375307 , n27702 );
buf ( n375308 , n372556 );
buf ( n375309 , n358424 );
nand ( n27706 , n375308 , n375309 );
buf ( n375311 , n27706 );
nand ( n27708 , n24943 , n358417 );
nand ( n27709 , n375307 , n375311 , n27708 );
buf ( n375314 , n27709 );
xor ( n27711 , n375025 , n375045 );
and ( n27712 , n27711 , n375056 );
and ( n27713 , n375025 , n375045 );
or ( n27714 , n27712 , n27713 );
buf ( n375319 , n27714 );
buf ( n375320 , n375319 );
xor ( n27717 , n375314 , n375320 );
buf ( n375322 , n9814 );
buf ( n375323 , n592 );
and ( n27720 , n375322 , n375323 );
buf ( n375325 , n27720 );
buf ( n375326 , n375325 );
buf ( n375327 , n348946 );
not ( n27724 , n375327 );
buf ( n375329 , n592 );
not ( n27726 , n375329 );
buf ( n375331 , n7360 );
not ( n27728 , n375331 );
or ( n27729 , n27726 , n27728 );
buf ( n375334 , n7359 );
buf ( n375335 , n348910 );
nand ( n27732 , n375334 , n375335 );
buf ( n375337 , n27732 );
buf ( n375338 , n375337 );
nand ( n27735 , n27729 , n375338 );
buf ( n375340 , n27735 );
buf ( n375341 , n375340 );
not ( n27738 , n375341 );
or ( n27739 , n27724 , n27738 );
buf ( n375344 , n375031 );
buf ( n375345 , n375038 );
nand ( n27742 , n375344 , n375345 );
buf ( n375347 , n27742 );
buf ( n375348 , n375347 );
nand ( n27745 , n27739 , n375348 );
buf ( n375350 , n27745 );
buf ( n375351 , n375350 );
xor ( n27748 , n375326 , n375351 );
buf ( n375353 , n349035 );
not ( n27750 , n375353 );
and ( n27751 , n594 , n357355 );
not ( n27752 , n594 );
and ( n27753 , n27752 , n9664 );
or ( n27754 , n27751 , n27753 );
buf ( n375359 , n27754 );
not ( n27756 , n375359 );
or ( n27757 , n27750 , n27756 );
not ( n27758 , n8330 );
buf ( n375363 , n27758 );
buf ( n375364 , n349153 );
and ( n27761 , n375363 , n375364 );
buf ( n375366 , n27758 );
buf ( n375367 , n349160 );
nor ( n27764 , n375366 , n375367 );
buf ( n375369 , n27764 );
buf ( n375370 , n375369 );
nor ( n27767 , n27761 , n375370 );
buf ( n375372 , n27767 );
buf ( n375373 , n375372 );
nand ( n27770 , n27757 , n375373 );
buf ( n375375 , n27770 );
buf ( n375376 , n375375 );
xor ( n27773 , n27748 , n375376 );
buf ( n375378 , n27773 );
buf ( n375379 , n375378 );
xor ( n27776 , n27717 , n375379 );
buf ( n375381 , n27776 );
buf ( n375382 , n375381 );
xor ( n27779 , n27693 , n375382 );
buf ( n375384 , n27779 );
buf ( n375385 , n375384 );
xor ( n27782 , n375098 , n375182 );
and ( n27783 , n27782 , n375189 );
and ( n27784 , n375098 , n375182 );
or ( n27785 , n27783 , n27784 );
buf ( n375390 , n27785 );
buf ( n375391 , n375390 );
xor ( n27788 , n375385 , n375391 );
xor ( n27789 , n375132 , n375138 );
and ( n27790 , n27789 , n375179 );
and ( n27791 , n375132 , n375138 );
or ( n27792 , n27790 , n27791 );
buf ( n375397 , n27792 );
buf ( n375398 , n375397 );
buf ( n375399 , n604 );
not ( n27796 , n375399 );
not ( n27797 , n27133 );
buf ( n375402 , n27797 );
not ( n27799 , n375402 );
or ( n27800 , n27796 , n27799 );
not ( n27801 , n604 );
nand ( n27802 , n27801 , n27133 );
buf ( n375407 , n27802 );
nand ( n27804 , n27800 , n375407 );
buf ( n375409 , n27804 );
not ( n27806 , n375409 );
not ( n27807 , n6600 );
or ( n27808 , n27806 , n27807 );
nand ( n27809 , n27464 , n355075 );
nand ( n27810 , n27808 , n27809 );
buf ( n375415 , n27810 );
xor ( n27812 , n374963 , n374980 );
and ( n27813 , n27812 , n374996 );
and ( n27814 , n374963 , n374980 );
or ( n27815 , n27813 , n27814 );
buf ( n375420 , n27815 );
buf ( n375421 , n375420 );
xor ( n27818 , n375415 , n375421 );
buf ( n375423 , n607 );
not ( n27820 , n375423 );
buf ( n375425 , n606 );
not ( n27822 , n375425 );
buf ( n27823 , n365892 );
not ( n27824 , n27823 );
not ( n27825 , n17014 );
or ( n27826 , n27824 , n27825 );
nand ( n27827 , n17015 , n370956 );
nand ( n27828 , n27826 , n27827 );
buf ( n375433 , n27828 );
not ( n27830 , n375433 );
buf ( n375435 , n27830 );
buf ( n375436 , n375435 );
not ( n27833 , n375436 );
or ( n27834 , n27822 , n27833 );
buf ( n375439 , n375435 );
not ( n27836 , n375439 );
buf ( n375441 , n27836 );
buf ( n375442 , n375441 );
buf ( n375443 , n9642 );
nand ( n27840 , n375442 , n375443 );
buf ( n375445 , n27840 );
buf ( n375446 , n375445 );
nand ( n27843 , n27834 , n375446 );
buf ( n375448 , n27843 );
buf ( n375449 , n375448 );
not ( n27846 , n375449 );
or ( n27847 , n27820 , n27846 );
buf ( n375452 , n375171 );
buf ( n375453 , n357376 );
nand ( n27850 , n375452 , n375453 );
buf ( n375455 , n27850 );
buf ( n375456 , n375455 );
nand ( n27853 , n27847 , n375456 );
buf ( n375458 , n27853 );
buf ( n375459 , n375458 );
xor ( n27856 , n27818 , n375459 );
buf ( n375461 , n27856 );
buf ( n375462 , n375461 );
xor ( n27859 , n375398 , n375462 );
xor ( n27860 , n374957 , n374999 );
and ( n27861 , n27860 , n375082 );
and ( n27862 , n374957 , n374999 );
or ( n27863 , n27861 , n27862 );
buf ( n375468 , n27863 );
buf ( n375469 , n375468 );
xor ( n27866 , n27859 , n375469 );
buf ( n375471 , n27866 );
buf ( n375472 , n375471 );
xor ( n27869 , n27788 , n375472 );
buf ( n375474 , n27869 );
xor ( n27871 , n375085 , n375091 );
and ( n27872 , n27871 , n375192 );
and ( n27873 , n375085 , n375091 );
or ( n27874 , n27872 , n27873 );
buf ( n375479 , n27874 );
or ( n27876 , n375474 , n375479 );
not ( n27877 , n27876 );
not ( n27878 , n26912 );
not ( n27879 , n374776 );
not ( n27880 , n374785 );
or ( n27881 , n27879 , n27880 );
not ( n27882 , n375194 );
nand ( n27883 , n27882 , n374947 );
nand ( n27884 , n27881 , n27883 );
nor ( n27885 , n27884 , n26476 );
not ( n27886 , n27885 );
or ( n27887 , n27878 , n27886 );
not ( n27888 , n27884 );
and ( n27889 , n27888 , n374530 );
buf ( n375494 , n374776 );
buf ( n375495 , n374785 );
nor ( n27892 , n375494 , n375495 );
buf ( n375497 , n27892 );
buf ( n375498 , n375497 );
not ( n27895 , n375498 );
buf ( n375500 , n375207 );
not ( n27897 , n375500 );
or ( n27898 , n27895 , n27897 );
buf ( n375503 , n375203 );
nand ( n27900 , n27898 , n375503 );
buf ( n375505 , n27900 );
nor ( n27902 , n27889 , n375505 );
nand ( n27903 , n27887 , n27902 );
not ( n27904 , n27903 );
or ( n27905 , n27877 , n27904 );
nand ( n27906 , n375474 , n375479 );
buf ( n27907 , n27906 );
nand ( n27908 , n27905 , n27907 );
not ( n27909 , n347319 );
or ( n27910 , n348865 , n25566 );
nand ( n27911 , n25566 , n348865 );
nand ( n27912 , n27910 , n27911 );
not ( n27913 , n27912 );
or ( n27914 , n27909 , n27913 );
buf ( n375519 , n360105 );
buf ( n375520 , n1651 );
and ( n27917 , n375519 , n375520 );
buf ( n375522 , n374281 );
buf ( n375523 , n1649 );
and ( n27920 , n375522 , n375523 );
nor ( n27921 , n27917 , n27920 );
buf ( n375526 , n27921 );
nand ( n27923 , n27914 , n375526 );
buf ( n375528 , n27923 );
buf ( n375529 , n374674 );
buf ( n375530 , n357731 );
nor ( n27927 , n375529 , n375530 );
buf ( n375532 , n27927 );
buf ( n375533 , n375532 );
buf ( n375534 , n25627 );
buf ( n375535 , n357742 );
and ( n27932 , n375534 , n375535 );
buf ( n375537 , n27932 );
buf ( n375538 , n375537 );
nor ( n27935 , n375533 , n375538 );
buf ( n375540 , n27935 );
buf ( n375541 , n375540 );
not ( n27938 , n598 );
not ( n27939 , n25676 );
or ( n27940 , n27938 , n27939 );
buf ( n375545 , n25672 );
buf ( n375546 , n347312 );
nand ( n27943 , n375545 , n375546 );
buf ( n375548 , n27943 );
nand ( n27945 , n27940 , n375548 );
buf ( n375550 , n27945 );
buf ( n375551 , n4362 );
nand ( n27948 , n375550 , n375551 );
buf ( n375553 , n27948 );
buf ( n375554 , n375553 );
nand ( n27951 , n375541 , n375554 );
buf ( n375556 , n27951 );
buf ( n375557 , n375556 );
xor ( n27954 , n375528 , n375557 );
not ( n27955 , n1722 );
not ( n27956 , n600 );
not ( n27957 , n372556 );
or ( n27958 , n27956 , n27957 );
nand ( n27959 , n24943 , n26117 );
nand ( n27960 , n27958 , n27959 );
not ( n27961 , n27960 );
or ( n27962 , n27955 , n27961 );
nand ( n27963 , n27678 , n351924 );
nand ( n27964 , n27962 , n27963 );
buf ( n375569 , n27964 );
xor ( n27966 , n27954 , n375569 );
buf ( n375571 , n27966 );
buf ( n375572 , n375571 );
xor ( n27969 , n375314 , n375320 );
and ( n27970 , n27969 , n375379 );
and ( n27971 , n375314 , n375320 );
or ( n27972 , n27970 , n27971 );
buf ( n375577 , n27972 );
buf ( n375578 , n375577 );
xor ( n27975 , n375572 , n375578 );
buf ( n375580 , n602 );
not ( n27977 , n375580 );
buf ( n375582 , n372582 );
not ( n27979 , n375582 );
or ( n27980 , n27977 , n27979 );
buf ( n375585 , n374705 );
buf ( n375586 , n349406 );
nand ( n27983 , n375585 , n375586 );
buf ( n375588 , n27983 );
buf ( n375589 , n375588 );
nand ( n27986 , n27980 , n375589 );
buf ( n375591 , n27986 );
not ( n27988 , n375591 );
not ( n27989 , n354113 );
or ( n27990 , n27988 , n27989 );
and ( n27991 , n17009 , n373187 );
not ( n27992 , n17009 );
and ( n27993 , n27992 , n373176 );
nor ( n27994 , n27991 , n27993 );
nand ( n27995 , n27990 , n27994 );
buf ( n375600 , n27995 );
and ( n27997 , n375028 , n375029 );
buf ( n375602 , n27997 );
buf ( n375603 , n375602 );
buf ( n375604 , n348946 );
not ( n28001 , n375604 );
and ( n28002 , n592 , n8330 );
not ( n28003 , n592 );
and ( n28004 , n28003 , n8333 );
or ( n28005 , n28002 , n28004 );
buf ( n375610 , n28005 );
not ( n28007 , n375610 );
or ( n28008 , n28001 , n28007 );
buf ( n375613 , n375340 );
buf ( n375614 , n375038 );
nand ( n28011 , n375613 , n375614 );
buf ( n375616 , n28011 );
buf ( n375617 , n375616 );
nand ( n28014 , n28008 , n375617 );
buf ( n375619 , n28014 );
buf ( n375620 , n375619 );
xor ( n28017 , n375603 , n375620 );
buf ( n375622 , n1397 );
not ( n28019 , n375622 );
buf ( n375624 , n27754 );
not ( n28021 , n375624 );
or ( n28022 , n28019 , n28021 );
buf ( n375627 , n9635 );
buf ( n375628 , n372871 );
and ( n28025 , n375627 , n375628 );
not ( n28026 , n375627 );
buf ( n375631 , n372880 );
and ( n28028 , n28026 , n375631 );
nor ( n28029 , n28025 , n28028 );
buf ( n375634 , n28029 );
buf ( n375635 , n375634 );
nand ( n28032 , n28022 , n375635 );
buf ( n375637 , n28032 );
buf ( n375638 , n375637 );
xor ( n28035 , n28017 , n375638 );
buf ( n375640 , n28035 );
buf ( n375641 , n375640 );
xor ( n28038 , n375600 , n375641 );
buf ( n375643 , n355075 );
not ( n28040 , n375643 );
buf ( n375645 , n375409 );
not ( n28042 , n375645 );
or ( n28043 , n28040 , n28042 );
xor ( n28044 , n604 , n27554 );
buf ( n375649 , n28044 );
buf ( n375650 , n6600 );
nand ( n28047 , n375649 , n375650 );
buf ( n375652 , n28047 );
buf ( n375653 , n375652 );
nand ( n28050 , n28043 , n375653 );
buf ( n375655 , n28050 );
buf ( n375656 , n375655 );
xor ( n28053 , n28038 , n375656 );
buf ( n375658 , n28053 );
buf ( n375659 , n375658 );
xor ( n28056 , n27975 , n375659 );
buf ( n375661 , n28056 );
buf ( n375662 , n375661 );
xor ( n28059 , n375415 , n375421 );
and ( n28060 , n28059 , n375459 );
and ( n28061 , n375415 , n375421 );
or ( n28062 , n28060 , n28061 );
buf ( n375667 , n28062 );
buf ( n375668 , n375667 );
xor ( n28065 , n375326 , n375351 );
and ( n28066 , n28065 , n375376 );
and ( n28067 , n375326 , n375351 );
or ( n28068 , n28066 , n28067 );
buf ( n375673 , n28068 );
buf ( n375674 , n375673 );
xor ( n28071 , n375252 , n375276 );
and ( n28072 , n28071 , n375287 );
and ( n28073 , n375252 , n375276 );
or ( n28074 , n28072 , n28073 );
buf ( n375679 , n28074 );
buf ( n375680 , n375679 );
xor ( n28077 , n375674 , n375680 );
buf ( n375682 , n357376 );
not ( n28079 , n375682 );
buf ( n375684 , n375448 );
not ( n28081 , n375684 );
or ( n28082 , n28079 , n28081 );
buf ( n375687 , n607 );
buf ( n375688 , n606 );
not ( n28085 , n375688 );
not ( n28086 , n16815 );
nand ( n28087 , n16957 , n16856 , n24940 );
not ( n28088 , n28087 );
or ( n28089 , n28086 , n28088 );
nand ( n28090 , n371006 , n16856 , n16957 , n24940 );
nand ( n28091 , n28089 , n28090 );
buf ( n28092 , n28091 );
not ( n28093 , n28092 );
buf ( n375698 , n28093 );
not ( n28095 , n375698 );
or ( n28096 , n28085 , n28095 );
buf ( n375701 , n28092 );
buf ( n375702 , n9642 );
nand ( n28099 , n375701 , n375702 );
buf ( n375704 , n28099 );
buf ( n375705 , n375704 );
nand ( n28102 , n28096 , n375705 );
buf ( n375707 , n28102 );
buf ( n375708 , n375707 );
nand ( n28105 , n375687 , n375708 );
buf ( n375710 , n28105 );
buf ( n375711 , n375710 );
nand ( n28108 , n28082 , n375711 );
buf ( n375713 , n28108 );
buf ( n375714 , n375713 );
xor ( n28111 , n28077 , n375714 );
buf ( n375716 , n28111 );
buf ( n375717 , n375716 );
xor ( n28114 , n375668 , n375717 );
xor ( n28115 , n375290 , n375296 );
and ( n28116 , n28115 , n375382 );
and ( n28117 , n375290 , n375296 );
or ( n28118 , n28116 , n28117 );
buf ( n375723 , n28118 );
buf ( n375724 , n375723 );
xor ( n28121 , n28114 , n375724 );
buf ( n375726 , n28121 );
buf ( n375727 , n375726 );
xor ( n28124 , n375662 , n375727 );
xor ( n28125 , n375398 , n375462 );
and ( n28126 , n28125 , n375469 );
and ( n28127 , n375398 , n375462 );
or ( n28128 , n28126 , n28127 );
buf ( n375733 , n28128 );
buf ( n375734 , n375733 );
xor ( n28131 , n28124 , n375734 );
buf ( n375736 , n28131 );
buf ( n375737 , n375736 );
xor ( n28134 , n375385 , n375391 );
and ( n28135 , n28134 , n375472 );
and ( n28136 , n375385 , n375391 );
or ( n28137 , n28135 , n28136 );
buf ( n375742 , n28137 );
buf ( n375743 , n375742 );
nor ( n28140 , n375737 , n375743 );
buf ( n375745 , n28140 );
buf ( n375746 , n375745 );
buf ( n28143 , n375746 );
buf ( n375748 , n28143 );
not ( n28145 , n375748 );
buf ( n375750 , n375736 );
buf ( n28147 , n375750 );
buf ( n375752 , n28147 );
buf ( n375753 , n375752 );
buf ( n375754 , n375742 );
nand ( n28151 , n375753 , n375754 );
buf ( n375756 , n28151 );
and ( n28153 , n28145 , n375756 );
and ( n28154 , n27908 , n28153 );
not ( n28155 , n27908 );
nand ( n28156 , n28145 , n375756 );
and ( n28157 , n28155 , n28156 );
nor ( n28158 , n28154 , n28157 );
buf ( n28159 , n28158 );
buf ( n28160 , n28159 );
buf ( n375765 , n28160 );
xor ( n28162 , n27635 , n375765 );
buf ( n375767 , n28162 );
buf ( n375768 , n375767 );
buf ( n375769 , n363763 );
buf ( n375770 , n16138 );
xor ( n28167 , n375769 , n375770 );
not ( n28168 , n27903 );
nand ( n28169 , n27906 , n27876 );
and ( n28170 , n28168 , n28169 );
not ( n28171 , n28168 );
not ( n28172 , n28169 );
and ( n28173 , n28171 , n28172 );
nor ( n28174 , n28170 , n28173 );
buf ( n375779 , n28174 );
buf ( n28176 , n375779 );
buf ( n375781 , n28176 );
buf ( n375782 , n375781 );
buf ( n28179 , n375782 );
buf ( n375784 , n28179 );
buf ( n28181 , n375784 );
buf ( n375786 , n28181 );
and ( n28183 , n28167 , n375786 );
and ( n28184 , n375769 , n375770 );
or ( n28185 , n28183 , n28184 );
buf ( n375790 , n28185 );
buf ( n375791 , n375790 );
xor ( n28188 , n375768 , n375791 );
buf ( n375793 , n375226 );
xor ( n28190 , n375769 , n375770 );
xor ( n28191 , n28190 , n375786 );
buf ( n375796 , n28191 );
buf ( n375797 , n375796 );
xor ( n28194 , n375793 , n375797 );
buf ( n375799 , n375221 );
buf ( n375800 , n374809 );
xor ( n28197 , n375799 , n375800 );
xor ( n28198 , n362813 , n362807 );
buf ( n375803 , n373615 );
buf ( n375804 , n373845 );
or ( n28201 , n375803 , n375804 );
buf ( n375806 , n28201 );
nand ( n28203 , n375806 , n373848 );
not ( n28204 , n28203 );
not ( n28205 , n26475 );
not ( n28206 , n26912 );
or ( n28207 , n28205 , n28206 );
nand ( n28208 , n373851 , n374077 );
nand ( n28209 , n28207 , n28208 );
not ( n28210 , n28209 );
not ( n28211 , n28210 );
or ( n28212 , n28204 , n28211 );
not ( n28213 , n28203 );
nand ( n28214 , n28209 , n28213 );
nand ( n28215 , n28212 , n28214 );
buf ( n375820 , n28215 );
not ( n28217 , n375820 );
buf ( n375822 , n28217 );
and ( n28219 , n28198 , n375822 );
and ( n28220 , n362813 , n362807 );
or ( n28221 , n28219 , n28220 );
buf ( n375826 , n28221 );
buf ( n375827 , n374804 );
xor ( n28224 , n375826 , n375827 );
buf ( n375829 , n362416 );
buf ( n375830 , n362431 );
xor ( n28227 , n375829 , n375830 );
buf ( n375832 , n26475 );
buf ( n375833 , n28208 );
nand ( n28230 , n375832 , n375833 );
buf ( n375835 , n28230 );
buf ( n375836 , n375835 );
not ( n28233 , n375836 );
buf ( n375838 , n28233 );
not ( n28235 , n375838 );
buf ( n375840 , n26912 );
buf ( n28237 , n375840 );
buf ( n375842 , n28237 );
buf ( n375843 , n375842 );
not ( n28240 , n375843 );
buf ( n375845 , n28240 );
not ( n28242 , n375845 );
or ( n28243 , n28235 , n28242 );
buf ( n375848 , n375842 );
buf ( n375849 , n375835 );
nand ( n28246 , n375848 , n375849 );
buf ( n375851 , n28246 );
nand ( n28248 , n28243 , n375851 );
not ( n28249 , n28248 );
not ( n28250 , n28249 );
buf ( n375855 , n28250 );
and ( n28252 , n28227 , n375855 );
and ( n28253 , n375829 , n375830 );
or ( n28254 , n28252 , n28253 );
buf ( n375859 , n28254 );
buf ( n375860 , n375859 );
xor ( n28257 , n362109 , n361993 );
not ( n28258 , n374888 );
not ( n28259 , n27279 );
or ( n28260 , n28258 , n28259 );
nand ( n28261 , n28260 , n374894 );
buf ( n375866 , n26905 );
buf ( n28263 , n375866 );
buf ( n375868 , n28263 );
nand ( n28265 , n375868 , n374504 );
not ( n28266 , n28265 );
and ( n28267 , n28261 , n28266 );
not ( n28268 , n28261 );
and ( n28269 , n28268 , n28265 );
nor ( n28270 , n28267 , n28269 );
and ( n28271 , n28257 , n28270 );
and ( n28272 , n362109 , n361993 );
or ( n28273 , n28271 , n28272 );
buf ( n375878 , n28273 );
xor ( n28275 , n375829 , n375830 );
xor ( n28276 , n28275 , n375855 );
buf ( n375881 , n28276 );
buf ( n375882 , n375881 );
xor ( n28279 , n375878 , n375882 );
buf ( n375884 , n374909 );
not ( n28281 , n375884 );
xor ( n28282 , n361201 , n361190 );
not ( n28283 , n374475 );
and ( n28284 , n28283 , n374486 );
not ( n28285 , n28284 );
not ( n28286 , n374461 );
not ( n28287 , n26657 );
or ( n28288 , n28286 , n28287 );
nand ( n28289 , n28288 , n374480 );
not ( n28290 , n28289 );
not ( n28291 , n28290 );
or ( n28292 , n28285 , n28291 );
not ( n28293 , n28284 );
nand ( n28294 , n28293 , n28289 );
nand ( n28295 , n28292 , n28294 );
not ( n28296 , n28295 );
not ( n28297 , n28296 );
and ( n28298 , n28282 , n28297 );
and ( n28299 , n361201 , n361190 );
or ( n28300 , n28298 , n28299 );
buf ( n375905 , n28300 );
not ( n28302 , n375905 );
buf ( n375907 , n28302 );
buf ( n375908 , n375907 );
nand ( n28305 , n28281 , n375908 );
buf ( n375910 , n28305 );
buf ( n375911 , n375910 );
not ( n28308 , n375911 );
xor ( n28309 , n361201 , n361190 );
xor ( n28310 , n28309 , n28297 );
buf ( n375915 , n28310 );
not ( n28312 , n375915 );
buf ( n375917 , n374871 );
not ( n28314 , n375917 );
buf ( n375919 , n28314 );
buf ( n375920 , n375919 );
nand ( n28317 , n28312 , n375920 );
buf ( n375922 , n28317 );
buf ( n375923 , n375922 );
not ( n28320 , n375923 );
buf ( n375925 , n374842 );
not ( n28322 , n375925 );
buf ( n375927 , n374820 );
not ( n28324 , n375927 );
buf ( n375929 , n28324 );
buf ( n375930 , n375929 );
nand ( n28327 , n28322 , n375930 );
buf ( n375932 , n28327 );
xor ( n28329 , n12504 , n357071 );
xor ( n28330 , n28329 , n12470 );
not ( n28331 , n28330 );
not ( n28332 , n374847 );
nand ( n28333 , n28331 , n28332 );
and ( n28334 , n375932 , n28333 );
not ( n28335 , n28334 );
buf ( n375940 , n12497 );
buf ( n28337 , n354819 );
buf ( n28338 , n28337 );
buf ( n375943 , n28338 );
xor ( n28340 , n375940 , n375943 );
not ( n28341 , n359288 );
not ( n28342 , n28341 );
not ( n28343 , n359282 );
not ( n28344 , n28343 );
or ( n28345 , n28342 , n28344 );
nand ( n28346 , n28345 , n359296 );
not ( n28347 , n28346 );
buf ( n28348 , n11584 );
not ( n28349 , n28348 );
or ( n28350 , n28347 , n28349 );
or ( n28351 , n28348 , n28346 );
nand ( n28352 , n28350 , n28351 );
buf ( n28353 , n28352 );
buf ( n375958 , n28353 );
xor ( n28355 , n28340 , n375958 );
buf ( n375960 , n28355 );
buf ( n375961 , n375960 );
not ( n28358 , n375961 );
buf ( n375963 , n374933 );
not ( n28360 , n375963 );
buf ( n375965 , n28360 );
buf ( n375966 , n375965 );
nand ( n28363 , n28358 , n375966 );
buf ( n375968 , n28363 );
buf ( n375969 , n375968 );
not ( n28366 , n375969 );
buf ( n375971 , n374928 );
buf ( n375972 , n352680 );
buf ( n375973 , n12486 );
xor ( n28370 , n375972 , n375973 );
buf ( n375975 , n358313 );
not ( n28372 , n375975 );
buf ( n375977 , n11576 );
nand ( n28374 , n28372 , n375977 );
buf ( n375979 , n28374 );
buf ( n375980 , n375979 );
buf ( n375981 , n11573 );
buf ( n28378 , n375981 );
buf ( n375983 , n28378 );
buf ( n375984 , n375983 );
not ( n28381 , n375984 );
buf ( n375986 , n28381 );
buf ( n375987 , n375986 );
and ( n28384 , n375980 , n375987 );
not ( n28385 , n375980 );
buf ( n375990 , n375983 );
and ( n28387 , n28385 , n375990 );
nor ( n28388 , n28384 , n28387 );
buf ( n375993 , n28388 );
buf ( n28390 , n375993 );
buf ( n375995 , n28390 );
and ( n28392 , n28370 , n375995 );
and ( n28393 , n375972 , n375973 );
or ( n28394 , n28392 , n28393 );
buf ( n375999 , n28394 );
buf ( n376000 , n375999 );
or ( n28397 , n375971 , n376000 );
xor ( n28398 , n375972 , n375973 );
xor ( n28399 , n28398 , n375995 );
buf ( n376004 , n28399 );
not ( n28401 , n376004 );
buf ( n376006 , n352445 );
buf ( n376007 , n12487 );
xor ( n28404 , n376006 , n376007 );
buf ( n376009 , n359239 );
not ( n28406 , n376009 );
buf ( n376011 , n359229 );
not ( n28408 , n376011 );
buf ( n376013 , n28408 );
buf ( n376014 , n376013 );
not ( n28411 , n376014 );
or ( n28412 , n28406 , n28411 );
buf ( n376017 , n359248 );
nand ( n28414 , n28412 , n376017 );
buf ( n376019 , n28414 );
buf ( n376020 , n376019 );
buf ( n28417 , n359225 );
not ( n28418 , n28417 );
buf ( n376023 , n28418 );
and ( n28420 , n376020 , n376023 );
not ( n28421 , n376020 );
buf ( n376026 , n28417 );
and ( n28423 , n28421 , n376026 );
nor ( n28424 , n28420 , n28423 );
buf ( n376029 , n28424 );
buf ( n376030 , n376029 );
xor ( n28427 , n28404 , n376030 );
buf ( n376032 , n28427 );
buf ( n376033 , n376032 );
buf ( n376034 , n372536 );
or ( n28431 , n376033 , n376034 );
buf ( n376036 , n28431 );
buf ( n376037 , n376036 );
not ( n28434 , n376037 );
buf ( n376039 , n372480 );
buf ( n376040 , n372495 );
xor ( n28437 , n376039 , n376040 );
buf ( n376042 , n372454 );
not ( n28439 , n376042 );
buf ( n376044 , n372475 );
not ( n28441 , n376044 );
or ( n28442 , n28439 , n28441 );
buf ( n376047 , n372454 );
buf ( n376048 , n372475 );
or ( n28445 , n376047 , n376048 );
buf ( n376050 , n372449 );
buf ( n376051 , n372441 );
or ( n28448 , n376050 , n376051 );
buf ( n376053 , n372436 );
buf ( n376054 , n372428 );
or ( n28451 , n376053 , n376054 );
buf ( n376056 , n372382 );
buf ( n376057 , n375232 );
buf ( n376058 , n347813 );
buf ( n376059 , n347906 );
not ( n28456 , n376059 );
buf ( n376061 , n28456 );
buf ( n376062 , n376061 );
xor ( n28459 , n376058 , n376062 );
buf ( n376064 , n347961 );
buf ( n376065 , n348033 );
xor ( n28462 , n376064 , n376065 );
buf ( n376067 , n347996 );
and ( n28464 , n28462 , n376067 );
or ( n28465 , n28464 , C0 );
buf ( n376070 , n28465 );
buf ( n376071 , n376070 );
and ( n28468 , n28459 , n376071 );
and ( n28469 , n376058 , n376062 );
or ( n28470 , n28468 , n28469 );
buf ( n376075 , n28470 );
buf ( n376076 , n376075 );
buf ( n376077 , n347906 );
xor ( n28474 , n376076 , n376077 );
buf ( n376079 , n375230 );
and ( n28476 , n28474 , n376079 );
and ( n28477 , n376076 , n376077 );
or ( n28478 , n28476 , n28477 );
buf ( n376083 , n28478 );
buf ( n376084 , n376083 );
xor ( n28481 , n376057 , n376084 );
buf ( n376086 , n372377 );
and ( n28483 , n28481 , n376086 );
and ( n28484 , n376057 , n376084 );
or ( n28485 , n28483 , n28484 );
buf ( n376090 , n28485 );
buf ( n376091 , n376090 );
xor ( n28488 , n376056 , n376091 );
buf ( n376093 , n372398 );
and ( n28490 , n28488 , n376093 );
and ( n28491 , n376056 , n376091 );
or ( n28492 , n28490 , n28491 );
buf ( n376097 , n28492 );
buf ( n376098 , n376097 );
not ( n28495 , n376098 );
buf ( n376100 , n28495 );
buf ( n376101 , n376100 );
buf ( n376102 , n372423 );
buf ( n376103 , n372403 );
nor ( n28500 , n376102 , n376103 );
buf ( n376105 , n28500 );
buf ( n376106 , n376105 );
or ( n28503 , n376101 , n376106 );
buf ( n376108 , n372423 );
buf ( n376109 , n372403 );
nand ( n28506 , n376108 , n376109 );
buf ( n376111 , n28506 );
buf ( n376112 , n376111 );
nand ( n28509 , n28503 , n376112 );
buf ( n376114 , n28509 );
buf ( n376115 , n376114 );
nand ( n28512 , n28451 , n376115 );
buf ( n376117 , n28512 );
buf ( n376118 , n376117 );
buf ( n376119 , n372436 );
buf ( n376120 , n372428 );
nand ( n28517 , n376119 , n376120 );
buf ( n376122 , n28517 );
buf ( n376123 , n376122 );
nand ( n28520 , n376118 , n376123 );
buf ( n376125 , n28520 );
buf ( n376126 , n376125 );
nand ( n28523 , n28448 , n376126 );
buf ( n376128 , n28523 );
buf ( n376129 , n376128 );
buf ( n376130 , n372441 );
buf ( n376131 , n372449 );
nand ( n28528 , n376130 , n376131 );
buf ( n376133 , n28528 );
buf ( n376134 , n376133 );
nand ( n28531 , n376129 , n376134 );
buf ( n376136 , n28531 );
buf ( n376137 , n376136 );
nand ( n28534 , n28445 , n376137 );
buf ( n376139 , n28534 );
buf ( n376140 , n376139 );
nand ( n28537 , n28442 , n376140 );
buf ( n376142 , n28537 );
buf ( n376143 , n376142 );
and ( n28540 , n28437 , n376143 );
and ( n28541 , n376039 , n376040 );
or ( n28542 , n28540 , n28541 );
buf ( n376147 , n28542 );
buf ( n376148 , n376147 );
not ( n28545 , n376148 );
buf ( n376150 , n28545 );
buf ( n376151 , n372531 );
buf ( n376152 , n372500 );
nor ( n28549 , n376151 , n376152 );
buf ( n376154 , n28549 );
or ( n28551 , n376150 , n376154 );
buf ( n376156 , n372531 );
buf ( n376157 , n372500 );
nand ( n28554 , n376156 , n376157 );
buf ( n376159 , n28554 );
nand ( n28556 , n28551 , n376159 );
buf ( n376161 , n28556 );
not ( n28558 , n376161 );
or ( n28559 , n28434 , n28558 );
buf ( n376164 , n376032 );
buf ( n376165 , n372536 );
nand ( n28562 , n376164 , n376165 );
buf ( n376167 , n28562 );
buf ( n376168 , n376167 );
nand ( n28565 , n28559 , n376168 );
buf ( n376170 , n28565 );
xor ( n28567 , n376006 , n376007 );
and ( n28568 , n28567 , n376030 );
and ( n28569 , n376006 , n376007 );
or ( n28570 , n28568 , n28569 );
buf ( n376175 , n28570 );
or ( n28572 , n376170 , n376175 );
not ( n28573 , n28572 );
or ( n28574 , n28401 , n28573 );
nand ( n28575 , n376170 , n376175 );
nand ( n28576 , n28574 , n28575 );
buf ( n376181 , n28576 );
nand ( n28578 , n28397 , n376181 );
buf ( n376183 , n28578 );
buf ( n376184 , n376183 );
buf ( n376185 , n374928 );
buf ( n376186 , n375999 );
nand ( n28583 , n376185 , n376186 );
buf ( n376188 , n28583 );
buf ( n376189 , n376188 );
nand ( n28586 , n376184 , n376189 );
buf ( n376191 , n28586 );
buf ( n376192 , n376191 );
not ( n28589 , n376192 );
or ( n28590 , n28366 , n28589 );
buf ( n376195 , n375960 );
buf ( n376196 , n374933 );
nand ( n28593 , n376195 , n376196 );
buf ( n376198 , n28593 );
buf ( n376199 , n376198 );
nand ( n28596 , n28590 , n376199 );
buf ( n376201 , n28596 );
buf ( n376202 , n376201 );
not ( n28599 , n376202 );
buf ( n376204 , n28599 );
buf ( n376205 , n376204 );
buf ( n376206 , n374815 );
xor ( n28603 , n375940 , n375943 );
and ( n28604 , n28603 , n375958 );
and ( n28605 , n375940 , n375943 );
or ( n28606 , n28604 , n28605 );
buf ( n376211 , n28606 );
buf ( n376212 , n376211 );
nor ( n28609 , n376206 , n376212 );
buf ( n376214 , n28609 );
buf ( n376215 , n376214 );
or ( n28612 , n376205 , n376215 );
buf ( n376217 , n374815 );
buf ( n376218 , n376211 );
nand ( n28615 , n376217 , n376218 );
buf ( n376220 , n28615 );
buf ( n376221 , n376220 );
nand ( n28618 , n28612 , n376221 );
buf ( n376223 , n28618 );
not ( n28620 , n376223 );
or ( n28621 , n28335 , n28620 );
buf ( n376226 , n374842 );
buf ( n376227 , n374820 );
nand ( n28624 , n376226 , n376227 );
buf ( n376229 , n28624 );
not ( n28626 , n376229 );
and ( n28627 , n28333 , n28626 );
and ( n28628 , n28330 , n374847 );
nor ( n28629 , n28627 , n28628 );
nand ( n28630 , n28621 , n28629 );
not ( n28631 , n28630 );
xor ( n28632 , n359909 , n359730 );
not ( n28633 , n12458 );
not ( n28634 , n11650 );
or ( n28635 , n28633 , n28634 );
buf ( n28636 , n360142 );
nand ( n28637 , n28635 , n28636 );
nand ( n28638 , n374241 , n374254 );
not ( n28639 , n28638 );
and ( n28640 , n28637 , n28639 );
not ( n28641 , n28637 );
and ( n28642 , n28641 , n28638 );
nor ( n28643 , n28640 , n28642 );
buf ( n28644 , n28643 );
and ( n28645 , n28632 , n28644 );
and ( n28646 , n359909 , n359730 );
or ( n28647 , n28645 , n28646 );
buf ( n376252 , n28647 );
not ( n28649 , n376252 );
buf ( n376254 , n28649 );
buf ( n376255 , n374866 );
not ( n28652 , n376255 );
buf ( n376257 , n28652 );
nand ( n28654 , n376254 , n376257 );
xor ( n28655 , n12504 , n357071 );
and ( n28656 , n28655 , n12470 );
and ( n28657 , n12504 , n357071 );
or ( n28658 , n28656 , n28657 );
not ( n28659 , n28658 );
xor ( n28660 , n359909 , n359730 );
xor ( n28661 , n28660 , n28644 );
buf ( n376266 , n28661 );
not ( n28663 , n376266 );
buf ( n376268 , n28663 );
nand ( n28665 , n28659 , n376268 );
and ( n28666 , n28654 , n28665 );
not ( n28667 , n28666 );
or ( n28668 , n28631 , n28667 );
nand ( n28669 , n28661 , n28658 );
not ( n28670 , n28669 );
and ( n28671 , n28654 , n28670 );
buf ( n376276 , n376257 );
not ( n28673 , n376276 );
buf ( n376278 , n28673 );
and ( n28675 , n28647 , n376278 );
nor ( n28676 , n28671 , n28675 );
nand ( n28677 , n28668 , n28676 );
buf ( n376282 , n28677 );
not ( n28679 , n376282 );
or ( n28680 , n28320 , n28679 );
buf ( n376285 , n28310 );
buf ( n376286 , n375919 );
not ( n28683 , n376286 );
buf ( n376288 , n28683 );
buf ( n376289 , n376288 );
nand ( n28686 , n376285 , n376289 );
buf ( n376291 , n28686 );
buf ( n376292 , n376291 );
nand ( n28689 , n28680 , n376292 );
buf ( n376294 , n28689 );
buf ( n376295 , n376294 );
not ( n28692 , n376295 );
or ( n28693 , n28308 , n28692 );
buf ( n376298 , n374909 );
buf ( n376299 , n28300 );
nand ( n28696 , n376298 , n376299 );
buf ( n376301 , n28696 );
buf ( n376302 , n376301 );
nand ( n28699 , n28693 , n376302 );
buf ( n376304 , n28699 );
buf ( n376305 , n376304 );
not ( n28702 , n376305 );
xor ( n28703 , n362109 , n361993 );
xor ( n28704 , n28703 , n28270 );
buf ( n376309 , n28704 );
not ( n28706 , n376309 );
buf ( n376311 , n374914 );
not ( n28708 , n376311 );
buf ( n376313 , n28708 );
buf ( n376314 , n376313 );
nand ( n28711 , n28706 , n376314 );
buf ( n376316 , n28711 );
buf ( n376317 , n376316 );
not ( n28714 , n376317 );
or ( n28715 , n28702 , n28714 );
buf ( n376320 , n374914 );
buf ( n376321 , n28704 );
nand ( n28718 , n376320 , n376321 );
buf ( n376323 , n28718 );
buf ( n376324 , n376323 );
nand ( n28721 , n28715 , n376324 );
buf ( n376326 , n28721 );
buf ( n376327 , n376326 );
and ( n28724 , n28279 , n376327 );
and ( n28725 , n375878 , n375882 );
or ( n28726 , n28724 , n28725 );
buf ( n376331 , n28726 );
buf ( n376332 , n376331 );
xor ( n28729 , n375860 , n376332 );
xor ( n28730 , n362813 , n362807 );
xor ( n28731 , n28730 , n375822 );
buf ( n376336 , n28731 );
and ( n28733 , n28729 , n376336 );
and ( n28734 , n375860 , n376332 );
or ( n28735 , n28733 , n28734 );
buf ( n376340 , n28735 );
buf ( n376341 , n376340 );
and ( n28738 , n28224 , n376341 );
and ( n28739 , n375826 , n375827 );
or ( n28740 , n28738 , n28739 );
buf ( n376345 , n28740 );
buf ( n376346 , n376345 );
and ( n28743 , n28197 , n376346 );
and ( n28744 , n375799 , n375800 );
or ( n28745 , n28743 , n28744 );
buf ( n376350 , n28745 );
buf ( n376351 , n376350 );
and ( n28748 , n28194 , n376351 );
and ( n28749 , n375793 , n375797 );
or ( n28750 , n28748 , n28749 );
buf ( n376355 , n28750 );
buf ( n376356 , n376355 );
and ( n28753 , n28188 , n376356 );
and ( n28754 , n375768 , n375791 );
or ( n28755 , n28753 , n28754 );
buf ( n376360 , n28755 );
buf ( n376361 , n376360 );
buf ( n376362 , n364157 );
buf ( n376363 , n364164 );
xor ( n28760 , n376362 , n376363 );
buf ( n376365 , n375745 );
buf ( n376366 , n375474 );
buf ( n376367 , n375479 );
nor ( n28764 , n376366 , n376367 );
buf ( n376369 , n28764 );
buf ( n376370 , n376369 );
nor ( n28767 , n376365 , n376370 );
buf ( n376372 , n28767 );
buf ( n376373 , n376372 );
buf ( n28770 , n376373 );
buf ( n376375 , n28770 );
not ( n28772 , n376375 );
not ( n28773 , n27903 );
or ( n28774 , n28772 , n28773 );
buf ( n376379 , n375748 );
not ( n28776 , n376379 );
buf ( n376381 , n27906 );
not ( n28778 , n376381 );
and ( n28779 , n28776 , n28778 );
buf ( n376384 , n375756 );
not ( n28781 , n376384 );
buf ( n376386 , n28781 );
buf ( n376387 , n376386 );
nor ( n28784 , n28779 , n376387 );
buf ( n376389 , n28784 );
nand ( n28786 , n28774 , n376389 );
not ( n28787 , n4362 );
not ( n28788 , n598 );
not ( n28789 , n25741 );
or ( n28790 , n28788 , n28789 );
nand ( n28791 , n25700 , n347312 );
nand ( n28792 , n28790 , n28791 );
not ( n28793 , n28792 );
or ( n28794 , n28787 , n28793 );
nand ( n28795 , n27945 , n4443 );
nand ( n28796 , n28794 , n28795 );
buf ( n376401 , n28796 );
buf ( n376402 , n349035 );
not ( n28799 , n376402 );
buf ( n376404 , n594 );
not ( n28801 , n376404 );
buf ( n376406 , n360099 );
not ( n28803 , n376406 );
or ( n28804 , n28801 , n28803 );
buf ( n376409 , n12420 );
buf ( n376410 , n348975 );
nand ( n28807 , n376409 , n376410 );
buf ( n376412 , n28807 );
buf ( n376413 , n376412 );
nand ( n28810 , n28804 , n376413 );
buf ( n376415 , n28810 );
buf ( n376416 , n376415 );
not ( n28813 , n376416 );
or ( n28814 , n28799 , n28813 );
and ( n28815 , n9636 , n349153 );
buf ( n376420 , n9636 );
buf ( n376421 , n349160 );
nor ( n28818 , n376420 , n376421 );
buf ( n376423 , n28818 );
nor ( n28820 , n28815 , n376423 );
buf ( n376425 , n28820 );
nand ( n28822 , n28814 , n376425 );
buf ( n376427 , n28822 );
buf ( n376428 , n376427 );
xor ( n28825 , n376401 , n376428 );
buf ( n376430 , n351924 );
not ( n28827 , n376430 );
buf ( n376432 , n27960 );
not ( n28829 , n376432 );
or ( n28830 , n28827 , n28829 );
buf ( n376435 , n600 );
not ( n28832 , n376435 );
buf ( n376437 , n372582 );
not ( n28834 , n376437 );
or ( n28835 , n28832 , n28834 );
buf ( n376440 , n374705 );
buf ( n376441 , n6460 );
nand ( n28838 , n376440 , n376441 );
buf ( n376443 , n28838 );
buf ( n376444 , n376443 );
nand ( n28841 , n28835 , n376444 );
buf ( n376446 , n28841 );
buf ( n376447 , n376446 );
buf ( n376448 , n1722 );
nand ( n28845 , n376447 , n376448 );
buf ( n376450 , n28845 );
buf ( n376451 , n376450 );
nand ( n28848 , n28830 , n376451 );
buf ( n376453 , n28848 );
buf ( n376454 , n376453 );
xor ( n28851 , n28825 , n376454 );
buf ( n376456 , n28851 );
buf ( n376457 , n376456 );
xor ( n28854 , n375600 , n375641 );
and ( n28855 , n28854 , n375656 );
and ( n28856 , n375600 , n375641 );
or ( n28857 , n28855 , n28856 );
buf ( n376462 , n28857 );
buf ( n376463 , n376462 );
xor ( n28860 , n376457 , n376463 );
buf ( n376465 , n354113 );
not ( n28862 , n376465 );
buf ( n376467 , n602 );
buf ( n376468 , n17009 );
and ( n28865 , n376467 , n376468 );
not ( n28866 , n376467 );
buf ( n376471 , n373494 );
and ( n28868 , n28866 , n376471 );
nor ( n28869 , n28865 , n28868 );
buf ( n376474 , n28869 );
buf ( n376475 , n376474 );
not ( n28872 , n376475 );
or ( n28873 , n28862 , n28872 );
buf ( n376478 , n27137 );
buf ( n376479 , n373187 );
and ( n28876 , n376478 , n376479 );
buf ( n376481 , n27134 );
buf ( n376482 , n373176 );
and ( n28879 , n376481 , n376482 );
nor ( n28880 , n28876 , n28879 );
buf ( n376485 , n28880 );
buf ( n376486 , n376485 );
nand ( n28883 , n28873 , n376486 );
buf ( n376488 , n28883 );
buf ( n376489 , n376488 );
xor ( n28886 , n375603 , n375620 );
and ( n28887 , n28886 , n375638 );
and ( n28888 , n375603 , n375620 );
or ( n28889 , n28887 , n28888 );
buf ( n376494 , n28889 );
buf ( n376495 , n376494 );
xor ( n28892 , n376489 , n376495 );
buf ( n376497 , n607 );
not ( n28894 , n376497 );
buf ( n376499 , n606 );
not ( n28896 , n14501 );
not ( n28897 , n16814 );
not ( n28898 , n16855 );
and ( n28899 , n28896 , n28897 , n28898 );
nand ( n28900 , n16957 , n16958 );
not ( n28901 , n28900 );
and ( n28902 , n23381 , n23383 );
not ( n28903 , n23381 );
and ( n28904 , n28903 , n23382 );
nor ( n28905 , n28902 , n28904 );
not ( n28906 , n28905 );
nand ( n28907 , n28899 , n28901 , n28906 );
or ( n28908 , n14501 , n16855 );
not ( n28909 , n28897 );
or ( n28910 , n28908 , n28909 );
nand ( n28911 , n28910 , n28905 );
nand ( n28912 , n28900 , n28905 );
nand ( n28913 , n28907 , n28911 , n28912 );
buf ( n376518 , n28913 );
buf ( n28915 , n376518 );
buf ( n376520 , n28915 );
buf ( n376521 , n376520 );
and ( n28918 , n376499 , n376521 );
not ( n28919 , n376499 );
buf ( n376524 , n376520 );
not ( n28921 , n376524 );
buf ( n376526 , n28921 );
buf ( n376527 , n376526 );
and ( n28924 , n28919 , n376527 );
nor ( n28925 , n28918 , n28924 );
buf ( n376530 , n28925 );
buf ( n376531 , n376530 );
not ( n28928 , n376531 );
or ( n28929 , n28894 , n28928 );
buf ( n376534 , n375707 );
buf ( n376535 , n357376 );
nand ( n28932 , n376534 , n376535 );
buf ( n376537 , n28932 );
buf ( n376538 , n376537 );
nand ( n28935 , n28929 , n376538 );
buf ( n376540 , n28935 );
buf ( n376541 , n376540 );
xor ( n28938 , n28892 , n376541 );
buf ( n376543 , n28938 );
buf ( n376544 , n376543 );
xor ( n28941 , n28860 , n376544 );
buf ( n376546 , n28941 );
buf ( n376547 , n376546 );
xor ( n28944 , n375668 , n375717 );
and ( n28945 , n28944 , n375724 );
and ( n28946 , n375668 , n375717 );
or ( n28947 , n28945 , n28946 );
buf ( n376552 , n28947 );
buf ( n376553 , n376552 );
xor ( n28950 , n376547 , n376553 );
xor ( n28951 , n375674 , n375680 );
and ( n28952 , n28951 , n375714 );
and ( n28953 , n375674 , n375680 );
or ( n28954 , n28952 , n28953 );
buf ( n376559 , n28954 );
buf ( n376560 , n376559 );
buf ( n376561 , n6600 );
not ( n28958 , n376561 );
and ( n28959 , n604 , n375435 );
not ( n28960 , n604 );
buf ( n376565 , n27828 );
buf ( n28962 , n376565 );
buf ( n376567 , n28962 );
and ( n28964 , n28960 , n376567 );
or ( n28965 , n28959 , n28964 );
buf ( n376570 , n28965 );
not ( n28967 , n376570 );
or ( n28968 , n28958 , n28967 );
buf ( n376573 , n28044 );
buf ( n376574 , n355075 );
nand ( n28971 , n376573 , n376574 );
buf ( n376576 , n28971 );
buf ( n376577 , n376576 );
nand ( n28974 , n28968 , n376577 );
buf ( n376579 , n28974 );
buf ( n376580 , n376579 );
buf ( n376581 , n7359 );
buf ( n376582 , n592 );
and ( n28979 , n376581 , n376582 );
buf ( n376584 , n28979 );
buf ( n376585 , n376584 );
buf ( n376586 , n348946 );
not ( n28983 , n376586 );
buf ( n376588 , n592 );
not ( n28985 , n376588 );
buf ( n376590 , n357355 );
not ( n28987 , n376590 );
or ( n28988 , n28985 , n28987 );
buf ( n376593 , n9664 );
buf ( n376594 , n348910 );
nand ( n28991 , n376593 , n376594 );
buf ( n376596 , n28991 );
buf ( n376597 , n376596 );
nand ( n28994 , n28988 , n376597 );
buf ( n376599 , n28994 );
buf ( n376600 , n376599 );
not ( n28997 , n376600 );
or ( n28998 , n28983 , n28997 );
buf ( n376603 , n375038 );
buf ( n376604 , n28005 );
nand ( n29001 , n376603 , n376604 );
buf ( n376606 , n29001 );
buf ( n376607 , n376606 );
nand ( n29004 , n28998 , n376607 );
buf ( n376609 , n29004 );
buf ( n376610 , n376609 );
xor ( n29007 , n376585 , n376610 );
buf ( n376612 , n347319 );
not ( n29009 , n376612 );
not ( n29010 , n596 );
not ( n29011 , n25863 );
or ( n29012 , n29010 , n29011 );
buf ( n376617 , n25627 );
buf ( n376618 , n348865 );
nand ( n29015 , n376617 , n376618 );
buf ( n376620 , n29015 );
nand ( n29017 , n29012 , n376620 );
buf ( n376622 , n29017 );
not ( n29019 , n376622 );
or ( n29020 , n29009 , n29019 );
nand ( n29021 , n27912 , n372772 );
buf ( n376626 , n29021 );
nand ( n29023 , n29020 , n376626 );
buf ( n376628 , n29023 );
buf ( n376629 , n376628 );
xor ( n29026 , n29007 , n376629 );
buf ( n376631 , n29026 );
buf ( n376632 , n376631 );
xor ( n29029 , n376580 , n376632 );
xor ( n29030 , n375528 , n375557 );
and ( n29031 , n29030 , n375569 );
and ( n29032 , n375528 , n375557 );
or ( n29033 , n29031 , n29032 );
buf ( n376638 , n29033 );
buf ( n376639 , n376638 );
xor ( n29036 , n29029 , n376639 );
buf ( n376641 , n29036 );
buf ( n376642 , n376641 );
xor ( n29039 , n376560 , n376642 );
xor ( n29040 , n375572 , n375578 );
and ( n29041 , n29040 , n375659 );
and ( n29042 , n375572 , n375578 );
or ( n29043 , n29041 , n29042 );
buf ( n376648 , n29043 );
buf ( n376649 , n376648 );
xor ( n29046 , n29039 , n376649 );
buf ( n376651 , n29046 );
buf ( n376652 , n376651 );
xor ( n29049 , n28950 , n376652 );
buf ( n376654 , n29049 );
buf ( n376655 , n376654 );
not ( n29052 , n376655 );
xor ( n29053 , n375662 , n375727 );
and ( n29054 , n29053 , n375734 );
and ( n29055 , n375662 , n375727 );
or ( n29056 , n29054 , n29055 );
buf ( n376661 , n29056 );
buf ( n376662 , n376661 );
not ( n29059 , n376662 );
buf ( n376664 , n29059 );
buf ( n376665 , n376664 );
nand ( n29062 , n29052 , n376665 );
buf ( n376667 , n29062 );
buf ( n376668 , n376667 );
buf ( n29065 , n376668 );
buf ( n376670 , n29065 );
buf ( n376671 , n376654 );
buf ( n376672 , n376661 );
nand ( n29069 , n376671 , n376672 );
buf ( n376674 , n29069 );
nand ( n29071 , n376670 , n376674 );
not ( n29072 , n29071 );
and ( n29073 , n28786 , n29072 );
not ( n29074 , n28786 );
and ( n29075 , n29074 , n29071 );
nor ( n29076 , n29073 , n29075 );
buf ( n29077 , n29076 );
buf ( n29078 , n29077 );
buf ( n376683 , n29078 );
xor ( n29080 , n28760 , n376683 );
buf ( n376685 , n29080 );
buf ( n376686 , n376685 );
not ( n29083 , n376686 );
buf ( n376688 , n29083 );
buf ( n376689 , n376688 );
xor ( n29086 , n375237 , n375238 );
and ( n29087 , n29086 , n375765 );
and ( n29088 , n375237 , n375238 );
or ( n29089 , n29087 , n29088 );
buf ( n376694 , n29089 );
buf ( n376695 , n376694 );
not ( n29092 , n376695 );
buf ( n376697 , n29092 );
buf ( n376698 , n376697 );
nand ( n29095 , n376689 , n376698 );
buf ( n376700 , n29095 );
buf ( n376701 , n376700 );
and ( n29098 , n376361 , n376701 );
buf ( n376703 , n376688 );
buf ( n376704 , n376697 );
nor ( n29101 , n376703 , n376704 );
buf ( n376706 , n29101 );
buf ( n376707 , n376706 );
nor ( n29104 , n29098 , n376707 );
buf ( n376709 , n29104 );
buf ( n376710 , n376709 );
buf ( n376711 , n376360 );
buf ( n376712 , n376706 );
or ( n29109 , n376711 , n376712 );
buf ( n376714 , n376700 );
nand ( n29111 , n29109 , n376714 );
buf ( n376716 , n29111 );
buf ( n376717 , n376716 );
not ( n29114 , n376717 );
buf ( n376719 , n29114 );
buf ( n376720 , n376719 );
xor ( n29117 , n376362 , n376363 );
and ( n29118 , n29117 , n376683 );
and ( n29119 , n376362 , n376363 );
or ( n29120 , n29118 , n29119 );
buf ( n376725 , n29120 );
buf ( n376726 , n376725 );
buf ( n376727 , n375236 );
xor ( n29124 , n376726 , n376727 );
buf ( n376729 , n29124 );
buf ( n376730 , n376729 );
and ( n29127 , n376730 , n376720 );
not ( n29128 , n376730 );
and ( n29129 , n29128 , n376710 );
nor ( n29130 , n29127 , n29129 );
buf ( n376735 , n29130 );
buf ( n376736 , n376697 );
buf ( n376737 , n376685 );
and ( n29134 , n376736 , n376737 );
not ( n29135 , n376736 );
buf ( n376740 , n376688 );
and ( n29137 , n29135 , n376740 );
nor ( n29138 , n29134 , n29137 );
buf ( n376743 , n29138 );
buf ( n376744 , n376743 );
buf ( n376745 , n376360 );
buf ( n376746 , n376743 );
buf ( n376747 , n376360 );
not ( n29144 , n376744 );
not ( n29145 , n376745 );
or ( n29146 , n29144 , n29145 );
or ( n29147 , n376746 , n376747 );
nand ( n29148 , n29146 , n29147 );
buf ( n376753 , n29148 );
xor ( n29150 , n375768 , n375791 );
xor ( n29151 , n29150 , n376356 );
buf ( n376756 , n29151 );
xor ( n29153 , n375793 , n375797 );
xor ( n29154 , n29153 , n376351 );
buf ( n376759 , n29154 );
xor ( n29156 , n375799 , n375800 );
xor ( n29157 , n29156 , n376346 );
buf ( n376762 , n29157 );
xor ( n29159 , n375826 , n375827 );
xor ( n29160 , n29159 , n376341 );
buf ( n376765 , n29160 );
buf ( n376766 , n376223 );
buf ( n376767 , n374842 );
buf ( n376768 , n375929 );
and ( n29165 , n376767 , n376768 );
not ( n29166 , n376767 );
buf ( n376771 , n374820 );
and ( n29168 , n29166 , n376771 );
nor ( n29169 , n29165 , n29168 );
buf ( n376774 , n29169 );
buf ( n376775 , n376774 );
buf ( n376776 , n376774 );
buf ( n376777 , n376223 );
not ( n29174 , n376766 );
not ( n29175 , n376775 );
or ( n29176 , n29174 , n29175 );
or ( n29177 , n376776 , n376777 );
nand ( n29178 , n29176 , n29177 );
buf ( n376783 , n29178 );
buf ( n376784 , n376204 );
buf ( n376785 , n376201 );
buf ( n376786 , n374815 );
buf ( n376787 , n376211 );
xor ( n29184 , n376786 , n376787 );
buf ( n376789 , n29184 );
buf ( n376790 , n376789 );
and ( n29187 , n376790 , n376785 );
not ( n29188 , n376790 );
and ( n29189 , n29188 , n376784 );
nor ( n29190 , n29187 , n29189 );
buf ( n376795 , n29190 );
buf ( n376796 , n375960 );
buf ( n376797 , n375965 );
and ( n29194 , n376796 , n376797 );
not ( n29195 , n376796 );
buf ( n376800 , n374933 );
and ( n29197 , n29195 , n376800 );
nor ( n29198 , n29194 , n29197 );
buf ( n376803 , n29198 );
buf ( n376804 , n376803 );
buf ( n376805 , n376191 );
buf ( n376806 , n376803 );
buf ( n376807 , n376191 );
not ( n29204 , n376804 );
not ( n29205 , n376805 );
or ( n29206 , n29204 , n29205 );
or ( n29207 , n376806 , n376807 );
nand ( n29208 , n29206 , n29207 );
buf ( n376813 , n29208 );
buf ( n376814 , n28576 );
buf ( n376815 , n374928 );
buf ( n376816 , n375999 );
xnor ( n29213 , n376815 , n376816 );
buf ( n376818 , n29213 );
buf ( n376819 , n376818 );
buf ( n376820 , n376818 );
buf ( n376821 , n28576 );
not ( n29218 , n376814 );
not ( n29219 , n376819 );
or ( n29220 , n29218 , n29219 );
or ( n29221 , n376820 , n376821 );
nand ( n29222 , n29220 , n29221 );
buf ( n376827 , n29222 );
buf ( n376828 , n376004 );
buf ( n376829 , n376175 );
xnor ( n29226 , n376828 , n376829 );
buf ( n376831 , n29226 );
buf ( n376832 , n376831 );
buf ( n376833 , n376170 );
buf ( n376834 , n376170 );
buf ( n376835 , n376831 );
not ( n29232 , n376832 );
not ( n29233 , n376833 );
or ( n29234 , n29232 , n29233 );
or ( n29235 , n376834 , n376835 );
nand ( n29236 , n29234 , n29235 );
buf ( n376841 , n29236 );
buf ( n376842 , n376150 );
buf ( n376843 , n376147 );
buf ( n376844 , n372531 );
buf ( n376845 , n372500 );
xor ( n29242 , n376844 , n376845 );
buf ( n376847 , n29242 );
buf ( n376848 , n376847 );
and ( n29245 , n376848 , n376843 );
not ( n29246 , n376848 );
and ( n29247 , n29246 , n376842 );
nor ( n29248 , n29245 , n29247 );
buf ( n376853 , n29248 );
xor ( n29250 , n376039 , n376040 );
xor ( n29251 , n29250 , n376143 );
buf ( n376856 , n29251 );
buf ( n376857 , n372475 );
buf ( n376858 , n372454 );
xor ( n29255 , n376857 , n376858 );
buf ( n376860 , n29255 );
buf ( n376861 , n376860 );
buf ( n376862 , n376136 );
xor ( n29259 , n376861 , n376862 );
buf ( n376864 , n29259 );
buf ( n376865 , n372449 );
buf ( n376866 , n372441 );
xor ( n29263 , n376865 , n376866 );
buf ( n376868 , n29263 );
buf ( n376869 , n376868 );
buf ( n376870 , n376125 );
xor ( n29267 , n376869 , n376870 );
buf ( n376872 , n29267 );
buf ( n376873 , n372436 );
buf ( n376874 , n372428 );
xor ( n29271 , n376873 , n376874 );
buf ( n376876 , n29271 );
buf ( n376877 , n376876 );
buf ( n376878 , n376114 );
xor ( n29275 , n376877 , n376878 );
buf ( n376880 , n29275 );
buf ( n376881 , n376100 );
buf ( n376882 , n376097 );
buf ( n376883 , n372423 );
buf ( n376884 , n372403 );
xor ( n29281 , n376883 , n376884 );
buf ( n376886 , n29281 );
buf ( n376887 , n376886 );
and ( n29284 , n376887 , n376882 );
not ( n29285 , n376887 );
and ( n29286 , n29285 , n376881 );
nor ( n29287 , n29284 , n29286 );
buf ( n376892 , n29287 );
xor ( n29289 , n376056 , n376091 );
xor ( n29290 , n29289 , n376093 );
buf ( n376895 , n29290 );
xor ( n29292 , n376057 , n376084 );
xor ( n29293 , n29292 , n376086 );
buf ( n376898 , n29293 );
xor ( n29295 , n376076 , n376077 );
xor ( n29296 , n29295 , n376079 );
buf ( n376901 , n29296 );
xor ( n29298 , n376058 , n376062 );
xor ( n29299 , n29298 , n376071 );
buf ( n376904 , n29299 );
buf ( n376905 , n28332 );
buf ( n376906 , n374847 );
buf ( n376907 , n28330 );
and ( n29304 , n376907 , n376906 );
not ( n29305 , n376907 );
and ( n29306 , n29305 , n376905 );
nor ( n29307 , n29304 , n29306 );
buf ( n376912 , n29307 );
buf ( n376913 , n376268 );
buf ( n376914 , n28661 );
buf ( n376915 , n28658 );
and ( n29312 , n376915 , n376914 );
not ( n29313 , n376915 );
and ( n29314 , n29313 , n376913 );
nor ( n29315 , n29312 , n29314 );
buf ( n376920 , n29315 );
buf ( n376921 , n376313 );
buf ( n376922 , n374914 );
buf ( n376923 , n28704 );
and ( n29320 , n376923 , n376922 );
not ( n29321 , n376923 );
and ( n29322 , n29321 , n376921 );
nor ( n29323 , n29320 , n29322 );
buf ( n376928 , n29323 );
buf ( n376929 , n375907 );
buf ( n376930 , n28300 );
buf ( n376931 , n374909 );
and ( n29328 , n376931 , n376930 );
not ( n29329 , n376931 );
and ( n29330 , n29329 , n376929 );
nor ( n29331 , n29328 , n29330 );
buf ( n376936 , n29331 );
buf ( n376937 , n375919 );
buf ( n376938 , n376288 );
buf ( n376939 , n28310 );
and ( n29336 , n376939 , n376938 );
not ( n29337 , n376939 );
and ( n29338 , n29337 , n376937 );
nor ( n29339 , n29336 , n29338 );
buf ( n376944 , n29339 );
buf ( n376945 , n376254 );
buf ( n376946 , n28647 );
buf ( n376947 , n376278 );
and ( n29344 , n376947 , n376946 );
not ( n29345 , n376947 );
and ( n29346 , n29345 , n376945 );
nor ( n29347 , n29344 , n29346 );
buf ( n376952 , n29347 );
not ( n29349 , n375932 );
not ( n29350 , n376223 );
or ( n29351 , n29349 , n29350 );
nand ( n29352 , n29351 , n376229 );
buf ( n376957 , n29352 );
buf ( n376958 , n376912 );
xor ( n29355 , n376957 , n376958 );
buf ( n376960 , n29355 );
buf ( n376961 , n28630 );
buf ( n376962 , n376920 );
xor ( n29359 , n376961 , n376962 );
buf ( n376964 , n29359 );
not ( n29361 , n28665 );
not ( n29362 , n28630 );
or ( n29363 , n29361 , n29362 );
nand ( n29364 , n29363 , n28669 );
buf ( n376969 , n29364 );
buf ( n376970 , n376952 );
xor ( n29367 , n376969 , n376970 );
buf ( n376972 , n29367 );
buf ( n376973 , n28677 );
buf ( n376974 , n376944 );
xor ( n29371 , n376973 , n376974 );
buf ( n376976 , n29371 );
buf ( n376977 , n376294 );
buf ( n376978 , n376936 );
xor ( n29375 , n376977 , n376978 );
buf ( n376980 , n29375 );
buf ( n376981 , n376304 );
buf ( n376982 , n376928 );
xor ( n29379 , n376981 , n376982 );
buf ( n376984 , n29379 );
buf ( n376985 , n364834 );
not ( n29382 , n376985 );
buf ( n376987 , n576 );
not ( n29384 , n376987 );
buf ( n376989 , n365897 );
buf ( n29386 , n376989 );
buf ( n376991 , n29386 );
buf ( n376992 , n376991 );
not ( n29389 , n376992 );
buf ( n376994 , n29389 );
buf ( n376995 , n376994 );
not ( n29392 , n376995 );
or ( n29393 , n29384 , n29392 );
buf ( n376998 , n376991 );
buf ( n376999 , n354303 );
nand ( n29396 , n376998 , n376999 );
buf ( n377001 , n29396 );
buf ( n377002 , n377001 );
nand ( n29399 , n29393 , n377002 );
buf ( n377004 , n29399 );
buf ( n377005 , n377004 );
not ( n29402 , n377005 );
or ( n29403 , n29382 , n29402 );
buf ( n377008 , n576 );
not ( n29405 , n377008 );
buf ( n377010 , n27128 );
not ( n29407 , n377010 );
or ( n29408 , n29405 , n29407 );
buf ( n377013 , n17933 );
buf ( n377014 , n354303 );
nand ( n29411 , n377013 , n377014 );
buf ( n377016 , n29411 );
buf ( n377017 , n377016 );
nand ( n29414 , n29408 , n377017 );
buf ( n377019 , n29414 );
buf ( n377020 , n377019 );
buf ( n377021 , n17182 );
buf ( n29418 , n377021 );
buf ( n377023 , n29418 );
buf ( n377024 , n377023 );
nand ( n29421 , n377020 , n377024 );
buf ( n377026 , n29421 );
buf ( n377027 , n377026 );
nand ( n29424 , n29403 , n377027 );
buf ( n377029 , n29424 );
buf ( n377030 , n377029 );
buf ( n377031 , n17082 );
buf ( n377032 , n578 );
not ( n29429 , n377032 );
buf ( n377034 , n365892 );
not ( n29431 , n377034 );
buf ( n377036 , n29431 );
buf ( n377037 , n377036 );
not ( n29434 , n377037 );
or ( n29435 , n29429 , n29434 );
buf ( n377040 , n377036 );
not ( n29437 , n377040 );
buf ( n377042 , n29437 );
buf ( n377043 , n377042 );
buf ( n377044 , n364727 );
nand ( n29441 , n377043 , n377044 );
buf ( n377046 , n29441 );
buf ( n377047 , n377046 );
nand ( n29444 , n29435 , n377047 );
buf ( n377049 , n29444 );
buf ( n377050 , n377049 );
nand ( n29447 , n377031 , n377050 );
buf ( n377052 , n29447 );
not ( n29449 , n578 );
buf ( n377054 , n16815 );
buf ( n29451 , n377054 );
buf ( n377056 , n29451 );
buf ( n377057 , n377056 );
not ( n29454 , n377057 );
buf ( n377059 , n29454 );
not ( n29456 , n377059 );
or ( n29457 , n29449 , n29456 );
buf ( n377062 , n377056 );
buf ( n377063 , n364727 );
nand ( n29460 , n377062 , n377063 );
buf ( n377065 , n29460 );
nand ( n29462 , n29457 , n377065 );
nand ( n29463 , n29462 , n17037 );
nand ( n29464 , n377052 , n29463 );
buf ( n377069 , n29464 );
xor ( n29466 , n377030 , n377069 );
buf ( n377071 , n17905 );
buf ( n29468 , n377071 );
buf ( n377073 , n29468 );
buf ( n377074 , n377073 );
not ( n29471 , n377074 );
buf ( n377076 , n29471 );
buf ( n377077 , n377076 );
not ( n29474 , n377077 );
buf ( n377079 , n576 );
nand ( n29476 , n29474 , n377079 );
buf ( n377081 , n29476 );
buf ( n377082 , n377081 );
xor ( n29479 , n29466 , n377082 );
buf ( n377084 , n29479 );
buf ( n377085 , n377084 );
buf ( n377086 , n17209 );
not ( n29483 , n377086 );
buf ( n377088 , n580 );
not ( n29485 , n377088 );
not ( n29486 , n16799 );
not ( n29487 , n29486 );
not ( n29488 , n29487 );
buf ( n377093 , n29488 );
not ( n29490 , n377093 );
or ( n29491 , n29485 , n29490 );
buf ( n377096 , n29487 );
buf ( n377097 , n364896 );
nand ( n29494 , n377096 , n377097 );
buf ( n377099 , n29494 );
buf ( n377100 , n377099 );
nand ( n29497 , n29491 , n377100 );
buf ( n377102 , n29497 );
buf ( n377103 , n377102 );
not ( n29500 , n377103 );
or ( n29501 , n29483 , n29500 );
buf ( n377106 , n580 );
not ( n29503 , n377106 );
buf ( n377108 , n364664 );
not ( n29505 , n377108 );
or ( n29506 , n29503 , n29505 );
buf ( n377111 , n364661 );
buf ( n377112 , n364896 );
nand ( n29509 , n377111 , n377112 );
buf ( n377114 , n29509 );
buf ( n377115 , n377114 );
nand ( n29512 , n29506 , n377115 );
buf ( n377117 , n29512 );
buf ( n377118 , n377117 );
buf ( n377119 , n17230 );
nand ( n29516 , n377118 , n377119 );
buf ( n377121 , n29516 );
buf ( n377122 , n377121 );
nand ( n29519 , n29501 , n377122 );
buf ( n377124 , n29519 );
buf ( n377125 , n377124 );
buf ( n377126 , n364834 );
not ( n29523 , n377126 );
buf ( n377128 , n377019 );
not ( n29525 , n377128 );
or ( n29526 , n29523 , n29525 );
and ( n377131 , n377076 , n576 );
not ( n29528 , n377076 );
and ( n377133 , n29528 , n354303 );
or ( n29530 , n377131 , n377133 );
buf ( n377135 , n29530 );
buf ( n377136 , n377023 );
nand ( n377137 , n377135 , n377136 );
buf ( n377138 , n377137 );
buf ( n377139 , n377138 );
nand ( n29536 , n29526 , n377139 );
buf ( n377141 , n29536 );
buf ( n377142 , n377141 );
buf ( n377143 , n365661 );
buf ( n377144 , n576 );
and ( n377145 , n377143 , n377144 );
buf ( n377146 , n377145 );
buf ( n377147 , n377146 );
xor ( n29544 , n377142 , n377147 );
or ( n377149 , n17133 , n365151 );
buf ( n377150 , n582 );
not ( n377151 , n377150 );
buf ( n377152 , n364664 );
not ( n377153 , n377152 );
or ( n29550 , n377151 , n377153 );
buf ( n377155 , n364661 );
buf ( n377156 , n364797 );
nand ( n377157 , n377155 , n377156 );
buf ( n377158 , n377157 );
buf ( n377159 , n377158 );
nand ( n29556 , n29550 , n377159 );
buf ( n377161 , n29556 );
nand ( n29558 , n377149 , n377161 );
buf ( n377163 , n29558 );
and ( n29560 , n29544 , n377163 );
and ( n377165 , n377142 , n377147 );
or ( n29562 , n29560 , n377165 );
buf ( n377167 , n29562 );
buf ( n377168 , n377167 );
xor ( n377169 , n377125 , n377168 );
buf ( n377170 , n17037 );
not ( n377171 , n377170 );
buf ( n377172 , n377049 );
not ( n377173 , n377172 );
or ( n29570 , n377171 , n377173 );
buf ( n377175 , n578 );
not ( n29572 , n377175 );
buf ( n377177 , n375155 );
not ( n29574 , n377177 );
or ( n377179 , n29572 , n29574 );
buf ( n377180 , n376991 );
buf ( n377181 , n364727 );
nand ( n29578 , n377180 , n377181 );
buf ( n377183 , n29578 );
buf ( n377184 , n377183 );
nand ( n377185 , n377179 , n377184 );
buf ( n377186 , n377185 );
buf ( n377187 , n377186 );
buf ( n377188 , n17082 );
nand ( n377189 , n377187 , n377188 );
buf ( n377190 , n377189 );
buf ( n377191 , n377190 );
nand ( n29588 , n29570 , n377191 );
buf ( n377193 , n29588 );
buf ( n377194 , n377193 );
buf ( n377195 , n17230 );
not ( n29592 , n377195 );
buf ( n377197 , n377102 );
not ( n29594 , n377197 );
or ( n377199 , n29592 , n29594 );
buf ( n377200 , n580 );
not ( n377201 , n377200 );
buf ( n377202 , n28909 );
not ( n377203 , n377202 );
or ( n29600 , n377201 , n377203 );
buf ( n377205 , n377056 );
buf ( n377206 , n364896 );
nand ( n377207 , n377205 , n377206 );
buf ( n377208 , n377207 );
buf ( n377209 , n377208 );
nand ( n29606 , n29600 , n377209 );
buf ( n377211 , n29606 );
buf ( n377212 , n377211 );
buf ( n377213 , n17209 );
nand ( n29610 , n377212 , n377213 );
buf ( n377215 , n29610 );
buf ( n377216 , n377215 );
nand ( n377217 , n377199 , n377216 );
buf ( n377218 , n377217 );
buf ( n377219 , n377218 );
xor ( n29616 , n377194 , n377219 );
not ( n377221 , n23108 );
nand ( n29618 , n377221 , n576 );
buf ( n377223 , n29618 );
not ( n29620 , n377223 );
buf ( n377225 , n29620 );
buf ( n377226 , n377225 );
and ( n377227 , n29616 , n377226 );
and ( n29624 , n377194 , n377219 );
or ( n377229 , n377227 , n29624 );
buf ( n377230 , n377229 );
buf ( n377231 , n377230 );
xor ( n29628 , n377169 , n377231 );
buf ( n377233 , n29628 );
buf ( n377234 , n377233 );
xor ( n377235 , n377085 , n377234 );
xor ( n29632 , n377142 , n377147 );
xor ( n377237 , n29632 , n377163 );
buf ( n377238 , n377237 );
buf ( n377239 , n377238 );
buf ( n377240 , n377023 );
not ( n377241 , n377240 );
buf ( n377242 , n576 );
not ( n377243 , n377242 );
buf ( n377244 , n370818 );
not ( n377245 , n377244 );
or ( n29642 , n377243 , n377245 );
buf ( n377247 , n365661 );
buf ( n377248 , n354303 );
nand ( n377249 , n377247 , n377248 );
buf ( n377250 , n377249 );
buf ( n377251 , n377250 );
nand ( n29648 , n29642 , n377251 );
buf ( n377253 , n29648 );
buf ( n377254 , n377253 );
not ( n377255 , n377254 );
or ( n29652 , n377241 , n377255 );
buf ( n377257 , n29530 );
buf ( n377258 , n364834 );
nand ( n377259 , n377257 , n377258 );
buf ( n377260 , n377259 );
buf ( n377261 , n377260 );
nand ( n29658 , n29652 , n377261 );
buf ( n377263 , n29658 );
buf ( n377264 , n377263 );
buf ( n377265 , n17037 );
not ( n29662 , n377265 );
buf ( n377267 , n377186 );
not ( n29664 , n377267 );
or ( n377269 , n29662 , n29664 );
buf ( n377270 , n578 );
not ( n377271 , n377270 );
buf ( n377272 , n23236 );
not ( n377273 , n377272 );
or ( n29670 , n377271 , n377273 );
buf ( n377275 , n17933 );
buf ( n377276 , n364727 );
nand ( n377277 , n377275 , n377276 );
buf ( n377278 , n377277 );
buf ( n377279 , n377278 );
nand ( n29676 , n29670 , n377279 );
buf ( n377281 , n29676 );
buf ( n377282 , n377281 );
buf ( n377283 , n17082 );
nand ( n29680 , n377282 , n377283 );
buf ( n377285 , n29680 );
buf ( n377286 , n377285 );
nand ( n377287 , n377269 , n377286 );
buf ( n377288 , n377287 );
buf ( n377289 , n377288 );
xor ( n29686 , n377264 , n377289 );
buf ( n377291 , n17133 );
not ( n29688 , n377291 );
buf ( n377293 , n582 );
not ( n29690 , n377293 );
buf ( n377295 , n28906 );
not ( n29692 , n377295 );
or ( n377297 , n29690 , n29692 );
buf ( n377298 , n364797 );
buf ( n377299 , n28905 );
nand ( n29696 , n377298 , n377299 );
buf ( n377301 , n29696 );
buf ( n377302 , n377301 );
nand ( n377303 , n377297 , n377302 );
buf ( n377304 , n377303 );
buf ( n377305 , n377304 );
not ( n29702 , n377305 );
or ( n377307 , n29688 , n29702 );
buf ( n377308 , n377161 );
buf ( n377309 , n365151 );
nand ( n29706 , n377308 , n377309 );
buf ( n377311 , n29706 );
buf ( n377312 , n377311 );
nand ( n377313 , n377307 , n377312 );
buf ( n377314 , n377313 );
buf ( n377315 , n377314 );
and ( n29712 , n29686 , n377315 );
and ( n377317 , n377264 , n377289 );
or ( n29714 , n29712 , n377317 );
buf ( n377319 , n29714 );
buf ( n377320 , n377319 );
xor ( n377321 , n377239 , n377320 );
buf ( n377322 , n17230 );
not ( n377323 , n377322 );
buf ( n377324 , n377211 );
not ( n377325 , n377324 );
or ( n29722 , n377323 , n377325 );
buf ( n377327 , n580 );
not ( n29724 , n377327 );
buf ( n377329 , n370956 );
not ( n29726 , n377329 );
or ( n377331 , n29724 , n29726 );
buf ( n377332 , n365892 );
buf ( n377333 , n364896 );
nand ( n29730 , n377332 , n377333 );
buf ( n377335 , n29730 );
buf ( n377336 , n377335 );
nand ( n377337 , n377331 , n377336 );
buf ( n377338 , n377337 );
buf ( n377339 , n377338 );
buf ( n377340 , n17209 );
nand ( n377341 , n377339 , n377340 );
buf ( n377342 , n377341 );
buf ( n377343 , n377342 );
nand ( n29740 , n29722 , n377343 );
buf ( n377345 , n29740 );
buf ( n377346 , n377345 );
buf ( n377347 , n29618 );
xor ( n29744 , n377346 , n377347 );
buf ( n377349 , n19106 );
buf ( n377350 , n576 );
and ( n377351 , n377349 , n377350 );
buf ( n377352 , n377351 );
buf ( n377353 , n377352 );
buf ( n377354 , n365355 );
buf ( n377355 , n576 );
nand ( n29752 , n377354 , n377355 );
buf ( n377357 , n29752 );
buf ( n377358 , n377357 );
not ( n377359 , n377358 );
buf ( n377360 , n377359 );
buf ( n377361 , n377360 );
xor ( n29758 , n377353 , n377361 );
buf ( n377363 , n17037 );
not ( n29760 , n377363 );
buf ( n377365 , n377281 );
not ( n29762 , n377365 );
or ( n377367 , n29760 , n29762 );
buf ( n377368 , n578 );
not ( n377369 , n377368 );
buf ( n377370 , n377076 );
not ( n377371 , n377370 );
or ( n29768 , n377369 , n377371 );
buf ( n377373 , n377073 );
buf ( n377374 , n364727 );
nand ( n377375 , n377373 , n377374 );
buf ( n377376 , n377375 );
buf ( n377377 , n377376 );
nand ( n29774 , n29768 , n377377 );
buf ( n377379 , n29774 );
buf ( n377380 , n377379 );
buf ( n377381 , n17082 );
nand ( n29778 , n377380 , n377381 );
buf ( n377383 , n29778 );
buf ( n377384 , n377383 );
nand ( n377385 , n377367 , n377384 );
buf ( n377386 , n377385 );
buf ( n377387 , n377386 );
and ( n377388 , n29758 , n377387 );
and ( n377389 , n377353 , n377361 );
or ( n29783 , n377388 , n377389 );
buf ( n377391 , n29783 );
buf ( n377392 , n377391 );
and ( n29786 , n29744 , n377392 );
and ( n29787 , n377346 , n377347 );
or ( n29788 , n29786 , n29787 );
buf ( n377396 , n29788 );
buf ( n377397 , n377396 );
and ( n29791 , n377321 , n377397 );
and ( n29792 , n377239 , n377320 );
or ( n29793 , n29791 , n29792 );
buf ( n377401 , n29793 );
buf ( n377402 , n377401 );
xor ( n29796 , n377235 , n377402 );
buf ( n377404 , n29796 );
not ( n29798 , n377404 );
xor ( n377406 , n377194 , n377219 );
xor ( n29800 , n377406 , n377226 );
buf ( n377408 , n29800 );
buf ( n377409 , n377408 );
xor ( n29803 , n377239 , n377320 );
xor ( n377411 , n29803 , n377397 );
buf ( n377412 , n377411 );
buf ( n377413 , n377412 );
xor ( n29807 , n377409 , n377413 );
buf ( n377415 , n377023 );
not ( n377416 , n377415 );
buf ( n377417 , n576 );
not ( n29811 , n377417 );
buf ( n377419 , n365748 );
not ( n29813 , n377419 );
or ( n377421 , n29811 , n29813 );
nand ( n29815 , n18854 , n354303 );
buf ( n377423 , n29815 );
nand ( n29817 , n377421 , n377423 );
buf ( n377425 , n29817 );
buf ( n377426 , n377425 );
not ( n29820 , n377426 );
or ( n29821 , n377416 , n29820 );
buf ( n377429 , n377253 );
buf ( n377430 , n364834 );
nand ( n377431 , n377429 , n377430 );
buf ( n377432 , n377431 );
buf ( n377433 , n377432 );
nand ( n29827 , n29821 , n377433 );
buf ( n377435 , n29827 );
buf ( n377436 , n377435 );
buf ( n377437 , n17209 );
not ( n29831 , n377437 );
buf ( n377439 , n580 );
not ( n29833 , n377439 );
buf ( n377441 , n376994 );
not ( n29835 , n377441 );
or ( n29836 , n29833 , n29835 );
buf ( n377444 , n375155 );
not ( n29838 , n377444 );
buf ( n377446 , n364896 );
nand ( n29840 , n29838 , n377446 );
buf ( n377448 , n29840 );
buf ( n377449 , n377448 );
nand ( n29843 , n29836 , n377449 );
buf ( n377451 , n29843 );
buf ( n377452 , n377451 );
not ( n29846 , n377452 );
or ( n29847 , n29831 , n29846 );
buf ( n377455 , n377338 );
buf ( n377456 , n17230 );
nand ( n29850 , n377455 , n377456 );
buf ( n377458 , n29850 );
buf ( n377459 , n377458 );
nand ( n29853 , n29847 , n377459 );
buf ( n377461 , n29853 );
buf ( n377462 , n377461 );
xor ( n29856 , n377436 , n377462 );
not ( n29857 , n584 );
not ( n29858 , n364664 );
or ( n377466 , n29857 , n29858 );
buf ( n377467 , n364661 );
buf ( n377468 , n364771 );
nand ( n29862 , n377467 , n377468 );
buf ( n377470 , n29862 );
nand ( n377471 , n377466 , n377470 );
not ( n29865 , n364973 );
nand ( n29866 , n29865 , n365406 );
nand ( n29867 , n377471 , n29866 );
buf ( n377475 , n29867 );
and ( n377476 , n29856 , n377475 );
and ( n29870 , n377436 , n377462 );
or ( n29871 , n377476 , n29870 );
buf ( n377479 , n29871 );
buf ( n377480 , n377479 );
xor ( n377481 , n377264 , n377289 );
xor ( n29875 , n377481 , n377315 );
buf ( n377483 , n29875 );
buf ( n377484 , n377483 );
xor ( n29878 , n377480 , n377484 );
buf ( n377486 , n17133 );
not ( n29880 , n377486 );
buf ( n377488 , n582 );
not ( n29882 , n377488 );
buf ( n377490 , n377059 );
not ( n377491 , n377490 );
or ( n29885 , n29882 , n377491 );
buf ( n377493 , n28909 );
not ( n29887 , n377493 );
buf ( n377495 , n364797 );
nand ( n377496 , n29887 , n377495 );
buf ( n377497 , n377496 );
buf ( n377498 , n377497 );
nand ( n29892 , n29885 , n377498 );
buf ( n377500 , n29892 );
buf ( n377501 , n377500 );
not ( n29895 , n377501 );
or ( n29896 , n29880 , n29895 );
buf ( n377504 , n377304 );
buf ( n377505 , n365151 );
nand ( n377506 , n377504 , n377505 );
buf ( n377507 , n377506 );
buf ( n377508 , n377507 );
nand ( n29902 , n29896 , n377508 );
buf ( n377510 , n29902 );
buf ( n377511 , n377510 );
buf ( n377512 , n377357 );
buf ( n377513 , n17082 );
not ( n29907 , n377513 );
buf ( n377515 , n364727 );
not ( n377516 , n377515 );
buf ( n377517 , n366277 );
not ( n29911 , n377517 );
or ( n29912 , n377516 , n29911 );
buf ( n377520 , n370818 );
buf ( n377521 , n578 );
nand ( n29915 , n377520 , n377521 );
buf ( n377523 , n29915 );
buf ( n377524 , n377523 );
nand ( n29918 , n29912 , n377524 );
buf ( n377526 , n29918 );
buf ( n377527 , n377526 );
not ( n29921 , n377527 );
or ( n29922 , n29907 , n29921 );
buf ( n377530 , n377379 );
buf ( n377531 , n17037 );
nand ( n29925 , n377530 , n377531 );
buf ( n377533 , n29925 );
buf ( n377534 , n377533 );
nand ( n29928 , n29922 , n377534 );
buf ( n377536 , n29928 );
buf ( n377537 , n377536 );
xor ( n29931 , n377512 , n377537 );
buf ( n377539 , n364834 );
not ( n29933 , n377539 );
buf ( n377541 , n377425 );
not ( n29935 , n377541 );
or ( n29936 , n29933 , n29935 );
buf ( n377544 , n576 );
not ( n29938 , n377544 );
buf ( n377546 , n23025 );
not ( n29940 , n377546 );
or ( n29941 , n29938 , n29940 );
buf ( n377549 , n17519 );
buf ( n377550 , n354303 );
nand ( n377551 , n377549 , n377550 );
buf ( n377552 , n377551 );
buf ( n377553 , n377552 );
nand ( n29947 , n29941 , n377553 );
buf ( n377555 , n29947 );
buf ( n377556 , n377555 );
buf ( n377557 , n377556 );
buf ( n377558 , n377023 );
nand ( n29952 , n377557 , n377558 );
buf ( n377560 , n29952 );
buf ( n377561 , n377560 );
nand ( n29955 , n29936 , n377561 );
buf ( n377563 , n29955 );
buf ( n377564 , n377563 );
and ( n29958 , n29931 , n377564 );
and ( n377566 , n377512 , n377537 );
or ( n29960 , n29958 , n377566 );
buf ( n377568 , n29960 );
buf ( n377569 , n377568 );
xor ( n29963 , n377511 , n377569 );
xor ( n377571 , n377353 , n377361 );
xor ( n29965 , n377571 , n377387 );
buf ( n377573 , n29965 );
buf ( n377574 , n377573 );
and ( n29968 , n29963 , n377574 );
and ( n377576 , n377511 , n377569 );
or ( n29970 , n29968 , n377576 );
buf ( n377578 , n29970 );
buf ( n377579 , n377578 );
and ( n29973 , n29878 , n377579 );
and ( n377581 , n377480 , n377484 );
or ( n29975 , n29973 , n377581 );
buf ( n377583 , n29975 );
buf ( n377584 , n377583 );
and ( n29978 , n29807 , n377584 );
and ( n377586 , n377409 , n377413 );
or ( n29980 , n29978 , n377586 );
buf ( n377588 , n29980 );
not ( n29982 , n377588 );
and ( n29983 , n29798 , n29982 );
xor ( n377591 , n377346 , n377347 );
xor ( n29985 , n377591 , n377392 );
buf ( n377593 , n29985 );
buf ( n377594 , n377593 );
xor ( n29988 , n377480 , n377484 );
xor ( n377596 , n29988 , n377579 );
buf ( n377597 , n377596 );
buf ( n377598 , n377597 );
xor ( n29992 , n377594 , n377598 );
and ( n29993 , n576 , n366654 );
buf ( n377601 , n29993 );
not ( n29995 , n364834 );
not ( n29996 , n377555 );
or ( n29997 , n29995 , n29996 );
buf ( n377605 , n576 );
not ( n377606 , n377605 );
buf ( n377607 , n364936 );
not ( n30001 , n377607 );
or ( n30002 , n377606 , n30001 );
buf ( n377610 , n365355 );
buf ( n377611 , n354303 );
nand ( n30005 , n377610 , n377611 );
buf ( n377613 , n30005 );
buf ( n377614 , n377613 );
nand ( n30008 , n30002 , n377614 );
buf ( n377616 , n30008 );
nand ( n30010 , n377616 , n17182 );
nand ( n30011 , n29997 , n30010 );
buf ( n377619 , n30011 );
xor ( n30013 , n377601 , n377619 );
buf ( n377621 , n365403 );
buf ( n377622 , n377621 );
buf ( n377623 , n576 );
nand ( n30017 , n377622 , n377623 );
buf ( n377625 , n30017 );
buf ( n377626 , n377625 );
not ( n30020 , n377626 );
buf ( n377628 , n30020 );
buf ( n377629 , n377628 );
and ( n30023 , n30013 , n377629 );
and ( n377631 , n377601 , n377619 );
or ( n30025 , n30023 , n377631 );
buf ( n377633 , n30025 );
buf ( n377634 , n377633 );
buf ( n377635 , n17230 );
not ( n377636 , n377635 );
buf ( n377637 , n377451 );
not ( n30031 , n377637 );
or ( n30032 , n377636 , n30031 );
not ( n30033 , n580 );
not ( n377641 , n23236 );
or ( n30035 , n30033 , n377641 );
buf ( n377643 , n17933 );
buf ( n377644 , n364896 );
nand ( n30038 , n377643 , n377644 );
buf ( n377646 , n30038 );
nand ( n30040 , n30035 , n377646 );
buf ( n377648 , n30040 );
buf ( n377649 , n17209 );
nand ( n30043 , n377648 , n377649 );
buf ( n377651 , n30043 );
buf ( n377652 , n377651 );
nand ( n30046 , n30032 , n377652 );
buf ( n377654 , n30046 );
buf ( n377655 , n377654 );
xor ( n377656 , n377634 , n377655 );
not ( n30050 , n364925 );
not ( n30051 , n377471 );
or ( n30052 , n30050 , n30051 );
not ( n30053 , n584 );
not ( n377661 , n23388 );
or ( n30055 , n30053 , n377661 );
not ( n30056 , n29486 );
nand ( n30057 , n30056 , n364771 );
nand ( n30058 , n30055 , n30057 );
buf ( n377666 , n30058 );
buf ( n377667 , n364973 );
nand ( n30061 , n377666 , n377667 );
buf ( n377669 , n30061 );
nand ( n30063 , n30052 , n377669 );
buf ( n377671 , n30063 );
and ( n30065 , n377656 , n377671 );
and ( n30066 , n377634 , n377655 );
or ( n30067 , n30065 , n30066 );
buf ( n377675 , n30067 );
buf ( n377676 , n377675 );
xor ( n30070 , n377436 , n377462 );
xor ( n30071 , n30070 , n377475 );
buf ( n377679 , n30071 );
buf ( n377680 , n377679 );
xor ( n377681 , n377676 , n377680 );
xor ( n30075 , n377511 , n377569 );
xor ( n30076 , n30075 , n377574 );
buf ( n377684 , n30076 );
buf ( n377685 , n377684 );
and ( n377686 , n377681 , n377685 );
and ( n30080 , n377676 , n377680 );
or ( n30081 , n377686 , n30080 );
buf ( n377689 , n30081 );
buf ( n377690 , n377689 );
and ( n377691 , n29992 , n377690 );
and ( n30085 , n377594 , n377598 );
or ( n30086 , n377691 , n30085 );
buf ( n377694 , n30086 );
xor ( n30088 , n377409 , n377413 );
xor ( n377696 , n30088 , n377584 );
buf ( n377697 , n377696 );
nor ( n30091 , n377694 , n377697 );
nor ( n30092 , n29983 , n30091 );
buf ( n377700 , n30092 );
xor ( n377701 , n377085 , n377234 );
and ( n30095 , n377701 , n377402 );
and ( n30096 , n377085 , n377234 );
or ( n30097 , n30095 , n30096 );
buf ( n377705 , n30097 );
buf ( n377706 , n377705 );
not ( n30100 , n377706 );
buf ( n377708 , n30100 );
buf ( n377709 , n377708 );
xor ( n30103 , n377030 , n377069 );
and ( n377711 , n30103 , n377082 );
and ( n30105 , n377030 , n377069 );
or ( n30106 , n377711 , n30105 );
buf ( n377714 , n30106 );
buf ( n377715 , n377714 );
buf ( n377716 , n17082 );
not ( n30110 , n377716 );
buf ( n377718 , n29462 );
not ( n30112 , n377718 );
or ( n30113 , n30110 , n30112 );
buf ( n377721 , n578 );
not ( n30115 , n377721 );
buf ( n377723 , n29488 );
not ( n30117 , n377723 );
or ( n30118 , n30115 , n30117 );
buf ( n377726 , n29487 );
buf ( n377727 , n377726 );
buf ( n377728 , n364727 );
nand ( n30122 , n377727 , n377728 );
buf ( n377730 , n30122 );
buf ( n377731 , n377730 );
nand ( n30125 , n30118 , n377731 );
buf ( n377733 , n30125 );
buf ( n377734 , n377733 );
buf ( n377735 , n17037 );
nand ( n377736 , n377734 , n377735 );
buf ( n377737 , n377736 );
buf ( n377738 , n377737 );
nand ( n30132 , n30113 , n377738 );
buf ( n377740 , n30132 );
buf ( n377741 , n377740 );
buf ( n377742 , n377081 );
not ( n30136 , n377742 );
buf ( n377744 , n30136 );
buf ( n377745 , n377744 );
xor ( n377746 , n377741 , n377745 );
not ( n30140 , n27128 );
buf ( n377748 , n30140 );
buf ( n377749 , n576 );
and ( n30143 , n377748 , n377749 );
buf ( n377751 , n30143 );
buf ( n377752 , n377751 );
buf ( n377753 , n365019 );
not ( n30147 , n377753 );
buf ( n377755 , n17209 );
not ( n377756 , n377755 );
buf ( n377757 , n377756 );
buf ( n377758 , n377757 );
not ( n30152 , n377758 );
or ( n30153 , n30147 , n30152 );
buf ( n377761 , n377117 );
nand ( n30155 , n30153 , n377761 );
buf ( n377763 , n30155 );
buf ( n377764 , n377763 );
xor ( n30158 , n377752 , n377764 );
buf ( n377766 , n364834 );
not ( n30160 , n377766 );
buf ( n377768 , n576 );
buf ( n377769 , n365892 );
xor ( n30163 , n377768 , n377769 );
buf ( n377771 , n30163 );
buf ( n377772 , n377771 );
not ( n30166 , n377772 );
or ( n30167 , n30160 , n30166 );
buf ( n377775 , n377004 );
buf ( n377776 , n377023 );
nand ( n30170 , n377775 , n377776 );
buf ( n377778 , n30170 );
buf ( n377779 , n377778 );
nand ( n30173 , n30167 , n377779 );
buf ( n377781 , n30173 );
buf ( n377782 , n377781 );
xor ( n30176 , n30158 , n377782 );
buf ( n377784 , n30176 );
buf ( n377785 , n377784 );
xor ( n377786 , n377746 , n377785 );
buf ( n377787 , n377786 );
buf ( n377788 , n377787 );
xor ( n30182 , n377715 , n377788 );
xor ( n30183 , n377125 , n377168 );
and ( n377791 , n30183 , n377231 );
and ( n30185 , n377125 , n377168 );
or ( n30186 , n377791 , n30185 );
buf ( n377794 , n30186 );
buf ( n377795 , n377794 );
xor ( n377796 , n30182 , n377795 );
buf ( n377797 , n377796 );
buf ( n377798 , n377797 );
not ( n30192 , n377798 );
buf ( n377800 , n30192 );
buf ( n377801 , n377800 );
nand ( n30195 , n377709 , n377801 );
buf ( n377803 , n30195 );
buf ( n377804 , n377803 );
nand ( n30198 , n377700 , n377804 );
buf ( n377806 , n30198 );
buf ( n377807 , n377806 );
not ( n30201 , n377807 );
buf ( n377809 , n30201 );
not ( n30203 , n377809 );
buf ( n377811 , n365151 );
not ( n30205 , n377811 );
buf ( n377813 , n377500 );
not ( n30207 , n377813 );
or ( n30208 , n30205 , n30207 );
buf ( n377816 , n582 );
not ( n30210 , n377816 );
buf ( n377818 , n377036 );
not ( n30212 , n377818 );
or ( n30213 , n30210 , n30212 );
buf ( n377821 , n377042 );
buf ( n377822 , n364797 );
nand ( n30216 , n377821 , n377822 );
buf ( n377824 , n30216 );
buf ( n377825 , n377824 );
nand ( n377826 , n30213 , n377825 );
buf ( n377827 , n377826 );
buf ( n377828 , n377827 );
buf ( n377829 , n17133 );
nand ( n30223 , n377828 , n377829 );
buf ( n377831 , n30223 );
buf ( n377832 , n377831 );
nand ( n30226 , n30208 , n377832 );
buf ( n377834 , n30226 );
buf ( n377835 , n377834 );
buf ( n377836 , n17230 );
not ( n30230 , n377836 );
buf ( n377838 , n30040 );
not ( n30232 , n377838 );
or ( n30233 , n30230 , n30232 );
buf ( n377841 , n377073 );
buf ( n377842 , n364896 );
nand ( n30236 , n377841 , n377842 );
buf ( n377844 , n30236 );
not ( n30238 , n377844 );
nand ( n377846 , n377076 , n580 );
not ( n30240 , n377846 );
or ( n30241 , n30238 , n30240 );
nand ( n30242 , n30241 , n17209 );
buf ( n377850 , n30242 );
nand ( n377851 , n30233 , n377850 );
buf ( n377852 , n377851 );
buf ( n377853 , n377852 );
buf ( n377854 , n17082 );
not ( n30248 , n377854 );
buf ( n377856 , n578 );
not ( n30250 , n377856 );
buf ( n377858 , n23108 );
not ( n30252 , n377858 );
or ( n30253 , n30250 , n30252 );
buf ( n377861 , n365748 );
not ( n30255 , n377861 );
buf ( n377863 , n364727 );
nand ( n30257 , n30255 , n377863 );
buf ( n377865 , n30257 );
buf ( n377866 , n377865 );
nand ( n30260 , n30253 , n377866 );
buf ( n377868 , n30260 );
buf ( n377869 , n377868 );
not ( n30263 , n377869 );
or ( n377871 , n30248 , n30263 );
buf ( n377872 , n377526 );
buf ( n377873 , n17037 );
nand ( n30267 , n377872 , n377873 );
buf ( n377875 , n30267 );
buf ( n377876 , n377875 );
nand ( n30270 , n377871 , n377876 );
buf ( n377878 , n30270 );
buf ( n377879 , n377878 );
xor ( n30273 , n377853 , n377879 );
buf ( n377881 , n17133 );
not ( n30275 , n377881 );
buf ( n377883 , n582 );
not ( n30277 , n377883 );
buf ( n377885 , n375155 );
not ( n377886 , n377885 );
or ( n30280 , n30277 , n377886 );
buf ( n377888 , n370944 );
not ( n30282 , n377888 );
buf ( n377890 , n364797 );
nand ( n377891 , n30282 , n377890 );
buf ( n377892 , n377891 );
buf ( n377893 , n377892 );
nand ( n30287 , n30280 , n377893 );
buf ( n377895 , n30287 );
buf ( n377896 , n377895 );
not ( n30290 , n377896 );
or ( n30291 , n30275 , n30290 );
buf ( n377899 , n377827 );
buf ( n377900 , n365151 );
nand ( n377901 , n377899 , n377900 );
buf ( n377902 , n377901 );
buf ( n377903 , n377902 );
nand ( n30297 , n30291 , n377903 );
buf ( n377905 , n30297 );
buf ( n377906 , n377905 );
and ( n30300 , n30273 , n377906 );
and ( n30301 , n377853 , n377879 );
or ( n30302 , n30300 , n30301 );
buf ( n377910 , n30302 );
buf ( n377911 , n377910 );
xor ( n30305 , n377835 , n377911 );
xor ( n30306 , n377512 , n377537 );
xor ( n30307 , n30306 , n377564 );
buf ( n377915 , n30307 );
buf ( n377916 , n377915 );
xor ( n30310 , n30305 , n377916 );
buf ( n377918 , n30310 );
buf ( n377919 , n377918 );
buf ( n377920 , n586 );
not ( n377921 , n377920 );
buf ( n377922 , n16981 );
not ( n30316 , n377922 );
or ( n30317 , n377921 , n30316 );
buf ( n377925 , n16982 );
buf ( n377926 , n365334 );
nand ( n30320 , n377925 , n377926 );
buf ( n377928 , n30320 );
buf ( n377929 , n377928 );
nand ( n30323 , n30317 , n377929 );
buf ( n377931 , n30323 );
nand ( n30325 , n365350 , n369743 );
nand ( n30326 , n377931 , n30325 );
buf ( n377934 , n30326 );
buf ( n377935 , n364973 );
not ( n377936 , n377935 );
not ( n30330 , n584 );
not ( n30331 , n371006 );
or ( n30332 , n30330 , n30331 );
buf ( n377940 , n28897 );
buf ( n377941 , n364771 );
nand ( n30335 , n377940 , n377941 );
buf ( n377943 , n30335 );
nand ( n30337 , n30332 , n377943 );
buf ( n377945 , n30337 );
not ( n377946 , n377945 );
or ( n30340 , n377936 , n377946 );
buf ( n377948 , n30058 );
buf ( n377949 , n364925 );
nand ( n30343 , n377948 , n377949 );
buf ( n377951 , n30343 );
buf ( n377952 , n377951 );
nand ( n30346 , n30340 , n377952 );
buf ( n377954 , n30346 );
buf ( n377955 , n377954 );
xor ( n377956 , n377934 , n377955 );
xor ( n30350 , n377601 , n377619 );
xor ( n30351 , n30350 , n377629 );
buf ( n377959 , n30351 );
buf ( n377960 , n377959 );
and ( n377961 , n377956 , n377960 );
and ( n30355 , n377934 , n377955 );
or ( n30356 , n377961 , n30355 );
buf ( n377964 , n30356 );
buf ( n377965 , n377964 );
xor ( n377966 , n377634 , n377655 );
xor ( n30360 , n377966 , n377671 );
buf ( n377968 , n30360 );
buf ( n377969 , n377968 );
xor ( n30363 , n377965 , n377969 );
buf ( n377971 , n364834 );
not ( n30365 , n377971 );
buf ( n377973 , n377616 );
not ( n30367 , n377973 );
or ( n30368 , n30365 , n30367 );
xor ( n377976 , n576 , n366654 );
nand ( n30370 , n377976 , n377023 );
buf ( n377978 , n30370 );
nand ( n30372 , n30368 , n377978 );
buf ( n377980 , n30372 );
buf ( n377981 , n377980 );
buf ( n377982 , n377625 );
xor ( n30376 , n377981 , n377982 );
and ( n30377 , n576 , n360086 );
buf ( n377985 , n30377 );
buf ( n377986 , n364834 );
not ( n30380 , n377986 );
buf ( n377988 , n30380 );
buf ( n377989 , n377988 );
buf ( n377990 , n354303 );
nor ( n377991 , n377989 , n377990 );
buf ( n377992 , n377991 );
nand ( n30386 , n366657 , n377992 );
buf ( n377994 , n377988 );
buf ( n377995 , n576 );
nor ( n377996 , n377994 , n377995 );
buf ( n377997 , n377996 );
nand ( n30391 , n366654 , n377997 );
xor ( n30392 , n576 , n17021 );
nand ( n30393 , n30392 , n17182 );
nand ( n378001 , n30386 , n30391 , n30393 );
buf ( n378002 , n378001 );
xor ( n30396 , n377985 , n378002 );
buf ( n378004 , n357316 );
buf ( n378005 , n576 );
nand ( n378006 , n378004 , n378005 );
buf ( n378007 , n378006 );
buf ( n378008 , n378007 );
not ( n30402 , n378008 );
buf ( n378010 , n30402 );
buf ( n378011 , n378010 );
and ( n30405 , n30396 , n378011 );
and ( n30406 , n377985 , n378002 );
or ( n30407 , n30405 , n30406 );
buf ( n378015 , n30407 );
buf ( n378016 , n378015 );
and ( n30410 , n30376 , n378016 );
and ( n30411 , n377981 , n377982 );
or ( n30412 , n30410 , n30411 );
buf ( n378020 , n30412 );
buf ( n378021 , n378020 );
xor ( n30415 , n377853 , n377879 );
xor ( n30416 , n30415 , n377906 );
buf ( n378024 , n30416 );
buf ( n378025 , n378024 );
xor ( n30419 , n378021 , n378025 );
buf ( n378027 , n17209 );
not ( n30421 , n378027 );
buf ( n378029 , n364896 );
not ( n30423 , n378029 );
buf ( n378031 , n366277 );
not ( n30425 , n378031 );
or ( n30426 , n30423 , n30425 );
buf ( n378034 , n370818 );
buf ( n378035 , n580 );
nand ( n30429 , n378034 , n378035 );
buf ( n378037 , n30429 );
buf ( n378038 , n378037 );
nand ( n30432 , n30426 , n378038 );
buf ( n378040 , n30432 );
buf ( n378041 , n378040 );
not ( n30435 , n378041 );
or ( n30436 , n30421 , n30435 );
buf ( n378044 , n580 );
not ( n30438 , n378044 );
buf ( n378046 , n377076 );
not ( n30440 , n378046 );
or ( n30441 , n30438 , n30440 );
buf ( n378049 , n377844 );
nand ( n30443 , n30441 , n378049 );
buf ( n378051 , n30443 );
buf ( n378052 , n378051 );
buf ( n378053 , n17230 );
nand ( n30447 , n378052 , n378053 );
buf ( n378055 , n30447 );
buf ( n378056 , n378055 );
nand ( n30450 , n30436 , n378056 );
buf ( n378058 , n30450 );
buf ( n378059 , n378058 );
buf ( n378060 , n17037 );
not ( n30454 , n378060 );
buf ( n378062 , n377868 );
not ( n30456 , n378062 );
or ( n30457 , n30454 , n30456 );
buf ( n378065 , n578 );
not ( n30459 , n378065 );
buf ( n378067 , n17520 );
not ( n30461 , n378067 );
or ( n30462 , n30459 , n30461 );
buf ( n378070 , n17519 );
buf ( n378071 , n364727 );
nand ( n30465 , n378070 , n378071 );
buf ( n378073 , n30465 );
buf ( n378074 , n378073 );
nand ( n30468 , n30462 , n378074 );
buf ( n378076 , n30468 );
buf ( n378077 , n378076 );
buf ( n378078 , n17082 );
nand ( n30472 , n378077 , n378078 );
buf ( n378080 , n30472 );
buf ( n378081 , n378080 );
nand ( n30475 , n30457 , n378081 );
buf ( n378083 , n30475 );
buf ( n378084 , n378083 );
xor ( n30478 , n378059 , n378084 );
buf ( n378086 , n17133 );
not ( n30480 , n378086 );
buf ( n378088 , n582 );
not ( n30482 , n378088 );
buf ( n378090 , n23236 );
not ( n30484 , n378090 );
or ( n30485 , n30482 , n30484 );
buf ( n378093 , n17933 );
buf ( n378094 , n364797 );
nand ( n30488 , n378093 , n378094 );
buf ( n378096 , n30488 );
buf ( n378097 , n378096 );
nand ( n30491 , n30485 , n378097 );
buf ( n378099 , n30491 );
buf ( n378100 , n378099 );
not ( n30494 , n378100 );
or ( n30495 , n30480 , n30494 );
buf ( n378103 , n377895 );
buf ( n378104 , n365151 );
nand ( n30498 , n378103 , n378104 );
buf ( n378106 , n30498 );
buf ( n378107 , n378106 );
nand ( n30501 , n30495 , n378107 );
buf ( n378109 , n30501 );
buf ( n378110 , n378109 );
and ( n30504 , n30478 , n378110 );
and ( n30505 , n378059 , n378084 );
or ( n30506 , n30504 , n30505 );
buf ( n378114 , n30506 );
buf ( n378115 , n378114 );
and ( n30509 , n30419 , n378115 );
and ( n30510 , n378021 , n378025 );
or ( n30511 , n30509 , n30510 );
buf ( n378119 , n30511 );
buf ( n378120 , n378119 );
xor ( n30514 , n30363 , n378120 );
buf ( n378122 , n30514 );
buf ( n378123 , n378122 );
xor ( n30517 , n377919 , n378123 );
xor ( n30518 , n377934 , n377955 );
xor ( n30519 , n30518 , n377960 );
buf ( n378127 , n30519 );
buf ( n378128 , n378127 );
buf ( n378129 , n365375 );
not ( n30523 , n378129 );
buf ( n378131 , n586 );
not ( n30525 , n378131 );
buf ( n378133 , n29486 );
not ( n30527 , n378133 );
or ( n30528 , n30525 , n30527 );
buf ( n378136 , n23387 );
buf ( n378137 , n365334 );
nand ( n30531 , n378136 , n378137 );
buf ( n378139 , n30531 );
buf ( n378140 , n378139 );
nand ( n30534 , n30528 , n378140 );
buf ( n378142 , n30534 );
buf ( n378143 , n378142 );
not ( n30537 , n378143 );
or ( n30538 , n30523 , n30537 );
buf ( n378146 , n377931 );
buf ( n378147 , n365351 );
nand ( n30541 , n378146 , n378147 );
buf ( n378149 , n30541 );
buf ( n378150 , n378149 );
nand ( n30544 , n30538 , n378150 );
buf ( n378152 , n30544 );
buf ( n378153 , n378152 );
buf ( n378154 , n364925 );
not ( n30548 , n378154 );
buf ( n378156 , n30337 );
not ( n30550 , n378156 );
or ( n30551 , n30548 , n30550 );
buf ( n378159 , n584 );
not ( n30553 , n378159 );
buf ( n378161 , n377036 );
not ( n30555 , n378161 );
or ( n30556 , n30553 , n30555 );
buf ( n378164 , n377042 );
buf ( n378165 , n364771 );
nand ( n30559 , n378164 , n378165 );
buf ( n378167 , n30559 );
buf ( n378168 , n378167 );
nand ( n30562 , n30556 , n378168 );
buf ( n378170 , n30562 );
buf ( n378171 , n378170 );
buf ( n378172 , n364973 );
nand ( n30566 , n378171 , n378172 );
buf ( n378174 , n30566 );
buf ( n378175 , n378174 );
nand ( n30569 , n30551 , n378175 );
buf ( n378177 , n30569 );
buf ( n378178 , n378177 );
xor ( n30572 , n378153 , n378178 );
buf ( n378180 , n17037 );
not ( n30574 , n378180 );
buf ( n378182 , n378076 );
not ( n30576 , n378182 );
or ( n30577 , n30574 , n30576 );
buf ( n378185 , n578 );
not ( n30579 , n378185 );
buf ( n378187 , n364936 );
not ( n30581 , n378187 );
or ( n30582 , n30579 , n30581 );
buf ( n378190 , n367123 );
buf ( n378191 , n364727 );
nand ( n30585 , n378190 , n378191 );
buf ( n378193 , n30585 );
buf ( n378194 , n378193 );
nand ( n30588 , n30582 , n378194 );
buf ( n378196 , n30588 );
buf ( n378197 , n378196 );
buf ( n378198 , n17082 );
nand ( n30592 , n378197 , n378198 );
buf ( n378200 , n30592 );
buf ( n378201 , n378200 );
nand ( n30595 , n30577 , n378201 );
buf ( n378203 , n30595 );
buf ( n378204 , n378203 );
buf ( n378205 , n17209 );
not ( n30599 , n378205 );
and ( n30600 , n16900 , n364896 );
not ( n30601 , n16900 );
and ( n30602 , n30601 , n580 );
or ( n30603 , n30600 , n30602 );
buf ( n378211 , n30603 );
not ( n30605 , n378211 );
or ( n30606 , n30599 , n30605 );
buf ( n378214 , n378040 );
buf ( n378215 , n17230 );
nand ( n30609 , n378214 , n378215 );
buf ( n378217 , n30609 );
buf ( n378218 , n378217 );
nand ( n30612 , n30606 , n378218 );
buf ( n378220 , n30612 );
buf ( n378221 , n378220 );
xor ( n30615 , n378204 , n378221 );
buf ( n378223 , n365151 );
not ( n30617 , n378223 );
buf ( n378225 , n378099 );
not ( n30619 , n378225 );
or ( n30620 , n30617 , n30619 );
buf ( n378228 , n582 );
not ( n30622 , n378228 );
not ( n30623 , n17905 );
buf ( n378231 , n30623 );
not ( n30625 , n378231 );
or ( n30626 , n30622 , n30625 );
buf ( n378234 , n17002 );
buf ( n378235 , n364797 );
nand ( n30629 , n378234 , n378235 );
buf ( n378237 , n30629 );
buf ( n378238 , n378237 );
nand ( n30632 , n30626 , n378238 );
buf ( n378240 , n30632 );
buf ( n378241 , n378240 );
buf ( n378242 , n17133 );
nand ( n30636 , n378241 , n378242 );
buf ( n378244 , n30636 );
buf ( n378245 , n378244 );
nand ( n30639 , n30620 , n378245 );
buf ( n378247 , n30639 );
buf ( n378248 , n378247 );
and ( n30642 , n30615 , n378248 );
and ( n30643 , n378204 , n378221 );
or ( n30644 , n30642 , n30643 );
buf ( n378252 , n30644 );
buf ( n378253 , n378252 );
and ( n30647 , n30572 , n378253 );
and ( n30648 , n378153 , n378178 );
or ( n30649 , n30647 , n30648 );
buf ( n378257 , n30649 );
buf ( n378258 , n378257 );
xor ( n30652 , n378128 , n378258 );
xor ( n30653 , n377981 , n377982 );
xor ( n30654 , n30653 , n378016 );
buf ( n378262 , n30654 );
buf ( n378263 , n378262 );
not ( n30657 , n364834 );
not ( n30658 , n30392 );
or ( n30659 , n30657 , n30658 );
xor ( n30660 , n576 , n360086 );
nand ( n30661 , n30660 , n17182 );
nand ( n378269 , n30659 , n30661 );
buf ( n378270 , n378269 );
not ( n30664 , n17182 );
buf ( n378272 , n576 );
not ( n30666 , n378272 );
buf ( n378274 , n364891 );
not ( n30668 , n378274 );
or ( n30669 , n30666 , n30668 );
buf ( n378277 , n9625 );
buf ( n378278 , n354303 );
nand ( n30672 , n378277 , n378278 );
buf ( n378280 , n30672 );
buf ( n378281 , n378280 );
nand ( n30675 , n30669 , n378281 );
buf ( n378283 , n30675 );
not ( n30677 , n378283 );
or ( n30678 , n30664 , n30677 );
nand ( n30679 , n30660 , n364834 );
nand ( n30680 , n30678 , n30679 );
buf ( n378288 , n30680 );
xor ( n30682 , n378270 , n378288 );
buf ( n378290 , n378007 );
and ( n30684 , n30682 , n378290 );
and ( n30685 , n378270 , n378288 );
or ( n30686 , n30684 , n30685 );
buf ( n378294 , n30686 );
buf ( n378295 , n378294 );
xor ( n30689 , n377985 , n378002 );
xor ( n30690 , n30689 , n378011 );
buf ( n378298 , n30690 );
buf ( n378299 , n378298 );
xor ( n30693 , n378295 , n378299 );
buf ( n378301 , n364925 );
not ( n30695 , n378301 );
buf ( n378303 , n378170 );
not ( n30697 , n378303 );
or ( n30698 , n30695 , n30697 );
and ( n30699 , n365897 , n364771 );
not ( n30700 , n365897 );
and ( n30701 , n30700 , n584 );
or ( n30702 , n30699 , n30701 );
buf ( n378310 , n30702 );
buf ( n378311 , n364973 );
nand ( n30705 , n378310 , n378311 );
buf ( n378313 , n30705 );
buf ( n378314 , n378313 );
nand ( n30708 , n30698 , n378314 );
buf ( n378316 , n30708 );
buf ( n378317 , n378316 );
and ( n30711 , n30693 , n378317 );
and ( n30712 , n378295 , n378299 );
or ( n30713 , n30711 , n30712 );
buf ( n378321 , n30713 );
buf ( n378322 , n378321 );
xor ( n30716 , n378263 , n378322 );
xor ( n30717 , n378059 , n378084 );
xor ( n30718 , n30717 , n378110 );
buf ( n378326 , n30718 );
buf ( n378327 , n378326 );
and ( n30721 , n30716 , n378327 );
and ( n30722 , n378263 , n378322 );
or ( n30723 , n30721 , n30722 );
buf ( n378331 , n30723 );
buf ( n378332 , n378331 );
and ( n30726 , n30652 , n378332 );
and ( n30727 , n378128 , n378258 );
or ( n30728 , n30726 , n30727 );
buf ( n378336 , n30728 );
buf ( n378337 , n378336 );
xor ( n30731 , n30517 , n378337 );
buf ( n378339 , n30731 );
not ( n30733 , n378339 );
xor ( n30734 , n378021 , n378025 );
xor ( n30735 , n30734 , n378115 );
buf ( n378343 , n30735 );
buf ( n378344 , n378343 );
xor ( n30738 , n378128 , n378258 );
xor ( n30739 , n30738 , n378332 );
buf ( n378347 , n30739 );
buf ( n378348 , n378347 );
xor ( n30742 , n378344 , n378348 );
xor ( n30743 , n378153 , n378178 );
xor ( n30744 , n30743 , n378253 );
buf ( n378352 , n30744 );
buf ( n378353 , n378352 );
buf ( n378354 , n368307 );
not ( n30748 , n378354 );
buf ( n378356 , n17875 );
not ( n30750 , n378356 );
or ( n30751 , n30748 , n30750 );
buf ( n378359 , n588 );
not ( n30753 , n378359 );
buf ( n378361 , n16981 );
not ( n30755 , n378361 );
or ( n30756 , n30753 , n30755 );
buf ( n378364 , n588 );
not ( n30758 , n378364 );
buf ( n378366 , n16982 );
nand ( n30760 , n30758 , n378366 );
buf ( n378368 , n30760 );
buf ( n378369 , n378368 );
nand ( n30763 , n30756 , n378369 );
buf ( n378371 , n30763 );
buf ( n378372 , n378371 );
nand ( n30766 , n30751 , n378372 );
buf ( n378374 , n30766 );
buf ( n378375 , n378374 );
buf ( n378376 , n365375 );
not ( n30770 , n378376 );
buf ( n378378 , n586 );
not ( n30772 , n378378 );
buf ( n378380 , n28909 );
not ( n30774 , n378380 );
or ( n30775 , n30772 , n30774 );
buf ( n378383 , n28897 );
buf ( n378384 , n365334 );
nand ( n30778 , n378383 , n378384 );
buf ( n378386 , n30778 );
buf ( n378387 , n378386 );
nand ( n30781 , n30775 , n378387 );
buf ( n378389 , n30781 );
buf ( n378390 , n378389 );
not ( n30784 , n378390 );
or ( n30785 , n30770 , n30784 );
buf ( n378393 , n378142 );
buf ( n378394 , n365351 );
nand ( n30788 , n378393 , n378394 );
buf ( n378396 , n30788 );
buf ( n378397 , n378396 );
nand ( n30791 , n30785 , n378397 );
buf ( n378399 , n30791 );
buf ( n378400 , n378399 );
xor ( n30794 , n378375 , n378400 );
buf ( n378402 , n17037 );
not ( n30796 , n378402 );
buf ( n378404 , n378196 );
not ( n30798 , n378404 );
or ( n30799 , n30796 , n30798 );
and ( n30800 , n14498 , n364727 );
not ( n30801 , n14498 );
and ( n30802 , n30801 , n578 );
or ( n30803 , n30800 , n30802 );
buf ( n378411 , n30803 );
buf ( n378412 , n17082 );
nand ( n30806 , n378411 , n378412 );
buf ( n378414 , n30806 );
buf ( n378415 , n378414 );
nand ( n30809 , n30799 , n378415 );
buf ( n378417 , n30809 );
buf ( n378418 , n378417 );
buf ( n378419 , n17230 );
not ( n30813 , n378419 );
buf ( n378421 , n30603 );
not ( n30815 , n378421 );
or ( n30816 , n30813 , n30815 );
buf ( n378424 , n580 );
not ( n30818 , n378424 );
buf ( n378426 , n366255 );
not ( n30820 , n378426 );
or ( n30821 , n30818 , n30820 );
buf ( n378429 , n17519 );
buf ( n378430 , n364896 );
nand ( n30824 , n378429 , n378430 );
buf ( n378432 , n30824 );
buf ( n378433 , n378432 );
nand ( n30827 , n30821 , n378433 );
buf ( n378435 , n30827 );
buf ( n378436 , n378435 );
buf ( n378437 , n17209 );
nand ( n30831 , n378436 , n378437 );
buf ( n378439 , n30831 );
buf ( n378440 , n378439 );
nand ( n30834 , n30816 , n378440 );
buf ( n378442 , n30834 );
buf ( n378443 , n378442 );
xor ( n30837 , n378418 , n378443 );
buf ( n378445 , n357348 );
buf ( n378446 , n576 );
and ( n30840 , n378445 , n378446 );
buf ( n378448 , n30840 );
buf ( n378449 , n378448 );
not ( n30843 , n30680 );
buf ( n378451 , n30843 );
xor ( n30845 , n378449 , n378451 );
buf ( n378453 , n17037 );
not ( n30847 , n378453 );
buf ( n378455 , n30803 );
not ( n30849 , n378455 );
or ( n30850 , n30847 , n30849 );
buf ( n378458 , n578 );
not ( n30852 , n378458 );
buf ( n378460 , n364790 );
not ( n30854 , n378460 );
or ( n30855 , n30852 , n30854 );
buf ( n378463 , n17021 );
buf ( n378464 , n364727 );
nand ( n30858 , n378463 , n378464 );
buf ( n378466 , n30858 );
buf ( n378467 , n378466 );
nand ( n30861 , n30855 , n378467 );
buf ( n378469 , n30861 );
buf ( n378470 , n378469 );
buf ( n378471 , n17082 );
nand ( n30865 , n378470 , n378471 );
buf ( n378473 , n30865 );
buf ( n378474 , n378473 );
nand ( n30868 , n30850 , n378474 );
buf ( n378476 , n30868 );
buf ( n378477 , n378476 );
and ( n30871 , n30845 , n378477 );
and ( n30872 , n378449 , n378451 );
or ( n30873 , n30871 , n30872 );
buf ( n378481 , n30873 );
buf ( n378482 , n378481 );
and ( n30876 , n30837 , n378482 );
and ( n30877 , n378418 , n378443 );
or ( n30878 , n30876 , n30877 );
buf ( n378486 , n30878 );
buf ( n378487 , n378486 );
and ( n30881 , n30794 , n378487 );
and ( n30882 , n378375 , n378400 );
or ( n30883 , n30881 , n30882 );
buf ( n378491 , n30883 );
buf ( n378492 , n378491 );
xor ( n30886 , n378353 , n378492 );
not ( n30887 , n17133 );
buf ( n378495 , n364797 );
not ( n30889 , n378495 );
buf ( n378497 , n16955 );
not ( n30891 , n378497 );
or ( n30892 , n30889 , n30891 );
buf ( n378500 , n370818 );
buf ( n378501 , n582 );
nand ( n30895 , n378500 , n378501 );
buf ( n378503 , n30895 );
buf ( n378504 , n378503 );
nand ( n30898 , n30892 , n378504 );
buf ( n378506 , n30898 );
not ( n30900 , n378506 );
or ( n30901 , n30887 , n30900 );
not ( n30902 , n378237 );
nand ( n30903 , n30623 , n582 );
not ( n30904 , n30903 );
or ( n30905 , n30902 , n30904 );
nand ( n30906 , n30905 , n365151 );
nand ( n30907 , n30901 , n30906 );
buf ( n378515 , n30907 );
xor ( n30909 , n378270 , n378288 );
xor ( n30910 , n30909 , n378290 );
buf ( n378518 , n30910 );
buf ( n378519 , n378518 );
xor ( n30913 , n378515 , n378519 );
buf ( n378521 , n364925 );
not ( n30915 , n378521 );
buf ( n378523 , n30702 );
not ( n30917 , n378523 );
or ( n30918 , n30915 , n30917 );
buf ( n378526 , n17933 );
not ( n30920 , n378526 );
buf ( n378528 , n584 );
nand ( n30922 , n30920 , n378528 );
buf ( n378530 , n30922 );
buf ( n378531 , n378530 );
not ( n30925 , n378531 );
buf ( n378533 , n23236 );
not ( n30927 , n378533 );
buf ( n378535 , n364771 );
nand ( n30929 , n30927 , n378535 );
buf ( n378537 , n30929 );
buf ( n378538 , n378537 );
not ( n30932 , n378538 );
or ( n30933 , n30925 , n30932 );
buf ( n378541 , n364973 );
nand ( n30935 , n30933 , n378541 );
buf ( n378543 , n30935 );
buf ( n378544 , n378543 );
nand ( n30938 , n30918 , n378544 );
buf ( n378546 , n30938 );
buf ( n378547 , n378546 );
and ( n30941 , n30913 , n378547 );
and ( n30942 , n378515 , n378519 );
or ( n30943 , n30941 , n30942 );
buf ( n378551 , n30943 );
buf ( n378552 , n378551 );
xor ( n30946 , n378204 , n378221 );
xor ( n30947 , n30946 , n378248 );
buf ( n378555 , n30947 );
buf ( n378556 , n378555 );
xor ( n30950 , n378552 , n378556 );
xor ( n30951 , n378295 , n378299 );
xor ( n30952 , n30951 , n378317 );
buf ( n378560 , n30952 );
buf ( n378561 , n378560 );
and ( n30955 , n30950 , n378561 );
and ( n30956 , n378552 , n378556 );
or ( n30957 , n30955 , n30956 );
buf ( n378565 , n30957 );
buf ( n378566 , n378565 );
and ( n30960 , n30886 , n378566 );
and ( n30961 , n378353 , n378492 );
or ( n30962 , n30960 , n30961 );
buf ( n378570 , n30962 );
buf ( n378571 , n378570 );
and ( n30965 , n30742 , n378571 );
and ( n30966 , n378344 , n378348 );
or ( n30967 , n30965 , n30966 );
buf ( n378575 , n30967 );
not ( n30969 , n378575 );
and ( n30970 , n30733 , n30969 );
xor ( n30971 , n378344 , n378348 );
xor ( n30972 , n30971 , n378571 );
buf ( n378580 , n30972 );
xor ( n30974 , n378263 , n378322 );
xor ( n30975 , n30974 , n378327 );
buf ( n378583 , n30975 );
buf ( n378584 , n378583 );
xor ( n30978 , n378353 , n378492 );
xor ( n30979 , n30978 , n378566 );
buf ( n378587 , n30979 );
buf ( n378588 , n378587 );
xor ( n30982 , n378584 , n378588 );
xor ( n30983 , n378375 , n378400 );
xor ( n30984 , n30983 , n378487 );
buf ( n378592 , n30984 );
buf ( n378593 , n378592 );
buf ( n378594 , n365646 );
not ( n30988 , n378594 );
and ( n30989 , n588 , n29486 );
not ( n30990 , n588 );
and ( n30991 , n30990 , n23387 );
or ( n30992 , n30989 , n30991 );
buf ( n378600 , n30992 );
not ( n30994 , n378600 );
or ( n30995 , n30988 , n30994 );
buf ( n378603 , n378371 );
buf ( n378604 , n17867 );
nand ( n30998 , n378603 , n378604 );
buf ( n378606 , n30998 );
buf ( n378607 , n378606 );
nand ( n31001 , n30995 , n378607 );
buf ( n378609 , n31001 );
buf ( n378610 , n378609 );
buf ( n378611 , n365351 );
not ( n31005 , n378611 );
buf ( n378613 , n378389 );
not ( n31007 , n378613 );
or ( n31008 , n31005 , n31007 );
buf ( n378616 , n365892 );
not ( n31010 , n378616 );
buf ( n378618 , n365334 );
not ( n31012 , n378618 );
and ( n31013 , n31010 , n31012 );
buf ( n378621 , n370956 );
not ( n31015 , n378621 );
buf ( n378623 , n31015 );
buf ( n378624 , n378623 );
buf ( n378625 , n365334 );
and ( n31019 , n378624 , n378625 );
nor ( n31020 , n31013 , n31019 );
buf ( n378628 , n31020 );
buf ( n378629 , n378628 );
not ( n31023 , n378629 );
buf ( n378631 , n365375 );
nand ( n31025 , n31023 , n378631 );
buf ( n378633 , n31025 );
buf ( n378634 , n378633 );
nand ( n31028 , n31008 , n378634 );
buf ( n378636 , n31028 );
buf ( n378637 , n378636 );
xor ( n31031 , n378610 , n378637 );
buf ( n378639 , n17230 );
not ( n31033 , n378639 );
buf ( n378641 , n378435 );
not ( n31035 , n378641 );
or ( n31036 , n31033 , n31035 );
buf ( n378644 , n580 );
not ( n31038 , n378644 );
buf ( n378646 , n364936 );
not ( n31040 , n378646 );
or ( n31041 , n31038 , n31040 );
buf ( n378649 , n365355 );
buf ( n378650 , n364896 );
nand ( n31044 , n378649 , n378650 );
buf ( n378652 , n31044 );
buf ( n378653 , n378652 );
nand ( n31047 , n31041 , n378653 );
buf ( n378655 , n31047 );
buf ( n378656 , n378655 );
buf ( n378657 , n17209 );
nand ( n31051 , n378656 , n378657 );
buf ( n378659 , n31051 );
buf ( n378660 , n378659 );
nand ( n31054 , n31036 , n378660 );
buf ( n378662 , n31054 );
buf ( n378663 , n378662 );
buf ( n378664 , n364834 );
not ( n31058 , n378664 );
buf ( n378666 , n378283 );
not ( n31060 , n378666 );
or ( n31061 , n31058 , n31060 );
nand ( n31062 , n23185 , n17182 );
buf ( n378670 , n31062 );
nand ( n31064 , n31061 , n378670 );
buf ( n378672 , n31064 );
buf ( n378673 , n378672 );
and ( n31067 , n370682 , n370683 );
buf ( n378675 , n31067 );
buf ( n378676 , n378675 );
xor ( n31070 , n378673 , n378676 );
buf ( n378678 , n17037 );
not ( n31072 , n378678 );
buf ( n378680 , n378469 );
not ( n31074 , n378680 );
or ( n31075 , n31072 , n31074 );
not ( n31076 , n370772 );
not ( n31077 , n23163 );
or ( n31078 , n31076 , n31077 );
nand ( n31079 , n31078 , n17082 );
buf ( n378687 , n31079 );
nand ( n31081 , n31075 , n378687 );
buf ( n378689 , n31081 );
buf ( n378690 , n378689 );
and ( n31084 , n31070 , n378690 );
and ( n31085 , n378673 , n378676 );
or ( n31086 , n31084 , n31085 );
buf ( n378694 , n31086 );
buf ( n378695 , n378694 );
xor ( n31089 , n378663 , n378695 );
buf ( n378697 , n17133 );
not ( n31091 , n378697 );
nand ( n31092 , n582 , n23108 );
buf ( n378700 , n364797 );
buf ( n378701 , n16900 );
nand ( n31095 , n378700 , n378701 );
buf ( n378703 , n31095 );
nand ( n31097 , n31092 , n378703 );
buf ( n378705 , n31097 );
not ( n31099 , n378705 );
or ( n31100 , n31091 , n31099 );
buf ( n378708 , n378506 );
buf ( n378709 , n365151 );
nand ( n31103 , n378708 , n378709 );
buf ( n378711 , n31103 );
buf ( n378712 , n378711 );
nand ( n31106 , n31100 , n378712 );
buf ( n378714 , n31106 );
buf ( n378715 , n378714 );
and ( n31109 , n31089 , n378715 );
and ( n31110 , n378663 , n378695 );
or ( n31111 , n31109 , n31110 );
buf ( n378719 , n31111 );
buf ( n378720 , n378719 );
and ( n31114 , n31031 , n378720 );
and ( n31115 , n378610 , n378637 );
or ( n31116 , n31114 , n31115 );
buf ( n378724 , n31116 );
buf ( n378725 , n378724 );
xor ( n31119 , n378593 , n378725 );
buf ( n378727 , n365881 );
not ( n31121 , n378727 );
buf ( n378729 , n365410 );
nand ( n31123 , n31121 , n378729 );
buf ( n378731 , n31123 );
buf ( n378732 , n378731 );
buf ( n378733 , n17905 );
not ( n31127 , n378733 );
buf ( n378735 , n369554 );
nand ( n31129 , n31127 , n378735 );
buf ( n378737 , n31129 );
buf ( n378738 , n378737 );
buf ( n378739 , n17905 );
buf ( n378740 , n370806 );
nand ( n31134 , n378739 , n378740 );
buf ( n378742 , n31134 );
buf ( n378743 , n378742 );
buf ( n378744 , n365881 );
buf ( n378745 , n365430 );
nand ( n31139 , n378744 , n378745 );
buf ( n378747 , n31139 );
buf ( n378748 , n378747 );
nand ( n31142 , n378732 , n378738 , n378743 , n378748 );
buf ( n378750 , n31142 );
buf ( n378751 , n378750 );
xor ( n31145 , n378449 , n378451 );
xor ( n31146 , n31145 , n378477 );
buf ( n378754 , n31146 );
buf ( n378755 , n378754 );
xor ( n31149 , n378751 , n378755 );
buf ( n378757 , n365375 );
not ( n31151 , n378757 );
buf ( n378759 , n365897 );
buf ( n378760 , n586 );
and ( n31154 , n378759 , n378760 );
not ( n31155 , n378759 );
buf ( n378763 , n365334 );
and ( n31157 , n31155 , n378763 );
nor ( n31158 , n31154 , n31157 );
buf ( n378766 , n31158 );
buf ( n378767 , n378766 );
not ( n31161 , n378767 );
or ( n31162 , n31151 , n31161 );
buf ( n378770 , n378628 );
buf ( n378771 , n365350 );
or ( n31165 , n378770 , n378771 );
nand ( n31166 , n31162 , n31165 );
buf ( n378774 , n31166 );
buf ( n378775 , n378774 );
and ( n31169 , n31149 , n378775 );
and ( n31170 , n378751 , n378755 );
or ( n31171 , n31169 , n31170 );
buf ( n378779 , n31171 );
buf ( n378780 , n378779 );
xor ( n31174 , n378418 , n378443 );
xor ( n31175 , n31174 , n378482 );
buf ( n378783 , n31175 );
buf ( n378784 , n378783 );
xor ( n31178 , n378780 , n378784 );
xor ( n31179 , n378515 , n378519 );
xor ( n31180 , n31179 , n378547 );
buf ( n378788 , n31180 );
buf ( n378789 , n378788 );
and ( n31183 , n31178 , n378789 );
and ( n31184 , n378780 , n378784 );
or ( n31185 , n31183 , n31184 );
buf ( n378793 , n31185 );
buf ( n378794 , n378793 );
and ( n31188 , n31119 , n378794 );
and ( n31189 , n378593 , n378725 );
or ( n31190 , n31188 , n31189 );
buf ( n378798 , n31190 );
buf ( n378799 , n378798 );
and ( n31193 , n30982 , n378799 );
and ( n31194 , n378584 , n378588 );
or ( n31195 , n31193 , n31194 );
buf ( n378803 , n31195 );
nor ( n31197 , n378580 , n378803 );
nor ( n31198 , n30970 , n31197 );
xor ( n31199 , n377835 , n377911 );
and ( n31200 , n31199 , n377916 );
and ( n31201 , n377835 , n377911 );
or ( n31202 , n31200 , n31201 );
buf ( n378810 , n31202 );
buf ( n378811 , n378810 );
xor ( n31205 , n377676 , n377680 );
xor ( n31206 , n31205 , n377685 );
buf ( n378814 , n31206 );
buf ( n378815 , n378814 );
xor ( n31209 , n378811 , n378815 );
xor ( n31210 , n377965 , n377969 );
and ( n31211 , n31210 , n378120 );
and ( n31212 , n377965 , n377969 );
or ( n31213 , n31211 , n31212 );
buf ( n378821 , n31213 );
buf ( n378822 , n378821 );
xor ( n31216 , n31209 , n378822 );
buf ( n378824 , n31216 );
not ( n31218 , n378824 );
xor ( n31219 , n377919 , n378123 );
and ( n31220 , n31219 , n378337 );
and ( n31221 , n377919 , n378123 );
or ( n31222 , n31220 , n31221 );
buf ( n378830 , n31222 );
not ( n31224 , n378830 );
and ( n31225 , n31218 , n31224 );
xor ( n31226 , n377594 , n377598 );
xor ( n31227 , n31226 , n377690 );
buf ( n378835 , n31227 );
not ( n31229 , n378835 );
xor ( n31230 , n378811 , n378815 );
and ( n31231 , n31230 , n378822 );
and ( n31232 , n378811 , n378815 );
or ( n31233 , n31231 , n31232 );
buf ( n378841 , n31233 );
not ( n31235 , n378841 );
and ( n31236 , n31229 , n31235 );
nor ( n31237 , n31225 , n31236 );
nand ( n31238 , n31198 , n31237 );
buf ( n378846 , n31238 );
not ( n31240 , n378846 );
buf ( n378848 , n31240 );
not ( n31242 , n378848 );
xor ( n31243 , n378780 , n378784 );
xor ( n31244 , n31243 , n378789 );
buf ( n378852 , n31244 );
buf ( n378853 , n378852 );
buf ( n378854 , n365351 );
not ( n31248 , n378854 );
buf ( n378856 , n378766 );
not ( n31250 , n378856 );
or ( n31251 , n31248 , n31250 );
buf ( n378859 , n370850 );
buf ( n378860 , n365375 );
nand ( n31254 , n378859 , n378860 );
buf ( n378862 , n31254 );
buf ( n378863 , n378862 );
nand ( n31257 , n31251 , n378863 );
buf ( n378865 , n31257 );
buf ( n378866 , n378865 );
buf ( n378867 , n17867 );
not ( n31261 , n378867 );
xor ( n31262 , n588 , n28897 );
buf ( n378870 , n31262 );
not ( n31264 , n378870 );
or ( n31265 , n31261 , n31264 );
buf ( n378873 , n370967 );
buf ( n378874 , n365646 );
nand ( n31268 , n378873 , n378874 );
buf ( n378876 , n31268 );
buf ( n378877 , n378876 );
nand ( n31271 , n31265 , n378877 );
buf ( n378879 , n31271 );
buf ( n378880 , n378879 );
xor ( n31274 , n378866 , n378880 );
buf ( n378882 , n365738 );
not ( n31276 , n378882 );
buf ( n378884 , n371000 );
not ( n31278 , n378884 );
or ( n31279 , n31276 , n31278 );
xor ( n31280 , n590 , n16982 );
buf ( n378888 , n31280 );
buf ( n378889 , n591 );
nand ( n31283 , n378888 , n378889 );
buf ( n378891 , n31283 );
buf ( n378892 , n378891 );
nand ( n31286 , n31279 , n378892 );
buf ( n378894 , n31286 );
buf ( n378895 , n378894 );
and ( n31289 , n31274 , n378895 );
and ( n31290 , n378866 , n378880 );
or ( n31291 , n31289 , n31290 );
buf ( n378899 , n31291 );
buf ( n378900 , n378899 );
buf ( n378901 , n370062 );
not ( n31295 , n378901 );
buf ( n378903 , n367116 );
not ( n31297 , n378903 );
or ( n31298 , n31295 , n31297 );
buf ( n378906 , n31280 );
nand ( n31300 , n31298 , n378906 );
buf ( n378908 , n31300 );
buf ( n378909 , n378908 );
buf ( n378910 , n17230 );
not ( n31304 , n378910 );
buf ( n378912 , n378655 );
not ( n31306 , n378912 );
or ( n31307 , n31304 , n31306 );
buf ( n378915 , n22996 );
buf ( n378916 , n17209 );
nand ( n31310 , n378915 , n378916 );
buf ( n378918 , n31310 );
buf ( n378919 , n378918 );
nand ( n31313 , n31307 , n378919 );
buf ( n378921 , n31313 );
buf ( n378922 , n378921 );
xor ( n31316 , n370761 , n370779 );
and ( n31317 , n31316 , n370797 );
and ( n31318 , n370761 , n370779 );
or ( n31319 , n31317 , n31318 );
buf ( n378927 , n31319 );
buf ( n378928 , n378927 );
xor ( n31322 , n378922 , n378928 );
xor ( n31323 , n378673 , n378676 );
xor ( n31324 , n31323 , n378690 );
buf ( n378932 , n31324 );
buf ( n378933 , n378932 );
and ( n31327 , n31322 , n378933 );
and ( n31328 , n378922 , n378928 );
or ( n31329 , n31327 , n31328 );
buf ( n378937 , n31329 );
buf ( n378938 , n378937 );
xor ( n31332 , n378909 , n378938 );
buf ( n378940 , n17867 );
not ( n31334 , n378940 );
buf ( n378942 , n30992 );
not ( n31336 , n378942 );
or ( n31337 , n31334 , n31336 );
buf ( n378945 , n31262 );
buf ( n378946 , n365646 );
nand ( n31340 , n378945 , n378946 );
buf ( n378948 , n31340 );
buf ( n378949 , n378948 );
nand ( n31343 , n31337 , n378949 );
buf ( n378951 , n31343 );
buf ( n378952 , n378951 );
xor ( n31346 , n31332 , n378952 );
buf ( n378954 , n31346 );
buf ( n378955 , n378954 );
xor ( n31349 , n378900 , n378955 );
xor ( n31350 , n378922 , n378928 );
xor ( n31351 , n31350 , n378933 );
buf ( n378959 , n31351 );
buf ( n378960 , n378959 );
xor ( n31354 , n370800 , n370832 );
and ( n31355 , n31354 , n370853 );
and ( n31356 , n370800 , n370832 );
or ( n31357 , n31355 , n31356 );
buf ( n378965 , n31357 );
buf ( n378966 , n378965 );
xor ( n31360 , n378960 , n378966 );
buf ( n378968 , n364973 );
not ( n31362 , n378968 );
buf ( n378970 , n364771 );
buf ( n378971 , n370818 );
and ( n31365 , n378970 , n378971 );
not ( n31366 , n378970 );
buf ( n378974 , n366277 );
and ( n31368 , n31366 , n378974 );
nor ( n31369 , n31365 , n31368 );
buf ( n378977 , n31369 );
buf ( n378978 , n378977 );
not ( n31372 , n378978 );
or ( n31373 , n31362 , n31372 );
buf ( n378981 , n584 );
not ( n31375 , n378981 );
buf ( n378983 , n30623 );
not ( n31377 , n378983 );
or ( n31378 , n31375 , n31377 );
buf ( n378986 , n364771 );
buf ( n378987 , n17002 );
nand ( n31381 , n378986 , n378987 );
buf ( n378989 , n31381 );
buf ( n378990 , n378989 );
nand ( n31384 , n31378 , n378990 );
buf ( n378992 , n31384 );
buf ( n378993 , n378992 );
buf ( n378994 , n364925 );
nand ( n31388 , n378993 , n378994 );
buf ( n378996 , n31388 );
buf ( n378997 , n378996 );
nand ( n31391 , n31373 , n378997 );
buf ( n378999 , n31391 );
buf ( n379000 , n378999 );
not ( n31394 , n365151 );
not ( n31395 , n31097 );
or ( n31396 , n31394 , n31395 );
and ( n31397 , n25697 , n364797 );
not ( n31398 , n25697 );
and ( n31399 , n31398 , n582 );
or ( n31400 , n31397 , n31399 );
nand ( n31401 , n31400 , n17133 );
nand ( n31402 , n31396 , n31401 );
buf ( n379010 , n31402 );
xor ( n31404 , n379000 , n379010 );
xor ( n31405 , n370616 , n370657 );
and ( n31406 , n31405 , n370701 );
and ( n31407 , n370616 , n370657 );
or ( n379015 , n31406 , n31407 );
buf ( n379016 , n379015 );
buf ( n379017 , n379016 );
xor ( n31411 , n31404 , n379017 );
buf ( n379019 , n31411 );
buf ( n379020 , n379019 );
and ( n31414 , n31360 , n379020 );
and ( n31415 , n378960 , n378966 );
or ( n31416 , n31414 , n31415 );
buf ( n379024 , n31416 );
buf ( n379025 , n379024 );
and ( n31419 , n31349 , n379025 );
and ( n31420 , n378900 , n378955 );
or ( n31421 , n31419 , n31420 );
buf ( n379029 , n31421 );
buf ( n379030 , n379029 );
xor ( n31424 , n378853 , n379030 );
xor ( n31425 , n378909 , n378938 );
and ( n31426 , n31425 , n378952 );
and ( n31427 , n378909 , n378938 );
or ( n31428 , n31426 , n31427 );
buf ( n379036 , n31428 );
buf ( n379037 , n379036 );
xor ( n31431 , n378610 , n378637 );
xor ( n31432 , n31431 , n378720 );
buf ( n379040 , n31432 );
buf ( n379041 , n379040 );
xor ( n31435 , n379037 , n379041 );
xor ( n31436 , n378663 , n378695 );
xor ( n31437 , n31436 , n378715 );
buf ( n379045 , n31437 );
buf ( n379046 , n379045 );
xor ( n31440 , n379000 , n379010 );
and ( n31441 , n31440 , n379017 );
and ( n31442 , n379000 , n379010 );
or ( n31443 , n31441 , n31442 );
buf ( n379051 , n31443 );
buf ( n379052 , n379051 );
xor ( n31446 , n379046 , n379052 );
xor ( n31447 , n378751 , n378755 );
xor ( n31448 , n31447 , n378775 );
buf ( n379056 , n31448 );
buf ( n379057 , n379056 );
and ( n31451 , n31446 , n379057 );
and ( n31452 , n379046 , n379052 );
or ( n31453 , n31451 , n31452 );
buf ( n379061 , n31453 );
buf ( n379062 , n379061 );
xor ( n31456 , n31435 , n379062 );
buf ( n379064 , n31456 );
buf ( n379065 , n379064 );
xor ( n31459 , n31424 , n379065 );
buf ( n379067 , n31459 );
buf ( n379068 , n379067 );
xor ( n31462 , n379046 , n379052 );
xor ( n31463 , n31462 , n379057 );
buf ( n379071 , n31463 );
buf ( n379072 , n379071 );
xor ( n31466 , n378900 , n378955 );
xor ( n31467 , n31466 , n379025 );
buf ( n379075 , n31467 );
buf ( n379076 , n379075 );
xor ( n31470 , n379072 , n379076 );
xor ( n31471 , n370975 , n370981 );
and ( n31472 , n31471 , n371016 );
and ( n31473 , n370975 , n370981 );
or ( n31474 , n31472 , n31473 );
buf ( n379082 , n31474 );
buf ( n379083 , n379082 );
xor ( n31477 , n378866 , n378880 );
xor ( n31478 , n31477 , n378895 );
buf ( n379086 , n31478 );
buf ( n379087 , n379086 );
xor ( n31481 , n379083 , n379087 );
xor ( n31482 , n370704 , n370757 );
and ( n31483 , n31482 , n370856 );
and ( n31484 , n370704 , n370757 );
or ( n31485 , n31483 , n31484 );
buf ( n379093 , n31485 );
buf ( n379094 , n379093 );
and ( n31488 , n31481 , n379094 );
and ( n31489 , n379083 , n379087 );
or ( n31490 , n31488 , n31489 );
buf ( n379098 , n31490 );
buf ( n379099 , n379098 );
and ( n31493 , n31470 , n379099 );
and ( n31494 , n379072 , n379076 );
or ( n31495 , n31493 , n31494 );
buf ( n379103 , n31495 );
buf ( n379104 , n379103 );
nor ( n31498 , n379068 , n379104 );
buf ( n379106 , n31498 );
xor ( n31500 , n379072 , n379076 );
xor ( n31501 , n31500 , n379099 );
buf ( n379109 , n31501 );
buf ( n379110 , n379109 );
xor ( n31504 , n378960 , n378966 );
xor ( n31505 , n31504 , n379020 );
buf ( n379113 , n31505 );
buf ( n379114 , n379113 );
xor ( n31508 , n379083 , n379087 );
xor ( n31509 , n31508 , n379094 );
buf ( n379117 , n31509 );
buf ( n379118 , n379117 );
xor ( n31512 , n379114 , n379118 );
xor ( n31513 , n370935 , n371019 );
and ( n31514 , n31513 , n371049 );
and ( n31515 , n370935 , n371019 );
or ( n31516 , n31514 , n31515 );
buf ( n379124 , n31516 );
buf ( n379125 , n379124 );
and ( n31519 , n31512 , n379125 );
and ( n31520 , n379114 , n379118 );
or ( n31521 , n31519 , n31520 );
buf ( n379129 , n31521 );
buf ( n379130 , n379129 );
nand ( n31524 , n379110 , n379130 );
buf ( n379132 , n31524 );
or ( n31526 , n379106 , n379132 );
buf ( n379134 , n379103 );
buf ( n379135 , n379067 );
nand ( n31529 , n379134 , n379135 );
buf ( n379137 , n31529 );
nand ( n31531 , n31526 , n379137 );
xor ( n31532 , n378552 , n378556 );
xor ( n31533 , n31532 , n378561 );
buf ( n379141 , n31533 );
buf ( n379142 , n379141 );
xor ( n31536 , n378593 , n378725 );
xor ( n31537 , n31536 , n378794 );
buf ( n379145 , n31537 );
buf ( n379146 , n379145 );
xor ( n31540 , n379142 , n379146 );
xor ( n31541 , n379037 , n379041 );
and ( n31542 , n31541 , n379062 );
and ( n31543 , n379037 , n379041 );
or ( n31544 , n31542 , n31543 );
buf ( n379152 , n31544 );
buf ( n379153 , n379152 );
xor ( n31547 , n31540 , n379153 );
buf ( n379155 , n31547 );
not ( n31549 , n379155 );
xor ( n31550 , n378853 , n379030 );
and ( n31551 , n31550 , n379065 );
and ( n31552 , n378853 , n379030 );
or ( n31553 , n31551 , n31552 );
buf ( n379161 , n31553 );
buf ( n379162 , n379161 );
not ( n31556 , n379162 );
buf ( n379164 , n31556 );
nand ( n31558 , n31549 , n379164 );
xor ( n31559 , n378584 , n378588 );
xor ( n31560 , n31559 , n378799 );
buf ( n379168 , n31560 );
not ( n31562 , n379168 );
xor ( n31563 , n379142 , n379146 );
and ( n31564 , n31563 , n379153 );
and ( n31565 , n379142 , n379146 );
or ( n31566 , n31564 , n31565 );
buf ( n379174 , n31566 );
not ( n31568 , n379174 );
nand ( n31569 , n31562 , n31568 );
nand ( n31570 , n31531 , n31558 , n31569 );
nor ( n31571 , n379168 , n379174 );
not ( n31572 , n31571 );
nand ( n31573 , n379155 , n379161 );
not ( n31574 , n31573 );
and ( n31575 , n31572 , n31574 );
buf ( n379183 , n31568 );
not ( n31577 , n379183 );
buf ( n379185 , n31577 );
not ( n31579 , n31562 );
and ( n31580 , n379185 , n31579 );
nor ( n31581 , n31575 , n31580 );
nand ( n31582 , n31570 , n31581 );
not ( n31583 , n31582 );
or ( n31584 , n31242 , n31583 );
buf ( n379192 , n379155 );
not ( n31586 , n379192 );
buf ( n379194 , n31586 );
nand ( n31588 , n379164 , n379194 );
not ( n31589 , n379109 );
not ( n31590 , n379129 );
and ( n31591 , n31589 , n31590 );
nor ( n31592 , n379067 , n379103 );
nor ( n31593 , n31591 , n31592 );
nand ( n31594 , n31568 , n31562 );
nand ( n31595 , n31588 , n31593 , n31594 );
nor ( n31596 , n31238 , n31595 );
not ( n31597 , n371054 );
not ( n31598 , n371074 );
and ( n31599 , n31597 , n31598 );
xor ( n31600 , n379114 , n379118 );
xor ( n31601 , n31600 , n379125 );
buf ( n379209 , n31601 );
buf ( n379210 , n379209 );
xor ( n31604 , n370859 , n370928 );
and ( n31605 , n31604 , n371052 );
and ( n31606 , n370859 , n370928 );
or ( n31607 , n31605 , n31606 );
buf ( n379215 , n31607 );
buf ( n379216 , n379215 );
nor ( n31610 , n379210 , n379216 );
buf ( n379218 , n31610 );
nor ( n31612 , n31599 , n379218 );
not ( n31613 , n31612 );
not ( n31614 , n371128 );
or ( n31615 , n31613 , n31614 );
buf ( n379223 , n379218 );
not ( n31617 , n379223 );
buf ( n379225 , n371081 );
not ( n31619 , n379225 );
and ( n31620 , n31617 , n31619 );
buf ( n379228 , n379209 );
buf ( n379229 , n379215 );
and ( n31623 , n379228 , n379229 );
buf ( n379231 , n31623 );
buf ( n379232 , n379231 );
nor ( n31626 , n31620 , n379232 );
buf ( n379234 , n31626 );
nand ( n31628 , n31615 , n379234 );
nand ( n31629 , n31596 , n31628 );
nand ( n31630 , n31584 , n31629 );
buf ( n379238 , n31630 );
not ( n31632 , n379238 );
buf ( n379240 , n31632 );
buf ( n379241 , n379240 );
not ( n31635 , n31237 );
buf ( n379243 , n378339 );
buf ( n31637 , n379243 );
buf ( n379245 , n31637 );
buf ( n379246 , n379245 );
buf ( n379247 , n378575 );
buf ( n31641 , n379247 );
buf ( n379249 , n31641 );
buf ( n379250 , n379249 );
nor ( n31644 , n379246 , n379250 );
buf ( n379252 , n31644 );
buf ( n379253 , n378580 );
buf ( n31647 , n379253 );
buf ( n379255 , n31647 );
nand ( n31649 , n379255 , n378803 );
or ( n31650 , n379252 , n31649 );
buf ( n379258 , n379245 );
buf ( n379259 , n379249 );
nand ( n31653 , n379258 , n379259 );
buf ( n379261 , n31653 );
nand ( n31655 , n31650 , n379261 );
not ( n31656 , n31655 );
or ( n31657 , n31635 , n31656 );
buf ( n379265 , n378835 );
buf ( n31659 , n379265 );
buf ( n379267 , n31659 );
buf ( n379268 , n379267 );
not ( n31662 , n379268 );
buf ( n379270 , n31662 );
not ( n31664 , n379270 );
buf ( n379272 , n378841 );
buf ( n31666 , n379272 );
buf ( n379274 , n31666 );
buf ( n379275 , n379274 );
not ( n31669 , n379275 );
buf ( n379277 , n31669 );
not ( n31671 , n379277 );
and ( n31672 , n31664 , n31671 );
buf ( n379280 , n378824 );
buf ( n31674 , n379280 );
buf ( n379282 , n31674 );
buf ( n379283 , n379282 );
buf ( n31677 , n378830 );
buf ( n379285 , n31677 );
nand ( n31679 , n379283 , n379285 );
buf ( n379287 , n31679 );
buf ( n379288 , n379287 );
not ( n31682 , n379288 );
buf ( n379290 , n31682 );
buf ( n379291 , n379270 );
buf ( n379292 , n379277 );
nand ( n31686 , n379291 , n379292 );
buf ( n379294 , n31686 );
and ( n31688 , n379290 , n379294 );
nor ( n31689 , n31672 , n31688 );
nand ( n31690 , n31657 , n31689 );
buf ( n379298 , n31690 );
not ( n31692 , n379298 );
buf ( n379300 , n31692 );
buf ( n379301 , n379300 );
nand ( n31695 , n379241 , n379301 );
buf ( n379303 , n31695 );
not ( n31697 , n379303 );
or ( n31698 , n30203 , n31697 );
buf ( n379306 , n377708 );
buf ( n379307 , n377800 );
nand ( n31701 , n379306 , n379307 );
buf ( n379309 , n31701 );
buf ( n379310 , n379309 );
not ( n31704 , n379310 );
buf ( n379312 , n377588 );
buf ( n379313 , n377404 );
nor ( n31707 , n379312 , n379313 );
buf ( n379315 , n31707 );
buf ( n379316 , n377694 );
buf ( n379317 , n377697 );
nand ( n31711 , n379316 , n379317 );
buf ( n379319 , n31711 );
or ( n31713 , n379315 , n379319 );
buf ( n379321 , n377588 );
buf ( n379322 , n377404 );
nand ( n31716 , n379321 , n379322 );
buf ( n379324 , n31716 );
nand ( n31718 , n31713 , n379324 );
buf ( n379326 , n31718 );
not ( n31720 , n379326 );
or ( n31721 , n31704 , n31720 );
buf ( n379329 , n377800 );
not ( n31723 , n379329 );
buf ( n379331 , n377705 );
nand ( n31725 , n31723 , n379331 );
buf ( n379333 , n31725 );
buf ( n379334 , n379333 );
nand ( n31728 , n31721 , n379334 );
buf ( n379336 , n31728 );
buf ( n379337 , n379336 );
not ( n31731 , n379337 );
buf ( n379339 , n31731 );
nand ( n31733 , n31698 , n379339 );
xor ( n31734 , n377715 , n377788 );
and ( n31735 , n31734 , n377795 );
and ( n31736 , n377715 , n377788 );
or ( n31737 , n31735 , n31736 );
buf ( n379345 , n31737 );
buf ( n379346 , n379345 );
xor ( n31740 , n377752 , n377764 );
and ( n31741 , n31740 , n377782 );
and ( n31742 , n377752 , n377764 );
or ( n31743 , n31741 , n31742 );
buf ( n379351 , n31743 );
buf ( n379352 , n379351 );
buf ( n379353 , n364834 );
not ( n31747 , n379353 );
buf ( n379355 , n576 );
not ( n31749 , n379355 );
buf ( n379357 , n377059 );
not ( n31751 , n379357 );
or ( n31752 , n31749 , n31751 );
buf ( n379360 , n377056 );
buf ( n379361 , n354303 );
nand ( n31755 , n379360 , n379361 );
buf ( n379363 , n31755 );
buf ( n379364 , n379363 );
nand ( n31758 , n31752 , n379364 );
buf ( n379366 , n31758 );
buf ( n379367 , n379366 );
not ( n31761 , n379367 );
or ( n31762 , n31747 , n31761 );
buf ( n379370 , n377771 );
buf ( n379371 , n377023 );
nand ( n31765 , n379370 , n379371 );
buf ( n379373 , n31765 );
buf ( n379374 , n379373 );
nand ( n31768 , n31762 , n379374 );
buf ( n379376 , n31768 );
buf ( n379377 , n379376 );
buf ( n379378 , n17082 );
not ( n31772 , n379378 );
buf ( n379380 , n377733 );
not ( n31774 , n379380 );
or ( n31775 , n31772 , n31774 );
buf ( n379383 , n578 );
not ( n31777 , n379383 );
buf ( n379385 , n364664 );
not ( n31779 , n379385 );
or ( n31780 , n31777 , n31779 );
buf ( n379388 , n364661 );
buf ( n379389 , n364727 );
nand ( n31783 , n379388 , n379389 );
buf ( n379391 , n31783 );
buf ( n379392 , n379391 );
nand ( n31786 , n31780 , n379392 );
buf ( n379394 , n31786 );
buf ( n379395 , n379394 );
buf ( n379396 , n17037 );
nand ( n31790 , n379395 , n379396 );
buf ( n379398 , n31790 );
buf ( n379399 , n379398 );
nand ( n31793 , n31775 , n379399 );
buf ( n379401 , n31793 );
buf ( n379402 , n379401 );
xor ( n31796 , n379377 , n379402 );
buf ( n379404 , n376991 );
buf ( n379405 , n576 );
nand ( n31799 , n379404 , n379405 );
buf ( n379407 , n31799 );
buf ( n379408 , n379407 );
xor ( n31802 , n31796 , n379408 );
buf ( n379410 , n31802 );
buf ( n379411 , n379410 );
xor ( n31805 , n379352 , n379411 );
xor ( n31806 , n377741 , n377745 );
and ( n31807 , n31806 , n377785 );
and ( n31808 , n377741 , n377745 );
or ( n31809 , n31807 , n31808 );
buf ( n379417 , n31809 );
buf ( n379418 , n379417 );
xor ( n31812 , n31805 , n379418 );
buf ( n379420 , n31812 );
buf ( n379421 , n379420 );
nor ( n31815 , n379346 , n379421 );
buf ( n379423 , n31815 );
buf ( n379424 , n379423 );
not ( n31818 , n379424 );
buf ( n379426 , n31818 );
not ( n31820 , n379426 );
buf ( n379428 , n379345 );
buf ( n379429 , n379420 );
and ( n31823 , n379428 , n379429 );
buf ( n379431 , n31823 );
nor ( n31825 , n31820 , n379431 );
and ( n31826 , n31733 , n31825 );
not ( n31827 , n31733 );
not ( n31828 , n31825 );
and ( n31829 , n31827 , n31828 );
nor ( n31830 , n31826 , n31829 );
not ( n31831 , n31830 );
not ( n31832 , n30092 );
nand ( n31833 , n379240 , n379300 );
not ( n31834 , n31833 );
or ( n31835 , n31832 , n31834 );
not ( n31836 , n31718 );
nand ( n31837 , n31835 , n31836 );
buf ( n31838 , n379333 );
nand ( n31839 , n31838 , n377803 );
not ( n31840 , n31839 );
and ( n31841 , n31837 , n31840 );
not ( n31842 , n31837 );
and ( n31843 , n31842 , n31839 );
nor ( n31844 , n31841 , n31843 );
not ( n31845 , n31844 );
or ( n31846 , n31831 , n31845 );
not ( n31847 , n31844 );
not ( n31848 , n31830 );
nand ( n31849 , n31847 , n31848 );
nand ( n31850 , n31846 , n31849 );
buf ( n379458 , n31850 );
buf ( n31852 , n379458 );
buf ( n379460 , n31852 );
buf ( n379461 , n379460 );
not ( n31855 , n379461 );
buf ( n379463 , n31855 );
buf ( n379464 , n379463 );
buf ( n31858 , n379464 );
buf ( n379466 , n31858 );
buf ( n379467 , n379466 );
not ( n31861 , n379467 );
buf ( n379469 , n379407 );
not ( n31863 , n379469 );
buf ( n379471 , n31863 );
buf ( n379472 , n379471 );
buf ( n379473 , n17037 );
not ( n31867 , n379473 );
buf ( n379475 , n31867 );
buf ( n379476 , n379475 );
not ( n31870 , n379476 );
buf ( n379478 , n17081 );
not ( n31872 , n379478 );
or ( n31873 , n31870 , n31872 );
buf ( n379481 , n379394 );
nand ( n31875 , n31873 , n379481 );
buf ( n379483 , n31875 );
buf ( n379484 , n379483 );
and ( n31878 , n377768 , n377769 );
buf ( n379486 , n31878 );
buf ( n379487 , n379486 );
xor ( n31881 , n379484 , n379487 );
buf ( n379489 , n364834 );
not ( n31883 , n379489 );
buf ( n379491 , n576 );
buf ( n379492 , n29487 );
xor ( n31886 , n379491 , n379492 );
buf ( n379494 , n31886 );
buf ( n379495 , n379494 );
not ( n31889 , n379495 );
or ( n31890 , n31883 , n31889 );
buf ( n379498 , n379366 );
buf ( n379499 , n377023 );
nand ( n31893 , n379498 , n379499 );
buf ( n379501 , n31893 );
buf ( n379502 , n379501 );
nand ( n31896 , n31890 , n379502 );
buf ( n379504 , n31896 );
buf ( n379505 , n379504 );
xor ( n31899 , n31881 , n379505 );
buf ( n379507 , n31899 );
buf ( n379508 , n379507 );
xor ( n31902 , n379472 , n379508 );
xor ( n31903 , n379377 , n379402 );
and ( n31904 , n31903 , n379408 );
and ( n31905 , n379377 , n379402 );
or ( n31906 , n31904 , n31905 );
buf ( n379514 , n31906 );
buf ( n379515 , n379514 );
xor ( n31909 , n31902 , n379515 );
buf ( n379517 , n31909 );
xor ( n31911 , n379352 , n379411 );
and ( n31912 , n31911 , n379418 );
and ( n31913 , n379352 , n379411 );
or ( n31914 , n31912 , n31913 );
buf ( n379522 , n31914 );
or ( n31916 , n379517 , n379522 );
buf ( n379524 , n379522 );
buf ( n379525 , n379517 );
nand ( n31919 , n379524 , n379525 );
buf ( n379527 , n31919 );
nand ( n31921 , n31916 , n379527 );
buf ( n379529 , n31921 );
not ( n31923 , n379529 );
buf ( n379531 , n31923 );
not ( n31925 , n379531 );
buf ( n379533 , n31630 );
buf ( n379534 , n31690 );
or ( n31928 , n379533 , n379534 );
buf ( n379536 , n377806 );
buf ( n379537 , n379423 );
nor ( n31931 , n379536 , n379537 );
buf ( n379539 , n31931 );
buf ( n379540 , n379539 );
buf ( n31934 , n379540 );
buf ( n379542 , n31934 );
buf ( n379543 , n379542 );
nand ( n31937 , n31928 , n379543 );
buf ( n379545 , n31937 );
buf ( n379546 , n379545 );
buf ( n379547 , n379336 );
buf ( n379548 , n379431 );
or ( n31942 , n379547 , n379548 );
buf ( n379550 , n379426 );
nand ( n31944 , n31942 , n379550 );
buf ( n379552 , n31944 );
buf ( n379553 , n379552 );
buf ( n31947 , n379553 );
buf ( n379555 , n31947 );
buf ( n379556 , n379555 );
nand ( n31950 , n379546 , n379556 );
buf ( n379558 , n31950 );
buf ( n379559 , n379558 );
not ( n31953 , n379559 );
buf ( n379561 , n31953 );
not ( n31955 , n379561 );
or ( n31956 , n31925 , n31955 );
buf ( n379564 , n379558 );
buf ( n379565 , n31921 );
nand ( n31959 , n379564 , n379565 );
buf ( n379567 , n31959 );
nand ( n31961 , n31956 , n379567 );
not ( n31962 , n31961 );
not ( n31963 , n31962 );
buf ( n31964 , n31963 );
buf ( n379572 , n31964 );
not ( n31966 , n379572 );
buf ( n379574 , n31966 );
buf ( n379575 , n379574 );
not ( n31969 , n379575 );
buf ( n379577 , n31969 );
buf ( n379578 , n379577 );
not ( n31972 , n379578 );
buf ( n379580 , n351924 );
not ( n31974 , n379580 );
buf ( n379582 , n600 );
not ( n31976 , n379582 );
buf ( n379584 , n16993 );
not ( n31978 , n379584 );
buf ( n379586 , n31978 );
buf ( n379587 , n379586 );
not ( n31981 , n379587 );
or ( n31982 , n31976 , n31981 );
buf ( n379590 , n16993 );
buf ( n379591 , n4193 );
nand ( n31985 , n379590 , n379591 );
buf ( n379593 , n31985 );
buf ( n379594 , n379593 );
nand ( n31988 , n31982 , n379594 );
buf ( n379596 , n31988 );
buf ( n379597 , n379596 );
not ( n31991 , n379597 );
or ( n31992 , n31974 , n31991 );
buf ( n379600 , n600 );
not ( n31994 , n379600 );
buf ( n379602 , n16995 );
buf ( n31996 , n379602 );
buf ( n379604 , n31996 );
buf ( n379605 , n379604 );
not ( n31999 , n379605 );
buf ( n379607 , n31999 );
buf ( n379608 , n379607 );
not ( n32002 , n379608 );
or ( n32003 , n31994 , n32002 );
buf ( n379611 , n379604 );
buf ( n379612 , n4193 );
nand ( n32006 , n379611 , n379612 );
buf ( n379614 , n32006 );
buf ( n379615 , n379614 );
nand ( n32009 , n32003 , n379615 );
buf ( n379617 , n32009 );
buf ( n379618 , n379617 );
buf ( n379619 , n9751 );
nand ( n32013 , n379618 , n379619 );
buf ( n379621 , n32013 );
buf ( n379622 , n379621 );
nand ( n32016 , n31992 , n379622 );
buf ( n379624 , n32016 );
buf ( n379625 , n379624 );
buf ( n379626 , n372772 );
not ( n32020 , n379626 );
buf ( n379628 , n596 );
not ( n32022 , n379628 );
buf ( n379630 , n27797 );
not ( n32024 , n379630 );
or ( n32025 , n32022 , n32024 );
buf ( n379633 , n27137 );
buf ( n379634 , n348865 );
nand ( n32028 , n379633 , n379634 );
buf ( n379636 , n32028 );
buf ( n379637 , n379636 );
nand ( n32031 , n32025 , n379637 );
buf ( n379639 , n32031 );
buf ( n379640 , n379639 );
not ( n32034 , n379640 );
or ( n32035 , n32020 , n32034 );
buf ( n379643 , n596 );
not ( n32037 , n379643 );
buf ( n379645 , n27554 );
not ( n32039 , n379645 );
buf ( n379647 , n32039 );
buf ( n379648 , n379647 );
not ( n32042 , n379648 );
or ( n32043 , n32037 , n32042 );
buf ( n379651 , n27554 );
buf ( n379652 , n348865 );
nand ( n32046 , n379651 , n379652 );
buf ( n379654 , n32046 );
buf ( n379655 , n379654 );
nand ( n32049 , n32043 , n379655 );
buf ( n379657 , n32049 );
buf ( n379658 , n379657 );
buf ( n379659 , n347319 );
nand ( n32053 , n379658 , n379659 );
buf ( n379661 , n32053 );
buf ( n379662 , n379661 );
nand ( n32056 , n32035 , n379662 );
buf ( n379664 , n32056 );
buf ( n379665 , n379664 );
buf ( n379666 , n374674 );
buf ( n379667 , n592 );
nand ( n32061 , n379666 , n379667 );
buf ( n379669 , n32061 );
buf ( n379670 , n379669 );
not ( n32064 , n379670 );
buf ( n379672 , n32064 );
buf ( n379673 , n379672 );
xor ( n32067 , n379665 , n379673 );
buf ( n379675 , n602 );
not ( n32069 , n379675 );
buf ( n379677 , n16995 );
not ( n32071 , n379677 );
buf ( n379679 , n32071 );
buf ( n379680 , n379679 );
not ( n32074 , n379680 );
or ( n32075 , n32069 , n32074 );
buf ( n379683 , n16995 );
buf ( n379684 , n349406 );
nand ( n32078 , n379683 , n379684 );
buf ( n379686 , n32078 );
buf ( n379687 , n379686 );
nand ( n32081 , n32075 , n379687 );
buf ( n379689 , n32081 );
buf ( n379690 , n379689 );
buf ( n379691 , n354113 );
not ( n32085 , n379691 );
buf ( n379693 , n4464 );
nand ( n32087 , n32085 , n379693 );
buf ( n379695 , n32087 );
buf ( n379696 , n379695 );
nand ( n32090 , n379690 , n379696 );
buf ( n379698 , n32090 );
buf ( n379699 , n379698 );
and ( n32093 , n32067 , n379699 );
and ( n32094 , n379665 , n379673 );
or ( n32095 , n32093 , n32094 );
buf ( n379703 , n32095 );
buf ( n379704 , n379703 );
xor ( n32098 , n379625 , n379704 );
not ( n32099 , n348946 );
buf ( n379707 , n592 );
not ( n32101 , n379707 );
buf ( n379709 , n372582 );
not ( n32103 , n379709 );
or ( n32104 , n32101 , n32103 );
buf ( n379712 , n372582 );
not ( n32106 , n379712 );
buf ( n379714 , n32106 );
buf ( n379715 , n379714 );
buf ( n379716 , n348910 );
nand ( n32110 , n379715 , n379716 );
buf ( n379718 , n32110 );
buf ( n379719 , n379718 );
nand ( n32113 , n32104 , n379719 );
buf ( n379721 , n32113 );
not ( n32115 , n379721 );
or ( n32116 , n32099 , n32115 );
buf ( n379724 , n592 );
not ( n32118 , n379724 );
buf ( n379726 , n375105 );
not ( n32120 , n379726 );
or ( n32121 , n32118 , n32120 );
buf ( n379729 , n375105 );
not ( n32123 , n379729 );
buf ( n379731 , n32123 );
buf ( n379732 , n379731 );
buf ( n379733 , n348910 );
nand ( n32127 , n379732 , n379733 );
buf ( n379735 , n32127 );
buf ( n379736 , n379735 );
nand ( n32130 , n32121 , n379736 );
buf ( n379738 , n32130 );
nand ( n32132 , n379738 , n375038 );
nand ( n32133 , n32116 , n32132 );
buf ( n379741 , n32133 );
buf ( n379742 , n1397 );
not ( n32136 , n379742 );
buf ( n379744 , n594 );
not ( n32138 , n379744 );
buf ( n379746 , n17009 );
not ( n32140 , n379746 );
buf ( n379748 , n32140 );
buf ( n379749 , n379748 );
not ( n32143 , n379749 );
or ( n32144 , n32138 , n32143 );
buf ( n379752 , n17009 );
buf ( n379753 , n348975 );
nand ( n32147 , n379752 , n379753 );
buf ( n379755 , n32147 );
buf ( n379756 , n379755 );
nand ( n32150 , n32144 , n379756 );
buf ( n379758 , n32150 );
buf ( n379759 , n379758 );
not ( n32153 , n379759 );
or ( n32154 , n32136 , n32153 );
not ( n32155 , n594 );
not ( n32156 , n27797 );
or ( n32157 , n32155 , n32156 );
buf ( n379765 , n27137 );
buf ( n379766 , n348975 );
nand ( n32160 , n379765 , n379766 );
buf ( n379768 , n32160 );
nand ( n32162 , n32157 , n379768 );
nand ( n32163 , n32162 , n349035 );
buf ( n379771 , n32163 );
nand ( n32165 , n32154 , n379771 );
buf ( n379773 , n32165 );
buf ( n379774 , n379773 );
xor ( n32168 , n379741 , n379774 );
buf ( n379776 , n27516 );
buf ( n379777 , n592 );
nand ( n32171 , n379776 , n379777 );
buf ( n379779 , n32171 );
buf ( n379780 , n379779 );
xor ( n32174 , n32168 , n379780 );
buf ( n379782 , n32174 );
buf ( n379783 , n379782 );
xor ( n32177 , n32098 , n379783 );
buf ( n379785 , n32177 );
buf ( n379786 , n379785 );
buf ( n379787 , n4362 );
not ( n32181 , n379787 );
buf ( n379789 , n598 );
not ( n32183 , n379789 );
buf ( n379791 , n376520 );
not ( n32185 , n379791 );
buf ( n379793 , n32185 );
buf ( n379794 , n379793 );
not ( n32188 , n379794 );
or ( n32189 , n32183 , n32188 );
buf ( n379797 , n376526 );
not ( n32191 , n379797 );
buf ( n379799 , n32191 );
buf ( n379800 , n379799 );
buf ( n379801 , n347312 );
nand ( n32195 , n379800 , n379801 );
buf ( n379803 , n32195 );
buf ( n379804 , n379803 );
nand ( n32198 , n32189 , n379804 );
buf ( n379806 , n32198 );
buf ( n379807 , n379806 );
not ( n32201 , n379807 );
or ( n32202 , n32181 , n32201 );
buf ( n379810 , n598 );
not ( n32204 , n379810 );
not ( n32205 , n28092 );
buf ( n379813 , n32205 );
not ( n32207 , n379813 );
or ( n32208 , n32204 , n32207 );
buf ( n379816 , n28092 );
buf ( n379817 , n347312 );
nand ( n32211 , n379816 , n379817 );
buf ( n379819 , n32211 );
buf ( n379820 , n379819 );
nand ( n32214 , n32208 , n379820 );
buf ( n379822 , n32214 );
buf ( n379823 , n379822 );
buf ( n379824 , n4443 );
nand ( n32218 , n379823 , n379824 );
buf ( n379826 , n32218 );
buf ( n379827 , n379826 );
nand ( n32221 , n32202 , n379827 );
buf ( n379829 , n32221 );
buf ( n379830 , n379829 );
not ( n32224 , n347319 );
nand ( n32225 , n375441 , n348865 );
nand ( n32226 , n596 , n375435 );
nand ( n32227 , n32225 , n32226 );
not ( n32228 , n32227 );
or ( n32229 , n32224 , n32228 );
buf ( n379837 , n379657 );
buf ( n379838 , n372772 );
nand ( n32232 , n379837 , n379838 );
buf ( n379840 , n32232 );
nand ( n32234 , n32229 , n379840 );
buf ( n379842 , n32234 );
xor ( n32236 , n379830 , n379842 );
buf ( n379844 , n373283 );
buf ( n379845 , n592 );
and ( n32239 , n379844 , n379845 );
buf ( n379847 , n32239 );
buf ( n379848 , n379847 );
buf ( n379849 , n348946 );
not ( n32243 , n379849 );
buf ( n379851 , n379738 );
not ( n32245 , n379851 );
or ( n32246 , n32243 , n32245 );
buf ( n379854 , n592 );
not ( n32248 , n379854 );
buf ( n379856 , n25703 );
not ( n32250 , n379856 );
or ( n32251 , n32248 , n32250 );
buf ( n379859 , n25700 );
buf ( n379860 , n348910 );
nand ( n32254 , n379859 , n379860 );
buf ( n379862 , n32254 );
buf ( n379863 , n379862 );
nand ( n32257 , n32251 , n379863 );
buf ( n379865 , n32257 );
buf ( n379866 , n379865 );
buf ( n379867 , n375038 );
nand ( n32261 , n379866 , n379867 );
buf ( n379869 , n32261 );
buf ( n379870 , n379869 );
nand ( n32264 , n32246 , n379870 );
buf ( n379872 , n32264 );
buf ( n379873 , n379872 );
xor ( n32267 , n379848 , n379873 );
buf ( n379875 , n349035 );
not ( n32269 , n379875 );
buf ( n379877 , n379758 );
not ( n32271 , n379877 );
or ( n32272 , n32269 , n32271 );
buf ( n379880 , n594 );
not ( n32274 , n379880 );
buf ( n379882 , n372588 );
not ( n32276 , n379882 );
buf ( n379884 , n32276 );
buf ( n379885 , n379884 );
not ( n32279 , n379885 );
or ( n32280 , n32274 , n32279 );
buf ( n379888 , n372588 );
buf ( n379889 , n348975 );
nand ( n32283 , n379888 , n379889 );
buf ( n379891 , n32283 );
buf ( n379892 , n379891 );
nand ( n32286 , n32280 , n379892 );
buf ( n379894 , n32286 );
buf ( n379895 , n379894 );
buf ( n379896 , n1397 );
nand ( n32290 , n379895 , n379896 );
buf ( n379898 , n32290 );
buf ( n379899 , n379898 );
nand ( n32293 , n32272 , n379899 );
buf ( n379901 , n32293 );
buf ( n379902 , n379901 );
and ( n32296 , n32267 , n379902 );
and ( n32297 , n379848 , n379873 );
or ( n32298 , n32296 , n32297 );
buf ( n379906 , n32298 );
buf ( n379907 , n379906 );
xor ( n32301 , n32236 , n379907 );
buf ( n379909 , n32301 );
buf ( n379910 , n379909 );
buf ( n379911 , n4362 );
not ( n32305 , n379911 );
buf ( n379913 , n379822 );
not ( n32307 , n379913 );
or ( n32308 , n32305 , n32307 );
buf ( n379916 , n598 );
not ( n32310 , n379916 );
buf ( n379918 , n375435 );
not ( n32312 , n379918 );
or ( n32313 , n32310 , n32312 );
buf ( n379921 , n375441 );
buf ( n379922 , n347312 );
nand ( n32316 , n379921 , n379922 );
buf ( n379924 , n32316 );
buf ( n379925 , n379924 );
nand ( n32319 , n32313 , n379925 );
buf ( n379927 , n32319 );
buf ( n379928 , n379927 );
buf ( n379929 , n4443 );
nand ( n32323 , n379928 , n379929 );
buf ( n379931 , n32323 );
buf ( n379932 , n379931 );
nand ( n32326 , n32308 , n379932 );
buf ( n379934 , n32326 );
buf ( n379935 , n379934 );
buf ( n379936 , n9751 );
not ( n32330 , n379936 );
buf ( n379938 , n379596 );
not ( n32332 , n379938 );
or ( n32333 , n32330 , n32332 );
buf ( n379941 , n379793 );
not ( n32335 , n379941 );
buf ( n379943 , n32335 );
buf ( n379944 , n379943 );
buf ( n379945 , n358055 );
and ( n32339 , n379944 , n379945 );
buf ( n379947 , n379799 );
not ( n32341 , n379947 );
buf ( n379949 , n32341 );
buf ( n379950 , n379949 );
buf ( n379951 , n358065 );
and ( n32345 , n379950 , n379951 );
nor ( n32346 , n32339 , n32345 );
buf ( n379954 , n32346 );
buf ( n379955 , n379954 );
nand ( n32349 , n32333 , n379955 );
buf ( n379957 , n32349 );
buf ( n379958 , n379957 );
xor ( n32352 , n379935 , n379958 );
not ( n32353 , n348946 );
not ( n32354 , n379865 );
or ( n32355 , n32353 , n32354 );
buf ( n379963 , n592 );
not ( n32357 , n379963 );
buf ( n379965 , n25676 );
not ( n32359 , n379965 );
or ( n32360 , n32357 , n32359 );
buf ( n379968 , n25672 );
buf ( n379969 , n348910 );
nand ( n32363 , n379968 , n379969 );
buf ( n379971 , n32363 );
buf ( n379972 , n379971 );
nand ( n32366 , n32360 , n379972 );
buf ( n379974 , n32366 );
buf ( n379975 , n379974 );
buf ( n379976 , n375038 );
nand ( n32370 , n379975 , n379976 );
buf ( n379978 , n32370 );
nand ( n32372 , n32355 , n379978 );
buf ( n379980 , n32372 );
buf ( n379981 , n1397 );
not ( n32375 , n379981 );
buf ( n379983 , n594 );
not ( n32377 , n379983 );
buf ( n379985 , n375105 );
not ( n32379 , n379985 );
or ( n32380 , n32377 , n32379 );
buf ( n379988 , n24943 );
buf ( n379989 , n348975 );
nand ( n32383 , n379988 , n379989 );
buf ( n379991 , n32383 );
buf ( n379992 , n379991 );
nand ( n32386 , n32380 , n379992 );
buf ( n379994 , n32386 );
buf ( n379995 , n379994 );
not ( n32389 , n379995 );
or ( n32390 , n32375 , n32389 );
buf ( n379998 , n379894 );
buf ( n379999 , n349035 );
nand ( n32393 , n379998 , n379999 );
buf ( n380001 , n32393 );
buf ( n380002 , n380001 );
nand ( n32396 , n32390 , n380002 );
buf ( n380004 , n32396 );
buf ( n380005 , n380004 );
xor ( n32399 , n379980 , n380005 );
buf ( n380007 , n372772 );
not ( n32401 , n380007 );
buf ( n380009 , n596 );
not ( n32403 , n380009 );
buf ( n380011 , n379748 );
not ( n32405 , n380011 );
or ( n32406 , n32403 , n32405 );
buf ( n380014 , n17009 );
buf ( n380015 , n348865 );
nand ( n32409 , n380014 , n380015 );
buf ( n380017 , n32409 );
buf ( n380018 , n380017 );
nand ( n32412 , n32406 , n380018 );
buf ( n380020 , n32412 );
buf ( n380021 , n380020 );
not ( n32415 , n380021 );
or ( n32416 , n32401 , n32415 );
buf ( n380024 , n379639 );
buf ( n380025 , n347319 );
nand ( n32419 , n380024 , n380025 );
buf ( n380027 , n32419 );
buf ( n380028 , n380027 );
nand ( n32422 , n32416 , n380028 );
buf ( n380030 , n32422 );
buf ( n380031 , n380030 );
and ( n32425 , n32399 , n380031 );
and ( n32426 , n379980 , n380005 );
or ( n32427 , n32425 , n32426 );
buf ( n380035 , n32427 );
buf ( n380036 , n380035 );
and ( n32430 , n32352 , n380036 );
and ( n32431 , n379935 , n379958 );
or ( n32432 , n32430 , n32431 );
buf ( n380040 , n32432 );
buf ( n380041 , n380040 );
xor ( n32435 , n379910 , n380041 );
xor ( n32436 , n379848 , n379873 );
xor ( n32437 , n32436 , n379902 );
buf ( n380045 , n32437 );
buf ( n380046 , n380045 );
xor ( n32440 , n379665 , n379673 );
xor ( n32441 , n32440 , n379699 );
buf ( n380049 , n32441 );
buf ( n380050 , n380049 );
xor ( n32444 , n380046 , n380050 );
buf ( n380052 , n379669 );
buf ( n380053 , n600 );
not ( n32447 , n380053 );
buf ( n380055 , n28093 );
not ( n32449 , n380055 );
or ( n32450 , n32447 , n32449 );
buf ( n380058 , n600 );
not ( n32452 , n380058 );
buf ( n380060 , n28092 );
nand ( n32454 , n32452 , n380060 );
buf ( n380062 , n32454 );
buf ( n380063 , n380062 );
nand ( n32457 , n32450 , n380063 );
buf ( n380065 , n32457 );
buf ( n380066 , n380065 );
buf ( n380067 , n351924 );
nand ( n32461 , n380066 , n380067 );
buf ( n380069 , n32461 );
buf ( n380070 , n380069 );
buf ( n380071 , n379793 );
buf ( n380072 , n373257 );
nand ( n32466 , n380071 , n380072 );
buf ( n380074 , n32466 );
buf ( n380075 , n380074 );
buf ( n380076 , n379943 );
buf ( n380077 , n373251 );
nand ( n32471 , n380076 , n380077 );
buf ( n380079 , n32471 );
buf ( n380080 , n380079 );
nand ( n32474 , n380070 , n380075 , n380080 );
buf ( n380082 , n32474 );
buf ( n380083 , n380082 );
xor ( n32477 , n380052 , n380083 );
buf ( n380085 , n4362 );
not ( n32479 , n380085 );
buf ( n380087 , n379927 );
not ( n32481 , n380087 );
or ( n32482 , n32479 , n32481 );
buf ( n380090 , n598 );
not ( n32484 , n380090 );
buf ( n380092 , n379647 );
not ( n32486 , n380092 );
or ( n32487 , n32484 , n32486 );
buf ( n380095 , n27554 );
buf ( n380096 , n347312 );
nand ( n32490 , n380095 , n380096 );
buf ( n380098 , n32490 );
buf ( n380099 , n380098 );
nand ( n32493 , n32487 , n380099 );
buf ( n380101 , n32493 );
buf ( n380102 , n380101 );
buf ( n380103 , n4443 );
nand ( n32497 , n380102 , n380103 );
buf ( n380105 , n32497 );
buf ( n380106 , n380105 );
nand ( n32500 , n32482 , n380106 );
buf ( n380108 , n32500 );
buf ( n380109 , n380108 );
and ( n32503 , n32477 , n380109 );
and ( n32504 , n380052 , n380083 );
or ( n32505 , n32503 , n32504 );
buf ( n380113 , n32505 );
buf ( n380114 , n380113 );
and ( n32508 , n32444 , n380114 );
and ( n32509 , n380046 , n380050 );
or ( n32510 , n32508 , n32509 );
buf ( n380118 , n32510 );
buf ( n380119 , n380118 );
xor ( n32513 , n32435 , n380119 );
buf ( n380121 , n32513 );
buf ( n380122 , n380121 );
xor ( n32516 , n379786 , n380122 );
xor ( n32517 , n379935 , n379958 );
xor ( n32518 , n32517 , n380036 );
buf ( n380126 , n32518 );
buf ( n380127 , n380126 );
not ( n32521 , n379689 );
not ( n32522 , n352149 );
or ( n32523 , n32521 , n32522 );
and ( n32524 , n379586 , n358424 );
not ( n32525 , n379586 );
and ( n32526 , n32525 , n358417 );
nor ( n32527 , n32524 , n32526 );
nand ( n32528 , n32523 , n32527 );
buf ( n380136 , n32528 );
buf ( n380137 , n348946 );
not ( n32531 , n380137 );
buf ( n380139 , n379974 );
not ( n32533 , n380139 );
or ( n32534 , n32531 , n32533 );
not ( n32535 , n592 );
not ( n32536 , n25863 );
or ( n32537 , n32535 , n32536 );
buf ( n380145 , n25627 );
buf ( n380146 , n348910 );
nand ( n32540 , n380145 , n380146 );
buf ( n380148 , n32540 );
nand ( n32542 , n32537 , n380148 );
buf ( n380150 , n32542 );
buf ( n380151 , n375038 );
nand ( n32545 , n380150 , n380151 );
buf ( n380153 , n32545 );
buf ( n380154 , n380153 );
nand ( n32548 , n32534 , n380154 );
buf ( n380156 , n32548 );
buf ( n380157 , n380156 );
buf ( n380158 , n592 );
buf ( n380159 , n373806 );
and ( n32553 , n380158 , n380159 );
buf ( n380161 , n32553 );
buf ( n380162 , n380161 );
xor ( n32556 , n380157 , n380162 );
buf ( n380164 , n349035 );
not ( n32558 , n380164 );
buf ( n380166 , n379994 );
not ( n32560 , n380166 );
or ( n32561 , n32558 , n32560 );
buf ( n380169 , n594 );
not ( n32563 , n380169 );
buf ( n380171 , n25703 );
not ( n32565 , n380171 );
or ( n32566 , n32563 , n32565 );
buf ( n380174 , n25700 );
buf ( n380175 , n348975 );
nand ( n32569 , n380174 , n380175 );
buf ( n380177 , n32569 );
buf ( n380178 , n380177 );
nand ( n32572 , n32566 , n380178 );
buf ( n380180 , n32572 );
buf ( n380181 , n380180 );
buf ( n380182 , n1397 );
nand ( n32576 , n380181 , n380182 );
buf ( n380184 , n32576 );
buf ( n380185 , n380184 );
nand ( n32579 , n32561 , n380185 );
buf ( n380187 , n32579 );
buf ( n380188 , n380187 );
and ( n32582 , n32556 , n380188 );
and ( n32583 , n380157 , n380162 );
or ( n32584 , n32582 , n32583 );
buf ( n380192 , n32584 );
buf ( n380193 , n380192 );
xor ( n32587 , n380136 , n380193 );
buf ( n380195 , n347319 );
not ( n32589 , n380195 );
buf ( n380197 , n380020 );
not ( n32591 , n380197 );
or ( n32592 , n32589 , n32591 );
buf ( n380200 , n596 );
not ( n32594 , n380200 );
buf ( n380202 , n372582 );
not ( n32596 , n380202 );
or ( n32597 , n32594 , n32596 );
buf ( n380205 , n379714 );
buf ( n380206 , n348865 );
nand ( n32600 , n380205 , n380206 );
buf ( n380208 , n32600 );
buf ( n380209 , n380208 );
nand ( n32603 , n32597 , n380209 );
buf ( n380211 , n32603 );
buf ( n380212 , n380211 );
buf ( n380213 , n372772 );
nand ( n32607 , n380212 , n380213 );
buf ( n380215 , n32607 );
buf ( n380216 , n380215 );
nand ( n32610 , n32592 , n380216 );
buf ( n380218 , n32610 );
buf ( n380219 , n380218 );
not ( n32613 , n1397 );
not ( n32614 , n594 );
not ( n32615 , n25676 );
or ( n32616 , n32614 , n32615 );
buf ( n380224 , n25672 );
buf ( n380225 , n348975 );
nand ( n32619 , n380224 , n380225 );
buf ( n380227 , n32619 );
nand ( n32621 , n32616 , n380227 );
not ( n32622 , n32621 );
or ( n32623 , n32613 , n32622 );
buf ( n380231 , n380180 );
buf ( n380232 , n349035 );
nand ( n32626 , n380231 , n380232 );
buf ( n380234 , n32626 );
nand ( n32628 , n32623 , n380234 );
buf ( n380236 , n32628 );
xor ( n32630 , n380219 , n380236 );
not ( n32631 , n4362 );
not ( n32632 , n380101 );
or ( n32633 , n32631 , n32632 );
buf ( n380241 , n27137 );
buf ( n380242 , n347312 );
nand ( n32636 , n380241 , n380242 );
buf ( n380244 , n32636 );
nand ( n32638 , n27797 , n598 );
nand ( n32639 , n380244 , n32638 );
nand ( n32640 , n32639 , n4443 );
nand ( n32641 , n32633 , n32640 );
buf ( n380249 , n32641 );
and ( n32643 , n32630 , n380249 );
and ( n32644 , n380219 , n380236 );
or ( n32645 , n32643 , n32644 );
buf ( n380253 , n32645 );
buf ( n380254 , n380253 );
and ( n32648 , n32587 , n380254 );
and ( n32649 , n380136 , n380193 );
or ( n32650 , n32648 , n32649 );
buf ( n380258 , n32650 );
buf ( n380259 , n380258 );
xor ( n32653 , n380127 , n380259 );
xor ( n32654 , n379980 , n380005 );
xor ( n32655 , n32654 , n380031 );
buf ( n380263 , n32655 );
buf ( n380264 , n380263 );
xor ( n32658 , n380052 , n380083 );
xor ( n32659 , n32658 , n380109 );
buf ( n380267 , n32659 );
buf ( n380268 , n380267 );
xor ( n32662 , n380264 , n380268 );
buf ( n380270 , n351924 );
not ( n32664 , n380270 );
and ( n32665 , n600 , n375435 );
not ( n32666 , n600 );
and ( n32667 , n32666 , n376567 );
or ( n32668 , n32665 , n32667 );
buf ( n380276 , n32668 );
not ( n32670 , n380276 );
or ( n32671 , n32664 , n32670 );
and ( n32672 , n28092 , n373251 );
not ( n32673 , n28092 );
and ( n32674 , n32673 , n373257 );
nor ( n32675 , n32672 , n32674 );
buf ( n380283 , n32675 );
nand ( n32677 , n32671 , n380283 );
buf ( n380285 , n32677 );
buf ( n380286 , n380285 );
xor ( n32680 , n604 , n16995 );
buf ( n380288 , n32680 );
buf ( n380289 , n355075 );
not ( n32683 , n380289 );
buf ( n380291 , n358937 );
nand ( n32685 , n32683 , n380291 );
buf ( n380293 , n32685 );
buf ( n380294 , n380293 );
nand ( n32688 , n380288 , n380294 );
buf ( n380296 , n32688 );
buf ( n380297 , n380296 );
xor ( n32691 , n380286 , n380297 );
xor ( n32692 , n380157 , n380162 );
xor ( n32693 , n32692 , n380188 );
buf ( n380301 , n32693 );
buf ( n380302 , n380301 );
and ( n32696 , n32691 , n380302 );
and ( n32697 , n380286 , n380297 );
or ( n32698 , n32696 , n32697 );
buf ( n380306 , n32698 );
buf ( n380307 , n380306 );
and ( n32701 , n32662 , n380307 );
and ( n32702 , n380264 , n380268 );
or ( n32703 , n32701 , n32702 );
buf ( n380311 , n32703 );
buf ( n380312 , n380311 );
and ( n32706 , n32653 , n380312 );
and ( n32707 , n380127 , n380259 );
or ( n32708 , n32706 , n32707 );
buf ( n380316 , n32708 );
buf ( n380317 , n380316 );
xor ( n32711 , n32516 , n380317 );
buf ( n380319 , n32711 );
not ( n32713 , n380319 );
xor ( n32714 , n380046 , n380050 );
xor ( n32715 , n32714 , n380114 );
buf ( n380323 , n32715 );
buf ( n380324 , n380323 );
xor ( n32718 , n380127 , n380259 );
xor ( n32719 , n32718 , n380312 );
buf ( n380327 , n32719 );
buf ( n380328 , n380327 );
xor ( n32722 , n380324 , n380328 );
xor ( n32723 , n380136 , n380193 );
xor ( n32724 , n32723 , n380254 );
buf ( n380332 , n32724 );
buf ( n380333 , n380332 );
buf ( n380334 , n602 );
not ( n32728 , n380334 );
buf ( n380336 , n379793 );
not ( n32730 , n380336 );
or ( n32731 , n32728 , n32730 );
buf ( n380339 , n376520 );
buf ( n380340 , n349406 );
nand ( n32734 , n380339 , n380340 );
buf ( n380342 , n32734 );
buf ( n380343 , n380342 );
nand ( n32737 , n32731 , n380343 );
buf ( n380345 , n32737 );
buf ( n380346 , n380345 );
buf ( n380347 , n354113 );
nand ( n32741 , n380346 , n380347 );
buf ( n380349 , n32741 );
buf ( n380350 , n380349 );
buf ( n380351 , n16993 );
not ( n32745 , n380351 );
buf ( n380353 , n32745 );
buf ( n380354 , n380353 );
buf ( n380355 , n373176 );
nand ( n32749 , n380354 , n380355 );
buf ( n380357 , n32749 );
buf ( n380358 , n380357 );
buf ( n380359 , n16993 );
not ( n32753 , n380359 );
buf ( n380361 , n32753 );
buf ( n380362 , n380361 );
not ( n32756 , n380362 );
buf ( n380364 , n32756 );
buf ( n380365 , n380364 );
buf ( n380366 , n373187 );
nand ( n32760 , n380365 , n380366 );
buf ( n380368 , n32760 );
buf ( n380369 , n380368 );
nand ( n32763 , n380350 , n380358 , n380369 );
buf ( n380371 , n32763 );
buf ( n380372 , n380371 );
buf ( n380373 , n375038 );
not ( n32767 , n380373 );
xor ( n32768 , n380158 , n380159 );
buf ( n380376 , n32768 );
buf ( n380377 , n380376 );
not ( n32771 , n380377 );
or ( n32772 , n32767 , n32771 );
buf ( n380380 , n32542 );
buf ( n380381 , n348946 );
nand ( n32775 , n380380 , n380381 );
buf ( n380383 , n32775 );
buf ( n380384 , n380383 );
nand ( n32778 , n32772 , n380384 );
buf ( n380386 , n32778 );
buf ( n380387 , n380386 );
buf ( n380388 , n592 );
buf ( n380389 , n374656 );
and ( n32783 , n380388 , n380389 );
buf ( n380391 , n32783 );
buf ( n380392 , n380391 );
xor ( n32786 , n380387 , n380392 );
buf ( n380394 , n372772 );
not ( n32788 , n380394 );
and ( n32789 , n372550 , n596 );
not ( n32790 , n372550 );
and ( n32791 , n32790 , n348865 );
or ( n32792 , n32789 , n32791 );
buf ( n380400 , n32792 );
not ( n32794 , n380400 );
or ( n32795 , n32788 , n32794 );
buf ( n380403 , n380211 );
buf ( n380404 , n347319 );
nand ( n32798 , n380403 , n380404 );
buf ( n380406 , n32798 );
buf ( n380407 , n380406 );
nand ( n32801 , n32795 , n380407 );
buf ( n380409 , n32801 );
buf ( n380410 , n380409 );
and ( n32804 , n32786 , n380410 );
and ( n32805 , n380387 , n380392 );
or ( n32806 , n32804 , n32805 );
buf ( n380414 , n32806 );
buf ( n380415 , n380414 );
xor ( n32809 , n380372 , n380415 );
not ( n32810 , n9637 );
nand ( n32811 , n32810 , n592 );
buf ( n380419 , n32811 );
not ( n32813 , n380419 );
buf ( n380421 , n32813 );
buf ( n380422 , n380421 );
buf ( n380423 , n32628 );
not ( n32817 , n380423 );
buf ( n380425 , n32817 );
buf ( n380426 , n380425 );
xor ( n32820 , n380422 , n380426 );
buf ( n380428 , n4362 );
not ( n32822 , n380428 );
buf ( n380430 , n32639 );
not ( n32824 , n380430 );
or ( n32825 , n32822 , n32824 );
buf ( n380433 , n598 );
not ( n32827 , n380433 );
buf ( n380435 , n379748 );
not ( n32829 , n380435 );
or ( n32830 , n32827 , n32829 );
buf ( n380438 , n17009 );
buf ( n380439 , n347312 );
nand ( n32833 , n380438 , n380439 );
buf ( n380441 , n32833 );
buf ( n380442 , n380441 );
nand ( n32836 , n32830 , n380442 );
buf ( n380444 , n32836 );
buf ( n380445 , n380444 );
buf ( n380446 , n4443 );
nand ( n32840 , n380445 , n380446 );
buf ( n380448 , n32840 );
buf ( n380449 , n380448 );
nand ( n32843 , n32825 , n380449 );
buf ( n380451 , n32843 );
buf ( n380452 , n380451 );
and ( n32846 , n32820 , n380452 );
and ( n32847 , n380422 , n380426 );
or ( n32848 , n32846 , n32847 );
buf ( n380456 , n32848 );
buf ( n380457 , n380456 );
and ( n32851 , n32809 , n380457 );
and ( n32852 , n380372 , n380415 );
or ( n32853 , n32851 , n32852 );
buf ( n380461 , n32853 );
buf ( n380462 , n380461 );
xor ( n32856 , n380333 , n380462 );
xor ( n32857 , n380219 , n380236 );
xor ( n32858 , n32857 , n380249 );
buf ( n380466 , n32858 );
buf ( n380467 , n380466 );
xor ( n32861 , n380286 , n380297 );
xor ( n32862 , n32861 , n380302 );
buf ( n380470 , n32862 );
buf ( n380471 , n380470 );
xor ( n32865 , n380467 , n380471 );
buf ( n380473 , n352149 );
not ( n32867 , n380473 );
buf ( n380475 , n380345 );
not ( n32869 , n380475 );
or ( n32870 , n32867 , n32869 );
buf ( n380478 , n602 );
not ( n32872 , n380478 );
buf ( n380480 , n32205 );
not ( n32874 , n380480 );
or ( n32875 , n32872 , n32874 );
buf ( n380483 , n28092 );
buf ( n380484 , n349406 );
nand ( n32878 , n380483 , n380484 );
buf ( n380486 , n32878 );
buf ( n380487 , n380486 );
nand ( n32881 , n32875 , n380487 );
buf ( n380489 , n32881 );
buf ( n380490 , n380489 );
buf ( n380491 , n354113 );
nand ( n32885 , n380490 , n380491 );
buf ( n380493 , n32885 );
buf ( n380494 , n380493 );
nand ( n32888 , n32870 , n380494 );
buf ( n380496 , n32888 );
buf ( n380497 , n380496 );
buf ( n380498 , n1722 );
not ( n32892 , n380498 );
buf ( n380500 , n32668 );
not ( n32894 , n380500 );
or ( n32895 , n32892 , n32894 );
buf ( n380503 , n600 );
not ( n32897 , n380503 );
buf ( n380505 , n375161 );
not ( n32899 , n380505 );
or ( n32900 , n32897 , n32899 );
buf ( n380508 , n27554 );
buf ( n380509 , n4193 );
nand ( n32903 , n380508 , n380509 );
buf ( n380511 , n32903 );
buf ( n380512 , n380511 );
nand ( n32906 , n32900 , n380512 );
buf ( n380514 , n32906 );
buf ( n380515 , n380514 );
buf ( n380516 , n351924 );
nand ( n32910 , n380515 , n380516 );
buf ( n380518 , n32910 );
buf ( n380519 , n380518 );
nand ( n32913 , n32895 , n380519 );
buf ( n380521 , n32913 );
buf ( n380522 , n380521 );
xor ( n32916 , n380497 , n380522 );
xor ( n32917 , n380387 , n380392 );
xor ( n32918 , n32917 , n380410 );
buf ( n380526 , n32918 );
buf ( n380527 , n380526 );
and ( n32921 , n32916 , n380527 );
and ( n32922 , n380497 , n380522 );
or ( n32923 , n32921 , n32922 );
buf ( n380531 , n32923 );
buf ( n380532 , n380531 );
and ( n32926 , n32865 , n380532 );
and ( n32927 , n380467 , n380471 );
or ( n32928 , n32926 , n32927 );
buf ( n380536 , n32928 );
buf ( n380537 , n380536 );
and ( n32931 , n32856 , n380537 );
and ( n32932 , n380333 , n380462 );
or ( n32933 , n32931 , n32932 );
buf ( n380541 , n32933 );
buf ( n380542 , n380541 );
and ( n32936 , n32722 , n380542 );
and ( n32937 , n380324 , n380328 );
or ( n32938 , n32936 , n32937 );
buf ( n380546 , n32938 );
not ( n32940 , n380546 );
and ( n32941 , n32713 , n32940 );
xor ( n32942 , n380264 , n380268 );
xor ( n32943 , n32942 , n380307 );
buf ( n380551 , n32943 );
buf ( n380552 , n380551 );
xor ( n32946 , n380333 , n380462 );
xor ( n32947 , n32946 , n380537 );
buf ( n380555 , n32947 );
buf ( n380556 , n380555 );
xor ( n32950 , n380552 , n380556 );
xor ( n32951 , n380372 , n380415 );
xor ( n32952 , n32951 , n380457 );
buf ( n380560 , n32952 );
buf ( n380561 , n380560 );
buf ( n380562 , n355075 );
not ( n32956 , n380562 );
buf ( n380564 , n604 );
buf ( n380565 , n16993 );
and ( n32959 , n380564 , n380565 );
not ( n32960 , n380564 );
buf ( n380568 , n380361 );
and ( n32962 , n32960 , n380568 );
nor ( n32963 , n32959 , n32962 );
buf ( n380571 , n32963 );
buf ( n380572 , n380571 );
not ( n32966 , n380572 );
or ( n32967 , n32956 , n32966 );
buf ( n380575 , n32680 );
buf ( n380576 , n6600 );
nand ( n32970 , n380575 , n380576 );
buf ( n380578 , n32970 );
buf ( n380579 , n380578 );
nand ( n32973 , n32967 , n380579 );
buf ( n380581 , n32973 );
buf ( n380582 , n380581 );
buf ( n380583 , n1397 );
not ( n32977 , n380583 );
buf ( n380585 , n594 );
not ( n32979 , n380585 );
buf ( n380587 , n374042 );
not ( n32981 , n380587 );
or ( n32982 , n32979 , n32981 );
buf ( n380590 , n25627 );
buf ( n380591 , n348975 );
nand ( n32985 , n380590 , n380591 );
buf ( n380593 , n32985 );
buf ( n380594 , n380593 );
nand ( n32988 , n32982 , n380594 );
buf ( n380596 , n32988 );
buf ( n380597 , n380596 );
not ( n32991 , n380597 );
or ( n32992 , n32977 , n32991 );
nand ( n32993 , n32621 , n349035 );
buf ( n380601 , n32993 );
nand ( n32995 , n32992 , n380601 );
buf ( n380603 , n32995 );
buf ( n380604 , n380603 );
buf ( n380605 , n348946 );
not ( n32999 , n380605 );
buf ( n380607 , n380376 );
not ( n33001 , n380607 );
or ( n33002 , n32999 , n33001 );
xor ( n33003 , n380388 , n380389 );
buf ( n380611 , n33003 );
buf ( n380612 , n380611 );
buf ( n380613 , n375038 );
nand ( n33007 , n380612 , n380613 );
buf ( n380615 , n33007 );
buf ( n380616 , n380615 );
nand ( n33010 , n33002 , n380616 );
buf ( n380618 , n33010 );
buf ( n380619 , n380618 );
xor ( n33013 , n380604 , n380619 );
buf ( n380621 , n347319 );
not ( n33015 , n380621 );
buf ( n380623 , n32792 );
not ( n33017 , n380623 );
or ( n33018 , n33015 , n33017 );
buf ( n380626 , n596 );
not ( n33020 , n380626 );
buf ( n380628 , n25741 );
not ( n33022 , n380628 );
or ( n33023 , n33020 , n33022 );
buf ( n380631 , n25700 );
buf ( n380632 , n348865 );
nand ( n33026 , n380631 , n380632 );
buf ( n380634 , n33026 );
buf ( n380635 , n380634 );
nand ( n33029 , n33023 , n380635 );
buf ( n380637 , n33029 );
buf ( n380638 , n380637 );
buf ( n380639 , n372772 );
nand ( n33033 , n380638 , n380639 );
buf ( n380641 , n33033 );
buf ( n380642 , n380641 );
nand ( n33036 , n33018 , n380642 );
buf ( n380644 , n33036 );
buf ( n380645 , n380644 );
and ( n33039 , n33013 , n380645 );
and ( n33040 , n380604 , n380619 );
or ( n33041 , n33039 , n33040 );
buf ( n380649 , n33041 );
buf ( n380650 , n380649 );
xor ( n33044 , n380582 , n380650 );
buf ( n380652 , n32811 );
buf ( n380653 , n4362 );
not ( n33047 , n380653 );
buf ( n380655 , n380444 );
not ( n33049 , n380655 );
or ( n33050 , n33047 , n33049 );
buf ( n380658 , n598 );
not ( n33052 , n380658 );
buf ( n380660 , n379884 );
not ( n33054 , n380660 );
or ( n33055 , n33052 , n33054 );
buf ( n380663 , n379714 );
buf ( n380664 , n347312 );
nand ( n33058 , n380663 , n380664 );
buf ( n380666 , n33058 );
buf ( n380667 , n380666 );
nand ( n33061 , n33055 , n380667 );
buf ( n380669 , n33061 );
buf ( n380670 , n380669 );
buf ( n380671 , n4443 );
nand ( n33065 , n380670 , n380671 );
buf ( n380673 , n33065 );
buf ( n380674 , n380673 );
nand ( n33068 , n33050 , n380674 );
buf ( n380676 , n33068 );
buf ( n380677 , n380676 );
xor ( n33071 , n380652 , n380677 );
buf ( n380679 , n351924 );
not ( n33073 , n380679 );
and ( n33074 , n600 , n27134 );
not ( n33075 , n600 );
and ( n33076 , n33075 , n27137 );
or ( n33077 , n33074 , n33076 );
buf ( n380685 , n33077 );
not ( n33079 , n380685 );
or ( n33080 , n33073 , n33079 );
buf ( n380688 , n380514 );
buf ( n380689 , n9751 );
nand ( n33083 , n380688 , n380689 );
buf ( n380691 , n33083 );
buf ( n380692 , n380691 );
nand ( n33086 , n33080 , n380692 );
buf ( n380694 , n33086 );
buf ( n380695 , n380694 );
and ( n33089 , n33071 , n380695 );
and ( n33090 , n380652 , n380677 );
or ( n33091 , n33089 , n33090 );
buf ( n380699 , n33091 );
buf ( n380700 , n380699 );
and ( n33094 , n33044 , n380700 );
and ( n33095 , n380582 , n380650 );
or ( n33096 , n33094 , n33095 );
buf ( n380704 , n33096 );
buf ( n380705 , n380704 );
xor ( n33099 , n380561 , n380705 );
xor ( n33100 , n380422 , n380426 );
xor ( n33101 , n33100 , n380452 );
buf ( n380709 , n33101 );
buf ( n380710 , n380709 );
buf ( n380711 , n354113 );
not ( n33105 , n380711 );
xor ( n33106 , n375435 , n349406 );
buf ( n380714 , n33106 );
not ( n33108 , n380714 );
or ( n33109 , n33105 , n33108 );
buf ( n380717 , n602 );
not ( n33111 , n380717 );
buf ( n380719 , n28093 );
not ( n33113 , n380719 );
or ( n33114 , n33111 , n33113 );
buf ( n380722 , n380486 );
nand ( n33116 , n33114 , n380722 );
buf ( n380724 , n33116 );
buf ( n380725 , n380724 );
buf ( n380726 , n352149 );
nand ( n33120 , n380725 , n380726 );
buf ( n380728 , n33120 );
buf ( n380729 , n380728 );
nand ( n33123 , n33109 , n380729 );
buf ( n380731 , n33123 );
buf ( n380732 , n380731 );
buf ( n380733 , n9664 );
buf ( n380734 , n592 );
and ( n33128 , n380733 , n380734 );
buf ( n380736 , n33128 );
buf ( n380737 , n380736 );
buf ( n380738 , n372772 );
not ( n33132 , n380738 );
buf ( n380740 , n596 );
not ( n33134 , n380740 );
buf ( n380742 , n25676 );
not ( n33136 , n380742 );
or ( n33137 , n33134 , n33136 );
buf ( n380745 , n25672 );
buf ( n380746 , n348865 );
nand ( n33140 , n380745 , n380746 );
buf ( n380748 , n33140 );
buf ( n380749 , n380748 );
nand ( n33143 , n33137 , n380749 );
buf ( n380751 , n33143 );
buf ( n380752 , n380751 );
not ( n33146 , n380752 );
or ( n33147 , n33132 , n33146 );
buf ( n380755 , n380637 );
buf ( n380756 , n347319 );
nand ( n33150 , n380755 , n380756 );
buf ( n380758 , n33150 );
buf ( n380759 , n380758 );
nand ( n33153 , n33147 , n380759 );
buf ( n380761 , n33153 );
buf ( n380762 , n380761 );
xor ( n33156 , n380737 , n380762 );
buf ( n380764 , n348946 );
not ( n33158 , n380764 );
buf ( n380766 , n380611 );
not ( n33160 , n380766 );
or ( n33161 , n33158 , n33160 );
buf ( n380769 , n592 );
not ( n33163 , n380769 );
buf ( n380771 , n9637 );
not ( n33165 , n380771 );
or ( n33166 , n33163 , n33165 );
buf ( n380774 , n9636 );
buf ( n380775 , n348910 );
nand ( n33169 , n380774 , n380775 );
buf ( n380777 , n33169 );
buf ( n380778 , n380777 );
nand ( n33172 , n33166 , n380778 );
buf ( n380780 , n33172 );
buf ( n380781 , n380780 );
buf ( n380782 , n375038 );
nand ( n33176 , n380781 , n380782 );
buf ( n380784 , n33176 );
buf ( n380785 , n380784 );
nand ( n33179 , n33161 , n380785 );
buf ( n380787 , n33179 );
buf ( n380788 , n380787 );
and ( n33182 , n33156 , n380788 );
and ( n33183 , n380737 , n380762 );
or ( n33184 , n33182 , n33183 );
buf ( n380792 , n33184 );
buf ( n380793 , n380792 );
xor ( n33187 , n380732 , n380793 );
buf ( n380795 , n606 );
not ( n33189 , n380795 );
buf ( n380797 , n379679 );
not ( n33191 , n380797 );
or ( n33192 , n33189 , n33191 );
buf ( n380800 , n16995 );
buf ( n380801 , n9642 );
nand ( n33195 , n380800 , n380801 );
buf ( n380803 , n33195 );
buf ( n380804 , n380803 );
nand ( n33198 , n33192 , n380804 );
buf ( n380806 , n33198 );
buf ( n380807 , n380806 );
buf ( n380808 , n357376 );
not ( n33202 , n380808 );
buf ( n380810 , n358969 );
nand ( n33204 , n33202 , n380810 );
buf ( n380812 , n33204 );
buf ( n380813 , n380812 );
nand ( n33207 , n380807 , n380813 );
buf ( n380815 , n33207 );
buf ( n380816 , n380815 );
and ( n33210 , n33187 , n380816 );
and ( n33211 , n380732 , n380793 );
or ( n33212 , n33210 , n33211 );
buf ( n380820 , n33212 );
buf ( n380821 , n380820 );
xor ( n33215 , n380710 , n380821 );
xor ( n33216 , n380497 , n380522 );
xor ( n33217 , n33216 , n380527 );
buf ( n380825 , n33217 );
buf ( n380826 , n380825 );
and ( n33220 , n33215 , n380826 );
and ( n33221 , n380710 , n380821 );
or ( n33222 , n33220 , n33221 );
buf ( n380830 , n33222 );
buf ( n380831 , n380830 );
and ( n33225 , n33099 , n380831 );
and ( n33226 , n380561 , n380705 );
or ( n33227 , n33225 , n33226 );
buf ( n380835 , n33227 );
buf ( n380836 , n380835 );
and ( n33230 , n32950 , n380836 );
and ( n33231 , n380552 , n380556 );
or ( n33232 , n33230 , n33231 );
buf ( n380840 , n33232 );
buf ( n380841 , n380840 );
xor ( n33235 , n380324 , n380328 );
xor ( n33236 , n33235 , n380542 );
buf ( n380844 , n33236 );
buf ( n380845 , n380844 );
nor ( n33239 , n380841 , n380845 );
buf ( n380847 , n33239 );
nor ( n33241 , n32941 , n380847 );
xor ( n33242 , n379625 , n379704 );
and ( n33243 , n33242 , n379783 );
and ( n33244 , n379625 , n379704 );
or ( n33245 , n33243 , n33244 );
buf ( n380853 , n33245 );
buf ( n380854 , n380853 );
xor ( n33248 , n379830 , n379842 );
and ( n33249 , n33248 , n379907 );
and ( n33250 , n379830 , n379842 );
or ( n33251 , n33249 , n33250 );
buf ( n380859 , n33251 );
buf ( n380860 , n380859 );
buf ( n380861 , n349035 );
not ( n33255 , n380861 );
buf ( n380863 , n594 );
not ( n33257 , n380863 );
buf ( n380865 , n379647 );
not ( n33259 , n380865 );
or ( n33260 , n33257 , n33259 );
buf ( n380868 , n27554 );
buf ( n380869 , n348975 );
nand ( n33263 , n380868 , n380869 );
buf ( n380871 , n33263 );
buf ( n380872 , n380871 );
nand ( n33266 , n33260 , n380872 );
buf ( n380874 , n33266 );
buf ( n380875 , n380874 );
not ( n33269 , n380875 );
or ( n33270 , n33255 , n33269 );
nand ( n33271 , n32162 , n1397 );
buf ( n380879 , n33271 );
nand ( n33273 , n33270 , n380879 );
buf ( n380881 , n33273 );
buf ( n380882 , n380881 );
buf ( n380883 , n358041 );
not ( n33277 , n380883 );
buf ( n380885 , n351924 );
not ( n33279 , n380885 );
buf ( n380887 , n33279 );
buf ( n380888 , n380887 );
not ( n33282 , n380888 );
or ( n33283 , n33277 , n33282 );
buf ( n380891 , n379617 );
nand ( n33285 , n33283 , n380891 );
buf ( n380893 , n33285 );
buf ( n380894 , n380893 );
xor ( n33288 , n380882 , n380894 );
buf ( n380896 , n372772 );
not ( n33290 , n380896 );
buf ( n380898 , n32227 );
not ( n33292 , n380898 );
or ( n33293 , n33290 , n33292 );
buf ( n380901 , n596 );
not ( n33295 , n380901 );
buf ( n380903 , n32205 );
not ( n33297 , n380903 );
or ( n33298 , n33295 , n33297 );
not ( n33299 , n32205 );
buf ( n380907 , n33299 );
buf ( n380908 , n348865 );
nand ( n33302 , n380907 , n380908 );
buf ( n380910 , n33302 );
buf ( n380911 , n380910 );
nand ( n33305 , n33298 , n380911 );
buf ( n380913 , n33305 );
buf ( n380914 , n380913 );
buf ( n380915 , n347319 );
nand ( n33309 , n380914 , n380915 );
buf ( n380917 , n33309 );
buf ( n380918 , n380917 );
nand ( n33312 , n33293 , n380918 );
buf ( n380920 , n33312 );
buf ( n380921 , n380920 );
xor ( n33315 , n33288 , n380921 );
buf ( n380923 , n33315 );
buf ( n380924 , n380923 );
xor ( n33318 , n380860 , n380924 );
buf ( n380926 , n4362 );
not ( n33320 , n380926 );
buf ( n380928 , n598 );
not ( n33322 , n380928 );
buf ( n380930 , n379586 );
not ( n33324 , n380930 );
or ( n33325 , n33322 , n33324 );
buf ( n380933 , n380364 );
buf ( n380934 , n347312 );
nand ( n33328 , n380933 , n380934 );
buf ( n380936 , n33328 );
buf ( n380937 , n380936 );
nand ( n33331 , n33325 , n380937 );
buf ( n380939 , n33331 );
buf ( n380940 , n380939 );
not ( n33334 , n380940 );
or ( n33335 , n33320 , n33334 );
buf ( n380943 , n379806 );
buf ( n380944 , n4443 );
nand ( n33338 , n380943 , n380944 );
buf ( n380946 , n33338 );
buf ( n380947 , n380946 );
nand ( n33341 , n33335 , n380947 );
buf ( n380949 , n33341 );
buf ( n380950 , n380949 );
xor ( n33344 , n379741 , n379774 );
and ( n33345 , n33344 , n379780 );
and ( n33346 , n379741 , n379774 );
or ( n33347 , n33345 , n33346 );
buf ( n380955 , n33347 );
buf ( n380956 , n380955 );
xor ( n33350 , n380950 , n380956 );
buf ( n380958 , n348946 );
not ( n33352 , n380958 );
buf ( n380960 , n592 );
buf ( n380961 , n379748 );
not ( n33355 , n380961 );
buf ( n380963 , n33355 );
buf ( n380964 , n380963 );
xor ( n33358 , n380960 , n380964 );
buf ( n380966 , n33358 );
buf ( n380967 , n380966 );
not ( n33361 , n380967 );
or ( n33362 , n33352 , n33361 );
buf ( n380970 , n379721 );
buf ( n380971 , n375038 );
nand ( n33365 , n380970 , n380971 );
buf ( n380973 , n33365 );
buf ( n380974 , n380973 );
nand ( n33368 , n33362 , n380974 );
buf ( n380976 , n33368 );
buf ( n380977 , n380976 );
buf ( n380978 , n379731 );
buf ( n380979 , n592 );
and ( n33373 , n380978 , n380979 );
buf ( n380981 , n33373 );
buf ( n380982 , n380981 );
xor ( n33376 , n380977 , n380982 );
buf ( n380984 , n379779 );
not ( n33378 , n380984 );
buf ( n380986 , n33378 );
buf ( n380987 , n380986 );
xor ( n33381 , n33376 , n380987 );
buf ( n380989 , n33381 );
buf ( n380990 , n380989 );
xor ( n33384 , n33350 , n380990 );
buf ( n380992 , n33384 );
buf ( n380993 , n380992 );
xor ( n33387 , n33318 , n380993 );
buf ( n380995 , n33387 );
buf ( n380996 , n380995 );
xor ( n33390 , n380854 , n380996 );
xor ( n33391 , n379910 , n380041 );
and ( n33392 , n33391 , n380119 );
and ( n33393 , n379910 , n380041 );
or ( n33394 , n33392 , n33393 );
buf ( n381002 , n33394 );
buf ( n381003 , n381002 );
xor ( n33397 , n33390 , n381003 );
buf ( n381005 , n33397 );
not ( n33399 , n381005 );
xor ( n33400 , n379786 , n380122 );
and ( n33401 , n33400 , n380317 );
and ( n33402 , n379786 , n380122 );
or ( n33403 , n33401 , n33402 );
buf ( n381011 , n33403 );
not ( n33405 , n381011 );
nand ( n33406 , n33399 , n33405 );
nand ( n33407 , n33241 , n33406 );
buf ( n381015 , n347319 );
not ( n33409 , n381015 );
buf ( n381017 , n596 );
not ( n33411 , n381017 );
buf ( n381019 , n379949 );
not ( n33413 , n381019 );
or ( n33414 , n33411 , n33413 );
buf ( n381022 , n379949 );
not ( n33416 , n381022 );
buf ( n381024 , n33416 );
buf ( n381025 , n381024 );
buf ( n381026 , n348865 );
nand ( n33420 , n381025 , n381026 );
buf ( n381028 , n33420 );
buf ( n381029 , n381028 );
nand ( n33423 , n33414 , n381029 );
buf ( n381031 , n33423 );
buf ( n381032 , n381031 );
not ( n33426 , n381032 );
or ( n33427 , n33409 , n33426 );
buf ( n381035 , n380913 );
buf ( n381036 , n372772 );
nand ( n33430 , n381035 , n381036 );
buf ( n381038 , n33430 );
buf ( n381039 , n381038 );
nand ( n33433 , n33427 , n381039 );
buf ( n381041 , n33433 );
buf ( n381042 , n381041 );
buf ( n381043 , n4443 );
not ( n33437 , n381043 );
buf ( n381045 , n380939 );
not ( n33439 , n381045 );
or ( n33440 , n33437 , n33439 );
buf ( n381048 , n598 );
not ( n33442 , n381048 );
buf ( n381050 , n379607 );
not ( n33444 , n381050 );
or ( n33445 , n33442 , n33444 );
buf ( n381053 , n379604 );
buf ( n381054 , n347312 );
nand ( n33448 , n381053 , n381054 );
buf ( n381056 , n33448 );
buf ( n381057 , n381056 );
nand ( n33451 , n33445 , n381057 );
buf ( n381059 , n33451 );
buf ( n381060 , n381059 );
buf ( n381061 , n4362 );
nand ( n33455 , n381060 , n381061 );
buf ( n381063 , n33455 );
buf ( n381064 , n381063 );
nand ( n33458 , n33440 , n381064 );
buf ( n381066 , n33458 );
buf ( n381067 , n381066 );
xor ( n33461 , n381042 , n381067 );
xor ( n33462 , n380977 , n380982 );
and ( n33463 , n33462 , n380987 );
and ( n33464 , n380977 , n380982 );
or ( n33465 , n33463 , n33464 );
buf ( n381073 , n33465 );
buf ( n381074 , n381073 );
xor ( n33468 , n33461 , n381074 );
buf ( n381076 , n33468 );
buf ( n381077 , n381076 );
xor ( n33471 , n380882 , n380894 );
and ( n33472 , n33471 , n380921 );
and ( n33473 , n380882 , n380894 );
or ( n33474 , n33472 , n33473 );
buf ( n381082 , n33474 );
buf ( n381083 , n381082 );
buf ( n381084 , n348946 );
not ( n33478 , n381084 );
buf ( n381086 , n592 );
not ( n33480 , n381086 );
buf ( n381088 , n27797 );
not ( n33482 , n381088 );
or ( n33483 , n33480 , n33482 );
buf ( n381091 , n27137 );
buf ( n381092 , n348910 );
nand ( n33486 , n381091 , n381092 );
buf ( n381094 , n33486 );
buf ( n381095 , n381094 );
nand ( n33489 , n33483 , n381095 );
buf ( n381097 , n33489 );
buf ( n381098 , n381097 );
not ( n33492 , n381098 );
or ( n33493 , n33478 , n33492 );
buf ( n381101 , n380966 );
buf ( n381102 , n375038 );
nand ( n33496 , n381101 , n381102 );
buf ( n381104 , n33496 );
buf ( n381105 , n381104 );
nand ( n33499 , n33493 , n381105 );
buf ( n381107 , n33499 );
buf ( n381108 , n381107 );
not ( n33502 , n349035 );
buf ( n381110 , n375441 );
buf ( n33504 , n381110 );
buf ( n381112 , n33504 );
and ( n33506 , n381112 , n594 );
not ( n33507 , n381112 );
and ( n33508 , n33507 , n348975 );
nor ( n33509 , n33506 , n33508 );
not ( n33510 , n33509 );
or ( n33511 , n33502 , n33510 );
nand ( n33512 , n380874 , n1397 );
nand ( n33513 , n33511 , n33512 );
buf ( n381121 , n33513 );
xor ( n33515 , n381108 , n381121 );
buf ( n381123 , n379714 );
buf ( n381124 , n592 );
and ( n33518 , n381123 , n381124 );
buf ( n381126 , n33518 );
buf ( n381127 , n381126 );
not ( n33521 , n381127 );
buf ( n381129 , n33521 );
buf ( n381130 , n381129 );
xor ( n33524 , n33515 , n381130 );
buf ( n381132 , n33524 );
buf ( n381133 , n381132 );
xor ( n33527 , n381083 , n381133 );
xor ( n33528 , n380950 , n380956 );
and ( n33529 , n33528 , n380990 );
and ( n33530 , n380950 , n380956 );
or ( n33531 , n33529 , n33530 );
buf ( n381139 , n33531 );
buf ( n381140 , n381139 );
xor ( n33534 , n33527 , n381140 );
buf ( n381142 , n33534 );
buf ( n381143 , n381142 );
xor ( n33537 , n381077 , n381143 );
xor ( n33538 , n380860 , n380924 );
and ( n33539 , n33538 , n380993 );
and ( n33540 , n380860 , n380924 );
or ( n33541 , n33539 , n33540 );
buf ( n381149 , n33541 );
buf ( n381150 , n381149 );
xor ( n33544 , n33537 , n381150 );
buf ( n381152 , n33544 );
xor ( n33546 , n380854 , n380996 );
and ( n33547 , n33546 , n381003 );
and ( n33548 , n380854 , n380996 );
or ( n33549 , n33547 , n33548 );
buf ( n381157 , n33549 );
nor ( n33551 , n381152 , n381157 );
buf ( n33552 , n33551 );
nor ( n33553 , n33407 , n33552 );
not ( n33554 , n33553 );
buf ( n381162 , n592 );
buf ( n381163 , n27554 );
and ( n33557 , n381162 , n381163 );
buf ( n381165 , n33557 );
buf ( n381166 , n381165 );
buf ( n381167 , n357712 );
not ( n33561 , n381167 );
buf ( n381169 , n372772 );
not ( n33563 , n381169 );
buf ( n381171 , n33563 );
buf ( n381172 , n381171 );
not ( n33566 , n381172 );
or ( n33567 , n33561 , n33566 );
buf ( n381175 , n596 );
not ( n33569 , n381175 );
buf ( n381177 , n379607 );
not ( n33571 , n381177 );
or ( n33572 , n33569 , n33571 );
buf ( n381180 , n379604 );
buf ( n381181 , n348865 );
nand ( n33575 , n381180 , n381181 );
buf ( n381183 , n33575 );
buf ( n381184 , n381183 );
nand ( n33578 , n33572 , n381184 );
buf ( n381186 , n33578 );
buf ( n381187 , n381186 );
nand ( n33581 , n33567 , n381187 );
buf ( n381189 , n33581 );
buf ( n381190 , n381189 );
xor ( n33584 , n381166 , n381190 );
buf ( n381192 , n348946 );
not ( n33586 , n381192 );
buf ( n381194 , n592 );
buf ( n381195 , n33299 );
xor ( n33589 , n381194 , n381195 );
buf ( n381197 , n33589 );
buf ( n381198 , n381197 );
not ( n33592 , n381198 );
or ( n33593 , n33586 , n33592 );
buf ( n381201 , n592 );
not ( n33595 , n381201 );
buf ( n381203 , n375435 );
not ( n33597 , n381203 );
or ( n33598 , n33595 , n33597 );
buf ( n381206 , n381112 );
buf ( n381207 , n348910 );
nand ( n33601 , n381206 , n381207 );
buf ( n381209 , n33601 );
buf ( n381210 , n381209 );
nand ( n33604 , n33598 , n381210 );
buf ( n381212 , n33604 );
buf ( n381213 , n381212 );
buf ( n381214 , n375038 );
nand ( n33608 , n381213 , n381214 );
buf ( n381216 , n33608 );
buf ( n381217 , n381216 );
nand ( n33611 , n33593 , n381217 );
buf ( n381219 , n33611 );
buf ( n381220 , n381219 );
and ( n33614 , n33584 , n381220 );
and ( n33615 , n381166 , n381190 );
or ( n33616 , n33614 , n33615 );
buf ( n381224 , n33616 );
buf ( n381225 , n381224 );
buf ( n381226 , n348946 );
not ( n33620 , n381226 );
and ( n33621 , n381024 , n348910 );
not ( n33622 , n381024 );
and ( n33623 , n33622 , n592 );
or ( n33624 , n33621 , n33623 );
buf ( n381232 , n33624 );
not ( n33626 , n381232 );
or ( n33627 , n33620 , n33626 );
buf ( n381235 , n381197 );
buf ( n381236 , n375038 );
nand ( n33630 , n381235 , n381236 );
buf ( n381238 , n33630 );
buf ( n381239 , n381238 );
nand ( n33633 , n33627 , n381239 );
buf ( n381241 , n33633 );
buf ( n381242 , n381241 );
buf ( n381243 , n1397 );
not ( n33637 , n381243 );
buf ( n381245 , n594 );
not ( n33639 , n381245 );
buf ( n381247 , n380353 );
not ( n33641 , n381247 );
or ( n33642 , n33639 , n33641 );
buf ( n381250 , n380353 );
not ( n33644 , n381250 );
buf ( n381252 , n33644 );
buf ( n381253 , n381252 );
buf ( n381254 , n348975 );
nand ( n33648 , n381253 , n381254 );
buf ( n381256 , n33648 );
buf ( n381257 , n381256 );
nand ( n33651 , n33642 , n381257 );
buf ( n381259 , n33651 );
buf ( n381260 , n381259 );
not ( n33654 , n381260 );
or ( n33655 , n33637 , n33654 );
buf ( n381263 , n594 );
not ( n33657 , n381263 );
buf ( n381265 , n379607 );
not ( n33659 , n381265 );
or ( n33660 , n33657 , n33659 );
buf ( n381268 , n379604 );
buf ( n381269 , n348975 );
nand ( n33663 , n381268 , n381269 );
buf ( n381271 , n33663 );
buf ( n381272 , n381271 );
nand ( n33666 , n33660 , n381272 );
buf ( n381274 , n33666 );
buf ( n381275 , n381274 );
buf ( n381276 , n349035 );
nand ( n33670 , n381275 , n381276 );
buf ( n381278 , n33670 );
buf ( n381279 , n381278 );
nand ( n33673 , n33655 , n381279 );
buf ( n381281 , n33673 );
buf ( n381282 , n381281 );
xor ( n33676 , n381242 , n381282 );
buf ( n381284 , n381112 );
buf ( n381285 , n592 );
nand ( n33679 , n381284 , n381285 );
buf ( n381287 , n33679 );
buf ( n381288 , n381287 );
xor ( n33682 , n33676 , n381288 );
buf ( n381290 , n33682 );
buf ( n381291 , n381290 );
xor ( n33685 , n381225 , n381291 );
buf ( n381293 , n349035 );
not ( n33687 , n381293 );
buf ( n381295 , n381259 );
not ( n33689 , n381295 );
or ( n33690 , n33687 , n33689 );
not ( n33691 , n594 );
not ( n33692 , n379793 );
or ( n33693 , n33691 , n33692 );
buf ( n381301 , n379799 );
buf ( n381302 , n348975 );
nand ( n33696 , n381301 , n381302 );
buf ( n381304 , n33696 );
nand ( n33698 , n33693 , n381304 );
nand ( n33699 , n33698 , n1397 );
buf ( n381307 , n33699 );
nand ( n33701 , n33690 , n381307 );
buf ( n381309 , n33701 );
buf ( n381310 , n381309 );
buf ( n381311 , n27137 );
buf ( n381312 , n592 );
nand ( n33706 , n381311 , n381312 );
buf ( n381314 , n33706 );
buf ( n381315 , n381314 );
not ( n33709 , n381315 );
buf ( n381317 , n33709 );
buf ( n381318 , n381317 );
xor ( n33712 , n381310 , n381318 );
xor ( n33713 , n381166 , n381190 );
xor ( n33714 , n33713 , n381220 );
buf ( n381322 , n33714 );
buf ( n381323 , n381322 );
and ( n33717 , n33712 , n381323 );
and ( n33718 , n381310 , n381318 );
or ( n33719 , n33717 , n33718 );
buf ( n381327 , n33719 );
buf ( n381328 , n381327 );
xor ( n33722 , n33685 , n381328 );
buf ( n381330 , n33722 );
not ( n33724 , n381330 );
buf ( n381332 , n348946 );
not ( n33726 , n381332 );
buf ( n381334 , n381212 );
not ( n33728 , n381334 );
or ( n33729 , n33726 , n33728 );
xor ( n33730 , n381162 , n381163 );
buf ( n381338 , n33730 );
buf ( n381339 , n381338 );
buf ( n381340 , n375038 );
nand ( n33734 , n381339 , n381340 );
buf ( n381342 , n33734 );
buf ( n381343 , n381342 );
nand ( n33737 , n33729 , n381343 );
buf ( n381345 , n33737 );
buf ( n381346 , n381345 );
buf ( n381347 , n594 );
not ( n33741 , n381347 );
buf ( n381349 , n32205 );
not ( n33743 , n381349 );
or ( n33744 , n33741 , n33743 );
buf ( n381352 , n28092 );
buf ( n381353 , n348975 );
nand ( n33747 , n381352 , n381353 );
buf ( n381355 , n33747 );
buf ( n381356 , n381355 );
nand ( n33750 , n33744 , n381356 );
buf ( n381358 , n33750 );
and ( n33752 , n381358 , n1397 );
not ( n33753 , n33752 );
nand ( n33754 , n349035 , n594 , n379793 );
not ( n33755 , n381304 );
nand ( n33756 , n33755 , n349035 );
nand ( n33757 , n33753 , n33754 , n33756 );
buf ( n381365 , n33757 );
xor ( n33759 , n381346 , n381365 );
buf ( n381367 , n372772 );
not ( n33761 , n381367 );
buf ( n381369 , n596 );
not ( n33763 , n381369 );
buf ( n381371 , n380353 );
not ( n33765 , n381371 );
or ( n33766 , n33763 , n33765 );
buf ( n381374 , n380364 );
buf ( n381375 , n348865 );
nand ( n33769 , n381374 , n381375 );
buf ( n381377 , n33769 );
buf ( n381378 , n381377 );
nand ( n33772 , n33766 , n381378 );
buf ( n381380 , n33772 );
buf ( n381381 , n381380 );
not ( n33775 , n381381 );
or ( n33776 , n33761 , n33775 );
buf ( n381384 , n381186 );
buf ( n381385 , n347319 );
nand ( n33779 , n381384 , n381385 );
buf ( n381387 , n33779 );
buf ( n381388 , n381387 );
nand ( n33782 , n33776 , n381388 );
buf ( n381390 , n33782 );
buf ( n381391 , n381390 );
and ( n33785 , n33759 , n381391 );
and ( n33786 , n381346 , n381365 );
or ( n33787 , n33785 , n33786 );
buf ( n381395 , n33787 );
buf ( n381396 , n381395 );
xor ( n33790 , n381310 , n381318 );
xor ( n33791 , n33790 , n381323 );
buf ( n381399 , n33791 );
buf ( n381400 , n381399 );
xor ( n33794 , n381396 , n381400 );
buf ( n381402 , n381314 );
and ( n33796 , n380960 , n380964 );
buf ( n381404 , n33796 );
buf ( n381405 , n381404 );
buf ( n381406 , n375038 );
not ( n33800 , n381406 );
buf ( n381408 , n381097 );
not ( n33802 , n381408 );
or ( n33803 , n33800 , n33802 );
buf ( n381411 , n381338 );
buf ( n381412 , n348946 );
nand ( n33806 , n381411 , n381412 );
buf ( n381414 , n33806 );
buf ( n381415 , n381414 );
nand ( n33809 , n33803 , n381415 );
buf ( n381417 , n33809 );
buf ( n381418 , n381417 );
xor ( n33812 , n381405 , n381418 );
buf ( n381420 , n381059 );
buf ( n381421 , n4443 );
not ( n33815 , n381421 );
buf ( n381423 , n352112 );
nand ( n33817 , n33815 , n381423 );
buf ( n381425 , n33817 );
buf ( n381426 , n381425 );
nand ( n33820 , n381420 , n381426 );
buf ( n381428 , n33820 );
buf ( n381429 , n381428 );
and ( n33823 , n33812 , n381429 );
and ( n33824 , n381405 , n381418 );
or ( n33825 , n33823 , n33824 );
buf ( n381433 , n33825 );
buf ( n381434 , n381433 );
xor ( n33828 , n381402 , n381434 );
xor ( n33829 , n381346 , n381365 );
xor ( n33830 , n33829 , n381391 );
buf ( n381438 , n33830 );
buf ( n381439 , n381438 );
and ( n33833 , n33828 , n381439 );
and ( n33834 , n381402 , n381434 );
or ( n33835 , n33833 , n33834 );
buf ( n381443 , n33835 );
buf ( n381444 , n381443 );
and ( n33838 , n33794 , n381444 );
and ( n33839 , n381396 , n381400 );
or ( n33840 , n33838 , n33839 );
buf ( n381448 , n33840 );
not ( n33842 , n381448 );
and ( n33843 , n33724 , n33842 );
xor ( n33844 , n381077 , n381143 );
and ( n33845 , n33844 , n381150 );
and ( n33846 , n381077 , n381143 );
or ( n33847 , n33845 , n33846 );
buf ( n381455 , n33847 );
xor ( n33849 , n381042 , n381067 );
and ( n33850 , n33849 , n381074 );
and ( n33851 , n381042 , n381067 );
or ( n33852 , n33850 , n33851 );
buf ( n381460 , n33852 );
buf ( n381461 , n381460 );
xor ( n33855 , n381405 , n381418 );
xor ( n33856 , n33855 , n381429 );
buf ( n381464 , n33856 );
buf ( n381465 , n381464 );
xor ( n33859 , n381108 , n381121 );
and ( n33860 , n33859 , n381130 );
and ( n33861 , n381108 , n381121 );
or ( n33862 , n33860 , n33861 );
buf ( n381470 , n33862 );
buf ( n381471 , n381470 );
xor ( n33865 , n381465 , n381471 );
buf ( n381473 , n381126 );
not ( n33867 , n1397 );
not ( n33868 , n33509 );
or ( n33869 , n33867 , n33868 );
buf ( n381477 , n381358 );
buf ( n381478 , n349035 );
nand ( n33872 , n381477 , n381478 );
buf ( n381480 , n33872 );
nand ( n33874 , n33869 , n381480 );
buf ( n381482 , n33874 );
xor ( n33876 , n381473 , n381482 );
buf ( n381484 , n347319 );
not ( n33878 , n381484 );
buf ( n381486 , n381380 );
not ( n33880 , n381486 );
or ( n33881 , n33878 , n33880 );
buf ( n381489 , n381031 );
buf ( n381490 , n372772 );
nand ( n33884 , n381489 , n381490 );
buf ( n381492 , n33884 );
buf ( n381493 , n381492 );
nand ( n33887 , n33881 , n381493 );
buf ( n381495 , n33887 );
buf ( n381496 , n381495 );
xor ( n33890 , n33876 , n381496 );
buf ( n381498 , n33890 );
buf ( n381499 , n381498 );
xor ( n33893 , n33865 , n381499 );
buf ( n381501 , n33893 );
buf ( n381502 , n381501 );
xor ( n33896 , n381461 , n381502 );
xor ( n33897 , n381083 , n381133 );
and ( n33898 , n33897 , n381140 );
and ( n33899 , n381083 , n381133 );
or ( n33900 , n33898 , n33899 );
buf ( n381508 , n33900 );
buf ( n381509 , n381508 );
xor ( n33903 , n33896 , n381509 );
buf ( n381511 , n33903 );
nor ( n33905 , n381455 , n381511 );
buf ( n381513 , n33905 );
xor ( n33907 , n381461 , n381502 );
and ( n33908 , n33907 , n381509 );
and ( n33909 , n381461 , n381502 );
or ( n33910 , n33908 , n33909 );
buf ( n381518 , n33910 );
buf ( n381519 , n381518 );
xor ( n33913 , n381473 , n381482 );
and ( n33914 , n33913 , n381496 );
and ( n33915 , n381473 , n381482 );
or ( n33916 , n33914 , n33915 );
buf ( n381524 , n33916 );
buf ( n381525 , n381524 );
xor ( n33919 , n381402 , n381434 );
xor ( n33920 , n33919 , n381439 );
buf ( n381528 , n33920 );
buf ( n381529 , n381528 );
xor ( n33923 , n381525 , n381529 );
xor ( n33924 , n381465 , n381471 );
and ( n33925 , n33924 , n381499 );
and ( n33926 , n381465 , n381471 );
or ( n33927 , n33925 , n33926 );
buf ( n381535 , n33927 );
buf ( n381536 , n381535 );
xor ( n33930 , n33923 , n381536 );
buf ( n381538 , n33930 );
buf ( n381539 , n381538 );
nor ( n33933 , n381519 , n381539 );
buf ( n381541 , n33933 );
buf ( n381542 , n381541 );
nor ( n33936 , n381513 , n381542 );
buf ( n381544 , n33936 );
buf ( n381545 , n381544 );
xor ( n33939 , n381525 , n381529 );
and ( n33940 , n33939 , n381536 );
and ( n33941 , n381525 , n381529 );
or ( n33942 , n33940 , n33941 );
buf ( n381550 , n33942 );
xor ( n33944 , n381396 , n381400 );
xor ( n33945 , n33944 , n381444 );
buf ( n381553 , n33945 );
or ( n33947 , n381550 , n381553 );
buf ( n381555 , n33947 );
nand ( n33949 , n381545 , n381555 );
buf ( n381557 , n33949 );
nor ( n33951 , n33843 , n381557 );
buf ( n381559 , n33951 );
not ( n33953 , n381559 );
buf ( n381561 , n33953 );
nor ( n33955 , n33554 , n381561 );
xor ( n33956 , n380552 , n380556 );
xor ( n33957 , n33956 , n380836 );
buf ( n381565 , n33957 );
buf ( n381566 , n381565 );
xor ( n33960 , n380467 , n380471 );
xor ( n33961 , n33960 , n380532 );
buf ( n381569 , n33961 );
buf ( n381570 , n381569 );
xor ( n33964 , n380561 , n380705 );
xor ( n33965 , n33964 , n380831 );
buf ( n381573 , n33965 );
buf ( n381574 , n381573 );
xor ( n33968 , n381570 , n381574 );
xor ( n33969 , n380582 , n380650 );
xor ( n33970 , n33969 , n380700 );
buf ( n381578 , n33970 );
buf ( n381579 , n381578 );
xor ( n33973 , n380604 , n380619 );
xor ( n33974 , n33973 , n380645 );
buf ( n381582 , n33974 );
buf ( n381583 , n381582 );
buf ( n381584 , n6600 );
not ( n33978 , n381584 );
buf ( n381586 , n380571 );
not ( n33980 , n381586 );
or ( n33981 , n33978 , n33980 );
buf ( n381589 , n604 );
not ( n33983 , n381589 );
buf ( n381591 , n376526 );
not ( n33985 , n381591 );
or ( n33986 , n33983 , n33985 );
buf ( n381594 , n376520 );
buf ( n381595 , n11145 );
nand ( n33989 , n381594 , n381595 );
buf ( n381597 , n33989 );
buf ( n381598 , n381597 );
nand ( n33992 , n33986 , n381598 );
buf ( n381600 , n33992 );
buf ( n381601 , n381600 );
buf ( n381602 , n355075 );
nand ( n33996 , n381601 , n381602 );
buf ( n381604 , n33996 );
buf ( n381605 , n381604 );
nand ( n33999 , n33981 , n381605 );
buf ( n381607 , n33999 );
buf ( n381608 , n381607 );
xor ( n34002 , n381583 , n381608 );
buf ( n381610 , n1397 );
not ( n34004 , n381610 );
buf ( n381612 , n594 );
not ( n34006 , n381612 );
buf ( n381614 , n25811 );
not ( n34008 , n381614 );
or ( n34009 , n34006 , n34008 );
buf ( n381617 , n25566 );
buf ( n381618 , n348975 );
nand ( n34012 , n381617 , n381618 );
buf ( n381620 , n34012 );
buf ( n381621 , n381620 );
nand ( n34015 , n34009 , n381621 );
buf ( n381623 , n34015 );
buf ( n381624 , n381623 );
not ( n34018 , n381624 );
or ( n34019 , n34004 , n34018 );
buf ( n381627 , n380596 );
buf ( n381628 , n349035 );
nand ( n34022 , n381627 , n381628 );
buf ( n381630 , n34022 );
buf ( n381631 , n381630 );
nand ( n34025 , n34019 , n381631 );
buf ( n381633 , n34025 );
buf ( n381634 , n381633 );
buf ( n381635 , n4443 );
not ( n34029 , n381635 );
and ( n34030 , n24943 , n347312 );
not ( n34031 , n24943 );
and ( n34032 , n34031 , n598 );
or ( n34033 , n34030 , n34032 );
buf ( n381641 , n34033 );
not ( n34035 , n381641 );
or ( n34036 , n34029 , n34035 );
buf ( n381644 , n380669 );
buf ( n381645 , n4362 );
nand ( n34039 , n381644 , n381645 );
buf ( n381647 , n34039 );
buf ( n381648 , n381647 );
nand ( n34042 , n34036 , n381648 );
buf ( n381650 , n34042 );
buf ( n381651 , n381650 );
xor ( n34045 , n381634 , n381651 );
buf ( n381653 , n351924 );
not ( n34047 , n381653 );
buf ( n381655 , n600 );
not ( n34049 , n381655 );
buf ( n381657 , n373494 );
not ( n34051 , n381657 );
or ( n34052 , n34049 , n34051 );
buf ( n381660 , n17009 );
buf ( n381661 , n6460 );
nand ( n34055 , n381660 , n381661 );
buf ( n381663 , n34055 );
buf ( n381664 , n381663 );
nand ( n34058 , n34052 , n381664 );
buf ( n381666 , n34058 );
buf ( n381667 , n381666 );
not ( n34061 , n381667 );
or ( n34062 , n34047 , n34061 );
buf ( n381670 , n33077 );
buf ( n381671 , n1722 );
nand ( n34065 , n381670 , n381671 );
buf ( n381673 , n34065 );
buf ( n381674 , n381673 );
nand ( n34068 , n34062 , n381674 );
buf ( n381676 , n34068 );
buf ( n381677 , n381676 );
and ( n34071 , n34045 , n381677 );
and ( n34072 , n381634 , n381651 );
or ( n34073 , n34071 , n34072 );
buf ( n381681 , n34073 );
buf ( n381682 , n381681 );
and ( n34076 , n34002 , n381682 );
and ( n34077 , n381583 , n381608 );
or ( n34078 , n34076 , n34077 );
buf ( n381686 , n34078 );
buf ( n381687 , n381686 );
xor ( n34081 , n381579 , n381687 );
xor ( n34082 , n380652 , n380677 );
xor ( n34083 , n34082 , n380695 );
buf ( n381691 , n34083 );
buf ( n381692 , n381691 );
buf ( n381693 , n27758 );
buf ( n381694 , n592 );
and ( n34088 , n381693 , n381694 );
buf ( n381696 , n34088 );
buf ( n381697 , n381696 );
buf ( n381698 , n375038 );
not ( n34092 , n381698 );
buf ( n381700 , n376599 );
not ( n34094 , n381700 );
or ( n34095 , n34092 , n34094 );
and ( n34096 , n9635 , n348910 );
not ( n34097 , n9635 );
and ( n34098 , n34097 , n592 );
or ( n34099 , n34096 , n34098 );
nand ( n34100 , n34099 , n348946 );
buf ( n381708 , n34100 );
nand ( n34102 , n34095 , n381708 );
buf ( n381710 , n34102 );
buf ( n381711 , n381710 );
xor ( n34105 , n381697 , n381711 );
not ( n34106 , n372772 );
not ( n34107 , n29017 );
or ( n34108 , n34106 , n34107 );
nand ( n34109 , n380751 , n347319 );
nand ( n34110 , n34108 , n34109 );
buf ( n381718 , n34110 );
and ( n34112 , n34105 , n381718 );
and ( n34113 , n381697 , n381711 );
or ( n34114 , n34112 , n34113 );
buf ( n381722 , n34114 );
buf ( n381723 , n381722 );
buf ( n381724 , n6600 );
not ( n34118 , n381724 );
buf ( n381726 , n381600 );
not ( n34120 , n381726 );
or ( n34121 , n34118 , n34120 );
and ( n34122 , n604 , n28093 );
not ( n34123 , n604 );
and ( n34124 , n34123 , n28092 );
or ( n34125 , n34122 , n34124 );
buf ( n381733 , n34125 );
buf ( n381734 , n355075 );
nand ( n34128 , n381733 , n381734 );
buf ( n381736 , n34128 );
buf ( n381737 , n381736 );
nand ( n34131 , n34121 , n381737 );
buf ( n381739 , n34131 );
buf ( n381740 , n381739 );
xor ( n34134 , n381723 , n381740 );
buf ( n381742 , n352149 );
not ( n34136 , n381742 );
buf ( n381744 , n33106 );
not ( n34138 , n381744 );
or ( n34139 , n34136 , n34138 );
buf ( n381747 , n27554 );
not ( n34141 , n381747 );
buf ( n381749 , n373465 );
not ( n34143 , n381749 );
and ( n34144 , n34141 , n34143 );
buf ( n381752 , n27554 );
buf ( n381753 , n358417 );
and ( n34147 , n381752 , n381753 );
nor ( n34148 , n34144 , n34147 );
buf ( n381756 , n34148 );
buf ( n381757 , n381756 );
nand ( n34151 , n34139 , n381757 );
buf ( n381759 , n34151 );
buf ( n381760 , n381759 );
and ( n34154 , n34134 , n381760 );
and ( n34155 , n381723 , n381740 );
or ( n34156 , n34154 , n34155 );
buf ( n381764 , n34156 );
buf ( n381765 , n381764 );
xor ( n34159 , n381692 , n381765 );
xor ( n34160 , n380732 , n380793 );
xor ( n34161 , n34160 , n380816 );
buf ( n381769 , n34161 );
buf ( n381770 , n381769 );
and ( n34164 , n34159 , n381770 );
and ( n34165 , n381692 , n381765 );
or ( n34166 , n34164 , n34165 );
buf ( n381774 , n34166 );
buf ( n381775 , n381774 );
and ( n34169 , n34081 , n381775 );
and ( n34170 , n381579 , n381687 );
or ( n34171 , n34169 , n34170 );
buf ( n381779 , n34171 );
buf ( n381780 , n381779 );
and ( n34174 , n33968 , n381780 );
and ( n34175 , n381570 , n381574 );
or ( n34176 , n34174 , n34175 );
buf ( n381784 , n34176 );
buf ( n381785 , n381784 );
nor ( n34179 , n381566 , n381785 );
buf ( n381787 , n34179 );
buf ( n381788 , n381787 );
xor ( n34182 , n381570 , n381574 );
xor ( n34183 , n34182 , n381780 );
buf ( n381791 , n34183 );
buf ( n381792 , n381791 );
xor ( n34186 , n380710 , n380821 );
xor ( n34187 , n34186 , n380826 );
buf ( n381795 , n34187 );
buf ( n381796 , n381795 );
xor ( n34190 , n381579 , n381687 );
xor ( n34191 , n34190 , n381775 );
buf ( n381799 , n34191 );
buf ( n381800 , n381799 );
xor ( n34194 , n381796 , n381800 );
xor ( n34195 , n380737 , n380762 );
xor ( n34196 , n34195 , n380788 );
buf ( n381804 , n34196 );
buf ( n381805 , n381804 );
buf ( n381806 , n357376 );
not ( n34200 , n381806 );
buf ( n381808 , n9642 );
buf ( n381809 , n379586 );
and ( n34203 , n381808 , n381809 );
not ( n34204 , n381808 );
buf ( n381812 , n16993 );
and ( n34206 , n34204 , n381812 );
nor ( n34207 , n34203 , n34206 );
buf ( n381815 , n34207 );
buf ( n381816 , n381815 );
not ( n34210 , n381816 );
or ( n34211 , n34200 , n34210 );
buf ( n381819 , n380806 );
buf ( n381820 , n607 );
nand ( n34214 , n381819 , n381820 );
buf ( n381822 , n34214 );
buf ( n381823 , n381822 );
nand ( n34217 , n34211 , n381823 );
buf ( n381825 , n34217 );
buf ( n381826 , n381825 );
xor ( n34220 , n381805 , n381826 );
buf ( n381828 , n349035 );
not ( n34222 , n381828 );
buf ( n381830 , n381623 );
not ( n34224 , n381830 );
or ( n34225 , n34222 , n34224 );
buf ( n381833 , n376415 );
buf ( n381834 , n1397 );
nand ( n34228 , n381833 , n381834 );
buf ( n381836 , n34228 );
buf ( n381837 , n381836 );
nand ( n34231 , n34225 , n381837 );
buf ( n381839 , n34231 );
buf ( n381840 , n381839 );
buf ( n381841 , n4362 );
not ( n34235 , n381841 );
buf ( n381843 , n34033 );
not ( n34237 , n381843 );
or ( n34238 , n34235 , n34237 );
nand ( n34239 , n28792 , n4443 );
buf ( n381847 , n34239 );
nand ( n34241 , n34238 , n381847 );
buf ( n381849 , n34241 );
buf ( n381850 , n381849 );
xor ( n34244 , n381840 , n381850 );
buf ( n381852 , n1722 );
not ( n34246 , n381852 );
buf ( n381854 , n381666 );
not ( n34248 , n381854 );
or ( n34249 , n34246 , n34248 );
buf ( n381857 , n376446 );
buf ( n381858 , n351924 );
nand ( n34252 , n381857 , n381858 );
buf ( n381860 , n34252 );
buf ( n381861 , n381860 );
nand ( n34255 , n34249 , n381861 );
buf ( n381863 , n34255 );
buf ( n381864 , n381863 );
and ( n34258 , n34244 , n381864 );
and ( n34259 , n381840 , n381850 );
or ( n34260 , n34258 , n34259 );
buf ( n381868 , n34260 );
buf ( n381869 , n381868 );
and ( n34263 , n34220 , n381869 );
and ( n34264 , n381805 , n381826 );
or ( n34265 , n34263 , n34264 );
buf ( n381873 , n34265 );
buf ( n381874 , n381873 );
xor ( n34268 , n381583 , n381608 );
xor ( n34269 , n34268 , n381682 );
buf ( n381877 , n34269 );
buf ( n381878 , n381877 );
xor ( n34272 , n381874 , n381878 );
xor ( n34273 , n381634 , n381651 );
xor ( n34274 , n34273 , n381677 );
buf ( n381882 , n34274 );
buf ( n381883 , n381882 );
buf ( n381884 , n354113 );
not ( n34278 , n381884 );
buf ( n381886 , n27137 );
buf ( n381887 , n602 );
and ( n34281 , n381886 , n381887 );
not ( n34282 , n381886 );
buf ( n381890 , n349406 );
and ( n34284 , n34282 , n381890 );
nor ( n34285 , n34281 , n34284 );
buf ( n381893 , n34285 );
buf ( n381894 , n381893 );
not ( n34288 , n381894 );
or ( n34289 , n34278 , n34288 );
buf ( n381897 , n27554 );
buf ( n381898 , n373187 );
and ( n34292 , n381897 , n381898 );
buf ( n381900 , n375161 );
buf ( n381901 , n373176 );
and ( n34295 , n381900 , n381901 );
nor ( n34296 , n34292 , n34295 );
buf ( n381904 , n34296 );
buf ( n381905 , n381904 );
nand ( n34299 , n34289 , n381905 );
buf ( n381907 , n34299 );
buf ( n381908 , n381907 );
xor ( n34302 , n381697 , n381711 );
xor ( n34303 , n34302 , n381718 );
buf ( n381911 , n34303 );
buf ( n381912 , n381911 );
xor ( n34306 , n381908 , n381912 );
buf ( n381914 , n355075 );
not ( n34308 , n381914 );
buf ( n381916 , n28965 );
not ( n34310 , n381916 );
or ( n34311 , n34308 , n34310 );
buf ( n381919 , n34125 );
buf ( n381920 , n6600 );
nand ( n34314 , n381919 , n381920 );
buf ( n381922 , n34314 );
buf ( n381923 , n381922 );
nand ( n34317 , n34311 , n381923 );
buf ( n381925 , n34317 );
buf ( n381926 , n381925 );
and ( n34320 , n34306 , n381926 );
and ( n34321 , n381908 , n381912 );
or ( n34322 , n34320 , n34321 );
buf ( n381930 , n34322 );
buf ( n381931 , n381930 );
xor ( n34325 , n381883 , n381931 );
xor ( n34326 , n381723 , n381740 );
xor ( n34327 , n34326 , n381760 );
buf ( n381935 , n34327 );
buf ( n381936 , n381935 );
and ( n34330 , n34325 , n381936 );
and ( n34331 , n381883 , n381931 );
or ( n381939 , n34330 , n34331 );
buf ( n381940 , n381939 );
buf ( n381941 , n381940 );
and ( n34335 , n34272 , n381941 );
and ( n34336 , n381874 , n381878 );
or ( n34337 , n34335 , n34336 );
buf ( n381945 , n34337 );
buf ( n381946 , n381945 );
and ( n34340 , n34194 , n381946 );
and ( n34341 , n381796 , n381800 );
or ( n34342 , n34340 , n34341 );
buf ( n381950 , n34342 );
buf ( n381951 , n381950 );
nor ( n34345 , n381792 , n381951 );
buf ( n381953 , n34345 );
buf ( n381954 , n381953 );
nor ( n34348 , n381788 , n381954 );
buf ( n381956 , n34348 );
not ( n34350 , n381956 );
xor ( n34351 , n381796 , n381800 );
xor ( n34352 , n34351 , n381946 );
buf ( n381960 , n34352 );
buf ( n381961 , n381960 );
xor ( n34355 , n381692 , n381765 );
xor ( n34356 , n34355 , n381770 );
buf ( n381964 , n34356 );
buf ( n381965 , n381964 );
xor ( n34359 , n381874 , n381878 );
xor ( n34360 , n34359 , n381941 );
buf ( n381968 , n34360 );
buf ( n381969 , n381968 );
xor ( n34363 , n381965 , n381969 );
xor ( n34364 , n376585 , n376610 );
and ( n34365 , n34364 , n376629 );
and ( n34366 , n376585 , n376610 );
or ( n34367 , n34365 , n34366 );
buf ( n381975 , n34367 );
buf ( n381976 , n381975 );
xor ( n34370 , n376401 , n376428 );
and ( n34371 , n34370 , n376454 );
and ( n34372 , n376401 , n376428 );
or ( n34373 , n34371 , n34372 );
buf ( n381981 , n34373 );
buf ( n381982 , n381981 );
xor ( n34376 , n381976 , n381982 );
buf ( n381984 , n607 );
not ( n34378 , n381984 );
buf ( n381986 , n381815 );
not ( n34380 , n381986 );
or ( n34381 , n34378 , n34380 );
buf ( n381989 , n379799 );
not ( n34383 , n381989 );
buf ( n381991 , n357376 );
nand ( n34385 , n34383 , n381991 );
buf ( n381993 , n34385 );
buf ( n381994 , n381993 );
nand ( n34388 , n34381 , n381994 );
buf ( n381996 , n34388 );
buf ( n381997 , n381996 );
and ( n34391 , n34376 , n381997 );
and ( n34392 , n381976 , n381982 );
or ( n34393 , n34391 , n34392 );
buf ( n382001 , n34393 );
buf ( n382002 , n382001 );
xor ( n34396 , n381805 , n381826 );
xor ( n34397 , n34396 , n381869 );
buf ( n382005 , n34397 );
buf ( n382006 , n382005 );
xor ( n34400 , n382002 , n382006 );
xor ( n34401 , n381840 , n381850 );
xor ( n34402 , n34401 , n381864 );
buf ( n382010 , n34402 );
buf ( n382011 , n382010 );
xor ( n34405 , n376489 , n376495 );
and ( n34406 , n34405 , n376541 );
and ( n34407 , n376489 , n376495 );
or ( n34408 , n34406 , n34407 );
buf ( n382016 , n34408 );
buf ( n382017 , n382016 );
xor ( n34411 , n382011 , n382017 );
xor ( n34412 , n381908 , n381912 );
xor ( n34413 , n34412 , n381926 );
buf ( n382021 , n34413 );
buf ( n382022 , n382021 );
and ( n34416 , n34411 , n382022 );
and ( n34417 , n382011 , n382017 );
or ( n34418 , n34416 , n34417 );
buf ( n382026 , n34418 );
buf ( n382027 , n382026 );
and ( n34421 , n34400 , n382027 );
and ( n34422 , n382002 , n382006 );
or ( n34423 , n34421 , n34422 );
buf ( n382031 , n34423 );
buf ( n382032 , n382031 );
and ( n34426 , n34363 , n382032 );
and ( n34427 , n381965 , n381969 );
or ( n34428 , n34426 , n34427 );
buf ( n382036 , n34428 );
buf ( n382037 , n382036 );
nand ( n34431 , n381961 , n382037 );
buf ( n382039 , n34431 );
buf ( n382040 , n382039 );
xor ( n34434 , n381965 , n381969 );
xor ( n34435 , n34434 , n382032 );
buf ( n382043 , n34435 );
buf ( n382044 , n382043 );
xor ( n34438 , n381883 , n381931 );
xor ( n34439 , n34438 , n381936 );
buf ( n382047 , n34439 );
buf ( n382048 , n382047 );
xor ( n34442 , n376580 , n376632 );
and ( n34443 , n34442 , n376639 );
and ( n34444 , n376580 , n376632 );
or ( n34445 , n34443 , n34444 );
buf ( n382053 , n34445 );
buf ( n382054 , n382053 );
xor ( n34448 , n381976 , n381982 );
xor ( n34449 , n34448 , n381997 );
buf ( n382057 , n34449 );
buf ( n382058 , n382057 );
xor ( n34452 , n382054 , n382058 );
xor ( n34453 , n376457 , n376463 );
and ( n34454 , n34453 , n376544 );
and ( n34455 , n376457 , n376463 );
or ( n34456 , n34454 , n34455 );
buf ( n382064 , n34456 );
buf ( n382065 , n382064 );
and ( n34459 , n34452 , n382065 );
and ( n34460 , n382054 , n382058 );
or ( n34461 , n34459 , n34460 );
buf ( n382069 , n34461 );
buf ( n382070 , n382069 );
xor ( n34464 , n382048 , n382070 );
xor ( n34465 , n382002 , n382006 );
xor ( n34466 , n34465 , n382027 );
buf ( n382074 , n34466 );
buf ( n382075 , n382074 );
and ( n34469 , n34464 , n382075 );
and ( n34470 , n382048 , n382070 );
or ( n34471 , n34469 , n34470 );
buf ( n382079 , n34471 );
buf ( n382080 , n382079 );
nand ( n34474 , n382044 , n382080 );
buf ( n382082 , n34474 );
buf ( n382083 , n382082 );
and ( n34477 , n382040 , n382083 );
buf ( n382085 , n381960 );
buf ( n382086 , n382036 );
nor ( n34480 , n382085 , n382086 );
buf ( n382088 , n34480 );
buf ( n382089 , n382088 );
nor ( n34483 , n34477 , n382089 );
buf ( n382091 , n34483 );
not ( n34485 , n382091 );
or ( n34486 , n34350 , n34485 );
buf ( n382094 , n381565 );
buf ( n382095 , n381784 );
nor ( n34489 , n382094 , n382095 );
buf ( n382097 , n34489 );
buf ( n382098 , n382097 );
not ( n34492 , n382098 );
nand ( n34493 , n381950 , n381791 );
buf ( n382101 , n34493 );
not ( n34495 , n382101 );
and ( n34496 , n34492 , n34495 );
buf ( n382104 , n381565 );
buf ( n382105 , n381784 );
and ( n34499 , n382104 , n382105 );
buf ( n382107 , n34499 );
buf ( n382108 , n382107 );
nor ( n34502 , n34496 , n382108 );
buf ( n382110 , n34502 );
nand ( n34504 , n34486 , n382110 );
not ( n34505 , n34504 );
nor ( n34506 , n382036 , n381960 );
buf ( n382114 , n382043 );
buf ( n382115 , n382079 );
nor ( n34509 , n382114 , n382115 );
buf ( n382117 , n34509 );
nor ( n34511 , n34506 , n382117 );
and ( n34512 , n381956 , n34511 );
xor ( n34513 , n382011 , n382017 );
xor ( n34514 , n34513 , n382022 );
buf ( n382122 , n34514 );
buf ( n382123 , n382122 );
xor ( n34517 , n382054 , n382058 );
xor ( n34518 , n34517 , n382065 );
buf ( n382126 , n34518 );
buf ( n382127 , n382126 );
xor ( n34521 , n382123 , n382127 );
xor ( n34522 , n376560 , n376642 );
and ( n34523 , n34522 , n376649 );
and ( n34524 , n376560 , n376642 );
or ( n34525 , n34523 , n34524 );
buf ( n382133 , n34525 );
buf ( n382134 , n382133 );
xor ( n34528 , n34521 , n382134 );
buf ( n382136 , n34528 );
buf ( n382137 , n382136 );
not ( n34531 , n382137 );
buf ( n382139 , n34531 );
buf ( n382140 , n382139 );
xor ( n34534 , n376547 , n376553 );
and ( n34535 , n34534 , n376652 );
and ( n34536 , n376547 , n376553 );
or ( n34537 , n34535 , n34536 );
buf ( n382145 , n34537 );
buf ( n382146 , n382145 );
not ( n34540 , n382146 );
buf ( n382148 , n34540 );
buf ( n382149 , n382148 );
nand ( n34543 , n382140 , n382149 );
buf ( n382151 , n34543 );
xor ( n34545 , n382048 , n382070 );
xor ( n34546 , n34545 , n382075 );
buf ( n382154 , n34546 );
buf ( n382155 , n382154 );
not ( n34549 , n382155 );
xor ( n34550 , n382123 , n382127 );
and ( n34551 , n34550 , n382134 );
and ( n34552 , n382123 , n382127 );
or ( n34553 , n34551 , n34552 );
buf ( n382161 , n34553 );
buf ( n382162 , n382161 );
not ( n34556 , n382162 );
buf ( n382164 , n34556 );
buf ( n382165 , n382164 );
nand ( n34559 , n34549 , n382165 );
buf ( n382167 , n34559 );
nand ( n34561 , n382151 , n382167 );
not ( n34562 , n34561 );
not ( n34563 , n375474 );
not ( n34564 , n375479 );
or ( n34565 , n34563 , n34564 );
buf ( n382173 , n375736 );
buf ( n382174 , n375742 );
nand ( n34568 , n382173 , n382174 );
buf ( n382176 , n34568 );
nand ( n34570 , n34565 , n382176 );
not ( n34571 , n34570 );
buf ( n382179 , n376654 );
buf ( n382180 , n376661 );
nor ( n34574 , n382179 , n382180 );
buf ( n382182 , n34574 );
buf ( n382183 , n382182 );
buf ( n382184 , n375745 );
nor ( n34578 , n382183 , n382184 );
buf ( n382186 , n34578 );
not ( n34580 , n382186 );
or ( n34581 , n34571 , n34580 );
buf ( n382189 , n382136 );
buf ( n382190 , n382145 );
nand ( n34584 , n382189 , n382190 );
buf ( n382192 , n34584 );
buf ( n382193 , n382192 );
buf ( n382194 , n376654 );
buf ( n382195 , n376661 );
nand ( n34589 , n382194 , n382195 );
buf ( n382197 , n34589 );
buf ( n382198 , n382197 );
and ( n34592 , n382193 , n382198 );
buf ( n382200 , n34592 );
nand ( n34594 , n34581 , n382200 );
nand ( n34595 , n34562 , n34594 );
not ( n34596 , n34561 );
and ( n34597 , n376372 , n376667 );
nand ( n34598 , n34596 , n27903 , n34597 );
buf ( n34599 , n382161 );
buf ( n382207 , n382154 );
buf ( n34601 , n382207 );
buf ( n382209 , n34601 );
nand ( n34603 , n34599 , n382209 );
nand ( n34604 , n34595 , n34598 , n34603 );
nand ( n34605 , n34512 , n34604 );
nand ( n34606 , n34505 , n34605 );
nand ( n34607 , n33955 , n34606 );
not ( n34608 , n34607 );
buf ( n382216 , n380319 );
buf ( n382217 , n380546 );
nand ( n34611 , n382216 , n382217 );
buf ( n382219 , n34611 );
not ( n34613 , n382219 );
buf ( n382221 , n380840 );
buf ( n382222 , n380844 );
nand ( n34616 , n382221 , n382222 );
buf ( n382224 , n34616 );
not ( n34618 , n382224 );
or ( n34619 , n34613 , n34618 );
not ( n34620 , n380319 );
buf ( n382228 , n380546 );
not ( n34622 , n382228 );
buf ( n382230 , n34622 );
nand ( n34624 , n34620 , n382230 );
nand ( n34625 , n34619 , n34624 );
not ( n34626 , n34625 );
nand ( n34627 , n381152 , n381157 );
nand ( n34628 , n381005 , n381011 );
and ( n34629 , n34627 , n34628 );
not ( n34630 , n34629 );
or ( n34631 , n34626 , n34630 );
not ( n34632 , n381005 );
nand ( n34633 , n34632 , n33405 );
not ( n34634 , n381152 );
not ( n34635 , n381157 );
nand ( n34636 , n34634 , n34635 );
nand ( n34637 , n34633 , n34636 );
nand ( n34638 , n34627 , n34637 );
nand ( n34639 , n34631 , n34638 );
not ( n34640 , n34639 );
buf ( n382248 , n381561 );
not ( n34642 , n382248 );
buf ( n382250 , n34642 );
and ( n34644 , n34640 , n382250 );
or ( n34645 , n381330 , n381448 );
nand ( n34646 , n381455 , n381511 );
nor ( n34647 , n381538 , n381518 );
or ( n34648 , n34646 , n34647 );
nand ( n34649 , n381538 , n381518 );
nand ( n34650 , n34648 , n34649 );
nand ( n34651 , n34645 , n34650 , n33947 );
nand ( n34652 , n381553 , n381550 );
not ( n34653 , n34652 );
nand ( n34654 , n34645 , n34653 );
nand ( n34655 , n381330 , n381448 );
nand ( n34656 , n34651 , n34654 , n34655 );
nor ( n34657 , n34644 , n34656 );
buf ( n382265 , n34657 );
not ( n34659 , n382265 );
buf ( n382267 , n375038 );
not ( n34661 , n382267 );
buf ( n382269 , n592 );
buf ( n382270 , n381252 );
xor ( n34664 , n382269 , n382270 );
buf ( n382272 , n34664 );
buf ( n382273 , n382272 );
not ( n34667 , n382273 );
or ( n34668 , n34661 , n34667 );
buf ( n382276 , n592 );
not ( n34670 , n382276 );
buf ( n382278 , n379607 );
not ( n34672 , n382278 );
or ( n34673 , n34670 , n34672 );
buf ( n382281 , n379604 );
buf ( n382282 , n348910 );
nand ( n34676 , n382281 , n382282 );
buf ( n382284 , n34676 );
buf ( n382285 , n382284 );
nand ( n34679 , n34673 , n382285 );
buf ( n382287 , n34679 );
buf ( n382288 , n382287 );
buf ( n382289 , n348946 );
nand ( n34683 , n382288 , n382289 );
buf ( n382291 , n34683 );
buf ( n382292 , n382291 );
nand ( n34686 , n34668 , n382292 );
buf ( n382294 , n34686 );
buf ( n382295 , n382294 );
buf ( n382296 , n381024 );
buf ( n382297 , n592 );
nand ( n34691 , n382296 , n382297 );
buf ( n382299 , n34691 );
buf ( n382300 , n382299 );
xor ( n34694 , n382295 , n382300 );
buf ( n382302 , n1335 );
not ( n34696 , n382302 );
buf ( n382304 , n1396 );
not ( n34698 , n382304 );
or ( n34699 , n34696 , n34698 );
buf ( n382307 , n381274 );
nand ( n34701 , n34699 , n382307 );
buf ( n382309 , n34701 );
buf ( n382310 , n382309 );
and ( n34704 , n381194 , n381195 );
buf ( n382312 , n34704 );
buf ( n382313 , n382312 );
xor ( n34707 , n382310 , n382313 );
buf ( n382315 , n348946 );
not ( n34709 , n382315 );
buf ( n382317 , n382272 );
not ( n34711 , n382317 );
or ( n34712 , n34709 , n34711 );
buf ( n382320 , n33624 );
buf ( n382321 , n375038 );
nand ( n34715 , n382320 , n382321 );
buf ( n382323 , n34715 );
buf ( n382324 , n382323 );
nand ( n34718 , n34712 , n382324 );
buf ( n382326 , n34718 );
buf ( n382327 , n382326 );
and ( n34721 , n34707 , n382327 );
and ( n34722 , n382310 , n382313 );
or ( n34723 , n34721 , n34722 );
buf ( n382331 , n34723 );
buf ( n382332 , n382331 );
and ( n34726 , n34694 , n382332 );
and ( n34727 , n382295 , n382300 );
or ( n34728 , n34726 , n34727 );
buf ( n382336 , n34728 );
buf ( n382337 , n349013 );
not ( n34731 , n382337 );
buf ( n382339 , n375038 );
not ( n34733 , n382339 );
buf ( n382341 , n34733 );
buf ( n382342 , n382341 );
not ( n34736 , n382342 );
or ( n34737 , n34731 , n34736 );
buf ( n382345 , n382287 );
nand ( n34739 , n34737 , n382345 );
buf ( n382347 , n34739 );
buf ( n382348 , n382347 );
and ( n34742 , n382269 , n382270 );
buf ( n382350 , n34742 );
buf ( n382351 , n382350 );
xor ( n34745 , n382348 , n382351 );
buf ( n382353 , n382299 );
not ( n34747 , n382353 );
buf ( n382355 , n34747 );
buf ( n382356 , n382355 );
xor ( n34750 , n34745 , n382356 );
buf ( n382358 , n34750 );
or ( n34752 , n382336 , n382358 );
not ( n34753 , n34752 );
buf ( n382361 , n34753 );
xor ( n34755 , n382348 , n382351 );
and ( n34756 , n34755 , n382356 );
and ( n34757 , n382348 , n382351 );
or ( n34758 , n34756 , n34757 );
buf ( n382366 , n34758 );
buf ( n382367 , n379604 );
buf ( n382368 , n592 );
nand ( n34763 , n382367 , n382368 );
buf ( n382370 , n34763 );
buf ( n382371 , C0 );
buf ( n382372 , n382371 );
nor ( n34769 , n382361 , n382372 );
buf ( n382374 , n34769 );
buf ( n382375 , n382374 );
not ( n34772 , n382375 );
buf ( n382377 , n381287 );
not ( n34774 , n382377 );
buf ( n382379 , n34774 );
buf ( n382380 , n382379 );
xor ( n34777 , n382310 , n382313 );
xor ( n34778 , n34777 , n382327 );
buf ( n382383 , n34778 );
buf ( n382384 , n382383 );
xor ( n34781 , n382380 , n382384 );
xor ( n34782 , n381242 , n381282 );
and ( n34783 , n34782 , n381288 );
and ( n34784 , n381242 , n381282 );
or ( n34785 , n34783 , n34784 );
buf ( n382390 , n34785 );
buf ( n382391 , n382390 );
xor ( n34788 , n34781 , n382391 );
buf ( n382393 , n34788 );
xor ( n34790 , n381225 , n381291 );
and ( n34791 , n34790 , n381328 );
and ( n34792 , n381225 , n381291 );
or ( n34793 , n34791 , n34792 );
buf ( n382398 , n34793 );
nand ( n34795 , n382393 , n382398 );
buf ( n382400 , n34795 );
xor ( n34797 , n382380 , n382384 );
and ( n34798 , n34797 , n382391 );
and ( n34799 , n382380 , n382384 );
or ( n34800 , n34798 , n34799 );
buf ( n382405 , n34800 );
buf ( n382406 , n382405 );
xor ( n34803 , n382295 , n382300 );
xor ( n34804 , n34803 , n382332 );
buf ( n382409 , n34804 );
buf ( n382410 , n382409 );
nor ( n34807 , n382406 , n382410 );
buf ( n382412 , n34807 );
buf ( n382413 , n382412 );
or ( n34810 , n382400 , n382413 );
buf ( n382415 , n382405 );
buf ( n382416 , n382409 );
nand ( n34813 , n382415 , n382416 );
buf ( n382418 , n34813 );
buf ( n382419 , n382418 );
nand ( n34816 , n34810 , n382419 );
buf ( n382421 , n34816 );
buf ( n382422 , n382421 );
not ( n34819 , n382422 );
or ( n34820 , n34772 , n34819 );
nand ( n34821 , n382336 , n382358 );
buf ( n382426 , n34821 );
buf ( n382427 , n382371 );
nor ( n34824 , n382426 , n382427 );
buf ( n382429 , n34824 );
buf ( n382430 , n382429 );
buf ( n382431 , n382366 );
buf ( n382432 , n382370 );
and ( n34829 , n382431 , n382432 );
buf ( n382434 , n34829 );
buf ( n382435 , n382434 );
nor ( n34832 , n382430 , n382435 );
buf ( n382437 , n34832 );
buf ( n382438 , n382437 );
nand ( n34835 , n34820 , n382438 );
buf ( n382440 , n34835 );
buf ( n382441 , n382440 );
nor ( n34838 , n34659 , n382441 );
buf ( n382443 , n34838 );
not ( n34840 , n382443 );
or ( n34841 , n34608 , n34840 );
buf ( n382446 , n382374 );
not ( n34843 , n382446 );
nor ( n34844 , n382398 , n382393 );
buf ( n382449 , n34844 );
buf ( n382450 , n382412 );
nor ( n34847 , n382449 , n382450 );
buf ( n382452 , n34847 );
buf ( n382453 , n382452 );
not ( n34850 , n382453 );
or ( n34851 , n34843 , n34850 );
buf ( n382456 , n382440 );
not ( n34853 , n382456 );
buf ( n382458 , n34853 );
buf ( n382459 , n382458 );
nand ( n34856 , n34851 , n382459 );
buf ( n382461 , n34856 );
nand ( n34858 , n34841 , n382461 );
not ( n34859 , n34858 );
not ( n34860 , n34859 );
not ( n34861 , n34860 );
not ( n34862 , n34861 );
not ( n34863 , n34862 );
buf ( n382468 , n34863 );
not ( n34865 , n382468 );
or ( n34866 , n31972 , n34865 );
buf ( n382471 , n34863 );
not ( n34868 , n382471 );
buf ( n382473 , n34868 );
buf ( n382474 , n382473 );
buf ( n382475 , n379574 );
nand ( n34872 , n382474 , n382475 );
buf ( n382477 , n34872 );
buf ( n382478 , n382477 );
nand ( n34875 , n34866 , n382478 );
buf ( n382480 , n34875 );
buf ( n382481 , n382480 );
not ( n34878 , n382481 );
or ( n34879 , n31861 , n34878 );
buf ( n382484 , n379577 );
not ( n34881 , n382484 );
not ( n34882 , n382452 );
not ( n34883 , n34656 );
or ( n34884 , n34882 , n34883 );
buf ( n382489 , n382421 );
not ( n34886 , n382489 );
buf ( n382491 , n34886 );
nand ( n34888 , n34884 , n382491 );
and ( n34889 , n34888 , n34752 );
not ( n34890 , n34821 );
nor ( n34891 , n34889 , n34890 );
nand ( n34892 , n33553 , n34512 , n34604 );
not ( n34893 , n34892 );
buf ( n382498 , n33951 );
buf ( n382499 , n382452 );
nand ( n34896 , n382498 , n382499 );
buf ( n382501 , n34896 );
nor ( n34898 , n34753 , n382501 );
nand ( n34899 , n34893 , n34898 );
not ( n34900 , n33241 );
not ( n34901 , n33551 );
nand ( n34902 , n34901 , n33406 );
nor ( n34903 , n34900 , n34902 );
not ( n34904 , n34903 );
not ( n34905 , n34504 );
or ( n34906 , n34904 , n34905 );
not ( n34907 , n34629 );
not ( n34908 , n34625 );
or ( n34909 , n34907 , n34908 );
nand ( n34910 , n34627 , n34637 );
nand ( n34911 , n34909 , n34910 );
nand ( n34912 , n34906 , n34911 );
nand ( n34913 , n34912 , n34898 );
nand ( n34914 , n34891 , n34899 , n34913 );
buf ( n382519 , n382371 );
buf ( n382520 , n382434 );
nor ( n34917 , n382519 , n382520 );
buf ( n382522 , n34917 );
xor ( n34919 , n34914 , n382522 );
buf ( n382524 , n34919 );
not ( n34921 , n382524 );
buf ( n382526 , n34921 );
buf ( n382527 , n382526 );
buf ( n34924 , n382527 );
buf ( n382529 , n34924 );
buf ( n382530 , n382529 );
not ( n34927 , n382530 );
buf ( n382532 , n34927 );
buf ( n382533 , n382532 );
not ( n34930 , n382533 );
buf ( n382535 , n34930 );
buf ( n382536 , n382535 );
buf ( n34933 , n382536 );
buf ( n382538 , n34933 );
buf ( n382539 , n382538 );
not ( n34936 , n382539 );
or ( n34937 , n34881 , n34936 );
buf ( n382542 , n379574 );
buf ( n382543 , n382526 );
not ( n34940 , n382543 );
buf ( n382545 , n34940 );
buf ( n382546 , n382545 );
not ( n34943 , n382546 );
buf ( n382548 , n34943 );
buf ( n382549 , n382548 );
not ( n34946 , n382549 );
buf ( n382551 , n34946 );
buf ( n382552 , n382551 );
nand ( n34949 , n382542 , n382552 );
buf ( n382554 , n34949 );
buf ( n382555 , n382554 );
nand ( n34952 , n34937 , n382555 );
buf ( n382557 , n34952 );
buf ( n382558 , n382557 );
buf ( n382559 , n31850 );
buf ( n382560 , n379531 );
not ( n34957 , n382560 );
buf ( n382562 , n379561 );
not ( n34959 , n382562 );
or ( n34960 , n34957 , n34959 );
buf ( n382565 , n379567 );
nand ( n34962 , n34960 , n382565 );
buf ( n382567 , n34962 );
buf ( n382568 , n382567 );
not ( n34965 , n382568 );
buf ( n382570 , n34965 );
buf ( n382571 , n382570 );
not ( n34968 , n382571 );
buf ( n382573 , n31830 );
not ( n34970 , n382573 );
or ( n34971 , n34968 , n34970 );
and ( n34972 , n31733 , n31825 );
not ( n34973 , n31733 );
and ( n34974 , n34973 , n31828 );
or ( n34975 , n34972 , n34974 );
buf ( n382580 , n34975 );
buf ( n382581 , n382567 );
nand ( n34978 , n382580 , n382581 );
buf ( n382583 , n34978 );
buf ( n382584 , n382583 );
nand ( n34981 , n34971 , n382584 );
buf ( n382586 , n34981 );
buf ( n382587 , n382586 );
nand ( n34984 , n382559 , n382587 );
buf ( n382589 , n34984 );
buf ( n382590 , n382589 );
buf ( n34987 , n382590 );
buf ( n382592 , n34987 );
buf ( n382593 , n382592 );
not ( n34990 , n382593 );
buf ( n382595 , n34990 );
buf ( n382596 , n382595 );
buf ( n34993 , n382596 );
buf ( n382598 , n34993 );
buf ( n382599 , n382598 );
buf ( n34996 , n382599 );
buf ( n382601 , n34996 );
buf ( n382602 , n382601 );
not ( n34999 , n382602 );
buf ( n382604 , n34999 );
buf ( n382605 , n382604 );
not ( n35002 , n382605 );
buf ( n382607 , n35002 );
buf ( n382608 , n382607 );
nand ( n35005 , n382558 , n382608 );
buf ( n382610 , n35005 );
buf ( n382611 , n382610 );
nand ( n35008 , n34879 , n382611 );
buf ( n382613 , n35008 );
buf ( n382614 , n382613 );
not ( n35011 , n382614 );
buf ( n382616 , n378848 );
not ( n35013 , n382616 );
buf ( n382618 , n379539 );
xor ( n35015 , n379472 , n379508 );
and ( n35016 , n35015 , n379515 );
and ( n35017 , n379472 , n379508 );
or ( n35018 , n35016 , n35017 );
buf ( n382623 , n35018 );
buf ( n382624 , n382623 );
buf ( n382625 , n377023 );
not ( n35022 , n382625 );
buf ( n382627 , n379494 );
not ( n35024 , n382627 );
or ( n35025 , n35022 , n35024 );
buf ( n382630 , n576 );
not ( n35027 , n382630 );
buf ( n382632 , n364664 );
not ( n35029 , n382632 );
or ( n35030 , n35027 , n35029 );
buf ( n382635 , n364661 );
buf ( n382636 , n354303 );
nand ( n35033 , n382635 , n382636 );
buf ( n382638 , n35033 );
buf ( n382639 , n382638 );
nand ( n35036 , n35030 , n382639 );
buf ( n382641 , n35036 );
buf ( n382642 , n382641 );
buf ( n382643 , n364834 );
nand ( n35040 , n382642 , n382643 );
buf ( n382645 , n35040 );
buf ( n382646 , n382645 );
nand ( n35043 , n35025 , n382646 );
buf ( n382648 , n35043 );
buf ( n382649 , n382648 );
buf ( n382650 , n377056 );
buf ( n382651 , n576 );
nand ( n382652 , n382650 , n382651 );
buf ( n382653 , n382652 );
buf ( n382654 , n382653 );
xor ( n35051 , n382649 , n382654 );
xor ( n35052 , n379484 , n379487 );
and ( n35053 , n35052 , n379505 );
and ( n35054 , n379484 , n379487 );
or ( n35055 , n35053 , n35054 );
buf ( n382660 , n35055 );
buf ( n382661 , n382660 );
xor ( n35058 , n35051 , n382661 );
buf ( n382663 , n35058 );
buf ( n382664 , n382663 );
or ( n35061 , n382624 , n382664 );
buf ( n382666 , n35061 );
nand ( n35063 , n382666 , n31916 );
buf ( n382668 , n35063 );
xor ( n35065 , n382649 , n382654 );
and ( n35066 , n35065 , n382661 );
and ( n35067 , n382649 , n382654 );
or ( n35068 , n35066 , n35067 );
buf ( n382673 , n35068 );
buf ( n382674 , n382673 );
buf ( n382675 , n377988 );
not ( n35072 , n382675 );
buf ( n382677 , n377023 );
not ( n35074 , n382677 );
buf ( n382679 , n35074 );
buf ( n382680 , n382679 );
not ( n35077 , n382680 );
or ( n35078 , n35072 , n35077 );
buf ( n382683 , n382641 );
nand ( n35080 , n35078 , n382683 );
buf ( n382685 , n35080 );
buf ( n382686 , n382685 );
and ( n35083 , n379491 , n379492 );
buf ( n382688 , n35083 );
buf ( n382689 , n382688 );
xor ( n35086 , n382686 , n382689 );
buf ( n382691 , n382653 );
not ( n35088 , n382691 );
buf ( n382693 , n35088 );
buf ( n382694 , n382693 );
xor ( n35091 , n35086 , n382694 );
buf ( n382696 , n35091 );
buf ( n382697 , n382696 );
nor ( n35094 , n382674 , n382697 );
buf ( n382699 , n35094 );
buf ( n382700 , n382699 );
nor ( n35097 , n382668 , n382700 );
buf ( n382702 , n35097 );
buf ( n382703 , n382702 );
nand ( n35100 , n382618 , n382703 );
buf ( n382705 , n35100 );
buf ( n382706 , n382705 );
nor ( n35103 , n35013 , n382706 );
buf ( n382708 , n35103 );
not ( n35105 , n382708 );
not ( n35106 , n31595 );
not ( n35107 , n35106 );
buf ( n382712 , n31612 );
not ( n35109 , n382712 );
buf ( n382714 , n371128 );
not ( n35111 , n382714 );
or ( n35112 , n35109 , n35111 );
buf ( n382717 , n379234 );
nand ( n35114 , n35112 , n382717 );
buf ( n382719 , n35114 );
not ( n35116 , n382719 );
or ( n35117 , n35107 , n35116 );
not ( n35118 , n31570 );
not ( n35119 , n31581 );
nor ( n35120 , n35118 , n35119 );
nand ( n35121 , n35117 , n35120 );
not ( n35122 , n35121 );
or ( n35123 , n35105 , n35122 );
not ( n35124 , n382705 );
nand ( n35125 , n35124 , n31690 );
nand ( n35126 , n35123 , n35125 );
not ( n35127 , n35126 );
not ( n35128 , n35127 );
buf ( n382733 , n382699 );
not ( n35130 , n382733 );
buf ( n382735 , n35130 );
buf ( n382736 , n382735 );
not ( n35133 , n382736 );
buf ( n382738 , n379552 );
buf ( n382739 , n35063 );
or ( n35136 , n382738 , n382739 );
buf ( n382741 , n382666 );
not ( n35138 , n382741 );
buf ( n382743 , n35138 );
buf ( n382744 , n382743 );
buf ( n382745 , n379527 );
or ( n35142 , n382744 , n382745 );
buf ( n382747 , n382623 );
buf ( n382748 , n382663 );
nand ( n35145 , n382747 , n382748 );
buf ( n382750 , n35145 );
buf ( n382751 , n382750 );
nand ( n35148 , n35142 , n382751 );
buf ( n382753 , n35148 );
buf ( n382754 , n382753 );
not ( n35151 , n382754 );
buf ( n382756 , n35151 );
buf ( n382757 , n382756 );
nand ( n35154 , n35136 , n382757 );
buf ( n382759 , n35154 );
buf ( n382760 , n382759 );
not ( n35157 , n382760 );
or ( n35158 , n35133 , n35157 );
buf ( n382763 , n382673 );
buf ( n382764 , n382696 );
nand ( n35161 , n382763 , n382764 );
buf ( n382766 , n35161 );
buf ( n382767 , n382766 );
nand ( n35164 , n35158 , n382767 );
buf ( n382769 , n35164 );
xor ( n35166 , n382686 , n382689 );
and ( n35167 , n35166 , n382694 );
and ( n35168 , n382686 , n382689 );
or ( n35169 , n35167 , n35168 );
buf ( n382774 , n35169 );
buf ( n382775 , n382774 );
buf ( n382776 , n364664 );
not ( n35173 , n382776 );
buf ( n382778 , n576 );
nand ( n35175 , n35173 , n382778 );
buf ( n382780 , n35175 );
buf ( n382781 , n382780 );
and ( n35178 , n382775 , n382781 );
buf ( n382783 , n35178 );
not ( n35180 , n382783 );
buf ( n382785 , n382774 );
buf ( n382786 , n382780 );
or ( n35183 , n382785 , n382786 );
buf ( n382788 , n35183 );
nand ( n35185 , n35180 , n382788 );
nor ( n35186 , n382769 , n35185 );
not ( n35187 , n35186 );
or ( n35188 , n35128 , n35187 );
or ( n35189 , n35126 , n382769 );
nand ( n35190 , n35189 , n35185 );
nand ( n35191 , n35188 , n35190 );
not ( n35192 , n35191 );
buf ( n382797 , n379542 );
not ( n35194 , n382797 );
buf ( n382799 , n35063 );
nor ( n35196 , n35194 , n382799 );
buf ( n382801 , n35196 );
buf ( n382802 , n382801 );
not ( n35199 , n382802 );
buf ( n382804 , n379303 );
not ( n35201 , n382804 );
or ( n35202 , n35199 , n35201 );
buf ( n382807 , n382759 );
not ( n35204 , n382807 );
buf ( n382809 , n35204 );
buf ( n382810 , n382809 );
nand ( n35207 , n35202 , n382810 );
buf ( n382812 , n35207 );
buf ( n382813 , n382735 );
buf ( n382814 , n382766 );
nand ( n35211 , n382813 , n382814 );
buf ( n382816 , n35211 );
buf ( n382817 , n382816 );
not ( n35214 , n382817 );
buf ( n382819 , n35214 );
and ( n35216 , n382812 , n382819 );
not ( n35217 , n382812 );
and ( n35218 , n35217 , n382816 );
nor ( n35219 , n35216 , n35218 );
buf ( n382824 , n35219 );
not ( n35221 , n382824 );
buf ( n382826 , n35221 );
not ( n35223 , n382826 );
or ( n35224 , n35192 , n35223 );
not ( n35225 , n35191 );
nand ( n35226 , n35219 , n35225 );
nand ( n35227 , n35224 , n35226 );
and ( n35231 , n382702 , n382788 );
not ( n35232 , n35231 );
not ( n35233 , n379558 );
or ( n35234 , n35232 , n35233 );
buf ( n382836 , n382735 );
not ( n35236 , n382836 );
buf ( n382838 , n382753 );
not ( n35238 , n382838 );
or ( n35239 , n35236 , n35238 );
buf ( n382841 , n382766 );
nand ( n35241 , n35239 , n382841 );
buf ( n382843 , n35241 );
buf ( n382844 , n382843 );
buf ( n382845 , n382788 );
and ( n35245 , n382844 , n382845 );
buf ( n382847 , n382783 );
nor ( n35247 , n35245 , n382847 );
buf ( n382849 , n35247 );
nand ( n35249 , n35234 , n382849 );
not ( n35262 , n35249 );
buf ( n382852 , n35262 );
buf ( n35264 , n382852 );
buf ( n382854 , n35264 );
buf ( n382855 , n382854 );
buf ( n35267 , n382855 );
buf ( n382857 , n35267 );
buf ( n382858 , n382857 );
not ( n35270 , n382858 );
not ( n35271 , n34912 );
nand ( n35272 , n35271 , n34892 );
buf ( n382862 , n35272 );
not ( n35274 , n382862 );
buf ( n382864 , n35274 );
buf ( n382865 , n382864 );
not ( n35277 , n382865 );
buf ( n382867 , n35277 );
not ( n35279 , n382867 );
buf ( n35280 , n34650 );
and ( n35281 , n35280 , n33947 );
nor ( n35282 , n35281 , n34653 );
not ( n35283 , n35282 );
nand ( n35284 , n34645 , n34655 );
nor ( n35285 , n35283 , n35284 );
nand ( n35286 , n35279 , n35285 );
buf ( n382876 , n381557 );
not ( n35288 , n382876 );
buf ( n382878 , n35288 );
not ( n35290 , n382878 );
not ( n35291 , n35284 );
nor ( n35292 , n35290 , n35291 );
nand ( n35293 , n382867 , n35292 );
not ( n35294 , n35291 );
not ( n35295 , n35282 );
and ( n35296 , n35294 , n35295 );
nor ( n35297 , n35284 , n382878 );
and ( n35298 , n35282 , n35297 );
nor ( n35299 , n35296 , n35298 );
nand ( n35300 , n35286 , n35293 , n35299 );
buf ( n35301 , n35300 );
buf ( n382891 , n35301 );
buf ( n35303 , n382891 );
buf ( n382893 , n35303 );
buf ( n382894 , n382893 );
not ( n35306 , n382894 );
buf ( n382896 , n35306 );
buf ( n382897 , n382896 );
not ( n35309 , n382897 );
or ( n35310 , n35270 , n35309 );
buf ( n382900 , n382893 );
buf ( n382901 , n382857 );
not ( n35313 , n382901 );
buf ( n382903 , n35313 );
buf ( n382904 , n382903 );
nand ( n35316 , n382900 , n382904 );
buf ( n382906 , n35316 );
buf ( n382907 , n382906 );
nand ( n35319 , n35310 , n382907 );
buf ( n382909 , n35319 );
buf ( n382910 , n382857 );
not ( n35325 , n382910 );
and ( n35326 , n382398 , n382393 );
nor ( n35327 , n35326 , n34844 );
not ( n35328 , n33955 );
not ( n35329 , n34606 );
or ( n35330 , n35328 , n35329 );
nand ( n35331 , n35330 , n34657 );
xor ( n35332 , n35327 , n35331 );
buf ( n382919 , n35332 );
buf ( n35334 , n382919 );
buf ( n382921 , n35334 );
buf ( n382922 , n382921 );
not ( n35337 , n382922 );
buf ( n382924 , n35337 );
buf ( n382925 , n382924 );
not ( n35340 , n382925 );
or ( n35341 , n35325 , n35340 );
buf ( n382928 , n382921 );
buf ( n382929 , n382903 );
nand ( n35344 , n382928 , n382929 );
buf ( n382931 , n35344 );
buf ( n382932 , n382931 );
nand ( n35347 , n35341 , n382932 );
buf ( n382934 , n35347 );
buf ( n382935 , n382934 );
buf ( n382936 , n35227 );
buf ( n35351 , n382936 );
buf ( n382938 , n35351 );
buf ( n382939 , n382938 );
not ( n35354 , n382939 );
buf ( n382941 , n35354 );
buf ( n382942 , n382941 );
buf ( n35357 , n382942 );
buf ( n382944 , n35357 );
buf ( n382945 , n382944 );
not ( n35360 , n382945 );
buf ( n382947 , n35360 );
buf ( n382948 , n382947 );
buf ( n35363 , n382948 );
buf ( n382950 , n35363 );
buf ( n382951 , n382950 );
nand ( n35366 , n382935 , n382951 );
buf ( n382953 , n35366 );
buf ( n382954 , n382953 );
nand ( n35369 , C1 , n382954 );
buf ( n382956 , n35369 );
buf ( n382957 , n382956 );
not ( n35372 , n382957 );
buf ( n382959 , n35372 );
buf ( n382960 , n382959 );
not ( n35375 , n382960 );
or ( n35376 , n35011 , n35375 );
buf ( n35377 , n35219 );
not ( n35378 , n31916 );
not ( n35379 , n379558 );
or ( n35380 , n35378 , n35379 );
nand ( n35381 , n35380 , n379527 );
buf ( n382968 , n382666 );
buf ( n382969 , n382750 );
nand ( n35384 , n382968 , n382969 );
buf ( n382971 , n35384 );
buf ( n382972 , n382971 );
not ( n35387 , n382972 );
buf ( n382974 , n35387 );
and ( n35389 , n35381 , n382974 );
not ( n35390 , n35381 );
and ( n35391 , n35390 , n382971 );
nor ( n35392 , n35389 , n35391 );
buf ( n382979 , n35392 );
not ( n35394 , n382979 );
buf ( n382981 , n35394 );
buf ( n382982 , n382981 );
not ( n35397 , n382982 );
buf ( n382984 , n35397 );
and ( n35399 , n35377 , n382984 );
buf ( n35400 , n35219 );
buf ( n382987 , n35400 );
not ( n35402 , n382987 );
buf ( n382989 , n35402 );
and ( n35404 , n382989 , n382981 );
nor ( n35405 , n35399 , n35404 );
buf ( n382992 , n31961 );
not ( n35407 , n382992 );
buf ( n382994 , n35407 );
buf ( n382995 , n382994 );
buf ( n382996 , n35381 );
buf ( n382997 , n382974 );
and ( n35412 , n382996 , n382997 );
not ( n35413 , n382996 );
buf ( n383000 , n382971 );
and ( n35415 , n35413 , n383000 );
nor ( n35416 , n35412 , n35415 );
buf ( n383003 , n35416 );
buf ( n383004 , n383003 );
and ( n35419 , n382995 , n383004 );
not ( n35420 , n382995 );
buf ( n383007 , n382981 );
and ( n35422 , n35420 , n383007 );
nor ( n35423 , n35419 , n35422 );
buf ( n383010 , n35423 );
nand ( n35425 , n35405 , n383010 );
buf ( n383012 , n35425 );
buf ( n35427 , n383012 );
buf ( n383014 , n35427 );
buf ( n383015 , n383014 );
not ( n35430 , n383015 );
buf ( n383017 , n35430 );
buf ( n35432 , n383017 );
buf ( n383019 , n35432 );
not ( n35434 , n383019 );
buf ( n35435 , n35400 );
buf ( n383022 , n35435 );
not ( n35437 , n383022 );
buf ( n383024 , n35437 );
buf ( n383025 , n383024 );
not ( n35440 , n383025 );
buf ( n383027 , n35440 );
buf ( n383028 , n383027 );
not ( n35443 , n383028 );
not ( n35444 , n34844 );
nand ( n35445 , n35331 , n35444 );
buf ( n383032 , n382412 );
not ( n35447 , n383032 );
buf ( n383034 , n382418 );
nand ( n35449 , n35447 , n383034 );
buf ( n383036 , n35449 );
not ( n35451 , n383036 );
or ( n35452 , n35445 , n35451 );
not ( n35453 , n34795 );
nand ( n35454 , n35453 , n383036 );
and ( n35455 , n35454 , n35444 );
not ( n35456 , n35455 );
not ( n35457 , n35331 );
or ( n35458 , n35456 , n35457 );
not ( n35459 , n34795 );
nor ( n35460 , n35459 , n383036 );
not ( n35461 , n35460 );
nand ( n35462 , n35461 , n35454 );
nand ( n35463 , n35458 , n35462 );
nand ( n35464 , n35452 , n35463 );
buf ( n383051 , n35464 );
buf ( n35466 , n383051 );
buf ( n383053 , n35466 );
buf ( n383054 , n383053 );
buf ( n35469 , n383054 );
buf ( n383056 , n35469 );
buf ( n383057 , n383056 );
not ( n35472 , n383057 );
buf ( n383059 , n35472 );
buf ( n383060 , n383059 );
buf ( n35475 , n383060 );
buf ( n383062 , n35475 );
buf ( n383063 , n383062 );
not ( n35478 , n383063 );
or ( n35479 , n35443 , n35478 );
buf ( n383066 , n383062 );
not ( n35481 , n383066 );
buf ( n383068 , n35481 );
buf ( n383069 , n383068 );
buf ( n383070 , n383027 );
not ( n35485 , n383070 );
buf ( n383072 , n35485 );
buf ( n383073 , n383072 );
nand ( n35488 , n383069 , n383073 );
buf ( n383075 , n35488 );
buf ( n383076 , n383075 );
nand ( n35491 , n35479 , n383076 );
buf ( n383078 , n35491 );
buf ( n383079 , n383078 );
not ( n35494 , n383079 );
or ( n35495 , n35434 , n35494 );
buf ( n383082 , n383027 );
not ( n35497 , n383082 );
not ( n35498 , n34892 );
nand ( n35499 , n34903 , n34504 );
not ( n35500 , n35499 );
or ( n35501 , n35498 , n35500 );
buf ( n383088 , n382501 );
not ( n35503 , n383088 );
buf ( n383090 , n35503 );
nand ( n35505 , n35501 , n383090 );
buf ( n383092 , n34640 );
buf ( n383093 , n383090 );
and ( n35508 , n383092 , n383093 );
buf ( n383095 , n34888 );
nor ( n35510 , n35508 , n383095 );
buf ( n383097 , n35510 );
nand ( n35512 , n35505 , n383097 );
nand ( n35513 , n34752 , n34821 );
not ( n35514 , n35513 );
and ( n35515 , n35512 , n35514 );
not ( n35516 , n35512 );
and ( n35517 , n35516 , n35513 );
nor ( n35518 , n35515 , n35517 );
buf ( n35519 , n35518 );
buf ( n383106 , n35519 );
not ( n35521 , n383106 );
buf ( n383108 , n35521 );
buf ( n383109 , n383108 );
not ( n35524 , n383109 );
buf ( n383111 , n35524 );
buf ( n383112 , n383111 );
not ( n35527 , n383112 );
buf ( n383114 , n35527 );
buf ( n383115 , n383114 );
buf ( n35530 , n383115 );
buf ( n383117 , n35530 );
buf ( n383118 , n383117 );
not ( n35533 , n383118 );
or ( n35534 , n35497 , n35533 );
buf ( n383121 , n383117 );
not ( n35536 , n383121 );
buf ( n383123 , n35536 );
buf ( n383124 , n383123 );
buf ( n383125 , n383072 );
nand ( n35540 , n383124 , n383125 );
buf ( n383127 , n35540 );
buf ( n383128 , n383127 );
nand ( n35543 , n35534 , n383128 );
buf ( n383130 , n35543 );
buf ( n383131 , n383130 );
buf ( n383132 , n383010 );
buf ( n35547 , n383132 );
buf ( n383134 , n35547 );
buf ( n383135 , n383134 );
not ( n35550 , n383135 );
buf ( n383137 , n35550 );
buf ( n383138 , n383137 );
nand ( n35553 , n383131 , n383138 );
buf ( n383140 , n35553 );
buf ( n383141 , n383140 );
nand ( n35556 , n35495 , n383141 );
buf ( n383143 , n35556 );
buf ( n383144 , n383143 );
nand ( n35559 , n35376 , n383144 );
buf ( n383146 , n35559 );
buf ( n383147 , n383146 );
buf ( n383148 , n382956 );
buf ( n383149 , n382613 );
not ( n35564 , n383149 );
buf ( n383151 , n35564 );
buf ( n383152 , n383151 );
nand ( n35567 , n383148 , n383152 );
buf ( n383154 , n35567 );
buf ( n383155 , n383154 );
and ( n35570 , n383147 , n383155 );
buf ( n383157 , n35570 );
buf ( n383158 , n383157 );
not ( n35573 , n383158 );
buf ( n383160 , n35573 );
buf ( n383161 , n383160 );
buf ( n383162 , n382613 );
nand ( n35577 , n383161 , n383162 );
buf ( n383164 , n35577 );
not ( n35579 , n383164 );
buf ( n383166 , n383027 );
not ( n35581 , n383166 );
buf ( n383168 , n382538 );
not ( n35583 , n383168 );
or ( n35584 , n35581 , n35583 );
buf ( n383171 , n382551 );
buf ( n383172 , n383072 );
nand ( n35587 , n383171 , n383172 );
buf ( n383174 , n35587 );
buf ( n383175 , n383174 );
nand ( n35590 , n35584 , n383175 );
buf ( n383177 , n35590 );
buf ( n383178 , n383177 );
not ( n35593 , n383178 );
buf ( n383180 , n383017 );
not ( n35595 , n383180 );
buf ( n383182 , n35595 );
buf ( n383183 , n383182 );
nor ( n35598 , n35593 , n383183 );
buf ( n383185 , n35598 );
buf ( n383186 , n383185 );
buf ( n383187 , n382473 );
not ( n35602 , n383187 );
buf ( n383189 , n383072 );
not ( n35604 , n383189 );
and ( n35605 , n35602 , n35604 );
buf ( n383192 , n382473 );
buf ( n383193 , n383072 );
and ( n35608 , n383192 , n383193 );
nor ( n35609 , n35605 , n35608 );
buf ( n383196 , n35609 );
buf ( n383197 , n383196 );
buf ( n383198 , n383137 );
not ( n35613 , n383198 );
buf ( n383200 , n35613 );
buf ( n383201 , n383200 );
nor ( n35616 , n383197 , n383201 );
buf ( n383203 , n35616 );
buf ( n383204 , n383203 );
nor ( n35619 , n383186 , n383204 );
buf ( n383206 , n35619 );
buf ( n383207 , n383206 );
buf ( n383208 , n382903 );
buf ( n383209 , n383062 );
xnor ( n35626 , n383208 , n383209 );
buf ( n383211 , n35626 );
buf ( n383212 , n382903 );
buf ( n383213 , n383117 );
and ( n35636 , n383212 , n383213 );
not ( n35637 , n383212 );
buf ( n383216 , n383123 );
and ( n35639 , n35637 , n383216 );
nor ( n35640 , n35636 , n35639 );
buf ( n383219 , n35640 );
buf ( n383220 , n383219 );
buf ( n383221 , n382950 );
nand ( n35644 , n383220 , n383221 );
buf ( n383223 , n35644 );
buf ( n383224 , n383223 );
nand ( n35647 , C1 , n383224 );
buf ( n383226 , n35647 );
buf ( n383227 , n383226 );
xor ( n35650 , n383207 , n383227 );
buf ( n383229 , n383137 );
not ( n35652 , n383229 );
buf ( n383231 , n383177 );
not ( n35654 , n383231 );
or ( n35655 , n35652 , n35654 );
buf ( n383234 , n383130 );
buf ( n383235 , n383017 );
nand ( n35658 , n383234 , n383235 );
buf ( n383237 , n35658 );
buf ( n383238 , n383237 );
nand ( n35661 , n35655 , n383238 );
buf ( n383240 , n35661 );
buf ( n383241 , n383240 );
not ( n35664 , n383241 );
buf ( n383243 , n379466 );
not ( n35666 , n383243 );
buf ( n383245 , n35666 );
buf ( n383246 , n383245 );
not ( n35669 , n383246 );
buf ( n383248 , n382604 );
not ( n35671 , n383248 );
or ( n35672 , n35669 , n35671 );
buf ( n383251 , n382480 );
nand ( n35674 , n35672 , n383251 );
buf ( n383253 , n35674 );
buf ( n383254 , n383253 );
not ( n35677 , n383254 );
buf ( n383256 , n35677 );
buf ( n383257 , n383256 );
nand ( n35680 , n35664 , n383257 );
buf ( n383259 , n35680 );
buf ( n383260 , n383259 );
not ( n35683 , n383260 );
buf ( n383262 , n383211 );
not ( n35685 , n383262 );
buf ( n383264 , n382950 );
not ( n35687 , n383264 );
buf ( n383266 , n35687 );
buf ( n383267 , n383266 );
not ( n35690 , n383267 );
and ( n35691 , n35685 , n35690 );
nor ( n35695 , n35691 , C0 );
buf ( n383271 , n35695 );
buf ( n383272 , n383271 );
not ( n35698 , n383272 );
buf ( n383274 , n35698 );
buf ( n383275 , n383274 );
not ( n35701 , n383275 );
or ( n35702 , n35683 , n35701 );
buf ( n383278 , n383253 );
buf ( n383279 , n383240 );
nand ( n35705 , n383278 , n383279 );
buf ( n383281 , n35705 );
buf ( n383282 , n383281 );
nand ( n35708 , n35702 , n383282 );
buf ( n383284 , n35708 );
buf ( n383285 , n383284 );
xor ( n35711 , n35650 , n383285 );
buf ( n383287 , n35711 );
not ( n35713 , n383287 );
buf ( n383289 , n383151 );
not ( n35715 , n383289 );
buf ( n383291 , n383157 );
not ( n35717 , n383291 );
or ( n35718 , n35715 , n35717 );
buf ( n383294 , n383271 );
not ( n35720 , n383294 );
buf ( n383296 , n383256 );
not ( n35722 , n383296 );
buf ( n383298 , n383240 );
not ( n35724 , n383298 );
or ( n35725 , n35722 , n35724 );
buf ( n383301 , n383240 );
buf ( n383302 , n383256 );
or ( n35728 , n383301 , n383302 );
nand ( n35729 , n35725 , n35728 );
buf ( n383305 , n35729 );
buf ( n383306 , n383305 );
not ( n35732 , n383306 );
and ( n35733 , n35720 , n35732 );
buf ( n383309 , n383271 );
buf ( n383310 , n383305 );
and ( n35736 , n383309 , n383310 );
nor ( n35737 , n35733 , n35736 );
buf ( n383313 , n35737 );
buf ( n383314 , n383313 );
not ( n35740 , n383314 );
buf ( n383316 , n35740 );
buf ( n383317 , n383316 );
nand ( n35743 , n35718 , n383317 );
buf ( n383319 , n35743 );
nand ( n35745 , n35713 , n383319 );
nor ( n35746 , n35579 , n35745 );
buf ( n383322 , n35746 );
not ( n35748 , n383322 );
nand ( n35749 , n383319 , n383164 );
buf ( n383325 , n35749 );
buf ( n383326 , n383287 );
nand ( n35752 , n383325 , n383326 );
buf ( n383328 , n35752 );
buf ( n383329 , n383328 );
nand ( n35755 , n35748 , n383329 );
buf ( n383331 , n35755 );
buf ( n383332 , n383331 );
buf ( n383333 , n383331 );
not ( n35759 , n383333 );
buf ( n383335 , n35759 );
buf ( n383336 , n383335 );
buf ( n383337 , n379466 );
not ( n35763 , n383337 );
buf ( n383339 , n382557 );
not ( n35765 , n383339 );
or ( n35766 , n35763 , n35765 );
buf ( n383342 , n383123 );
not ( n35768 , n383342 );
buf ( n383344 , n379574 );
not ( n35770 , n383344 );
and ( n35771 , n35768 , n35770 );
buf ( n383347 , n383123 );
buf ( n383348 , n379574 );
and ( n35774 , n383347 , n383348 );
nor ( n35775 , n35771 , n35774 );
buf ( n383351 , n35775 );
buf ( n383352 , n383351 );
not ( n35778 , n383352 );
buf ( n383354 , n382607 );
nand ( n35780 , n35778 , n383354 );
buf ( n383356 , n35780 );
buf ( n383357 , n383356 );
nand ( n35783 , n35766 , n383357 );
buf ( n383359 , n35783 );
buf ( n383360 , n383359 );
not ( n35786 , n383360 );
or ( n35787 , n377694 , n377697 );
buf ( n383363 , n379319 );
buf ( n35789 , n383363 );
buf ( n383365 , n35789 );
nand ( n35791 , n35787 , n383365 );
and ( n35792 , n31833 , n35791 );
not ( n35793 , n31833 );
not ( n35794 , n35791 );
and ( n35795 , n35793 , n35794 );
nor ( n35796 , n35792 , n35795 );
buf ( n35797 , n35796 );
not ( n35798 , n35797 );
not ( n35799 , n35798 );
nor ( n35800 , n377588 , n377404 );
buf ( n383376 , n35800 );
not ( n35802 , n383376 );
buf ( n383378 , n379324 );
nand ( n35804 , n35802 , n383378 );
buf ( n383380 , n35804 );
not ( n35806 , n383380 );
not ( n35807 , n35806 );
buf ( n383383 , n35787 );
not ( n35809 , n383383 );
buf ( n383385 , n31833 );
not ( n35811 , n383385 );
or ( n35812 , n35809 , n35811 );
buf ( n383388 , n383365 );
nand ( n35814 , n35812 , n383388 );
buf ( n383390 , n35814 );
not ( n35816 , n383390 );
not ( n35817 , n35816 );
or ( n35818 , n35807 , n35817 );
nand ( n35819 , n383390 , n383380 );
nand ( n35820 , n35818 , n35819 );
not ( n35821 , n35820 );
or ( n35822 , n35799 , n35821 );
not ( n35823 , n35820 );
nand ( n35824 , n35823 , n35797 );
nand ( n35825 , n35822 , n35824 );
buf ( n383401 , n35825 );
buf ( n35827 , n383401 );
buf ( n383403 , n35827 );
buf ( n383404 , n383403 );
not ( n35830 , n383404 );
buf ( n383406 , n35830 );
buf ( n383407 , n383406 );
buf ( n35833 , n383407 );
buf ( n383409 , n35833 );
buf ( n383410 , n383409 );
not ( n35836 , n383410 );
buf ( n383412 , n31844 );
buf ( n35838 , n383412 );
buf ( n383414 , n35838 );
buf ( n383415 , n383414 );
not ( n35841 , n383415 );
buf ( n383417 , n35841 );
buf ( n383418 , n383417 );
buf ( n35844 , n383418 );
buf ( n383420 , n35844 );
buf ( n383421 , n383420 );
not ( n35847 , n383421 );
buf ( n383423 , n35847 );
buf ( n383424 , n383423 );
not ( n35850 , n383424 );
buf ( n383426 , n35850 );
buf ( n383427 , n383426 );
not ( n35853 , n383427 );
buf ( n383429 , n35853 );
and ( n35855 , n383429 , n34863 );
not ( n35856 , n383429 );
and ( n35857 , n35856 , n382473 );
or ( n35858 , n35855 , n35857 );
buf ( n383434 , n35858 );
not ( n35860 , n383434 );
or ( n35861 , n35836 , n35860 );
buf ( n383437 , n383429 );
not ( n35863 , n383437 );
buf ( n383439 , n382538 );
not ( n35865 , n383439 );
or ( n35866 , n35863 , n35865 );
buf ( n383442 , n382551 );
buf ( n383443 , n383429 );
not ( n35869 , n383443 );
buf ( n383445 , n35869 );
buf ( n383446 , n383445 );
nand ( n35872 , n383442 , n383446 );
buf ( n383448 , n35872 );
buf ( n383449 , n383448 );
nand ( n35875 , n35866 , n383449 );
buf ( n383451 , n35875 );
buf ( n383452 , n383451 );
buf ( n383453 , n35825 );
buf ( n383454 , n35820 );
buf ( n383455 , n383414 );
and ( n35881 , n383454 , n383455 );
not ( n35882 , n383454 );
buf ( n383458 , n383414 );
not ( n35884 , n383458 );
buf ( n383460 , n35884 );
buf ( n383461 , n383460 );
and ( n35887 , n35882 , n383461 );
nor ( n35888 , n35881 , n35887 );
buf ( n383464 , n35888 );
buf ( n383465 , n383464 );
nand ( n35891 , n383453 , n383465 );
buf ( n383467 , n35891 );
buf ( n383468 , n383467 );
not ( n35894 , n383468 );
buf ( n383470 , n35894 );
buf ( n383471 , n383470 );
buf ( n35897 , n383471 );
buf ( n383473 , n35897 );
buf ( n383474 , n383473 );
not ( n35900 , n383474 );
buf ( n383476 , n35900 );
buf ( n383477 , n383476 );
buf ( n35903 , n383477 );
buf ( n383479 , n35903 );
buf ( n383480 , n383479 );
not ( n35906 , n383480 );
buf ( n383482 , n35906 );
buf ( n383483 , n383482 );
nand ( n35909 , n383452 , n383483 );
buf ( n383485 , n35909 );
buf ( n383486 , n383485 );
nand ( n35912 , n35861 , n383486 );
buf ( n383488 , n35912 );
buf ( n383489 , n383488 );
not ( n35915 , n383489 );
or ( n35916 , n35786 , n35915 );
buf ( n383492 , n383488 );
buf ( n383493 , n383359 );
or ( n35919 , n383492 , n383493 );
buf ( n383495 , n35858 );
buf ( n383496 , n383479 );
buf ( n383497 , n383409 );
not ( n35923 , n383497 );
buf ( n383499 , n35923 );
buf ( n383500 , n383499 );
nand ( n35926 , n383496 , n383500 );
buf ( n383502 , n35926 );
buf ( n383503 , n383502 );
and ( n35929 , n383495 , n383503 );
buf ( n383505 , n35929 );
buf ( n383506 , n383505 );
not ( n35932 , n383506 );
buf ( n383508 , n35932 );
buf ( n383509 , n383508 );
nand ( n35935 , n35919 , n383509 );
buf ( n383511 , n35935 );
buf ( n383512 , n383511 );
nand ( n35938 , n35916 , n383512 );
buf ( n383514 , n35938 );
buf ( n383515 , n383514 );
buf ( n383516 , n383143 );
not ( n35942 , n383516 );
buf ( n383518 , n382613 );
not ( n35944 , n383518 );
and ( n35945 , n35942 , n35944 );
buf ( n383521 , n383143 );
buf ( n383522 , n382613 );
and ( n35948 , n383521 , n383522 );
nor ( n35949 , n35945 , n35948 );
buf ( n383525 , n35949 );
and ( n35951 , n383525 , n382956 );
not ( n35952 , n383525 );
and ( n35953 , n35952 , n382959 );
or ( n35954 , n35951 , n35953 );
buf ( n383530 , n35954 );
xor ( n35956 , n383515 , n383530 );
buf ( n383532 , n35432 );
not ( n35958 , n383532 );
buf ( n383534 , n383027 );
not ( n35960 , n383534 );
buf ( n383536 , n382924 );
not ( n35962 , n383536 );
or ( n35963 , n35960 , n35962 );
buf ( n383539 , n382921 );
buf ( n383540 , n383072 );
nand ( n35966 , n383539 , n383540 );
buf ( n383542 , n35966 );
buf ( n383543 , n383542 );
nand ( n35969 , n35963 , n383543 );
buf ( n383545 , n35969 );
buf ( n383546 , n383545 );
not ( n35972 , n383546 );
or ( n35973 , n35958 , n35972 );
buf ( n383549 , n383078 );
buf ( n383550 , n383137 );
nand ( n35976 , n383549 , n383550 );
buf ( n383552 , n35976 );
buf ( n383553 , n383552 );
nand ( n35979 , n35973 , n383553 );
buf ( n383555 , n35979 );
buf ( n383556 , n383555 );
not ( n35982 , n383556 );
and ( n35983 , n382909 , n382950 );
buf ( n383559 , n382857 );
not ( n35985 , n383559 );
not ( n35986 , n35272 );
not ( n35987 , n381544 );
or ( n35988 , n35986 , n35987 );
not ( n35989 , n35280 );
nand ( n35990 , n35988 , n35989 );
nand ( n35991 , n33947 , n34652 );
not ( n35992 , n35991 );
and ( n35993 , n35990 , n35992 );
not ( n35994 , n35990 );
and ( n35995 , n35994 , n35991 );
nor ( n35996 , n35993 , n35995 );
buf ( n35997 , n35996 );
buf ( n383573 , n35997 );
not ( n35999 , n383573 );
buf ( n383575 , n35999 );
buf ( n383576 , n383575 );
buf ( n36002 , n383576 );
buf ( n383578 , n36002 );
buf ( n383579 , n383578 );
not ( n36005 , n383579 );
or ( n36006 , n35985 , n36005 );
buf ( n383582 , n383578 );
not ( n36008 , n383582 );
buf ( n383584 , n36008 );
buf ( n383585 , n383584 );
buf ( n383586 , n382903 );
nand ( n36012 , n383585 , n383586 );
buf ( n383588 , n36012 );
buf ( n383589 , n383588 );
nand ( n36015 , n36006 , n383589 );
buf ( n383591 , n36015 );
nor ( n36018 , n35983 , C0 );
buf ( n383593 , n36018 );
nand ( n36020 , n35982 , n383593 );
buf ( n383595 , n36020 );
buf ( n383596 , n383595 );
not ( n36023 , n383596 );
not ( n36024 , n383351 );
not ( n36025 , n383245 );
and ( n36026 , n36024 , n36025 );
buf ( n383601 , n379577 );
not ( n36028 , n383601 );
buf ( n383603 , n383062 );
not ( n36030 , n383603 );
or ( n36031 , n36028 , n36030 );
buf ( n383606 , n383068 );
buf ( n383607 , n379574 );
nand ( n36034 , n383606 , n383607 );
buf ( n383609 , n36034 );
buf ( n383610 , n383609 );
nand ( n36037 , n36031 , n383610 );
buf ( n383612 , n36037 );
and ( n36039 , n383612 , n382607 );
nor ( n36040 , n36026 , n36039 );
buf ( n383615 , n36040 );
not ( n36042 , n383615 );
buf ( n383617 , n36042 );
buf ( n383618 , n383617 );
not ( n36045 , n383618 );
buf ( n383620 , n382950 );
not ( n36047 , n383620 );
buf ( n383622 , n383591 );
not ( n36049 , n383622 );
or ( n36050 , n36047 , n36049 );
buf ( n383625 , n382857 );
not ( n36052 , n383625 );
not ( n36053 , n33905 );
not ( n36054 , n36053 );
not ( n36055 , n35272 );
or ( n36056 , n36054 , n36055 );
buf ( n36057 , n34646 );
nand ( n36058 , n36056 , n36057 );
not ( n36059 , n381541 );
nand ( n36060 , n36059 , n34649 );
not ( n36061 , n36060 );
and ( n36062 , n36058 , n36061 );
not ( n36063 , n36058 );
and ( n36064 , n36063 , n36060 );
nor ( n36065 , n36062 , n36064 );
buf ( n36066 , n36065 );
not ( n36067 , n36066 );
not ( n36068 , n36067 );
not ( n36069 , n36068 );
buf ( n383644 , n36069 );
not ( n36071 , n383644 );
or ( n36072 , n36052 , n36071 );
not ( n36073 , n36069 );
buf ( n383648 , n36073 );
buf ( n383649 , n382903 );
nand ( n36076 , n383648 , n383649 );
buf ( n383651 , n36076 );
buf ( n383652 , n383651 );
nand ( n36079 , n36072 , n383652 );
buf ( n383654 , n36079 );
buf ( n383655 , C1 );
buf ( n383656 , n383655 );
nand ( n36086 , n36050 , n383656 );
buf ( n383658 , n36086 );
buf ( n383659 , n383658 );
not ( n36089 , n383659 );
or ( n36090 , n36045 , n36089 );
buf ( n383662 , n383658 );
not ( n36092 , n383662 );
buf ( n383664 , n36092 );
buf ( n383665 , n383664 );
buf ( n383666 , n36040 );
nand ( n36096 , n383665 , n383666 );
buf ( n383668 , n36096 );
buf ( n383669 , n383668 );
buf ( n383670 , n383017 );
not ( n36100 , n383670 );
buf ( n383672 , n383027 );
not ( n36102 , n383672 );
buf ( n383674 , n382896 );
not ( n36104 , n383674 );
or ( n36105 , n36102 , n36104 );
buf ( n383677 , n382893 );
buf ( n383678 , n383072 );
nand ( n36108 , n383677 , n383678 );
buf ( n383680 , n36108 );
buf ( n383681 , n383680 );
nand ( n36111 , n36105 , n383681 );
buf ( n383683 , n36111 );
buf ( n383684 , n383683 );
not ( n36114 , n383684 );
or ( n36115 , n36100 , n36114 );
buf ( n383687 , n383545 );
buf ( n383688 , n383137 );
nand ( n36118 , n383687 , n383688 );
buf ( n383690 , n36118 );
buf ( n383691 , n383690 );
nand ( n36121 , n36115 , n383691 );
buf ( n383693 , n36121 );
buf ( n383694 , n383693 );
nand ( n36124 , n383669 , n383694 );
buf ( n383696 , n36124 );
buf ( n383697 , n383696 );
nand ( n36127 , n36090 , n383697 );
buf ( n383699 , n36127 );
buf ( n383700 , n383699 );
not ( n36130 , n383700 );
or ( n36131 , n36023 , n36130 );
buf ( n383703 , n36018 );
not ( n36133 , n383703 );
buf ( n383705 , n383555 );
nand ( n36135 , n36133 , n383705 );
buf ( n383707 , n36135 );
buf ( n383708 , n383707 );
nand ( n36138 , n36131 , n383708 );
buf ( n383710 , n36138 );
buf ( n383711 , n383710 );
and ( n36141 , n35956 , n383711 );
and ( n36142 , n383515 , n383530 );
or ( n36143 , n36141 , n36142 );
buf ( n383715 , n36143 );
not ( n36145 , n383715 );
buf ( n383717 , n383151 );
not ( n36147 , n383717 );
buf ( n383719 , n383316 );
not ( n36149 , n383719 );
or ( n36150 , n36147 , n36149 );
buf ( n383722 , n383313 );
buf ( n383723 , n382613 );
nand ( n36153 , n383722 , n383723 );
buf ( n383725 , n36153 );
buf ( n383726 , n383725 );
nand ( n36156 , n36150 , n383726 );
buf ( n383728 , n36156 );
buf ( n383729 , n383728 );
buf ( n383730 , n383157 );
and ( n36160 , n383729 , n383730 );
not ( n36161 , n383729 );
buf ( n383733 , n383160 );
and ( n36163 , n36161 , n383733 );
nor ( n36164 , n36160 , n36163 );
buf ( n383736 , n36164 );
nand ( n36166 , n36145 , n383736 );
not ( n36167 , n36166 );
buf ( n383739 , n383072 );
buf ( n383740 , n380847 );
not ( n36170 , n383740 );
buf ( n383742 , n36170 );
not ( n36172 , n383742 );
not ( n36173 , n34606 );
or ( n36174 , n36172 , n36173 );
buf ( n383746 , n380840 );
buf ( n383747 , n380844 );
nand ( n36177 , n383746 , n383747 );
buf ( n383749 , n36177 );
buf ( n36179 , n383749 );
nand ( n36180 , n36174 , n36179 );
xor ( n36181 , n34620 , n382230 );
not ( n36182 , n36181 );
and ( n36183 , n36180 , n36182 );
not ( n36184 , n36180 );
and ( n36185 , n36184 , n36181 );
nor ( n36186 , n36183 , n36185 );
not ( n36187 , n36186 );
buf ( n36188 , n36187 );
buf ( n383760 , n36188 );
not ( n36190 , n383760 );
buf ( n383762 , n36190 );
buf ( n383763 , n383762 );
not ( n36193 , n383763 );
buf ( n383765 , n36193 );
buf ( n383766 , n383765 );
and ( n36196 , n383739 , n383766 );
not ( n36197 , n383739 );
buf ( n383769 , n383762 );
and ( n36199 , n36197 , n383769 );
nor ( n36200 , n36196 , n36199 );
buf ( n383772 , n36200 );
or ( n36202 , n383772 , n383200 );
not ( n36203 , n383072 );
buf ( n383775 , n34606 );
not ( n36205 , n383775 );
buf ( n383777 , n36205 );
buf ( n383778 , n383742 );
buf ( n383779 , n383749 );
and ( n36209 , n383778 , n383779 );
buf ( n383781 , n36209 );
not ( n36211 , n383781 );
and ( n36212 , n383777 , n36211 );
not ( n36213 , n383777 );
and ( n36214 , n36213 , n383781 );
nor ( n36215 , n36212 , n36214 );
buf ( n36216 , n36215 );
buf ( n36217 , n36216 );
not ( n36218 , n36217 );
not ( n36219 , n36218 );
or ( n36220 , n36203 , n36219 );
not ( n36221 , n36218 );
nand ( n36222 , n383027 , n36221 );
nand ( n36223 , n36220 , n36222 );
not ( n36224 , n36223 );
nand ( n36225 , n36224 , n383017 );
nand ( n36226 , n36202 , n36225 );
not ( n36227 , n36226 );
not ( n36228 , n36227 );
buf ( n383800 , n31558 );
buf ( n383801 , n379194 );
not ( n36231 , n383801 );
buf ( n383803 , n379161 );
nand ( n36233 , n36231 , n383803 );
buf ( n383805 , n36233 );
buf ( n383806 , n383805 );
and ( n36236 , n383800 , n383806 );
buf ( n383808 , n36236 );
not ( n36238 , n383808 );
not ( n36239 , n36238 );
not ( n36240 , n31593 );
not ( n36241 , n31628 );
or ( n36242 , n36240 , n36241 );
not ( n36243 , n31531 );
nand ( n36244 , n36242 , n36243 );
not ( n36245 , n36244 );
not ( n36246 , n36245 );
or ( n36247 , n36239 , n36246 );
nand ( n36248 , n36244 , n383808 );
nand ( n36249 , n36247 , n36248 );
not ( n36250 , n36249 );
not ( n36251 , n36250 );
buf ( n36252 , n36251 );
not ( n36253 , n36252 );
not ( n36254 , n36253 );
not ( n36255 , n34861 );
or ( n36256 , n36254 , n36255 );
or ( n36257 , n34861 , n36253 );
nand ( n36258 , n36256 , n36257 );
not ( n36259 , n36249 );
buf ( n383831 , n36259 );
not ( n36261 , n383831 );
buf ( n383833 , n379109 );
buf ( n36263 , n383833 );
buf ( n383835 , n36263 );
buf ( n383836 , n383835 );
buf ( n383837 , n379129 );
buf ( n36267 , n383837 );
buf ( n383839 , n36267 );
buf ( n383840 , n383839 );
or ( n36270 , n383836 , n383840 );
buf ( n383842 , n36270 );
not ( n36272 , n383842 );
not ( n36273 , n31628 );
or ( n36274 , n36272 , n36273 );
buf ( n383846 , n383835 );
buf ( n383847 , n383839 );
nand ( n36277 , n383846 , n383847 );
buf ( n383849 , n36277 );
nand ( n36279 , n36274 , n383849 );
buf ( n383851 , n379106 );
not ( n36281 , n383851 );
buf ( n383853 , n379067 );
buf ( n383854 , n379103 );
nand ( n36284 , n383853 , n383854 );
buf ( n383856 , n36284 );
buf ( n383857 , n383856 );
nand ( n36287 , n36281 , n383857 );
buf ( n383859 , n36287 );
xnor ( n36289 , n36279 , n383859 );
buf ( n383861 , n36289 );
not ( n36291 , n383861 );
buf ( n383863 , n36291 );
buf ( n383864 , n383863 );
nand ( n36294 , n36261 , n383864 );
buf ( n383866 , n36294 );
and ( n36296 , n383842 , n383849 );
not ( n36297 , n36296 );
not ( n36298 , n31628 );
not ( n36299 , n36298 );
or ( n36300 , n36297 , n36299 );
not ( n36301 , n36298 );
xnor ( n36302 , n383835 , n383839 );
nand ( n36303 , n36301 , n36302 );
nand ( n36304 , n36300 , n36303 );
not ( n36305 , n36304 );
and ( n36306 , n36305 , n36289 );
not ( n36307 , n36305 );
not ( n36308 , n36289 );
and ( n36309 , n36307 , n36308 );
nor ( n36310 , n36306 , n36309 );
buf ( n383882 , n36259 );
xnor ( n36312 , n36279 , n383859 );
buf ( n383884 , n36312 );
nand ( n36314 , n383882 , n383884 );
buf ( n383886 , n36314 );
nand ( n36316 , n383866 , n36310 , n383886 );
not ( n36317 , n36316 );
buf ( n383889 , n36317 );
buf ( n36319 , n383889 );
buf ( n383891 , n36319 );
buf ( n383892 , n383891 );
buf ( n36322 , n383892 );
buf ( n383894 , n36322 );
buf ( n383895 , n383894 );
buf ( n36325 , n383895 );
buf ( n383897 , n36325 );
buf ( n383898 , n383897 );
not ( n36328 , n383898 );
buf ( n383900 , n36328 );
not ( n36330 , n36310 );
buf ( n383902 , n36330 );
buf ( n36332 , n383902 );
buf ( n383904 , n36332 );
buf ( n383905 , n383904 );
buf ( n36335 , n383905 );
buf ( n383907 , n36335 );
buf ( n383908 , n383907 );
not ( n36338 , n383908 );
buf ( n383910 , n36338 );
nand ( n36340 , n383900 , n383910 );
and ( n36341 , n36258 , n36340 );
buf ( n383913 , n36259 );
not ( n36343 , n383913 );
buf ( n383915 , n36343 );
not ( n36345 , n383915 );
buf ( n36346 , n31558 );
not ( n36347 , n36346 );
not ( n36348 , n36244 );
or ( n36349 , n36347 , n36348 );
nand ( n36350 , n36349 , n383805 );
nand ( n36351 , n379185 , n31579 );
nand ( n36352 , n36351 , n31594 );
not ( n36353 , n36352 );
and ( n36354 , n36350 , n36353 );
not ( n36355 , n36350 );
and ( n36356 , n36355 , n36352 );
nor ( n36357 , n36354 , n36356 );
not ( n36358 , n36357 );
or ( n36359 , n36345 , n36358 );
not ( n36360 , n36357 );
nand ( n36361 , n36360 , n36259 );
nand ( n36362 , n36359 , n36361 );
buf ( n36363 , n36362 );
buf ( n383935 , n36363 );
not ( n36365 , n383935 );
buf ( n383937 , n36365 );
buf ( n383938 , n383937 );
not ( n36368 , n383938 );
buf ( n383940 , n36368 );
buf ( n383941 , n383940 );
not ( n36371 , n383941 );
buf ( n383943 , n36371 );
buf ( n383944 , n383943 );
not ( n36374 , n383944 );
buf ( n383946 , n36374 );
not ( n36376 , n383946 );
or ( n36377 , n378580 , n378803 );
buf ( n383949 , n36377 );
buf ( n36379 , n31649 );
buf ( n383951 , n36379 );
nand ( n36381 , n383949 , n383951 );
buf ( n383953 , n36381 );
not ( n36383 , n383953 );
buf ( n383955 , n35121 );
buf ( n36385 , n383955 );
buf ( n383957 , n36385 );
not ( n36387 , n383957 );
or ( n36388 , n36383 , n36387 );
buf ( n383960 , n35121 );
buf ( n383961 , n383953 );
or ( n36391 , n383960 , n383961 );
buf ( n383963 , n36391 );
nand ( n36393 , n36388 , n383963 );
not ( n36394 , n36393 );
buf ( n36395 , n36394 );
not ( n36396 , n36395 );
buf ( n36397 , n36396 );
not ( n36398 , n36397 );
not ( n36399 , n36398 );
and ( n36400 , n36399 , n382535 );
not ( n36401 , n36399 );
buf ( n383973 , n382535 );
not ( n36403 , n383973 );
buf ( n383975 , n36403 );
and ( n36405 , n36401 , n383975 );
or ( n36406 , n36400 , n36405 );
not ( n36407 , n36406 );
or ( n36408 , n36376 , n36407 );
buf ( n383980 , n36399 );
not ( n36410 , n383980 );
buf ( n383982 , n383114 );
not ( n36412 , n383982 );
or ( n36413 , n36410 , n36412 );
buf ( n383985 , n383111 );
buf ( n383986 , n36398 );
nand ( n36416 , n383985 , n383986 );
buf ( n383988 , n36416 );
buf ( n383989 , n383988 );
nand ( n36419 , n36413 , n383989 );
buf ( n383991 , n36419 );
buf ( n383992 , n383991 );
not ( n36422 , n36360 );
not ( n36423 , n36422 );
buf ( n36424 , n36393 );
not ( n36425 , n36424 );
not ( n36426 , n36425 );
or ( n36427 , n36423 , n36426 );
nand ( n36428 , n36424 , n36360 );
nand ( n36429 , n36427 , n36428 );
buf ( n384001 , n36362 );
not ( n36431 , n384001 );
buf ( n384003 , n36431 );
nand ( n36433 , n36429 , n384003 );
buf ( n36434 , n36433 );
buf ( n384006 , n36434 );
buf ( n36436 , n384006 );
buf ( n384008 , n36436 );
buf ( n384009 , n384008 );
not ( n36439 , n384009 );
buf ( n384011 , n36439 );
buf ( n384012 , n384011 );
nand ( n36442 , n383992 , n384012 );
buf ( n384014 , n36442 );
nand ( n36444 , n36408 , n384014 );
xnor ( n36445 , n36341 , n36444 );
not ( n36446 , n36445 );
or ( n36447 , n36228 , n36446 );
not ( n36448 , n36444 );
nand ( n36449 , n36341 , n36448 );
not ( n36450 , n36449 );
not ( n36451 , n36341 );
and ( n36452 , n36444 , n36451 );
or ( n36453 , n36450 , n36452 );
nand ( n36454 , n36453 , n36226 );
nand ( n36455 , n36447 , n36454 );
not ( n36456 , n36455 );
buf ( n384028 , n384011 );
not ( n36458 , n384028 );
buf ( n384030 , n36399 );
not ( n36460 , n384030 );
buf ( n384032 , n383059 );
not ( n384033 , n384032 );
or ( n36463 , n36460 , n384033 );
buf ( n384035 , n383059 );
not ( n36465 , n384035 );
buf ( n384037 , n36465 );
buf ( n384038 , n384037 );
not ( n36468 , n36399 );
buf ( n384040 , n36468 );
nand ( n36470 , n384038 , n384040 );
buf ( n384042 , n36470 );
buf ( n384043 , n384042 );
nand ( n36473 , n36463 , n384043 );
buf ( n384045 , n36473 );
buf ( n384046 , n384045 );
not ( n36476 , n384046 );
or ( n36477 , n36458 , n36476 );
buf ( n384049 , n383991 );
buf ( n384050 , n383946 );
nand ( n36480 , n384049 , n384050 );
buf ( n384052 , n36480 );
buf ( n384053 , n384052 );
nand ( n36483 , n36477 , n384053 );
buf ( n384055 , n36483 );
buf ( n384056 , n384055 );
not ( n36486 , n382947 );
buf ( n384058 , n382854 );
not ( n36488 , n384058 );
buf ( n384060 , n382043 );
buf ( n384061 , n382079 );
nor ( n36491 , n384060 , n384061 );
buf ( n384063 , n36491 );
buf ( n384064 , n384063 );
not ( n36494 , n384064 );
buf ( n384066 , n382082 );
buf ( n36496 , n384066 );
buf ( n384068 , n36496 );
buf ( n384069 , n384068 );
nand ( n36499 , n36494 , n384069 );
buf ( n384071 , n36499 );
buf ( n384072 , n384071 );
not ( n36502 , n384072 );
buf ( n384074 , n36502 );
nand ( n36504 , n382209 , n382161 );
and ( n36505 , n34598 , n34595 , n36504 );
or ( n36506 , n384074 , n36505 );
nand ( n36507 , n384074 , n36505 );
nand ( n36508 , n36506 , n36507 );
buf ( n36509 , n36508 );
buf ( n384081 , n36509 );
not ( n36511 , n384081 );
buf ( n384083 , n36511 );
buf ( n384084 , n384083 );
not ( n36514 , n384084 );
or ( n36515 , n36488 , n36514 );
buf ( n384087 , n36509 );
not ( n36517 , n384087 );
buf ( n384089 , n36517 );
buf ( n384090 , n384089 );
not ( n36520 , n384090 );
buf ( n384092 , n36520 );
buf ( n384093 , n384092 );
buf ( n384094 , n382854 );
not ( n36524 , n384094 );
buf ( n384096 , n36524 );
buf ( n384097 , n384096 );
nand ( n36527 , n384093 , n384097 );
buf ( n384099 , n36527 );
buf ( n384100 , n384099 );
nand ( n36530 , n36515 , n384100 );
buf ( n384102 , n36530 );
not ( n36532 , n384102 );
or ( n36533 , n36486 , n36532 );
buf ( n384105 , n382854 );
not ( n36535 , n384105 );
buf ( n384107 , n382209 );
not ( n36537 , n384107 );
buf ( n384109 , n382164 );
nand ( n36539 , n36537 , n384109 );
buf ( n384111 , n36539 );
and ( n36541 , n384111 , n34603 );
buf ( n384113 , n382151 );
buf ( n36543 , n384113 );
buf ( n384115 , n36543 );
nand ( n36545 , n384115 , n34594 );
and ( n36546 , n36541 , n36545 );
not ( n36547 , n36546 );
not ( n36548 , n28168 );
buf ( n384120 , n384115 );
buf ( n384121 , n376670 );
nand ( n36551 , n384120 , n384121 );
buf ( n384123 , n36551 );
not ( n36553 , n384123 );
nand ( n36554 , n36548 , n36553 , n376375 );
buf ( n36555 , n36554 );
not ( n36556 , n36555 );
or ( n36557 , n36547 , n36556 );
not ( n36558 , n36545 );
not ( n36559 , n36554 );
or ( n36560 , n36558 , n36559 );
not ( n36561 , n36541 );
nand ( n36562 , n36560 , n36561 );
nand ( n36563 , n36557 , n36562 );
buf ( n36564 , n36563 );
not ( n36565 , n36564 );
buf ( n384137 , n36565 );
not ( n36567 , n384137 );
or ( n36568 , n36535 , n36567 );
buf ( n384140 , n36564 );
buf ( n384141 , n35262 );
not ( n36571 , n384141 );
buf ( n384143 , n36571 );
buf ( n384144 , n384143 );
nand ( n36574 , n384140 , n384144 );
buf ( n384146 , n36574 );
buf ( n384147 , n384146 );
nand ( n36577 , n36568 , n384147 );
buf ( n384149 , n36577 );
buf ( n384150 , C1 );
nand ( n36583 , n36533 , n384150 );
buf ( n384152 , n36583 );
buf ( n384153 , n383137 );
not ( n36586 , n384153 );
not ( n36587 , n383027 );
buf ( n36588 , n34511 );
or ( n36589 , n381791 , n381950 );
nand ( n36590 , n36588 , n36589 );
or ( n36591 , n36590 , n36505 );
buf ( n36592 , n382091 );
nand ( n36593 , n36592 , n36589 );
buf ( n36594 , n34493 );
nand ( n36595 , n36593 , n36594 );
not ( n36596 , n36595 );
nand ( n36597 , n36591 , n36596 );
buf ( n36598 , n382097 );
buf ( n36599 , n382107 );
nor ( n36600 , n36598 , n36599 );
not ( n36601 , n36600 );
nor ( n36602 , n36597 , n36601 );
buf ( n384171 , n36602 );
not ( n36604 , n384171 );
not ( n36605 , n36600 );
nand ( n36606 , n36605 , n36597 );
buf ( n384175 , n36606 );
nand ( n36608 , n36604 , n384175 );
buf ( n384177 , n36608 );
buf ( n384178 , n384177 );
buf ( n36611 , n384178 );
buf ( n384180 , n36611 );
buf ( n384181 , n384180 );
not ( n36614 , n384181 );
buf ( n384183 , n36614 );
buf ( n384184 , n384183 );
not ( n36617 , n384184 );
buf ( n384186 , n36617 );
buf ( n384187 , n384186 );
buf ( n36620 , n384187 );
buf ( n384189 , n36620 );
buf ( n384190 , n384189 );
not ( n36623 , n384190 );
buf ( n384192 , n36623 );
not ( n36625 , n384192 );
or ( n36626 , n36587 , n36625 );
buf ( n384195 , n36602 );
not ( n36628 , n384195 );
buf ( n384197 , n36606 );
nand ( n36630 , n36628 , n384197 );
buf ( n384199 , n36630 );
buf ( n384200 , n384199 );
not ( n36633 , n384200 );
buf ( n384202 , n36633 );
buf ( n384203 , n384202 );
not ( n36636 , n384203 );
buf ( n384205 , n36636 );
buf ( n384206 , n384205 );
not ( n36639 , n384206 );
buf ( n384208 , n36639 );
buf ( n384209 , n384208 );
buf ( n36642 , n384209 );
buf ( n384211 , n36642 );
buf ( n384212 , n384211 );
buf ( n384213 , n383027 );
or ( n36646 , n384212 , n384213 );
buf ( n384215 , n36646 );
nand ( n36648 , n36626 , n384215 );
buf ( n384217 , n36648 );
not ( n36650 , n384217 );
or ( n36651 , n36586 , n36650 );
buf ( n384220 , n383017 );
buf ( n384221 , n383027 );
not ( n36654 , n384221 );
and ( n36655 , n36594 , n36589 );
not ( n36656 , n36655 );
not ( n36657 , n36588 );
nand ( n36658 , n34598 , n34595 , n36504 );
not ( n36659 , n36658 );
or ( n36660 , n36657 , n36659 );
not ( n36661 , n36592 );
nand ( n36662 , n36660 , n36661 );
not ( n36663 , n36662 );
not ( n36664 , n36663 );
or ( n36665 , n36656 , n36664 );
not ( n36666 , n36655 );
nand ( n36667 , n36666 , n36662 );
nand ( n36668 , n36665 , n36667 );
buf ( n384237 , n36668 );
not ( n36670 , n384237 );
buf ( n384239 , n36670 );
buf ( n36672 , n384239 );
buf ( n384241 , n36672 );
not ( n36674 , n384241 );
or ( n36675 , n36654 , n36674 );
not ( n36676 , n36672 );
buf ( n384245 , n36676 );
buf ( n384246 , n383024 );
nand ( n36679 , n384245 , n384246 );
buf ( n384248 , n36679 );
buf ( n384249 , n384248 );
nand ( n36682 , n36675 , n384249 );
buf ( n384251 , n36682 );
buf ( n384252 , n384251 );
nand ( n36685 , n384220 , n384252 );
buf ( n384254 , n36685 );
buf ( n384255 , n384254 );
nand ( n36688 , n36651 , n384255 );
buf ( n384257 , n36688 );
buf ( n384258 , n384257 );
xor ( n36691 , n384152 , n384258 );
not ( n36692 , n382950 );
buf ( n384261 , n382854 );
not ( n36694 , n384261 );
not ( n36695 , n384063 );
not ( n36696 , n36695 );
not ( n36697 , n36658 );
or ( n36698 , n36696 , n36697 );
nand ( n36699 , n36698 , n384068 );
not ( n36700 , n382088 );
nand ( n36701 , n382036 , n381960 );
nand ( n36702 , n36700 , n36701 );
not ( n36703 , n36702 );
and ( n36704 , n36699 , n36703 );
not ( n36705 , n36699 );
and ( n36706 , n36705 , n36702 );
nor ( n36707 , n36704 , n36706 );
not ( n36708 , n36707 );
not ( n36709 , n36708 );
buf ( n384278 , n36709 );
not ( n36711 , n384278 );
buf ( n384280 , n36711 );
buf ( n384281 , n384280 );
not ( n36714 , n384281 );
or ( n36715 , n36694 , n36714 );
buf ( n384284 , n384280 );
not ( n36717 , n384284 );
buf ( n384286 , n36717 );
buf ( n384287 , n384286 );
buf ( n384288 , n384096 );
nand ( n36721 , n384287 , n384288 );
buf ( n384290 , n36721 );
buf ( n384291 , n384290 );
nand ( n36724 , n36715 , n384291 );
buf ( n384293 , n36724 );
not ( n36726 , n384293 );
or ( n36727 , n36692 , n36726 );
buf ( n384296 , C1 );
nand ( n36732 , n36727 , n384296 );
buf ( n384298 , n36732 );
and ( n36734 , n36691 , n384298 );
and ( n36735 , n384152 , n384258 );
or ( n36736 , n36734 , n36735 );
buf ( n384302 , n36736 );
buf ( n36738 , n384302 );
buf ( n384304 , n36738 );
xor ( n36740 , n384056 , n384304 );
not ( n36741 , n36377 );
not ( n36742 , n35121 );
or ( n36743 , n36741 , n36742 );
nand ( n36744 , n36743 , n36379 );
buf ( n384310 , n379245 );
buf ( n384311 , n379249 );
or ( n36747 , n384310 , n384311 );
buf ( n384313 , n36747 );
buf ( n384314 , n384313 );
buf ( n384315 , n379261 );
nand ( n36751 , n384314 , n384315 );
buf ( n384317 , n36751 );
and ( n36753 , n36744 , n384317 );
not ( n36754 , n36744 );
not ( n36755 , n384317 );
and ( n36756 , n36754 , n36755 );
nor ( n36757 , n36753 , n36756 );
not ( n36758 , n36757 );
not ( n36759 , n36758 );
nor ( n36760 , n378830 , n378824 );
buf ( n384326 , n36760 );
buf ( n36762 , n384326 );
buf ( n384328 , n36762 );
buf ( n384329 , n384328 );
not ( n36765 , n384329 );
buf ( n384331 , n379287 );
nand ( n36767 , n36765 , n384331 );
buf ( n384333 , n36767 );
not ( n36769 , n384333 );
not ( n36770 , n36769 );
not ( n36771 , n31198 );
not ( n36772 , n36771 );
not ( n36773 , n36772 );
not ( n36774 , n35121 );
or ( n36775 , n36773 , n36774 );
buf ( n384341 , n31655 );
not ( n36777 , n384341 );
buf ( n384343 , n36777 );
nand ( n36779 , n36775 , n384343 );
not ( n36780 , n36779 );
not ( n36781 , n36780 );
or ( n36782 , n36770 , n36781 );
buf ( n384348 , n36779 );
buf ( n384349 , n384333 );
nand ( n36785 , n384348 , n384349 );
buf ( n384351 , n36785 );
nand ( n36787 , n36782 , n384351 );
not ( n36788 , n36787 );
not ( n36789 , n36788 );
or ( n36790 , n36759 , n36789 );
nand ( n36791 , n36787 , n36757 );
nand ( n36792 , n36790 , n36791 );
not ( n36793 , n36757 );
not ( n36794 , n36393 );
or ( n36795 , n36793 , n36794 );
nand ( n36796 , n36394 , n36758 );
nand ( n36797 , n36795 , n36796 );
not ( n36798 , n36797 );
nand ( n36799 , n36792 , n36798 );
not ( n36800 , n36799 );
buf ( n36801 , n36800 );
buf ( n384367 , n36801 );
buf ( n36803 , n384367 );
buf ( n384369 , n36803 );
buf ( n384370 , n384369 );
not ( n36806 , n384370 );
or ( n36807 , n36779 , n384333 );
nand ( n36808 , n36807 , n384351 );
not ( n36809 , n36808 );
not ( n36810 , n36809 );
buf ( n36811 , n36810 );
buf ( n384377 , n36811 );
not ( n36813 , n384377 );
buf ( n384379 , n382893 );
not ( n36815 , n384379 );
buf ( n384381 , n36815 );
buf ( n384382 , n384381 );
not ( n36818 , n384382 );
or ( n36819 , n36813 , n36818 );
buf ( n384385 , n382893 );
not ( n36821 , n36809 );
not ( n36822 , n36821 );
buf ( n384388 , n36822 );
nand ( n36824 , n384385 , n384388 );
buf ( n384390 , n36824 );
buf ( n384391 , n384390 );
nand ( n36827 , n36819 , n384391 );
buf ( n384393 , n36827 );
buf ( n384394 , n384393 );
not ( n36830 , n384394 );
or ( n36831 , n36806 , n36830 );
buf ( n384397 , n36811 );
not ( n36833 , n384397 );
buf ( n384399 , n382924 );
not ( n36835 , n384399 );
or ( n36836 , n36833 , n36835 );
buf ( n384402 , n382921 );
buf ( n384403 , n36822 );
nand ( n36839 , n384402 , n384403 );
buf ( n384405 , n36839 );
buf ( n384406 , n384405 );
nand ( n36842 , n36836 , n384406 );
buf ( n384408 , n36842 );
buf ( n384409 , n384408 );
buf ( n36845 , n36798 );
buf ( n384411 , n36845 );
not ( n36847 , n384411 );
buf ( n384413 , n36847 );
buf ( n384414 , n384413 );
buf ( n36850 , n384414 );
buf ( n384416 , n36850 );
buf ( n384417 , n384416 );
nand ( n36853 , n384409 , n384417 );
buf ( n384419 , n36853 );
buf ( n384420 , n384419 );
nand ( n36856 , n36831 , n384420 );
buf ( n384422 , n36856 );
buf ( n384423 , n384422 );
and ( n36859 , n36740 , n384423 );
and ( n36860 , n384056 , n384304 );
or ( n36861 , n36859 , n36860 );
buf ( n384427 , n36861 );
xor ( n36863 , n36456 , n384427 );
buf ( n384429 , n383409 );
not ( n36865 , n384429 );
buf ( n384431 , n383429 );
not ( n36867 , n384431 );
buf ( n384433 , n36069 );
not ( n36869 , n384433 );
or ( n36870 , n36867 , n36869 );
buf ( n384436 , n36068 );
buf ( n384437 , n383445 );
nand ( n36873 , n384436 , n384437 );
buf ( n384439 , n36873 );
buf ( n384440 , n384439 );
nand ( n36876 , n36870 , n384440 );
buf ( n384442 , n36876 );
buf ( n384443 , n384442 );
not ( n36879 , n384443 );
or ( n36880 , n36865 , n36879 );
buf ( n384446 , n383429 );
not ( n36882 , n384446 );
buf ( n384448 , n36053 );
buf ( n384449 , n34646 );
nand ( n36885 , n384448 , n384449 );
buf ( n384451 , n36885 );
buf ( n384452 , n384451 );
not ( n36888 , n384452 );
buf ( n384454 , n36888 );
not ( n36890 , n384454 );
not ( n36891 , n382864 );
or ( n36892 , n36890 , n36891 );
buf ( n384458 , n35272 );
buf ( n384459 , n384451 );
nand ( n36895 , n384458 , n384459 );
buf ( n384461 , n36895 );
nand ( n36897 , n36892 , n384461 );
not ( n36898 , n36897 );
buf ( n36899 , n36898 );
buf ( n36900 , n36899 );
buf ( n384466 , n36900 );
not ( n36902 , n384466 );
or ( n36903 , n36882 , n36902 );
buf ( n384469 , n36900 );
not ( n36905 , n384469 );
buf ( n384471 , n36905 );
buf ( n384472 , n384471 );
buf ( n384473 , n383445 );
nand ( n36909 , n384472 , n384473 );
buf ( n384475 , n36909 );
buf ( n384476 , n384475 );
nand ( n36912 , n36903 , n384476 );
buf ( n384478 , n36912 );
buf ( n384479 , n384478 );
buf ( n384480 , n383482 );
nand ( n36916 , n384479 , n384480 );
buf ( n384482 , n36916 );
buf ( n384483 , n384482 );
nand ( n36919 , n36880 , n384483 );
buf ( n384485 , n36919 );
buf ( n384486 , n384485 );
buf ( n384487 , n384369 );
not ( n36923 , n384487 );
buf ( n384489 , n384408 );
not ( n36925 , n384489 );
or ( n36926 , n36923 , n36925 );
buf ( n384492 , n36811 );
not ( n36928 , n384492 );
buf ( n384494 , n383059 );
not ( n36930 , n384494 );
or ( n36931 , n36928 , n36930 );
buf ( n384497 , n384037 );
buf ( n384498 , n36822 );
nand ( n36934 , n384497 , n384498 );
buf ( n384500 , n36934 );
buf ( n384501 , n384500 );
nand ( n36937 , n36931 , n384501 );
buf ( n384503 , n36937 );
buf ( n384504 , n384503 );
buf ( n384505 , n384416 );
nand ( n36941 , n384504 , n384505 );
buf ( n384507 , n36941 );
buf ( n384508 , n384507 );
nand ( n36944 , n36926 , n384508 );
buf ( n384510 , n36944 );
buf ( n384511 , n384510 );
xor ( n36947 , n384486 , n384511 );
buf ( n384513 , n36787 );
nor ( n36949 , n384328 , n36771 );
nand ( n36950 , n36949 , n383957 );
not ( n36951 , n36950 );
or ( n36952 , n384343 , n384328 );
buf ( n36953 , n379287 );
nand ( n36954 , n36952 , n36953 );
buf ( n384520 , n379294 );
buf ( n384521 , n379267 );
buf ( n384522 , n379274 );
nand ( n36958 , n384521 , n384522 );
buf ( n384524 , n36958 );
buf ( n384525 , n384524 );
nand ( n36961 , n384520 , n384525 );
buf ( n384527 , n36961 );
nor ( n36963 , n36954 , n384527 );
not ( n36964 , n36963 );
or ( n36965 , n36951 , n36964 );
not ( n36966 , n36954 );
not ( n36967 , n36966 );
buf ( n384533 , n384527 );
not ( n36969 , n384533 );
buf ( n384535 , n36969 );
not ( n36971 , n384535 );
and ( n36972 , n36967 , n36971 );
not ( n36973 , n36949 );
nor ( n36974 , n36973 , n384535 );
and ( n36975 , n383957 , n36974 );
nor ( n36976 , n36972 , n36975 );
nand ( n36977 , n36965 , n36976 );
buf ( n384543 , n36977 );
xnor ( n36979 , n384513 , n384543 );
buf ( n384545 , n36979 );
buf ( n384546 , n384545 );
not ( n36982 , n384546 );
buf ( n384548 , n36982 );
buf ( n384549 , n384548 );
not ( n36985 , n384549 );
buf ( n384551 , n36985 );
buf ( n384552 , n384551 );
not ( n36988 , n384552 );
buf ( n384554 , n36988 );
buf ( n384555 , n384554 );
buf ( n36991 , n384555 );
buf ( n384557 , n36991 );
buf ( n384558 , n384557 );
not ( n36994 , n384558 );
buf ( n384560 , n35797 );
buf ( n36996 , n384560 );
buf ( n384562 , n36996 );
buf ( n384563 , n384562 );
buf ( n36999 , n384563 );
buf ( n384565 , n36999 );
buf ( n384566 , n384565 );
not ( n37002 , n384566 );
buf ( n384568 , n37002 );
buf ( n384569 , n384568 );
not ( n37005 , n384569 );
buf ( n384571 , n384381 );
not ( n37007 , n384571 );
or ( n37008 , n37005 , n37007 );
buf ( n384574 , n382893 );
buf ( n384575 , n384568 );
not ( n37011 , n384575 );
buf ( n384577 , n37011 );
buf ( n384578 , n384577 );
nand ( n37014 , n384574 , n384578 );
buf ( n384580 , n37014 );
buf ( n384581 , n384580 );
nand ( n37017 , n37008 , n384581 );
buf ( n384583 , n37017 );
buf ( n384584 , n384583 );
not ( n37020 , n384584 );
or ( n37021 , n36994 , n37020 );
buf ( n384587 , n384568 );
not ( n37023 , n384587 );
buf ( n384589 , n383578 );
not ( n37025 , n384589 );
or ( n37026 , n37023 , n37025 );
not ( n37027 , n35997 );
buf ( n384593 , n37027 );
not ( n37029 , n384593 );
buf ( n384595 , n384577 );
nand ( n37031 , n37029 , n384595 );
buf ( n384597 , n37031 );
buf ( n384598 , n384597 );
nand ( n37034 , n37026 , n384598 );
buf ( n384600 , n37034 );
buf ( n384601 , n384600 );
not ( n37037 , n35797 );
buf ( n384603 , n37037 );
buf ( n384604 , n36977 );
buf ( n37040 , n384604 );
buf ( n384606 , n37040 );
buf ( n384607 , n384606 );
nand ( n37043 , n384603 , n384607 );
buf ( n384609 , n37043 );
buf ( n384610 , n384609 );
buf ( n384611 , n384545 );
buf ( n384612 , n384606 );
not ( n37048 , n384612 );
buf ( n384614 , n37048 );
nand ( n37050 , n384614 , n35797 );
buf ( n384616 , n37050 );
nand ( n37052 , n384610 , n384611 , n384616 );
buf ( n384618 , n37052 );
buf ( n384619 , n384618 );
buf ( n37055 , n384619 );
buf ( n384621 , n37055 );
buf ( n384622 , n384621 );
not ( n37058 , n384622 );
buf ( n384624 , n37058 );
buf ( n384625 , n384624 );
buf ( n37061 , n384625 );
buf ( n384627 , n37061 );
buf ( n384628 , n384627 );
nand ( n37064 , n384601 , n384628 );
buf ( n384630 , n37064 );
buf ( n384631 , n384630 );
nand ( n37067 , n37021 , n384631 );
buf ( n384633 , n37067 );
buf ( n384634 , n384633 );
xnor ( n37070 , n36947 , n384634 );
buf ( n384636 , n37070 );
buf ( n384637 , n384636 );
not ( n37073 , n384637 );
buf ( n384639 , n37073 );
xor ( n37075 , n36863 , n384639 );
buf ( n384641 , n37075 );
buf ( n384642 , n383910 );
not ( n37078 , n384642 );
buf ( n384644 , n37078 );
buf ( n384645 , n384644 );
not ( n37081 , n384645 );
buf ( n384647 , n36253 );
not ( n37083 , n384647 );
buf ( n384649 , n382535 );
not ( n37085 , n384649 );
or ( n37086 , n37083 , n37085 );
buf ( n384652 , n382532 );
buf ( n384653 , n36252 );
nand ( n37089 , n384652 , n384653 );
buf ( n384655 , n37089 );
buf ( n384656 , n384655 );
nand ( n37092 , n37086 , n384656 );
buf ( n384658 , n37092 );
buf ( n384659 , n384658 );
not ( n37095 , n384659 );
or ( n37096 , n37081 , n37095 );
buf ( n384662 , n383900 );
not ( n37098 , n384662 );
buf ( n384664 , n36253 );
not ( n37100 , n384664 );
buf ( n384666 , n383114 );
not ( n37102 , n384666 );
or ( n37103 , n37100 , n37102 );
buf ( n384669 , n383111 );
buf ( n384670 , n36252 );
nand ( n37106 , n384669 , n384670 );
buf ( n384672 , n37106 );
buf ( n384673 , n384672 );
nand ( n37109 , n37103 , n384673 );
buf ( n384675 , n37109 );
buf ( n384676 , n384675 );
nand ( n37112 , n37098 , n384676 );
buf ( n384678 , n37112 );
buf ( n384679 , n384678 );
nand ( n37115 , n37096 , n384679 );
buf ( n384681 , n37115 );
buf ( n384682 , n384681 );
buf ( n384683 , n383409 );
not ( n37119 , n384683 );
buf ( n384685 , n383429 );
not ( n37121 , n384685 );
buf ( n384687 , n33241 );
buf ( n37123 , n384687 );
buf ( n384689 , n37123 );
not ( n37125 , n384689 );
not ( n37126 , n34504 );
or ( n37127 , n37125 , n37126 );
buf ( n384693 , n34625 );
buf ( n37129 , n384693 );
buf ( n384695 , n37129 );
nand ( n37131 , n37127 , n384695 );
buf ( n37132 , n34633 );
nand ( n37133 , n37131 , n37132 );
buf ( n384699 , n34605 );
buf ( n384700 , n33407 );
or ( n37136 , n384699 , n384700 );
buf ( n384702 , n37136 );
buf ( n37138 , n34627 );
nand ( n37139 , n37138 , n34636 );
and ( n37140 , n37139 , n34628 );
nand ( n37141 , n37133 , n384702 , n37140 );
or ( n37142 , n37133 , n37139 );
nor ( n37143 , n384702 , n37139 );
not ( n37144 , n37143 );
or ( n37145 , n37139 , n34628 );
nand ( n37146 , n37141 , n37142 , n37144 , n37145 );
buf ( n37147 , n37146 );
buf ( n384713 , n37147 );
buf ( n37149 , n384713 );
buf ( n384715 , n37149 );
buf ( n384716 , n384715 );
not ( n37152 , n384716 );
or ( n37153 , n37121 , n37152 );
buf ( n384719 , n384715 );
not ( n37155 , n384719 );
buf ( n384721 , n37155 );
buf ( n384722 , n384721 );
buf ( n384723 , n383445 );
nand ( n37159 , n384722 , n384723 );
buf ( n384725 , n37159 );
buf ( n384726 , n384725 );
nand ( n37162 , n37153 , n384726 );
buf ( n384728 , n37162 );
buf ( n384729 , n384728 );
not ( n37165 , n384729 );
or ( n37166 , n37119 , n37165 );
and ( n37167 , n37132 , n34628 );
not ( n37168 , n384689 );
not ( n37169 , n34606 );
or ( n37170 , n37168 , n37169 );
nand ( n37171 , n37170 , n384695 );
xor ( n37172 , n37167 , n37171 );
buf ( n37173 , n37172 );
buf ( n384739 , n37173 );
buf ( n37175 , n384739 );
buf ( n384741 , n37175 );
buf ( n384742 , n384741 );
not ( n37178 , n384742 );
buf ( n384744 , n37178 );
nand ( n37180 , n384744 , n383429 );
nand ( n37181 , n384741 , n383445 );
nand ( n37182 , n37180 , n37181 );
buf ( n384748 , n37182 );
buf ( n384749 , n383482 );
nand ( n37185 , n384748 , n384749 );
buf ( n384751 , n37185 );
buf ( n384752 , n384751 );
nand ( n37188 , n37166 , n384752 );
buf ( n384754 , n37188 );
buf ( n384755 , n384754 );
xor ( n37191 , n384682 , n384755 );
buf ( n384757 , n379466 );
not ( n37193 , n384757 );
buf ( n384759 , n31964 );
not ( n37195 , n384759 );
buf ( n384761 , n383762 );
not ( n37197 , n384761 );
or ( n37198 , n37195 , n37197 );
buf ( n384764 , n383765 );
buf ( n384765 , n379574 );
nand ( n37201 , n384764 , n384765 );
buf ( n384767 , n37201 );
buf ( n384768 , n384767 );
nand ( n37204 , n37198 , n384768 );
buf ( n384770 , n37204 );
buf ( n384771 , n384770 );
not ( n37207 , n384771 );
or ( n37208 , n37193 , n37207 );
buf ( n384774 , n31964 );
not ( n37210 , n384774 );
not ( n37211 , n36221 );
buf ( n384777 , n37211 );
not ( n37213 , n384777 );
or ( n37214 , n37210 , n37213 );
not ( n37215 , n36216 );
not ( n37216 , n37215 );
buf ( n384782 , n37216 );
buf ( n384783 , n379574 );
nand ( n37219 , n384782 , n384783 );
buf ( n384785 , n37219 );
buf ( n384786 , n384785 );
nand ( n37222 , n37214 , n384786 );
buf ( n384788 , n37222 );
buf ( n384789 , n384788 );
buf ( n384790 , n382601 );
nand ( n37226 , n384789 , n384790 );
buf ( n384792 , n37226 );
buf ( n384793 , n384792 );
nand ( n37229 , n37208 , n384793 );
buf ( n384795 , n37229 );
buf ( n384796 , n384795 );
and ( n37232 , n37191 , n384796 );
and ( n37233 , n384682 , n384755 );
or ( n37234 , n37232 , n37233 );
buf ( n384800 , n37234 );
buf ( n384801 , n384800 );
xnor ( n37242 , n382857 , n36672 );
buf ( n384803 , n37242 );
buf ( n384804 , n382950 );
nand ( n37245 , n384803 , n384804 );
buf ( n384806 , n37245 );
buf ( n384807 , n384806 );
nand ( n37248 , C1 , n384807 );
buf ( n384809 , n37248 );
buf ( n384810 , n384809 );
buf ( n384811 , n384644 );
not ( n37252 , n384811 );
buf ( n384813 , n36258 );
not ( n37254 , n384813 );
or ( n37255 , n37252 , n37254 );
buf ( n384816 , n384658 );
buf ( n384817 , n383897 );
nand ( n37258 , n384816 , n384817 );
buf ( n384819 , n37258 );
buf ( n384820 , n384819 );
nand ( n37261 , n37255 , n384820 );
buf ( n384822 , n37261 );
buf ( n384823 , n384822 );
xor ( n37264 , n384810 , n384823 );
buf ( n384825 , n383409 );
not ( n37266 , n384825 );
buf ( n384827 , n384478 );
not ( n37268 , n384827 );
or ( n37269 , n37266 , n37268 );
buf ( n384830 , n384728 );
buf ( n384831 , n383482 );
nand ( n37272 , n384830 , n384831 );
buf ( n384833 , n37272 );
buf ( n384834 , n384833 );
nand ( n37275 , n37269 , n384834 );
buf ( n384836 , n37275 );
buf ( n384837 , n384836 );
xor ( n37278 , n37264 , n384837 );
buf ( n384839 , n37278 );
buf ( n384840 , n384839 );
xor ( n37281 , n384801 , n384840 );
not ( n37282 , n23528 );
not ( n37283 , n37282 );
not ( n37284 , n37283 );
buf ( n384845 , n379218 );
buf ( n384846 , n379231 );
or ( n37287 , n384845 , n384846 );
buf ( n384848 , n37287 );
buf ( n384849 , n384848 );
not ( n37290 , n384849 );
buf ( n384851 , n37290 );
not ( n37292 , n384851 );
not ( n37293 , n37292 );
nand ( n37294 , n371131 , n371077 );
not ( n37295 , n37294 );
not ( n37296 , n37295 );
or ( n37297 , n37293 , n37296 );
not ( n37298 , n384851 );
not ( n37299 , n371081 );
and ( n37300 , n37298 , n37299 );
not ( n37301 , n371081 );
nor ( n37302 , n37301 , n384848 );
and ( n37303 , n37294 , n37302 );
nor ( n37304 , n37300 , n37303 );
nand ( n37305 , n37297 , n37304 );
buf ( n384866 , n37305 );
not ( n37307 , n384866 );
buf ( n384868 , n37307 );
not ( n37309 , n384868 );
not ( n37310 , n37309 );
or ( n37311 , n37284 , n37310 );
nand ( n37312 , n384868 , n37282 );
nand ( n37313 , n37311 , n37312 );
not ( n37314 , n37313 );
not ( n37315 , n37314 );
not ( n37316 , n37315 );
not ( n37317 , n37316 );
buf ( n384878 , n37317 );
not ( n37319 , n384878 );
buf ( n384880 , n36296 );
not ( n37321 , n384880 );
buf ( n384882 , n36298 );
not ( n37323 , n384882 );
or ( n37324 , n37321 , n37323 );
buf ( n384885 , n36303 );
nand ( n37326 , n37324 , n384885 );
buf ( n384887 , n37326 );
buf ( n384888 , n384887 );
buf ( n384889 , n37305 );
nand ( n37330 , n384888 , n384889 );
buf ( n384891 , n37330 );
not ( n37332 , n384891 );
nor ( n37333 , n36304 , n37305 );
nor ( n37334 , n37332 , n37333 );
or ( n37335 , n384868 , n37282 );
nand ( n37336 , n37335 , n37312 );
nand ( n37337 , n37334 , n37336 );
not ( n37338 , n37337 );
buf ( n384899 , n37338 );
not ( n37340 , n384899 );
buf ( n384901 , n37340 );
buf ( n384902 , n384901 );
not ( n37343 , n384902 );
or ( n37344 , n37319 , n37343 );
not ( n37345 , n36304 );
buf ( n37346 , n37345 );
not ( n37347 , n37346 );
buf ( n384908 , n37347 );
not ( n37349 , n384908 );
buf ( n384910 , n34863 );
not ( n37351 , n384910 );
or ( n37352 , n37349 , n37351 );
buf ( n384913 , n34862 );
not ( n37354 , n37347 );
buf ( n384915 , n37354 );
nand ( n37356 , n384913 , n384915 );
buf ( n384917 , n37356 );
buf ( n384918 , n384917 );
nand ( n37359 , n37352 , n384918 );
buf ( n384920 , n37359 );
buf ( n384921 , n384920 );
nand ( n37362 , n37344 , n384921 );
buf ( n384923 , n37362 );
buf ( n384924 , n384923 );
buf ( n384925 , n384557 );
not ( n37366 , n384925 );
and ( n37367 , n384568 , n36069 );
not ( n37368 , n384568 );
not ( n37369 , n36066 );
not ( n37370 , n37369 );
and ( n37371 , n37368 , n37370 );
or ( n37372 , n37367 , n37371 );
buf ( n384933 , n37372 );
not ( n37374 , n384933 );
or ( n37375 , n37366 , n37374 );
buf ( n384936 , n384568 );
not ( n37377 , n384936 );
buf ( n384938 , n36900 );
not ( n37379 , n384938 );
or ( n37380 , n37377 , n37379 );
not ( n37381 , n36899 );
buf ( n384942 , n37381 );
buf ( n384943 , n384565 );
nand ( n37384 , n384942 , n384943 );
buf ( n384945 , n37384 );
buf ( n384946 , n384945 );
nand ( n37387 , n37380 , n384946 );
buf ( n384948 , n37387 );
buf ( n384949 , n384948 );
buf ( n384950 , n384627 );
nand ( n37391 , n384949 , n384950 );
buf ( n384952 , n37391 );
buf ( n384953 , n384952 );
nand ( n37394 , n37375 , n384953 );
buf ( n384955 , n37394 );
buf ( n384956 , n384955 );
xor ( n37397 , n384924 , n384956 );
not ( n37398 , n36583 );
buf ( n384959 , n37398 );
buf ( n384960 , n383017 );
not ( n37401 , n384960 );
not ( n37402 , n35435 );
buf ( n384963 , n37402 );
not ( n37404 , n384963 );
buf ( n384965 , n37404 );
buf ( n384966 , n384965 );
not ( n37407 , n384966 );
buf ( n384968 , n384280 );
not ( n37409 , n384968 );
or ( n37410 , n37407 , n37409 );
not ( n37411 , n36708 );
buf ( n384972 , n37411 );
buf ( n37413 , n384972 );
buf ( n384974 , n37413 );
buf ( n384975 , n384974 );
buf ( n384976 , n383024 );
nand ( n37417 , n384975 , n384976 );
buf ( n384978 , n37417 );
buf ( n384979 , n384978 );
nand ( n37420 , n37410 , n384979 );
buf ( n384981 , n37420 );
buf ( n384982 , n384981 );
not ( n37423 , n384982 );
or ( n37424 , n37401 , n37423 );
buf ( n384985 , n384251 );
buf ( n384986 , n383137 );
nand ( n37427 , n384985 , n384986 );
buf ( n384988 , n37427 );
buf ( n384989 , n384988 );
nand ( n37430 , n37424 , n384989 );
buf ( n384991 , n37430 );
buf ( n384992 , n384991 );
xor ( n37433 , n384959 , n384992 );
buf ( n384994 , n379466 );
not ( n37435 , n384994 );
buf ( n384996 , n384788 );
not ( n37437 , n384996 );
or ( n37438 , n37435 , n37437 );
buf ( n384999 , n31964 );
buf ( n385000 , n384189 );
and ( n37441 , n384999 , n385000 );
not ( n37442 , n384999 );
buf ( n385003 , n384211 );
and ( n37444 , n37442 , n385003 );
nor ( n37445 , n37441 , n37444 );
buf ( n385006 , n37445 );
buf ( n385007 , n385006 );
buf ( n385008 , n382601 );
nand ( n37449 , n385007 , n385008 );
buf ( n385010 , n37449 );
buf ( n385011 , n385010 );
nand ( n37452 , n37438 , n385011 );
buf ( n385013 , n37452 );
buf ( n385014 , n385013 );
and ( n37455 , n37433 , n385014 );
and ( n37456 , n384959 , n384992 );
or ( n37457 , n37455 , n37456 );
buf ( n385018 , n37457 );
buf ( n385019 , n385018 );
and ( n37460 , n37397 , n385019 );
and ( n37461 , n384924 , n384956 );
or ( n37462 , n37460 , n37461 );
buf ( n385023 , n37462 );
buf ( n385024 , n385023 );
and ( n37465 , n37281 , n385024 );
and ( n37466 , n384801 , n384840 );
or ( n37467 , n37465 , n37466 );
buf ( n385028 , n37467 );
buf ( n385029 , n385028 );
not ( n37470 , n36223 );
not ( n37471 , n383200 );
and ( n37472 , n37470 , n37471 );
not ( n37473 , n383182 );
and ( n37474 , n36648 , n37473 );
nor ( n37475 , n37472 , n37474 );
buf ( n385036 , n37475 );
buf ( n385037 , n382601 );
not ( n37478 , n385037 );
buf ( n385039 , n384770 );
not ( n37480 , n385039 );
or ( n37481 , n37478 , n37480 );
buf ( n385042 , n31964 );
not ( n37483 , n385042 );
buf ( n385044 , n384744 );
not ( n37485 , n385044 );
or ( n37486 , n37483 , n37485 );
buf ( n385047 , n384741 );
buf ( n385048 , n379574 );
nand ( n37489 , n385047 , n385048 );
buf ( n385050 , n37489 );
buf ( n385051 , n385050 );
nand ( n37492 , n37486 , n385051 );
buf ( n385053 , n37492 );
buf ( n385054 , n385053 );
buf ( n385055 , n379466 );
nand ( n37496 , n385054 , n385055 );
buf ( n385057 , n37496 );
buf ( n385058 , n385057 );
nand ( n37499 , n37481 , n385058 );
buf ( n385060 , n37499 );
buf ( n385061 , n385060 );
xor ( n37502 , n385036 , n385061 );
buf ( n385063 , n384557 );
not ( n37504 , n385063 );
buf ( n385065 , n384600 );
not ( n37506 , n385065 );
or ( n37507 , n37504 , n37506 );
buf ( n385068 , n37372 );
buf ( n385069 , n384627 );
nand ( n37510 , n385068 , n385069 );
buf ( n385071 , n37510 );
buf ( n385072 , n385071 );
nand ( n37513 , n37507 , n385072 );
buf ( n385074 , n37513 );
buf ( n385075 , n385074 );
and ( n37516 , n37502 , n385075 );
and ( n37517 , n385036 , n385061 );
or ( n37518 , n37516 , n37517 );
buf ( n385079 , n37518 );
xor ( n37520 , n384810 , n384823 );
and ( n37521 , n37520 , n384837 );
and ( n37522 , n384810 , n384823 );
or ( n37523 , n37521 , n37522 );
buf ( n385084 , n37523 );
xor ( n37525 , n385079 , n385084 );
buf ( n385086 , n379466 );
not ( n37527 , n385086 );
buf ( n385088 , n31964 );
not ( n37529 , n385088 );
buf ( n385090 , n384715 );
not ( n37531 , n385090 );
or ( n37532 , n37529 , n37531 );
buf ( n385093 , n384721 );
buf ( n385094 , n379574 );
nand ( n37535 , n385093 , n385094 );
buf ( n385096 , n37535 );
buf ( n385097 , n385096 );
nand ( n37538 , n37532 , n385097 );
buf ( n385099 , n37538 );
buf ( n385100 , n385099 );
not ( n37541 , n385100 );
or ( n37542 , n37527 , n37541 );
buf ( n385103 , n385053 );
buf ( n385104 , n382601 );
nand ( n37545 , n385103 , n385104 );
buf ( n385106 , n37545 );
buf ( n385107 , n385106 );
nand ( n37548 , n37542 , n385107 );
buf ( n385109 , n37548 );
buf ( n385110 , n385109 );
buf ( n385111 , n37475 );
not ( n37552 , n385111 );
buf ( n385113 , n37552 );
buf ( n385114 , n385113 );
xor ( n37555 , n385110 , n385114 );
buf ( n385116 , n384192 );
buf ( n37557 , n385116 );
buf ( n385118 , n37557 );
not ( n37559 , n385118 );
xor ( n37560 , n382857 , n37559 );
not ( n37561 , n37560 );
not ( n37562 , n382950 );
or ( n37563 , n37561 , n37562 );
buf ( n385124 , C1 );
nand ( n37568 , n37563 , n385124 );
buf ( n385126 , n37568 );
xor ( n37570 , n37555 , n385126 );
buf ( n385128 , n37570 );
xor ( n37572 , n37525 , n385128 );
not ( n37573 , n37572 );
buf ( n385131 , n37573 );
and ( n37575 , n385029 , n385131 );
not ( n37576 , n385029 );
buf ( n385134 , n37572 );
and ( n37578 , n37576 , n385134 );
nor ( n37579 , n37575 , n37578 );
buf ( n385137 , n37579 );
buf ( n385138 , n385137 );
not ( n37582 , n385138 );
xor ( n37583 , n385036 , n385061 );
xor ( n37584 , n37583 , n385075 );
buf ( n385142 , n37584 );
buf ( n385143 , n385142 );
xor ( n37587 , n384056 , n384304 );
xor ( n37588 , n37587 , n384423 );
buf ( n385146 , n37588 );
buf ( n385147 , n385146 );
xor ( n37591 , n385143 , n385147 );
buf ( n385149 , n384416 );
not ( n37593 , n385149 );
buf ( n385151 , n384393 );
not ( n37595 , n385151 );
or ( n37596 , n37593 , n37595 );
not ( n37597 , n36811 );
not ( n37598 , n37597 );
not ( n37599 , n383584 );
or ( n37600 , n37598 , n37599 );
nand ( n37601 , n37027 , n36811 );
nand ( n37602 , n37600 , n37601 );
nand ( n37603 , n37602 , n384369 );
buf ( n385161 , n37603 );
nand ( n37605 , n37596 , n385161 );
buf ( n385163 , n37605 );
buf ( n385164 , n385163 );
buf ( n385165 , n384011 );
not ( n37609 , n385165 );
buf ( n385167 , n36399 );
not ( n37611 , n385167 );
buf ( n385169 , n382924 );
not ( n37613 , n385169 );
or ( n37614 , n37611 , n37613 );
buf ( n385172 , n382921 );
buf ( n385173 , n36468 );
nand ( n37617 , n385172 , n385173 );
buf ( n385175 , n37617 );
buf ( n385176 , n385175 );
nand ( n37620 , n37614 , n385176 );
buf ( n385178 , n37620 );
buf ( n385179 , n385178 );
not ( n37623 , n385179 );
or ( n37624 , n37609 , n37623 );
buf ( n385182 , n384045 );
buf ( n385183 , n383946 );
nand ( n37627 , n385182 , n385183 );
buf ( n385185 , n37627 );
buf ( n385186 , n385185 );
nand ( n37630 , n37624 , n385186 );
buf ( n385188 , n37630 );
buf ( n385189 , n385188 );
xor ( n37633 , n385164 , n385189 );
xor ( n37634 , n384152 , n384258 );
xor ( n37635 , n37634 , n384298 );
buf ( n385193 , n37635 );
buf ( n385194 , n385193 );
and ( n37638 , n37633 , n385194 );
and ( n37639 , n385164 , n385189 );
or ( n37640 , n37638 , n37639 );
buf ( n385198 , n37640 );
buf ( n385199 , n385198 );
and ( n37643 , n37591 , n385199 );
and ( n37644 , n385143 , n385147 );
or ( n37645 , n37643 , n37644 );
buf ( n385203 , n37645 );
buf ( n385204 , n385203 );
not ( n37648 , n385204 );
and ( n37649 , n37582 , n37648 );
buf ( n385207 , n385203 );
buf ( n385208 , n385137 );
and ( n37652 , n385207 , n385208 );
nor ( n37653 , n37649 , n37652 );
buf ( n385211 , n37653 );
buf ( n385212 , n385211 );
xor ( n37656 , n384641 , n385212 );
not ( n37657 , n384627 );
buf ( n385215 , n384565 );
buf ( n385216 , n384715 );
and ( n37660 , n385215 , n385216 );
not ( n37661 , n385215 );
buf ( n385219 , n384721 );
and ( n37663 , n37661 , n385219 );
nor ( n37664 , n37660 , n37663 );
buf ( n385222 , n37664 );
not ( n37666 , n385222 );
or ( n37667 , n37657 , n37666 );
buf ( n385225 , n384557 );
not ( n37669 , n385225 );
buf ( n385227 , n37669 );
not ( n37671 , n385227 );
nand ( n37672 , n37671 , n384948 );
nand ( n37673 , n37667 , n37672 );
buf ( n385231 , n37673 );
buf ( n385232 , n383482 );
not ( n37676 , n385232 );
and ( n37677 , n383429 , n383762 );
not ( n37678 , n383429 );
buf ( n37679 , n36186 );
not ( n37680 , n37679 );
and ( n37681 , n37678 , n37680 );
or ( n37682 , n37677 , n37681 );
buf ( n385240 , n37682 );
not ( n37684 , n385240 );
or ( n37685 , n37676 , n37684 );
buf ( n385243 , n37182 );
buf ( n385244 , n383409 );
nand ( n37688 , n385243 , n385244 );
buf ( n385246 , n37688 );
buf ( n385247 , n385246 );
nand ( n37691 , n37685 , n385247 );
buf ( n385249 , n37691 );
buf ( n385250 , n385249 );
xor ( n37694 , n385231 , n385250 );
not ( n37695 , n37317 );
buf ( n385253 , n37695 );
not ( n37697 , n385253 );
buf ( n385255 , n384920 );
not ( n37699 , n385255 );
or ( n37700 , n37697 , n37699 );
buf ( n385258 , n37347 );
buf ( n385259 , n383975 );
and ( n37703 , n385258 , n385259 );
not ( n37704 , n385258 );
buf ( n385262 , n382548 );
and ( n37706 , n37704 , n385262 );
nor ( n37707 , n37703 , n37706 );
buf ( n385265 , n37707 );
buf ( n385266 , n385265 );
buf ( n385267 , n384901 );
not ( n37711 , n385267 );
buf ( n385269 , n37711 );
buf ( n385270 , n385269 );
nand ( n37714 , n385266 , n385270 );
buf ( n385272 , n37714 );
buf ( n385273 , n385272 );
nand ( n37717 , n37700 , n385273 );
buf ( n385275 , n37717 );
buf ( n385276 , n385275 );
and ( n37720 , n37694 , n385276 );
and ( n37721 , n385231 , n385250 );
or ( n37722 , n37720 , n37721 );
buf ( n385280 , n37722 );
buf ( n385281 , n385280 );
xor ( n37725 , n384682 , n384755 );
xor ( n37726 , n37725 , n384796 );
buf ( n385284 , n37726 );
buf ( n385285 , n385284 );
xor ( n37729 , n385281 , n385285 );
not ( n37730 , n382947 );
not ( n37731 , n384149 );
or ( n37732 , n37730 , n37731 );
buf ( n385290 , n384143 );
not ( n37739 , n385290 );
buf ( n385292 , n37739 );
buf ( n385293 , n385292 );
not ( n37742 , n385293 );
not ( n37743 , n376674 );
nand ( n37744 , n28786 , n376670 );
not ( n37745 , n37744 );
or ( n37746 , n37743 , n37745 );
buf ( n385299 , n384115 );
buf ( n385300 , n382139 );
buf ( n385301 , n382148 );
or ( n37750 , n385300 , n385301 );
buf ( n385303 , n37750 );
buf ( n385304 , n385303 );
nand ( n37753 , n385299 , n385304 );
buf ( n385306 , n37753 );
nand ( n37755 , n37746 , n385306 );
not ( n37756 , n376670 );
not ( n37757 , n28786 );
or ( n37758 , n37756 , n37757 );
not ( n37759 , n376674 );
nor ( n37760 , n37759 , n385306 );
nand ( n37761 , n37758 , n37760 );
nand ( n37762 , n37755 , n37761 );
buf ( n37763 , n37762 );
buf ( n385316 , n37763 );
not ( n37765 , n385316 );
buf ( n385318 , n37765 );
buf ( n385319 , n385318 );
not ( n37768 , n385319 );
or ( n37769 , n37742 , n37768 );
buf ( n385322 , n37763 );
buf ( n37771 , n385322 );
buf ( n385324 , n37771 );
buf ( n385325 , n385324 );
buf ( n385326 , n35262 );
buf ( n37775 , n385326 );
buf ( n385328 , n37775 );
buf ( n385329 , n385328 );
not ( n37778 , n385329 );
buf ( n385331 , n37778 );
buf ( n385332 , n385331 );
nand ( n37781 , n385325 , n385332 );
buf ( n385334 , n37781 );
buf ( n385335 , n385334 );
nand ( n37784 , n37769 , n385335 );
buf ( n385337 , n37784 );
buf ( n385338 , C1 );
nand ( n37789 , n37732 , n385338 );
buf ( n385340 , n29077 );
buf ( n37791 , n385340 );
buf ( n385342 , n37791 );
buf ( n385343 , n385342 );
not ( n37794 , n385343 );
buf ( n385345 , n37794 );
buf ( n385346 , n385345 );
not ( n37797 , n385346 );
buf ( n385348 , n37797 );
buf ( n385349 , n385348 );
not ( n37800 , n385349 );
buf ( n385351 , n384143 );
not ( n37802 , n385351 );
and ( n37803 , n37800 , n37802 );
buf ( n385354 , n29077 );
not ( n37805 , n385354 );
buf ( n385356 , n37805 );
buf ( n385357 , n385356 );
not ( n37808 , n385357 );
buf ( n385359 , n37808 );
buf ( n385360 , n385359 );
buf ( n385361 , n384096 );
and ( n37812 , n385360 , n385361 );
nor ( n37813 , n37803 , n37812 );
buf ( n385364 , n37813 );
buf ( n385365 , n382947 );
buf ( n385366 , n385337 );
nand ( n37823 , n385365 , n385366 );
buf ( n385368 , n37823 );
nand ( n37825 , C1 , n385368 );
xor ( n37826 , n37789 , n37825 );
not ( n37827 , n384981 );
not ( n37828 , n383137 );
or ( n37829 , n37827 , n37828 );
buf ( n385374 , n383017 );
buf ( n385375 , n384965 );
not ( n37832 , n385375 );
buf ( n385377 , n384083 );
not ( n37834 , n385377 );
or ( n37835 , n37832 , n37834 );
buf ( n385380 , n36509 );
buf ( n385381 , n383024 );
nand ( n37838 , n385380 , n385381 );
buf ( n385383 , n37838 );
buf ( n385384 , n385383 );
nand ( n37841 , n37835 , n385384 );
buf ( n385386 , n37841 );
buf ( n385387 , n385386 );
nand ( n37844 , n385374 , n385387 );
buf ( n385389 , n37844 );
nand ( n37846 , n37829 , n385389 );
and ( n37847 , n37826 , n37846 );
and ( n37848 , n37789 , n37825 );
or ( n37849 , n37847 , n37848 );
not ( n37850 , n384416 );
not ( n37851 , n37602 );
or ( n385396 , n37850 , n37851 );
buf ( n385397 , n36811 );
not ( n37854 , n385397 );
buf ( n385399 , n36069 );
not ( n37856 , n385399 );
or ( n37857 , n37854 , n37856 );
buf ( n385402 , n37370 );
buf ( n385403 , n36822 );
nand ( n37860 , n385402 , n385403 );
buf ( n385405 , n37860 );
buf ( n385406 , n385405 );
nand ( n37863 , n37857 , n385406 );
buf ( n385408 , n37863 );
buf ( n385409 , n385408 );
buf ( n385410 , n384369 );
nand ( n37867 , n385409 , n385410 );
buf ( n385412 , n37867 );
nand ( n37869 , n385396 , n385412 );
xor ( n37870 , n37849 , n37869 );
not ( n37871 , n383897 );
buf ( n385416 , n36253 );
not ( n37873 , n385416 );
buf ( n385418 , n383059 );
not ( n37875 , n385418 );
or ( n37876 , n37873 , n37875 );
buf ( n385421 , n384037 );
buf ( n385422 , n36252 );
nand ( n37879 , n385421 , n385422 );
buf ( n385424 , n37879 );
buf ( n385425 , n385424 );
nand ( n37882 , n37876 , n385425 );
buf ( n385427 , n37882 );
not ( n37884 , n385427 );
or ( n37885 , n37871 , n37884 );
buf ( n385430 , n384675 );
buf ( n385431 , n384644 );
nand ( n37888 , n385430 , n385431 );
buf ( n385433 , n37888 );
nand ( n37890 , n37885 , n385433 );
and ( n37891 , n37870 , n37890 );
and ( n37892 , n37849 , n37869 );
or ( n37893 , n37891 , n37892 );
buf ( n385438 , n37893 );
and ( n37895 , n37729 , n385438 );
and ( n37896 , n385281 , n385285 );
or ( n37897 , n37895 , n37896 );
buf ( n385442 , n37897 );
buf ( n385443 , n385442 );
xor ( n37900 , n384801 , n384840 );
xor ( n37901 , n37900 , n385024 );
buf ( n385446 , n37901 );
buf ( n385447 , n385446 );
xor ( n37904 , n385443 , n385447 );
xor ( n37905 , n384924 , n384956 );
xor ( n37906 , n37905 , n385019 );
buf ( n385451 , n37906 );
buf ( n385452 , n385451 );
xor ( n37909 , n384959 , n384992 );
xor ( n37910 , n37909 , n385014 );
buf ( n385455 , n37910 );
buf ( n385456 , n385455 );
buf ( n37913 , n22981 );
or ( n37914 , n24029 , n37913 );
and ( n37915 , n24024 , n371623 );
not ( n37916 , n24024 );
not ( n37917 , n371623 );
and ( n37918 , n37916 , n37917 );
nor ( n37919 , n37915 , n37918 );
nand ( n37920 , n37919 , n37913 );
nand ( n37921 , n37914 , n37920 );
not ( n37922 , n37921 );
buf ( n37923 , n37922 );
buf ( n37924 , n37923 );
buf ( n385469 , n37924 );
not ( n37926 , n385469 );
buf ( n385471 , n23528 );
buf ( n37928 , n385471 );
buf ( n385473 , n37928 );
nand ( n37930 , n24030 , n385473 );
nand ( n37931 , n37919 , n37282 );
nand ( n37932 , n37930 , n37922 , n37931 );
buf ( n385477 , n37932 );
not ( n37934 , n385477 );
buf ( n385479 , n37934 );
buf ( n385480 , n385479 );
not ( n37937 , n385480 );
buf ( n385482 , n37937 );
buf ( n385483 , n385482 );
not ( n37940 , n385483 );
or ( n37941 , n37926 , n37940 );
buf ( n385486 , n385473 );
not ( n37943 , n385486 );
buf ( n385488 , n37943 );
buf ( n385489 , n385488 );
buf ( n37946 , n385489 );
buf ( n385491 , n37946 );
buf ( n385492 , n385491 );
not ( n37949 , n385492 );
buf ( n385494 , n37949 );
buf ( n385495 , n385494 );
not ( n37952 , n385495 );
buf ( n385497 , n34858 );
buf ( n37954 , n385497 );
buf ( n385499 , n37954 );
buf ( n385500 , n385499 );
not ( n37957 , n385500 );
buf ( n385502 , n37957 );
buf ( n385503 , n385502 );
not ( n37960 , n385503 );
or ( n37961 , n37952 , n37960 );
buf ( n385506 , n34860 );
buf ( n385507 , n385491 );
nand ( n37964 , n385506 , n385507 );
buf ( n385509 , n37964 );
buf ( n385510 , n385509 );
nand ( n37967 , n37961 , n385510 );
buf ( n385512 , n37967 );
buf ( n385513 , n385512 );
nand ( n37970 , n37941 , n385513 );
buf ( n385515 , n37970 );
not ( n37972 , n385006 );
not ( n37973 , n379466 );
or ( n37974 , n37972 , n37973 );
buf ( n385519 , n31964 );
not ( n37976 , n385519 );
buf ( n385521 , n36672 );
not ( n37978 , n385521 );
or ( n37979 , n37976 , n37978 );
buf ( n385524 , n36676 );
buf ( n385525 , n379574 );
nand ( n37982 , n385524 , n385525 );
buf ( n385527 , n37982 );
buf ( n385528 , n385527 );
nand ( n37985 , n37979 , n385528 );
buf ( n385530 , n37985 );
buf ( n385531 , n385530 );
buf ( n385532 , n382601 );
nand ( n37989 , n385531 , n385532 );
buf ( n385534 , n37989 );
nand ( n37991 , n37974 , n385534 );
xor ( n37992 , n385515 , n37991 );
buf ( n385537 , n384557 );
not ( n37994 , n385537 );
buf ( n385539 , n385222 );
not ( n37996 , n385539 );
or ( n37997 , n37994 , n37996 );
buf ( n385542 , n384568 );
buf ( n385543 , n384741 );
and ( n38000 , n385542 , n385543 );
not ( n38001 , n385542 );
buf ( n385546 , n384744 );
and ( n38003 , n38001 , n385546 );
nor ( n38004 , n38000 , n38003 );
buf ( n385549 , n38004 );
buf ( n385550 , n385549 );
buf ( n385551 , n384627 );
nand ( n38008 , n385550 , n385551 );
buf ( n385553 , n38008 );
buf ( n385554 , n385553 );
nand ( n38011 , n37997 , n385554 );
buf ( n385556 , n38011 );
and ( n38013 , n37992 , n385556 );
and ( n38014 , n385515 , n37991 );
or ( n38015 , n38013 , n38014 );
buf ( n385560 , n38015 );
xor ( n38017 , n385456 , n385560 );
not ( n38018 , n36399 );
not ( n38019 , n384381 );
or ( n38020 , n38018 , n38019 );
buf ( n385565 , n382893 );
buf ( n385566 , n36398 );
nand ( n38023 , n385565 , n385566 );
buf ( n385568 , n38023 );
nand ( n38025 , n38020 , n385568 );
not ( n38026 , n38025 );
not ( n38027 , n384011 );
or ( n38028 , n38026 , n38027 );
buf ( n385573 , n385178 );
buf ( n385574 , n383946 );
nand ( n38031 , n385573 , n385574 );
buf ( n385576 , n38031 );
nand ( n38033 , n38028 , n385576 );
buf ( n385578 , n38033 );
and ( n38035 , n38017 , n385578 );
and ( n38036 , n385456 , n385560 );
or ( n38037 , n38035 , n38036 );
buf ( n385582 , n38037 );
buf ( n385583 , n385582 );
xor ( n38040 , n385452 , n385583 );
xor ( n38041 , n385164 , n385189 );
xor ( n38042 , n38041 , n385194 );
buf ( n385587 , n38042 );
buf ( n385588 , n385587 );
and ( n38045 , n38040 , n385588 );
and ( n38046 , n385452 , n385583 );
or ( n38047 , n38045 , n38046 );
buf ( n385592 , n38047 );
buf ( n385593 , n385592 );
and ( n38050 , n37904 , n385593 );
and ( n38051 , n385443 , n385447 );
or ( n38052 , n38050 , n38051 );
buf ( n385597 , n38052 );
buf ( n385598 , n385597 );
not ( n38055 , n385598 );
buf ( n385600 , n38055 );
buf ( n385601 , n385600 );
xor ( n38058 , n37656 , n385601 );
buf ( n385603 , n38058 );
buf ( n385604 , n385603 );
xor ( n38061 , n385443 , n385447 );
xor ( n38062 , n38061 , n385593 );
buf ( n385607 , n38062 );
xor ( n38064 , n385143 , n385147 );
xor ( n38065 , n38064 , n385199 );
buf ( n385610 , n38065 );
nor ( n38067 , n385607 , n385610 );
not ( n38068 , n38067 );
xor ( n38069 , n385281 , n385285 );
xor ( n38070 , n38069 , n385438 );
buf ( n385615 , n38070 );
buf ( n385616 , n385615 );
buf ( n385617 , n383409 );
not ( n38074 , n385617 );
buf ( n385619 , n37682 );
not ( n38076 , n385619 );
or ( n38077 , n38074 , n38076 );
buf ( n385622 , n383429 );
not ( n38079 , n385622 );
buf ( n385624 , n36218 );
not ( n38081 , n385624 );
or ( n38082 , n38079 , n38081 );
buf ( n385627 , n36221 );
buf ( n385628 , n383460 );
not ( n38085 , n385628 );
buf ( n385630 , n38085 );
buf ( n385631 , n385630 );
not ( n38088 , n385631 );
buf ( n385633 , n38088 );
buf ( n385634 , n385633 );
nand ( n38091 , n385627 , n385634 );
buf ( n385636 , n38091 );
buf ( n385637 , n385636 );
nand ( n38094 , n38082 , n385637 );
buf ( n385639 , n38094 );
buf ( n385640 , n385639 );
buf ( n385641 , n383482 );
nand ( n38098 , n385640 , n385641 );
buf ( n385643 , n38098 );
buf ( n385644 , n385643 );
nand ( n38101 , n38077 , n385644 );
buf ( n385646 , n38101 );
buf ( n385647 , n385646 );
buf ( n385648 , n37695 );
not ( n38105 , n385648 );
buf ( n385650 , n385265 );
not ( n38107 , n385650 );
or ( n38108 , n38105 , n38107 );
buf ( n385653 , n37347 );
buf ( n385654 , n383111 );
and ( n38111 , n385653 , n385654 );
not ( n38112 , n385653 );
buf ( n385657 , n383108 );
and ( n38114 , n38112 , n385657 );
nor ( n38115 , n38111 , n38114 );
buf ( n385660 , n38115 );
buf ( n385661 , n385660 );
buf ( n385662 , n385269 );
nand ( n38119 , n385661 , n385662 );
buf ( n385664 , n38119 );
buf ( n385665 , n385664 );
nand ( n38122 , n38108 , n385665 );
buf ( n385667 , n38122 );
buf ( n385668 , n385667 );
xor ( n38125 , n385647 , n385668 );
xor ( n38126 , n37789 , n37825 );
xor ( n38127 , n38126 , n37846 );
buf ( n385672 , n38127 );
and ( n38129 , n38125 , n385672 );
and ( n38130 , n385647 , n385668 );
or ( n38131 , n38129 , n38130 );
buf ( n385676 , n38131 );
buf ( n385677 , n385676 );
xor ( n38134 , n385231 , n385250 );
xor ( n38135 , n38134 , n385276 );
buf ( n385680 , n38135 );
buf ( n385681 , n385680 );
xor ( n38138 , n385677 , n385681 );
xor ( n38139 , n37849 , n37869 );
xor ( n38140 , n38139 , n37890 );
buf ( n385685 , n38140 );
and ( n38142 , n38138 , n385685 );
and ( n38143 , n385677 , n385681 );
or ( n38144 , n38142 , n38143 );
buf ( n385689 , n38144 );
buf ( n385690 , n385689 );
xor ( n38147 , n385616 , n385690 );
buf ( n385692 , n37825 );
not ( n38149 , n385692 );
buf ( n385694 , n38149 );
buf ( n385695 , n385694 );
buf ( n385696 , n383027 );
nand ( n38153 , n36546 , n36555 );
nand ( n38154 , n36562 , n38153 );
buf ( n38155 , n38154 );
buf ( n385700 , n38155 );
and ( n38157 , n385696 , n385700 );
not ( n38158 , n385696 );
not ( n38159 , n38155 );
buf ( n385704 , n38159 );
and ( n38161 , n38158 , n385704 );
nor ( n38162 , n38157 , n38161 );
buf ( n385707 , n38162 );
buf ( n385708 , n385707 );
not ( n38165 , n385708 );
buf ( n385710 , n383017 );
not ( n38167 , n385710 );
or ( n38168 , n38165 , n38167 );
buf ( n385713 , n385386 );
buf ( n385714 , n383137 );
nand ( n38171 , n385713 , n385714 );
buf ( n385716 , n38171 );
buf ( n385717 , n385716 );
nand ( n38174 , n38168 , n385717 );
buf ( n385719 , n38174 );
buf ( n385720 , n385719 );
xor ( n38177 , n385695 , n385720 );
buf ( n385722 , n383409 );
not ( n38179 , n385722 );
buf ( n385724 , n385639 );
not ( n38181 , n385724 );
or ( n38182 , n38179 , n38181 );
buf ( n385727 , n385633 );
not ( n38184 , n385727 );
buf ( n385729 , n38184 );
buf ( n385730 , n385729 );
not ( n38187 , n385730 );
buf ( n385732 , n384202 );
buf ( n38189 , n385732 );
buf ( n385734 , n38189 );
buf ( n385735 , n385734 );
not ( n38192 , n385735 );
or ( n38193 , n38187 , n38192 );
buf ( n385738 , n385734 );
not ( n38195 , n385738 );
buf ( n385740 , n38195 );
buf ( n385741 , n385740 );
buf ( n385742 , n385633 );
nand ( n38199 , n385741 , n385742 );
buf ( n385744 , n38199 );
buf ( n385745 , n385744 );
nand ( n38202 , n38193 , n385745 );
buf ( n385747 , n38202 );
buf ( n385748 , n385747 );
buf ( n385749 , n383479 );
not ( n38206 , n385749 );
buf ( n385751 , n38206 );
buf ( n385752 , n385751 );
nand ( n38209 , n385748 , n385752 );
buf ( n385754 , n38209 );
buf ( n385755 , n385754 );
nand ( n38212 , n38182 , n385755 );
buf ( n385757 , n38212 );
buf ( n385758 , n385757 );
and ( n38215 , n38177 , n385758 );
and ( n38216 , n385695 , n385720 );
or ( n38217 , n38215 , n38216 );
buf ( n385762 , n38217 );
buf ( n385763 , n385762 );
buf ( n385764 , n384416 );
not ( n38221 , n385764 );
buf ( n385766 , n385408 );
not ( n38223 , n385766 );
or ( n38224 , n38221 , n38223 );
buf ( n385769 , n36811 );
not ( n38226 , n385769 );
not ( n38227 , n36898 );
buf ( n385772 , n38227 );
not ( n38229 , n385772 );
buf ( n385774 , n38229 );
buf ( n385775 , n385774 );
not ( n38232 , n385775 );
or ( n38233 , n38226 , n38232 );
buf ( n385778 , n37381 );
buf ( n385779 , n36822 );
nand ( n38236 , n385778 , n385779 );
buf ( n385781 , n38236 );
buf ( n385782 , n385781 );
nand ( n38239 , n38233 , n385782 );
buf ( n385784 , n38239 );
buf ( n385785 , n385784 );
buf ( n385786 , n384369 );
nand ( n38243 , n385785 , n385786 );
buf ( n385788 , n38243 );
buf ( n385789 , n385788 );
nand ( n38246 , n38224 , n385789 );
buf ( n385791 , n38246 );
buf ( n385792 , n385791 );
xor ( n38249 , n385763 , n385792 );
buf ( n385794 , n383897 );
not ( n38251 , n385794 );
buf ( n385796 , n36253 );
not ( n38253 , n385796 );
buf ( n385798 , n382924 );
not ( n38255 , n385798 );
or ( n38256 , n38253 , n38255 );
buf ( n385801 , n382921 );
buf ( n385802 , n36252 );
nand ( n38259 , n385801 , n385802 );
buf ( n385804 , n38259 );
buf ( n385805 , n385804 );
nand ( n38262 , n38256 , n385805 );
buf ( n385807 , n38262 );
buf ( n385808 , n385807 );
not ( n38265 , n385808 );
or ( n38266 , n38251 , n38265 );
buf ( n385811 , n385427 );
buf ( n385812 , n384644 );
nand ( n38269 , n385811 , n385812 );
buf ( n385814 , n38269 );
buf ( n385815 , n385814 );
nand ( n38272 , n38266 , n385815 );
buf ( n385817 , n38272 );
buf ( n385818 , n385817 );
and ( n38275 , n38249 , n385818 );
and ( n38276 , n385763 , n385792 );
or ( n38277 , n38275 , n38276 );
buf ( n385822 , n38277 );
buf ( n385823 , n385822 );
not ( n38280 , n383946 );
not ( n38281 , n38025 );
or ( n38282 , n38280 , n38281 );
buf ( n385827 , n36399 );
not ( n38284 , n385827 );
buf ( n385829 , n37027 );
not ( n38286 , n385829 );
or ( n38287 , n38284 , n38286 );
buf ( n385832 , n383575 );
not ( n38289 , n385832 );
buf ( n385834 , n38289 );
buf ( n385835 , n385834 );
buf ( n385836 , n36468 );
nand ( n38293 , n385835 , n385836 );
buf ( n385838 , n38293 );
buf ( n385839 , n385838 );
nand ( n38296 , n38287 , n385839 );
buf ( n385841 , n38296 );
buf ( n385842 , n385841 );
buf ( n385843 , n384011 );
nand ( n38300 , n385842 , n385843 );
buf ( n385845 , n38300 );
nand ( n38302 , n38282 , n385845 );
buf ( n385847 , n38302 );
buf ( n385848 , n382601 );
not ( n38305 , n385848 );
buf ( n385850 , n384974 );
not ( n38307 , n385850 );
buf ( n385852 , n38307 );
and ( n38309 , n31964 , n385852 );
not ( n38310 , n31964 );
and ( n38311 , n38310 , n384974 );
or ( n38312 , n38309 , n38311 );
buf ( n385857 , n38312 );
not ( n38314 , n385857 );
or ( n38315 , n38305 , n38314 );
buf ( n385860 , n385530 );
buf ( n385861 , n379466 );
nand ( n38318 , n385860 , n385861 );
buf ( n385863 , n38318 );
buf ( n385864 , n385863 );
nand ( n38321 , n38315 , n385864 );
buf ( n385866 , n38321 );
buf ( n385867 , n385866 );
not ( n38324 , n37924 );
buf ( n385869 , n38324 );
not ( n38326 , n385869 );
buf ( n385871 , n385512 );
not ( n38328 , n385871 );
or ( n38329 , n38326 , n38328 );
buf ( n385874 , n385494 );
not ( n38331 , n385874 );
buf ( n385876 , n382535 );
not ( n38333 , n385876 );
or ( n38334 , n38331 , n38333 );
buf ( n385879 , n382532 );
buf ( n385880 , n385491 );
nand ( n38337 , n385879 , n385880 );
buf ( n385882 , n38337 );
buf ( n385883 , n385882 );
nand ( n38340 , n38334 , n385883 );
buf ( n385885 , n38340 );
buf ( n385886 , n385885 );
buf ( n385887 , n385482 );
not ( n38344 , n385887 );
buf ( n385889 , n38344 );
buf ( n385890 , n385889 );
nand ( n38347 , n385886 , n385890 );
buf ( n385892 , n38347 );
buf ( n385893 , n385892 );
nand ( n38350 , n38329 , n385893 );
buf ( n385895 , n38350 );
buf ( n385896 , n385895 );
xor ( n38353 , n385867 , n385896 );
buf ( n385898 , n384369 );
not ( n38355 , n385898 );
buf ( n38356 , n37146 );
buf ( n38357 , n38356 );
and ( n38358 , n36821 , n38357 );
not ( n38359 , n36821 );
and ( n38360 , n38359 , n384721 );
or ( n38361 , n38358 , n38360 );
buf ( n385906 , n38361 );
not ( n38363 , n385906 );
or ( n38364 , n38355 , n38363 );
buf ( n385909 , n385784 );
buf ( n385910 , n384416 );
nand ( n38367 , n385909 , n385910 );
buf ( n385912 , n38367 );
buf ( n385913 , n385912 );
nand ( n38370 , n38364 , n385913 );
buf ( n385915 , n38370 );
buf ( n385916 , n385915 );
and ( n38373 , n38353 , n385916 );
and ( n38374 , n385867 , n385896 );
or ( n38375 , n38373 , n38374 );
buf ( n385920 , n38375 );
buf ( n385921 , n385920 );
xor ( n38378 , n385847 , n385921 );
xor ( n38379 , n385515 , n37991 );
xor ( n38380 , n38379 , n385556 );
buf ( n385925 , n38380 );
and ( n38382 , n38378 , n385925 );
and ( n38383 , n385847 , n385921 );
or ( n38384 , n38382 , n38383 );
buf ( n385929 , n38384 );
buf ( n385930 , n385929 );
xor ( n38387 , n385823 , n385930 );
xor ( n38388 , n385456 , n385560 );
xor ( n38389 , n38388 , n385578 );
buf ( n385934 , n38389 );
buf ( n385935 , n385934 );
and ( n38392 , n38387 , n385935 );
and ( n38393 , n385823 , n385930 );
or ( n38394 , n38392 , n38393 );
buf ( n385939 , n38394 );
buf ( n385940 , n385939 );
and ( n38397 , n38147 , n385940 );
and ( n38398 , n385616 , n385690 );
or ( n38399 , n38397 , n38398 );
buf ( n385944 , n38399 );
buf ( n385945 , n385944 );
not ( n38402 , n385945 );
buf ( n385947 , n38402 );
not ( n38404 , n385947 );
and ( n38405 , n38068 , n38404 );
buf ( n385950 , n385610 );
buf ( n385951 , n385607 );
and ( n38408 , n385950 , n385951 );
buf ( n385953 , n38408 );
nor ( n38410 , n38405 , n385953 );
buf ( n385955 , n38410 );
nand ( n38412 , n385604 , n385955 );
buf ( n385957 , n38412 );
buf ( n385958 , n385957 );
not ( n38415 , n385958 );
xor ( n38416 , n385763 , n385792 );
xor ( n38417 , n38416 , n385818 );
buf ( n385962 , n38417 );
buf ( n385963 , n385962 );
buf ( n385964 , n379466 );
not ( n38421 , n385964 );
buf ( n385966 , n38312 );
not ( n38423 , n385966 );
or ( n38424 , n38421 , n38423 );
not ( n38425 , n31962 );
buf ( n385970 , n38425 );
not ( n38427 , n385970 );
buf ( n385972 , n38427 );
buf ( n385973 , n385972 );
not ( n38430 , n385973 );
buf ( n385975 , n38430 );
buf ( n385976 , n385975 );
not ( n38433 , n385976 );
buf ( n385978 , n384089 );
not ( n38435 , n385978 );
or ( n38436 , n38433 , n38435 );
buf ( n385981 , n36509 );
buf ( n38438 , n385981 );
buf ( n385983 , n38438 );
buf ( n385984 , n385983 );
buf ( n385985 , n382570 );
buf ( n38442 , n385985 );
buf ( n385987 , n38442 );
buf ( n385988 , n385987 );
nand ( n38445 , n385984 , n385988 );
buf ( n385990 , n38445 );
buf ( n385991 , n385990 );
nand ( n38448 , n38436 , n385991 );
buf ( n385993 , n38448 );
buf ( n385994 , n385993 );
buf ( n385995 , n382598 );
nand ( n38452 , n385994 , n385995 );
buf ( n385997 , n38452 );
buf ( n385998 , n385997 );
nand ( n38455 , n38424 , n385998 );
buf ( n386000 , n38455 );
buf ( n386001 , n386000 );
buf ( n386002 , n383409 );
not ( n38459 , n386002 );
buf ( n386004 , n385747 );
not ( n38461 , n386004 );
or ( n38462 , n38459 , n38461 );
buf ( n386007 , n385751 );
buf ( n386008 , n383429 );
not ( n38465 , n386008 );
buf ( n386010 , n384239 );
buf ( n38467 , n386010 );
buf ( n386012 , n38467 );
buf ( n386013 , n386012 );
not ( n38470 , n386013 );
or ( n38471 , n38465 , n38470 );
not ( n38472 , n384239 );
buf ( n386017 , n38472 );
buf ( n386018 , n385633 );
nand ( n38475 , n386017 , n386018 );
buf ( n386020 , n38475 );
buf ( n386021 , n386020 );
nand ( n38478 , n38471 , n386021 );
buf ( n386023 , n38478 );
buf ( n386024 , n386023 );
nand ( n38481 , n386007 , n386024 );
buf ( n386026 , n38481 );
buf ( n386027 , n386026 );
nand ( n38484 , n38462 , n386027 );
buf ( n386029 , n38484 );
buf ( n386030 , n386029 );
xor ( n38487 , n386001 , n386030 );
buf ( n386032 , n384416 );
not ( n38489 , n386032 );
buf ( n386034 , n38361 );
not ( n38491 , n386034 );
or ( n38492 , n38489 , n38491 );
buf ( n386037 , n36821 );
not ( n38494 , n386037 );
buf ( n386039 , n384744 );
not ( n38496 , n386039 );
or ( n38497 , n38494 , n38496 );
nand ( n38498 , n37597 , n384741 );
buf ( n386043 , n38498 );
nand ( n38500 , n38497 , n386043 );
buf ( n386045 , n38500 );
buf ( n386046 , n386045 );
buf ( n386047 , n384369 );
nand ( n38504 , n386046 , n386047 );
buf ( n386049 , n38504 );
buf ( n386050 , n386049 );
nand ( n38507 , n38492 , n386050 );
buf ( n386052 , n38507 );
buf ( n386053 , n386052 );
and ( n38510 , n38487 , n386053 );
and ( n38511 , n386001 , n386030 );
or ( n38512 , n38510 , n38511 );
buf ( n386057 , n38512 );
buf ( n386058 , n386057 );
not ( n38515 , n386058 );
xor ( n38516 , n385867 , n385896 );
xor ( n38517 , n38516 , n385916 );
buf ( n386062 , n38517 );
buf ( n386063 , n386062 );
not ( n38520 , n386063 );
or ( n38521 , n38515 , n38520 );
buf ( n386066 , n386062 );
buf ( n386067 , n386057 );
or ( n38524 , n386066 , n386067 );
buf ( n386069 , n38324 );
not ( n38526 , n386069 );
buf ( n386071 , n385885 );
not ( n38528 , n386071 );
or ( n38529 , n38526 , n38528 );
buf ( n386074 , n385494 );
not ( n38531 , n386074 );
not ( n38532 , n35519 );
buf ( n386077 , n38532 );
not ( n38534 , n386077 );
or ( n38535 , n38531 , n38534 );
buf ( n386080 , n383111 );
buf ( n386081 , n385491 );
nand ( n386082 , n386080 , n386081 );
buf ( n386083 , n386082 );
buf ( n386084 , n386083 );
nand ( n38541 , n38535 , n386084 );
buf ( n386086 , n38541 );
buf ( n386087 , n386086 );
buf ( n386088 , n385889 );
nand ( n38545 , n386087 , n386088 );
buf ( n386090 , n38545 );
buf ( n386091 , n386090 );
nand ( n38548 , n38529 , n386091 );
buf ( n386093 , n38548 );
buf ( n386094 , n386093 );
not ( n38551 , n386094 );
buf ( n386096 , n384568 );
not ( n38553 , n386096 );
buf ( n386098 , n383762 );
not ( n38555 , n386098 );
or ( n38556 , n38553 , n38555 );
buf ( n386101 , n383765 );
buf ( n386102 , n384565 );
nand ( n38559 , n386101 , n386102 );
buf ( n386104 , n38559 );
buf ( n386105 , n386104 );
nand ( n38562 , n38556 , n386105 );
buf ( n386107 , n38562 );
buf ( n386108 , n386107 );
buf ( n386109 , n384557 );
and ( n38566 , n386108 , n386109 );
buf ( n386111 , n384568 );
not ( n38568 , n386111 );
buf ( n386113 , n36218 );
not ( n38570 , n386113 );
or ( n38571 , n38568 , n38570 );
buf ( n386116 , n37216 );
buf ( n386117 , n384565 );
nand ( n38574 , n386116 , n386117 );
buf ( n386119 , n38574 );
buf ( n386120 , n386119 );
nand ( n38577 , n38571 , n386120 );
buf ( n386122 , n38577 );
buf ( n386123 , n386122 );
not ( n38580 , n386123 );
buf ( n386125 , n384627 );
not ( n38582 , n386125 );
buf ( n386127 , n38582 );
buf ( n386128 , n386127 );
nor ( n38585 , n38580 , n386128 );
buf ( n386130 , n38585 );
buf ( n386131 , n386130 );
nor ( n38588 , n38566 , n386131 );
buf ( n386133 , n38588 );
buf ( n386134 , n386133 );
not ( n38591 , n386134 );
buf ( n386136 , n38591 );
buf ( n386137 , n386136 );
not ( n38594 , n386137 );
or ( n38595 , n38551 , n38594 );
buf ( n386140 , n386136 );
buf ( n386141 , n386093 );
or ( n38598 , n386140 , n386141 );
buf ( n386143 , n385292 );
not ( n38606 , n386143 );
buf ( n386145 , n375781 );
buf ( n38608 , n386145 );
buf ( n386147 , n38608 );
buf ( n386148 , n386147 );
not ( n38611 , n386148 );
buf ( n386150 , n38611 );
buf ( n386151 , n386150 );
not ( n38614 , n386151 );
and ( n38615 , n38606 , n38614 );
buf ( n386154 , n385292 );
buf ( n386155 , n386150 );
and ( n38618 , n386154 , n386155 );
nor ( n38619 , n38615 , n38618 );
buf ( n386158 , n38619 );
buf ( n386159 , n382938 );
not ( n38625 , n386159 );
buf ( n386161 , n38625 );
buf ( n386162 , n386161 );
buf ( n386163 , n385292 );
not ( n38629 , n386163 );
not ( n38630 , n28159 );
buf ( n38631 , n38630 );
buf ( n386167 , n38631 );
not ( n38633 , n386167 );
and ( n38634 , n38629 , n38633 );
buf ( n386170 , n384096 );
not ( n38636 , n386170 );
buf ( n386172 , n38636 );
buf ( n386173 , n386172 );
buf ( n386174 , n28159 );
not ( n38640 , n386174 );
buf ( n386176 , n38640 );
buf ( n386177 , n386176 );
buf ( n38643 , n386177 );
buf ( n386179 , n38643 );
buf ( n386180 , n386179 );
buf ( n38646 , n386180 );
buf ( n386182 , n38646 );
buf ( n386183 , n386182 );
and ( n38649 , n386173 , n386183 );
nor ( n38650 , n38634 , n38649 );
buf ( n386186 , n38650 );
buf ( n386187 , n386186 );
nor ( n38653 , n386162 , n386187 );
buf ( n386189 , n38653 );
buf ( n386190 , n386189 );
nor ( n38656 , C0 , n386190 );
buf ( n386192 , n38656 );
buf ( n386193 , n386192 );
not ( n38659 , n385975 );
not ( n38660 , n38155 );
not ( n38661 , n38660 );
or ( n38662 , n38659 , n38661 );
buf ( n386198 , n38155 );
buf ( n386199 , n385987 );
nand ( n38665 , n386198 , n386199 );
buf ( n386201 , n38665 );
nand ( n38667 , n38662 , n386201 );
not ( n38668 , n38667 );
not ( n38669 , n382598 );
or ( n38670 , n38668 , n38669 );
buf ( n386206 , n385993 );
buf ( n386207 , n379460 );
not ( n38673 , n386207 );
buf ( n386209 , n38673 );
buf ( n386210 , n386209 );
buf ( n38676 , n386210 );
buf ( n386212 , n38676 );
buf ( n386213 , n386212 );
nand ( n38679 , n386206 , n386213 );
buf ( n386215 , n38679 );
nand ( n38681 , n38670 , n386215 );
buf ( n386217 , n38681 );
xor ( n38683 , n386193 , n386217 );
buf ( n386219 , n383014 );
not ( n38685 , n35377 );
buf ( n386221 , n38685 );
not ( n38687 , n386221 );
buf ( n386223 , n38687 );
buf ( n386224 , n386223 );
buf ( n386225 , n385356 );
and ( n38691 , n386224 , n386225 );
not ( n38692 , n386224 );
buf ( n386228 , n385359 );
and ( n38694 , n38692 , n386228 );
nor ( n38695 , n38691 , n38694 );
buf ( n386231 , n38695 );
buf ( n386232 , n386231 );
or ( n38698 , n386219 , n386232 );
buf ( n386234 , n385324 );
not ( n38700 , n386234 );
buf ( n386236 , n38700 );
buf ( n386237 , n386236 );
buf ( n386238 , n386223 );
and ( n38704 , n386237 , n386238 );
buf ( n386240 , n385324 );
buf ( n386241 , n383024 );
and ( n38707 , n386240 , n386241 );
nor ( n38708 , n38704 , n38707 );
buf ( n386244 , n38708 );
buf ( n386245 , n386244 );
buf ( n386246 , n383134 );
or ( n38712 , n386245 , n386246 );
nand ( n38713 , n38698 , n38712 );
buf ( n386249 , n38713 );
buf ( n386250 , n386249 );
and ( n38716 , n38683 , n386250 );
and ( n38717 , n386193 , n386217 );
or ( n38718 , n38716 , n38717 );
buf ( n386254 , n38718 );
buf ( n386255 , n386254 );
nand ( n38721 , n38598 , n386255 );
buf ( n386257 , n38721 );
buf ( n386258 , n386257 );
nand ( n38724 , n38595 , n386258 );
buf ( n386260 , n38724 );
buf ( n386261 , n386260 );
nand ( n38727 , n38524 , n386261 );
buf ( n386263 , n38727 );
buf ( n386264 , n386263 );
nand ( n38730 , n38521 , n386264 );
buf ( n386266 , n38730 );
buf ( n386267 , n386266 );
xor ( n38733 , n385963 , n386267 );
xor ( n38734 , n385847 , n385921 );
xor ( n38735 , n38734 , n385925 );
buf ( n386271 , n38735 );
buf ( n386272 , n386271 );
xor ( n38738 , n38733 , n386272 );
buf ( n386274 , n38738 );
buf ( n386275 , n386274 );
not ( n38741 , n386275 );
xor ( n38742 , n385647 , n385668 );
xor ( n38743 , n38742 , n385672 );
buf ( n386279 , n38743 );
buf ( n386280 , n386279 );
buf ( n386281 , n382944 );
buf ( n386282 , n385364 );
or ( n38751 , n386281 , n386282 );
nand ( n38752 , C1 , n38751 );
buf ( n386285 , n38752 );
buf ( n386286 , n386285 );
buf ( n386287 , n386192 );
not ( n38756 , n386287 );
buf ( n386289 , n38756 );
buf ( n386290 , n386289 );
xor ( n38759 , n386286 , n386290 );
buf ( n386292 , n386244 );
not ( n38761 , n386292 );
buf ( n386294 , n38761 );
buf ( n386295 , n386294 );
not ( n38764 , n386295 );
not ( n38765 , n35425 );
buf ( n386298 , n38765 );
buf ( n38767 , n386298 );
buf ( n386300 , n38767 );
buf ( n386301 , n386300 );
not ( n38770 , n386301 );
or ( n38771 , n38764 , n38770 );
buf ( n386304 , n385707 );
buf ( n386305 , n383134 );
buf ( n38774 , n386305 );
buf ( n386307 , n38774 );
buf ( n386308 , n386307 );
not ( n38777 , n386308 );
buf ( n386310 , n38777 );
buf ( n386311 , n386310 );
nand ( n38780 , n386304 , n386311 );
buf ( n386313 , n38780 );
buf ( n386314 , n386313 );
nand ( n38783 , n38771 , n386314 );
buf ( n386316 , n38783 );
buf ( n386317 , n386316 );
and ( n38786 , n38759 , n386317 );
and ( n38787 , n386286 , n386290 );
or ( n38788 , n38786 , n38787 );
buf ( n386321 , n38788 );
buf ( n386322 , n386321 );
buf ( n386323 , n384627 );
not ( n38792 , n386323 );
buf ( n386325 , n386107 );
not ( n38794 , n386325 );
or ( n38795 , n38792 , n38794 );
buf ( n386328 , n385549 );
buf ( n386329 , n384557 );
nand ( n38798 , n386328 , n386329 );
buf ( n386331 , n38798 );
buf ( n386332 , n386331 );
nand ( n38801 , n38795 , n386332 );
buf ( n386334 , n38801 );
buf ( n386335 , n386334 );
xor ( n38804 , n386322 , n386335 );
xor ( n38805 , n385695 , n385720 );
xor ( n38806 , n38805 , n385758 );
buf ( n386339 , n38806 );
buf ( n386340 , n386339 );
and ( n38809 , n38804 , n386340 );
and ( n38810 , n386322 , n386335 );
or ( n38811 , n38809 , n38810 );
buf ( n386344 , n38811 );
buf ( n386345 , n386344 );
xor ( n38814 , n386280 , n386345 );
buf ( n386347 , n383946 );
not ( n38816 , n386347 );
buf ( n386349 , n385841 );
not ( n38818 , n386349 );
or ( n38819 , n38816 , n38818 );
buf ( n386352 , n36399 );
not ( n38821 , n386352 );
buf ( n38822 , n36066 );
not ( n38823 , n38822 );
buf ( n386356 , n38823 );
not ( n38825 , n386356 );
or ( n38826 , n38821 , n38825 );
buf ( n386359 , n37370 );
buf ( n386360 , n36398 );
nand ( n38829 , n386359 , n386360 );
buf ( n386362 , n38829 );
buf ( n386363 , n386362 );
nand ( n38832 , n38826 , n386363 );
buf ( n386365 , n38832 );
buf ( n386366 , n386365 );
buf ( n386367 , n384011 );
nand ( n38836 , n386366 , n386367 );
buf ( n386369 , n38836 );
buf ( n386370 , n386369 );
nand ( n38839 , n38819 , n386370 );
buf ( n386372 , n38839 );
buf ( n386373 , n386372 );
not ( n38842 , n386373 );
buf ( n386375 , n38842 );
buf ( n386376 , n386375 );
not ( n38845 , n386376 );
buf ( n386378 , n385807 );
buf ( n386379 , n384644 );
and ( n38848 , n386378 , n386379 );
buf ( n386381 , n36253 );
not ( n38850 , n386381 );
buf ( n386383 , n35301 );
not ( n38852 , n386383 );
buf ( n386385 , n38852 );
buf ( n386386 , n386385 );
not ( n38855 , n386386 );
or ( n38856 , n38850 , n38855 );
buf ( n386389 , n35301 );
not ( n38858 , n386389 );
buf ( n386391 , n38858 );
buf ( n386392 , n386391 );
not ( n38861 , n386392 );
buf ( n386394 , n36252 );
nand ( n38863 , n38861 , n386394 );
buf ( n386396 , n38863 );
buf ( n386397 , n386396 );
nand ( n38866 , n38856 , n386397 );
buf ( n386399 , n38866 );
buf ( n386400 , n386399 );
not ( n38869 , n386400 );
buf ( n386402 , n383900 );
nor ( n38871 , n38869 , n386402 );
buf ( n386404 , n38871 );
buf ( n386405 , n386404 );
nor ( n38874 , n38848 , n386405 );
buf ( n386407 , n38874 );
buf ( n386408 , n386407 );
not ( n38877 , n386408 );
or ( n38878 , n38845 , n38877 );
buf ( n386411 , n37347 );
not ( n38880 , n386411 );
buf ( n386413 , n383059 );
not ( n38882 , n386413 );
or ( n38883 , n38880 , n38882 );
buf ( n386416 , n383053 );
buf ( n38885 , n386416 );
buf ( n386418 , n38885 );
buf ( n386419 , n386418 );
not ( n38888 , n386419 );
buf ( n386421 , n38888 );
buf ( n386422 , n386421 );
buf ( n38891 , n386422 );
buf ( n386424 , n38891 );
buf ( n386425 , n386424 );
not ( n38894 , n386425 );
buf ( n386427 , n37354 );
nand ( n38896 , n38894 , n386427 );
buf ( n386429 , n38896 );
buf ( n386430 , n386429 );
nand ( n38899 , n38883 , n386430 );
buf ( n386432 , n38899 );
buf ( n386433 , n386432 );
buf ( n386434 , n385269 );
and ( n38903 , n386433 , n386434 );
buf ( n386436 , n385660 );
not ( n38905 , n386436 );
buf ( n386438 , n37317 );
nor ( n38907 , n38905 , n386438 );
buf ( n386440 , n38907 );
buf ( n386441 , n386440 );
nor ( n38910 , n38903 , n386441 );
buf ( n386443 , n38910 );
buf ( n386444 , n386443 );
not ( n38913 , n386444 );
buf ( n386446 , n38913 );
buf ( n386447 , n386446 );
nand ( n38916 , n38878 , n386447 );
buf ( n386449 , n38916 );
buf ( n386450 , n386449 );
buf ( n386451 , n386407 );
not ( n38920 , n386451 );
buf ( n386453 , n38920 );
buf ( n386454 , n386453 );
buf ( n386455 , n386372 );
nand ( n38924 , n386454 , n386455 );
buf ( n386457 , n38924 );
buf ( n386458 , n386457 );
nand ( n38927 , n386450 , n386458 );
buf ( n386460 , n38927 );
buf ( n386461 , n386460 );
xor ( n38930 , n38814 , n386461 );
buf ( n386463 , n38930 );
buf ( n386464 , n386463 );
not ( n38933 , n386464 );
not ( n38934 , n23988 );
buf ( n38935 , n24048 );
not ( n38936 , n38935 );
or ( n38937 , n38934 , n38936 );
or ( n38938 , n38935 , n23988 );
nand ( n38939 , n38937 , n38938 );
buf ( n386472 , n38939 );
buf ( n38941 , n386472 );
buf ( n386474 , n38941 );
buf ( n386475 , n386474 );
not ( n38944 , n386475 );
buf ( n386477 , n38944 );
buf ( n386478 , n386477 );
buf ( n38947 , n386478 );
buf ( n386480 , n38947 );
buf ( n386481 , n386480 );
not ( n38950 , n386481 );
buf ( n386483 , n38950 );
buf ( n386484 , n386483 );
not ( n38953 , n386484 );
and ( n38954 , n22981 , n23988 );
not ( n38955 , n22981 );
not ( n38956 , n23988 );
and ( n38957 , n38955 , n38956 );
nor ( n38958 , n38954 , n38957 );
nand ( n38959 , n38958 , n38939 );
buf ( n38960 , n38959 );
not ( n38961 , n38960 );
buf ( n386494 , n38961 );
buf ( n38963 , n386494 );
buf ( n386496 , n38963 );
buf ( n386497 , n386496 );
not ( n38966 , n386497 );
buf ( n386499 , n38966 );
buf ( n386500 , n386499 );
not ( n38969 , n386500 );
or ( n38970 , n38953 , n38969 );
not ( n38971 , n22982 );
not ( n38972 , n38971 );
buf ( n386505 , n38972 );
not ( n38974 , n386505 );
buf ( n386507 , n34861 );
not ( n38976 , n386507 );
or ( n38977 , n38974 , n38976 );
buf ( n386510 , n34860 );
buf ( n386511 , n38971 );
nand ( n38980 , n386510 , n386511 );
buf ( n386513 , n38980 );
buf ( n386514 , n386513 );
nand ( n38983 , n38977 , n386514 );
buf ( n386516 , n38983 );
buf ( n386517 , n386516 );
nand ( n38986 , n38970 , n386517 );
buf ( n386519 , n38986 );
buf ( n386520 , n386519 );
xor ( n38989 , n386286 , n386290 );
xor ( n38990 , n38989 , n386317 );
buf ( n386523 , n38990 );
buf ( n386524 , n386523 );
xor ( n38993 , n386520 , n386524 );
buf ( n386526 , n383946 );
not ( n38995 , n386526 );
buf ( n386528 , n386365 );
not ( n38997 , n386528 );
or ( n38998 , n38995 , n38997 );
buf ( n386531 , n36399 );
buf ( n386532 , n37381 );
and ( n39001 , n386531 , n386532 );
not ( n39002 , n386531 );
buf ( n386535 , n36900 );
and ( n39004 , n39002 , n386535 );
nor ( n39005 , n39001 , n39004 );
buf ( n386538 , n39005 );
buf ( n386539 , n386538 );
buf ( n386540 , n384011 );
nand ( n39009 , n386539 , n386540 );
buf ( n386542 , n39009 );
buf ( n386543 , n386542 );
nand ( n39012 , n38998 , n386543 );
buf ( n386545 , n39012 );
buf ( n386546 , n386545 );
and ( n39015 , n38993 , n386546 );
and ( n39016 , n386520 , n386524 );
or ( n39017 , n39015 , n39016 );
buf ( n386550 , n39017 );
buf ( n386551 , n386550 );
xor ( n39020 , n386322 , n386335 );
xor ( n39021 , n39020 , n386340 );
buf ( n386554 , n39021 );
buf ( n386555 , n386554 );
xor ( n39024 , n386551 , n386555 );
buf ( n386557 , n385269 );
not ( n39026 , n386557 );
buf ( n386559 , n382921 );
not ( n39028 , n386559 );
buf ( n386561 , n39028 );
and ( n39030 , n386561 , n37347 );
not ( n39031 , n386561 );
and ( n39032 , n39031 , n37354 );
or ( n39033 , n39030 , n39032 );
buf ( n386566 , n39033 );
not ( n39035 , n386566 );
or ( n39036 , n39026 , n39035 );
buf ( n386569 , n386432 );
buf ( n386570 , n37695 );
nand ( n39039 , n386569 , n386570 );
buf ( n386572 , n39039 );
buf ( n386573 , n386572 );
nand ( n39042 , n39036 , n386573 );
buf ( n386575 , n39042 );
buf ( n386576 , n386575 );
not ( n39045 , n386576 );
buf ( n386578 , n39045 );
buf ( n386579 , n386578 );
not ( n39048 , n386579 );
not ( n39049 , n383900 );
not ( n39050 , n36252 );
buf ( n39051 , n35997 );
not ( n39052 , n39051 );
or ( n39053 , n39050 , n39052 );
or ( n39054 , n39051 , n36252 );
nand ( n39055 , n39053 , n39054 );
not ( n39056 , n39055 );
not ( n39057 , n39056 );
and ( n39058 , n39049 , n39057 );
and ( n39059 , n386399 , n384644 );
nor ( n39060 , n39058 , n39059 );
buf ( n386593 , n39060 );
not ( n39062 , n386593 );
or ( n39063 , n39048 , n39062 );
xor ( n39064 , n386001 , n386030 );
xor ( n39065 , n39064 , n386053 );
buf ( n386598 , n39065 );
buf ( n386599 , n386598 );
nand ( n39068 , n39063 , n386599 );
buf ( n386601 , n39068 );
buf ( n386602 , n386601 );
not ( n39071 , n39060 );
buf ( n386604 , n39071 );
buf ( n386605 , n386575 );
nand ( n39074 , n386604 , n386605 );
buf ( n386607 , n39074 );
buf ( n386608 , n386607 );
nand ( n39077 , n386602 , n386608 );
buf ( n386610 , n39077 );
buf ( n386611 , n386610 );
and ( n39080 , n39024 , n386611 );
and ( n39081 , n386551 , n386555 );
or ( n39082 , n39080 , n39081 );
buf ( n386615 , n39082 );
buf ( n386616 , n386615 );
not ( n39085 , n386616 );
buf ( n386618 , n39085 );
buf ( n386619 , n386618 );
nand ( n39088 , n38933 , n386619 );
buf ( n386621 , n39088 );
buf ( n386622 , n386621 );
not ( n39091 , n386622 );
or ( n39092 , n38741 , n39091 );
buf ( n386625 , n386463 );
buf ( n386626 , n386615 );
nand ( n39095 , n386625 , n386626 );
buf ( n386628 , n39095 );
buf ( n386629 , n386628 );
nand ( n39098 , n39092 , n386629 );
buf ( n386631 , n39098 );
not ( n39100 , n386631 );
xor ( n39101 , n385677 , n385681 );
xor ( n39102 , n39101 , n385685 );
buf ( n386635 , n39102 );
buf ( n386636 , n386635 );
xor ( n39105 , n386280 , n386345 );
and ( n39106 , n39105 , n386461 );
and ( n39107 , n386280 , n386345 );
or ( n39108 , n39106 , n39107 );
buf ( n386641 , n39108 );
buf ( n386642 , n386641 );
xor ( n39111 , n386636 , n386642 );
xor ( n39112 , n385823 , n385930 );
xor ( n39113 , n39112 , n385935 );
buf ( n386646 , n39113 );
buf ( n386647 , n386646 );
xor ( n39116 , n39111 , n386647 );
buf ( n386649 , n39116 );
not ( n39118 , n386649 );
xor ( n39119 , n385963 , n386267 );
and ( n39120 , n39119 , n386272 );
and ( n39121 , n385963 , n386267 );
or ( n39122 , n39120 , n39121 );
buf ( n386655 , n39122 );
not ( n39124 , n386655 );
nand ( n39125 , n39118 , n39124 );
not ( n39126 , n39125 );
or ( n39127 , n39100 , n39126 );
buf ( n386660 , n386649 );
buf ( n386661 , n386655 );
nand ( n39130 , n386660 , n386661 );
buf ( n386663 , n39130 );
nand ( n39132 , n39127 , n386663 );
not ( n39133 , n39132 );
xor ( n39134 , n385452 , n385583 );
xor ( n39135 , n39134 , n385588 );
buf ( n386668 , n39135 );
xor ( n39137 , n386636 , n386642 );
and ( n39138 , n39137 , n386647 );
and ( n39139 , n386636 , n386642 );
or ( n39140 , n39138 , n39139 );
buf ( n386673 , n39140 );
xor ( n39142 , n386668 , n386673 );
xor ( n39143 , n385616 , n385690 );
xor ( n39144 , n39143 , n385940 );
buf ( n386677 , n39144 );
xor ( n39146 , n39142 , n386677 );
not ( n39147 , n39146 );
nand ( n39148 , n39133 , n39147 );
xor ( n39149 , n386668 , n386673 );
and ( n39150 , n39149 , n386677 );
and ( n39151 , n386668 , n386673 );
or ( n39152 , n39150 , n39151 );
xor ( n39153 , n385950 , n385951 );
buf ( n386686 , n39153 );
buf ( n386687 , n386686 );
buf ( n386688 , n385944 );
and ( n39157 , n386687 , n386688 );
not ( n39158 , n386687 );
buf ( n386691 , n385947 );
and ( n39160 , n39158 , n386691 );
nor ( n39161 , n39157 , n39160 );
buf ( n386694 , n39161 );
nor ( n39163 , n39152 , n386694 );
not ( n39164 , n39163 );
nand ( n39165 , n39148 , n39164 );
buf ( n386698 , n39165 );
nor ( n39167 , n38415 , n386698 );
buf ( n386700 , n39167 );
buf ( n386701 , n386700 );
buf ( n386702 , n385028 );
not ( n39171 , n386702 );
buf ( n386704 , n37573 );
nand ( n39173 , n39171 , n386704 );
buf ( n386706 , n39173 );
buf ( n386707 , n386706 );
not ( n39176 , n386707 );
buf ( n386709 , n385203 );
not ( n39178 , n386709 );
or ( n39179 , n39176 , n39178 );
buf ( n386712 , n37572 );
buf ( n386713 , n385028 );
nand ( n39182 , n386712 , n386713 );
buf ( n386715 , n39182 );
buf ( n386716 , n386715 );
nand ( n39185 , n39179 , n386716 );
buf ( n386718 , n39185 );
buf ( n386719 , n386718 );
not ( n39188 , n382950 );
and ( n39189 , n382857 , n36218 );
not ( n39190 , n382857 );
and ( n39191 , n39190 , n36221 );
or ( n39192 , n39189 , n39191 );
not ( n39193 , n39192 );
or ( n39194 , n39188 , n39193 );
buf ( n386727 , C1 );
nand ( n39211 , n39194 , n386727 );
not ( n39212 , n39211 );
buf ( n386730 , n383409 );
not ( n39214 , n386730 );
buf ( n386732 , n383429 );
not ( n39216 , n386732 );
buf ( n386734 , n383578 );
not ( n386735 , n386734 );
or ( n39219 , n39216 , n386735 );
buf ( n386737 , n383584 );
buf ( n386738 , n383445 );
nand ( n39222 , n386737 , n386738 );
buf ( n386740 , n39222 );
buf ( n386741 , n386740 );
nand ( n39225 , n39219 , n386741 );
buf ( n386743 , n39225 );
buf ( n386744 , n386743 );
not ( n39228 , n386744 );
or ( n39229 , n39214 , n39228 );
buf ( n386747 , n384442 );
buf ( n386748 , n383482 );
nand ( n39232 , n386747 , n386748 );
buf ( n386750 , n39232 );
buf ( n386751 , n386750 );
nand ( n39235 , n39229 , n386751 );
buf ( n386753 , n39235 );
and ( n39237 , n39212 , n386753 );
not ( n39238 , n39212 );
not ( n39239 , n386753 );
and ( n39240 , n39238 , n39239 );
nor ( n39241 , n39237 , n39240 );
buf ( n386759 , n384503 );
buf ( n386760 , n384369 );
and ( n39244 , n386759 , n386760 );
and ( n39245 , n383114 , n36811 );
not ( n39246 , n383114 );
and ( n39247 , n39246 , n36822 );
or ( n39248 , n39245 , n39247 );
buf ( n386766 , n39248 );
not ( n39250 , n386766 );
buf ( n386768 , n384416 );
not ( n39252 , n386768 );
buf ( n386770 , n39252 );
buf ( n386771 , n386770 );
nor ( n39255 , n39250 , n386771 );
buf ( n386773 , n39255 );
buf ( n386774 , n386773 );
nor ( n39258 , n39244 , n386774 );
buf ( n386776 , n39258 );
buf ( n386777 , n386776 );
not ( n39261 , n386777 );
buf ( n386779 , n39261 );
and ( n39263 , n39241 , n386779 );
not ( n39264 , n39241 );
and ( n39265 , n39264 , n386776 );
nor ( n39266 , n39263 , n39265 );
buf ( n386784 , n379466 );
not ( n39268 , n386784 );
buf ( n386786 , n31964 );
not ( n39270 , n386786 );
buf ( n386788 , n36900 );
not ( n39272 , n386788 );
or ( n39273 , n39270 , n39272 );
buf ( n386791 , n384471 );
buf ( n386792 , n379574 );
nand ( n39276 , n386791 , n386792 );
buf ( n386794 , n39276 );
buf ( n386795 , n386794 );
nand ( n39279 , n39273 , n386795 );
buf ( n386797 , n39279 );
buf ( n386798 , n386797 );
not ( n39282 , n386798 );
or ( n39283 , n39268 , n39282 );
buf ( n386801 , n385099 );
buf ( n386802 , n382601 );
nand ( n39286 , n386801 , n386802 );
buf ( n386804 , n39286 );
buf ( n386805 , n386804 );
nand ( n39289 , n39283 , n386805 );
buf ( n386807 , n39289 );
buf ( n386808 , n386807 );
not ( n39292 , n386808 );
buf ( n386810 , n383017 );
not ( n39294 , n386810 );
buf ( n386812 , n383772 );
not ( n39296 , n386812 );
buf ( n386814 , n39296 );
buf ( n386815 , n386814 );
not ( n39299 , n386815 );
or ( n39300 , n39294 , n39299 );
buf ( n386818 , n383027 );
not ( n39302 , n386818 );
buf ( n386820 , n384744 );
not ( n39304 , n386820 );
or ( n39305 , n39302 , n39304 );
buf ( n386823 , n384741 );
buf ( n386824 , n383072 );
nand ( n39308 , n386823 , n386824 );
buf ( n386826 , n39308 );
buf ( n386827 , n386826 );
nand ( n39311 , n39305 , n386827 );
buf ( n386829 , n39311 );
buf ( n386830 , n386829 );
buf ( n386831 , n383137 );
nand ( n39315 , n386830 , n386831 );
buf ( n386833 , n39315 );
buf ( n386834 , n386833 );
nand ( n39318 , n39300 , n386834 );
buf ( n386836 , n39318 );
buf ( n386837 , n386836 );
not ( n39321 , n386837 );
buf ( n386839 , n39321 );
buf ( n386840 , n386839 );
not ( n39324 , n386840 );
or ( n39325 , n39292 , n39324 );
buf ( n386843 , n386807 );
not ( n39327 , n386843 );
buf ( n386845 , n39327 );
buf ( n386846 , n386845 );
buf ( n386847 , n386836 );
nand ( n39331 , n386846 , n386847 );
buf ( n386849 , n39331 );
buf ( n386850 , n386849 );
nand ( n39334 , n39325 , n386850 );
buf ( n386852 , n39334 );
buf ( n386853 , n386852 );
buf ( n386854 , n384011 );
not ( n39338 , n386854 );
buf ( n386856 , n36406 );
not ( n39340 , n386856 );
or ( n39341 , n39338 , n39340 );
not ( n39342 , n36399 );
not ( n39343 , n34863 );
or ( n39344 , n39342 , n39343 );
buf ( n386862 , n34862 );
buf ( n386863 , n36468 );
nand ( n39347 , n386862 , n386863 );
buf ( n386865 , n39347 );
nand ( n39349 , n39344 , n386865 );
buf ( n386867 , n39349 );
buf ( n386868 , n383946 );
nand ( n39352 , n386867 , n386868 );
buf ( n386870 , n39352 );
buf ( n386871 , n386870 );
nand ( n39355 , n39341 , n386871 );
buf ( n386873 , n39355 );
buf ( n386874 , n386873 );
xor ( n39358 , n386853 , n386874 );
buf ( n386876 , n39358 );
xor ( n39360 , n39266 , n386876 );
buf ( n386878 , n384633 );
buf ( n386879 , n384510 );
or ( n39363 , n386878 , n386879 );
buf ( n386881 , n384485 );
nand ( n39365 , n39363 , n386881 );
buf ( n386883 , n39365 );
buf ( n386884 , n386883 );
buf ( n386885 , n384633 );
buf ( n386886 , n384510 );
nand ( n39370 , n386885 , n386886 );
buf ( n386888 , n39370 );
buf ( n386889 , n386888 );
nand ( n39373 , n386884 , n386889 );
buf ( n386891 , n39373 );
xnor ( n39375 , n39360 , n386891 );
buf ( n386893 , n39375 );
not ( n39377 , n386893 );
buf ( n386895 , n39377 );
buf ( n386896 , n386895 );
and ( n39380 , n386719 , n386896 );
not ( n39381 , n386719 );
buf ( n386899 , n39375 );
and ( n39383 , n39381 , n386899 );
nor ( n39384 , n39380 , n39383 );
buf ( n386902 , n39384 );
buf ( n386903 , n386902 );
buf ( n386904 , n36456 );
not ( n39388 , n386904 );
buf ( n386906 , n384636 );
not ( n39390 , n386906 );
or ( n39391 , n39388 , n39390 );
buf ( n386909 , n384427 );
nand ( n39393 , n39391 , n386909 );
buf ( n386911 , n39393 );
buf ( n386912 , n386911 );
nand ( n39396 , n384639 , n36455 );
buf ( n386914 , n39396 );
nand ( n39398 , n386912 , n386914 );
buf ( n386916 , n39398 );
not ( n39400 , n36449 );
not ( n39401 , n36226 );
or ( n39402 , n39400 , n39401 );
nand ( n39403 , n36444 , n36451 );
nand ( n39404 , n39402 , n39403 );
buf ( n386922 , n39404 );
buf ( n386923 , n384557 );
not ( n39407 , n386923 );
buf ( n386925 , n384568 );
not ( n39409 , n386925 );
buf ( n386927 , n382924 );
not ( n39411 , n386927 );
or ( n39412 , n39409 , n39411 );
buf ( n386930 , n382921 );
buf ( n386931 , n384577 );
nand ( n39415 , n386930 , n386931 );
buf ( n386933 , n39415 );
buf ( n386934 , n386933 );
nand ( n39418 , n39412 , n386934 );
buf ( n386936 , n39418 );
buf ( n386937 , n386936 );
not ( n39421 , n386937 );
or ( n39422 , n39407 , n39421 );
buf ( n386940 , n384583 );
buf ( n386941 , n384627 );
nand ( n39425 , n386940 , n386941 );
buf ( n386943 , n39425 );
buf ( n386944 , n386943 );
nand ( n39428 , n39422 , n386944 );
buf ( n386946 , n39428 );
buf ( n386947 , n386946 );
xor ( n39431 , n386922 , n386947 );
xor ( n39432 , n385110 , n385114 );
and ( n39433 , n39432 , n385126 );
and ( n39434 , n385110 , n385114 );
or ( n39435 , n39433 , n39434 );
buf ( n386953 , n39435 );
buf ( n386954 , n386953 );
xor ( n39438 , n39431 , n386954 );
buf ( n386956 , n39438 );
not ( n39440 , n386956 );
xor ( n39441 , n385079 , n385084 );
and ( n39442 , n39441 , n385128 );
and ( n39443 , n385079 , n385084 );
or ( n39444 , n39442 , n39443 );
buf ( n386962 , n39444 );
not ( n39446 , n386962 );
buf ( n386964 , n39446 );
not ( n39448 , n386964 );
or ( n39449 , n39440 , n39448 );
not ( n39450 , n386956 );
nand ( n39451 , n39450 , n39444 );
nand ( n39452 , n39449 , n39451 );
xnor ( n39453 , n386916 , n39452 );
buf ( n386971 , n39453 );
and ( n39455 , n386903 , n386971 );
not ( n39456 , n386903 );
buf ( n386974 , n39453 );
not ( n39458 , n386974 );
buf ( n386976 , n39458 );
buf ( n386977 , n386976 );
and ( n39461 , n39456 , n386977 );
nor ( n39462 , n39455 , n39461 );
buf ( n386980 , n39462 );
buf ( n386981 , n386980 );
xor ( n39465 , n384641 , n385212 );
and ( n39466 , n39465 , n385601 );
and ( n39467 , n384641 , n385212 );
or ( n39468 , n39466 , n39467 );
buf ( n386986 , n39468 );
buf ( n386987 , n386986 );
nand ( n39471 , n386981 , n386987 );
buf ( n386989 , n39471 );
buf ( n386990 , n386989 );
and ( n39474 , n386701 , n386990 );
buf ( n386992 , n39474 );
buf ( n386993 , n386992 );
buf ( n386994 , n379466 );
not ( n39478 , n386994 );
buf ( n386996 , n379577 );
not ( n39480 , n386996 );
buf ( n386998 , n382896 );
not ( n39482 , n386998 );
or ( n39483 , n39480 , n39482 );
buf ( n387001 , n382893 );
buf ( n387002 , n379574 );
nand ( n39486 , n387001 , n387002 );
buf ( n387004 , n39486 );
buf ( n387005 , n387004 );
nand ( n39489 , n39483 , n387005 );
buf ( n387007 , n39489 );
buf ( n387008 , n387007 );
not ( n39492 , n387008 );
or ( n39493 , n39478 , n39492 );
buf ( n387011 , n379577 );
not ( n39495 , n387011 );
buf ( n387013 , n383578 );
not ( n39497 , n387013 );
or ( n39498 , n39495 , n39497 );
buf ( n387016 , n383584 );
buf ( n387017 , n379574 );
nand ( n39501 , n387016 , n387017 );
buf ( n387019 , n39501 );
buf ( n387020 , n387019 );
nand ( n39504 , n39498 , n387020 );
buf ( n387022 , n39504 );
buf ( n387023 , n387022 );
buf ( n387024 , n382607 );
nand ( n39508 , n387023 , n387024 );
buf ( n387026 , n39508 );
buf ( n387027 , n387026 );
nand ( n39511 , n39493 , n387027 );
buf ( n387029 , n39511 );
buf ( n387030 , n387029 );
buf ( n387031 , n386770 );
not ( n39515 , n387031 );
buf ( n387033 , n384369 );
not ( n39517 , n387033 );
buf ( n387035 , n39517 );
buf ( n387036 , n387035 );
not ( n39520 , n387036 );
or ( n39521 , n39515 , n39520 );
buf ( n387039 , n36811 );
not ( n39523 , n387039 );
buf ( n387041 , n34863 );
not ( n39525 , n387041 );
or ( n39526 , n39523 , n39525 );
buf ( n387044 , n34862 );
buf ( n387045 , n36822 );
nand ( n39529 , n387044 , n387045 );
buf ( n387047 , n39529 );
buf ( n387048 , n387047 );
nand ( n39532 , n39526 , n387048 );
buf ( n387050 , n39532 );
buf ( n387051 , n387050 );
nand ( n39535 , n39521 , n387051 );
buf ( n387053 , n39535 );
buf ( n387054 , n387053 );
buf ( n387055 , n382950 );
not ( n39539 , n387055 );
buf ( n387057 , n382857 );
not ( n39541 , n387057 );
buf ( n387059 , n384715 );
not ( n39543 , n387059 );
or ( n39544 , n39541 , n39543 );
buf ( n387062 , n384721 );
buf ( n387063 , n382903 );
nand ( n39547 , n387062 , n387063 );
buf ( n387065 , n39547 );
buf ( n387066 , n387065 );
nand ( n39550 , n39544 , n387066 );
buf ( n387068 , n39550 );
buf ( n387069 , n387068 );
not ( n39553 , n387069 );
or ( n39554 , n39539 , n39553 );
and ( n39555 , n384744 , n382857 );
not ( n39556 , n384744 );
and ( n39557 , n39556 , n382903 );
or ( n39558 , n39555 , n39557 );
buf ( n387076 , C1 );
buf ( n387077 , n387076 );
nand ( n39564 , n39554 , n387077 );
buf ( n387079 , n39564 );
buf ( n387080 , n387079 );
xor ( n39567 , n387054 , n387080 );
buf ( n387082 , n384557 );
not ( n39569 , n387082 );
buf ( n387084 , n384568 );
not ( n39571 , n387084 );
buf ( n387086 , n382538 );
not ( n39573 , n387086 );
or ( n39574 , n39571 , n39573 );
buf ( n387089 , n384577 );
buf ( n387090 , n382551 );
nand ( n39577 , n387089 , n387090 );
buf ( n387092 , n39577 );
buf ( n387093 , n387092 );
nand ( n39580 , n39574 , n387093 );
buf ( n387095 , n39580 );
buf ( n387096 , n387095 );
not ( n39583 , n387096 );
or ( n39584 , n39569 , n39583 );
buf ( n387099 , n384568 );
not ( n39586 , n387099 );
buf ( n387101 , n383117 );
not ( n39588 , n387101 );
or ( n39589 , n39586 , n39588 );
buf ( n387104 , n383123 );
buf ( n387105 , n384577 );
nand ( n39592 , n387104 , n387105 );
buf ( n387107 , n39592 );
buf ( n387108 , n387107 );
nand ( n39595 , n39589 , n387108 );
buf ( n387110 , n39595 );
buf ( n387111 , n387110 );
buf ( n387112 , n384627 );
nand ( n39599 , n387111 , n387112 );
buf ( n387114 , n39599 );
buf ( n387115 , n387114 );
nand ( n39602 , n39584 , n387115 );
buf ( n387117 , n39602 );
buf ( n387118 , n387117 );
xor ( n39605 , n39567 , n387118 );
buf ( n387120 , n39605 );
buf ( n387121 , n387120 );
xor ( n39608 , n387030 , n387121 );
buf ( n387123 , n384369 );
not ( n39610 , n387123 );
buf ( n387125 , n36811 );
not ( n39612 , n387125 );
buf ( n387127 , n382535 );
not ( n39614 , n387127 );
or ( n39615 , n39612 , n39614 );
buf ( n387130 , n383975 );
buf ( n387131 , n36822 );
nand ( n39618 , n387130 , n387131 );
buf ( n387133 , n39618 );
buf ( n387134 , n387133 );
nand ( n39621 , n39615 , n387134 );
buf ( n387136 , n39621 );
buf ( n387137 , n387136 );
not ( n39624 , n387137 );
or ( n39625 , n39610 , n39624 );
buf ( n387140 , n387050 );
buf ( n387141 , n384416 );
nand ( n39628 , n387140 , n387141 );
buf ( n387143 , n39628 );
buf ( n387144 , n387143 );
nand ( n39631 , n39625 , n387144 );
buf ( n387146 , n39631 );
and ( n39635 , n383762 , n382857 );
not ( n39636 , n383762 );
and ( n39637 , n39636 , n382903 );
or ( n39638 , n39635 , n39637 );
buf ( n387151 , n39558 );
buf ( n387152 , n382950 );
nand ( n39644 , n387151 , n387152 );
buf ( n387154 , n39644 );
buf ( n387155 , n387154 );
nand ( n39647 , C1 , n387155 );
buf ( n387157 , n39647 );
xor ( n39649 , n387146 , n387157 );
buf ( n387159 , n31964 );
not ( n39651 , n387159 );
buf ( n387161 , n36069 );
not ( n39653 , n387161 );
or ( n39654 , n39651 , n39653 );
buf ( n387164 , n36073 );
buf ( n387165 , n379574 );
nand ( n39657 , n387164 , n387165 );
buf ( n387167 , n39657 );
buf ( n387168 , n387167 );
nand ( n39660 , n39654 , n387168 );
buf ( n387170 , n39660 );
buf ( n387171 , n387170 );
buf ( n387172 , n382607 );
nand ( n39664 , n387171 , n387172 );
buf ( n387174 , n39664 );
nand ( n39666 , n387022 , n379466 );
nand ( n39667 , n387174 , n39666 );
and ( n39668 , n39649 , n39667 );
and ( n39669 , n387146 , n387157 );
or ( n39670 , n39668 , n39669 );
buf ( n387180 , n39670 );
xnor ( n39672 , n39608 , n387180 );
buf ( n387182 , n39672 );
buf ( n387183 , n387182 );
not ( n39675 , n384008 );
not ( n39676 , n383943 );
or ( n39677 , n39675 , n39676 );
nand ( n39678 , n39677 , n39349 );
buf ( n387188 , n39678 );
not ( n39680 , n387188 );
buf ( n387190 , n384416 );
not ( n39682 , n387190 );
buf ( n387192 , n387136 );
not ( n39684 , n387192 );
or ( n39685 , n39682 , n39684 );
buf ( n387195 , n39248 );
buf ( n387196 , n384369 );
nand ( n39688 , n387195 , n387196 );
buf ( n387198 , n39688 );
buf ( n387199 , n387198 );
nand ( n39691 , n39685 , n387199 );
buf ( n387201 , n39691 );
buf ( n387202 , n387201 );
not ( n39694 , n387202 );
or ( n39695 , n39680 , n39694 );
buf ( n387205 , n387170 );
buf ( n387206 , n379466 );
and ( n39698 , n387205 , n387206 );
buf ( n387208 , n386797 );
not ( n39700 , n387208 );
buf ( n387210 , n382604 );
nor ( n39702 , n39700 , n387210 );
buf ( n387212 , n39702 );
buf ( n387213 , n387212 );
nor ( n39705 , n39698 , n387213 );
buf ( n387215 , n39705 );
buf ( n387216 , n387215 );
not ( n39708 , n387216 );
buf ( n387218 , n387201 );
not ( n39710 , n387218 );
buf ( n387220 , n39678 );
not ( n39712 , n387220 );
buf ( n387222 , n39712 );
buf ( n387223 , n387222 );
nand ( n39715 , n39710 , n387223 );
buf ( n387225 , n39715 );
buf ( n387226 , n387225 );
nand ( n39718 , n39708 , n387226 );
buf ( n387228 , n39718 );
buf ( n387229 , n387228 );
nand ( n39721 , n39695 , n387229 );
buf ( n387231 , n39721 );
not ( n39723 , n387231 );
xor ( n39724 , n387146 , n387157 );
xor ( n39725 , n39724 , n39667 );
not ( n39726 , n39725 );
nand ( n39727 , n39723 , n39726 );
buf ( n387237 , n39727 );
buf ( n387238 , n39211 );
buf ( n387239 , n383137 );
not ( n39731 , n387239 );
buf ( n387241 , n383072 );
buf ( n387242 , n384721 );
and ( n39734 , n387241 , n387242 );
not ( n39735 , n387241 );
buf ( n387245 , n384715 );
and ( n39737 , n39735 , n387245 );
nor ( n39738 , n39734 , n39737 );
buf ( n387248 , n39738 );
buf ( n387249 , n387248 );
not ( n39741 , n387249 );
buf ( n387251 , n39741 );
buf ( n387252 , n387251 );
not ( n39744 , n387252 );
or ( n39745 , n39731 , n39744 );
buf ( n387255 , n386829 );
buf ( n387256 , n383017 );
nand ( n39748 , n387255 , n387256 );
buf ( n387258 , n39748 );
buf ( n387259 , n387258 );
nand ( n39751 , n39745 , n387259 );
buf ( n387261 , n39751 );
buf ( n387262 , n387261 );
xor ( n39754 , n387238 , n387262 );
buf ( n387264 , n382950 );
not ( n39756 , n387264 );
buf ( n387266 , n39638 );
not ( n39758 , n387266 );
or ( n39759 , n39756 , n39758 );
buf ( n387269 , C1 );
buf ( n387270 , n387269 );
nand ( n39765 , n39759 , n387270 );
buf ( n387272 , n39765 );
buf ( n387273 , n387272 );
and ( n39768 , n39754 , n387273 );
and ( n39769 , n387238 , n387262 );
or ( n39770 , n39768 , n39769 );
buf ( n387277 , n39770 );
buf ( n387278 , n387277 );
and ( n39773 , n387237 , n387278 );
nor ( n39774 , n39726 , n39723 );
buf ( n387281 , n39774 );
nor ( n39776 , n39773 , n387281 );
buf ( n387283 , n39776 );
buf ( n387284 , n387283 );
not ( n39779 , n387284 );
buf ( n387286 , n383027 );
buf ( n387287 , n384471 );
and ( n39782 , n387286 , n387287 );
not ( n39783 , n387286 );
buf ( n387290 , n36900 );
and ( n39785 , n39783 , n387290 );
or ( n39786 , n39782 , n39785 );
buf ( n387293 , n39786 );
not ( n39788 , n387293 );
not ( n39789 , n383200 );
and ( n39790 , n39788 , n39789 );
buf ( n387297 , n387248 );
buf ( n387298 , n383182 );
nor ( n39793 , n387297 , n387298 );
buf ( n387300 , n39793 );
nor ( n39795 , n39790 , n387300 );
not ( n39796 , n39795 );
not ( n39797 , n387110 );
not ( n39798 , n384557 );
or ( n39799 , n39797 , n39798 );
buf ( n387306 , n383059 );
buf ( n387307 , n384568 );
and ( n39802 , n387306 , n387307 );
buf ( n387309 , n384037 );
buf ( n387310 , n384577 );
and ( n39805 , n387309 , n387310 );
nor ( n39806 , n39802 , n39805 );
buf ( n387313 , n39806 );
not ( n39808 , n387313 );
nand ( n39809 , n39808 , n384627 );
nand ( n39810 , n39799 , n39809 );
not ( n39811 , n39810 );
or ( n39812 , n39796 , n39811 );
or ( n39813 , n39810 , n39795 );
buf ( n387320 , n383482 );
not ( n39815 , n387320 );
and ( n39816 , n384381 , n383445 );
not ( n39817 , n384381 );
and ( n39818 , n39817 , n383429 );
nor ( n39819 , n39816 , n39818 );
buf ( n387326 , n39819 );
not ( n39821 , n387326 );
or ( n39822 , n39815 , n39821 );
and ( n39823 , n382924 , n383429 );
not ( n39824 , n382924 );
and ( n39825 , n39824 , n383445 );
or ( n39826 , n39823 , n39825 );
buf ( n387333 , n39826 );
buf ( n387334 , n383409 );
nand ( n39829 , n387333 , n387334 );
buf ( n387336 , n39829 );
buf ( n387337 , n387336 );
nand ( n39832 , n39822 , n387337 );
buf ( n387339 , n39832 );
not ( n39834 , n387339 );
not ( n39835 , n39834 );
nand ( n39836 , n39813 , n39835 );
nand ( n39837 , n39812 , n39836 );
not ( n39838 , n39837 );
buf ( n387345 , n383137 );
not ( n39840 , n387345 );
buf ( n387347 , n383027 );
not ( n39842 , n387347 );
buf ( n387349 , n36069 );
not ( n39844 , n387349 );
or ( n39845 , n39842 , n39844 );
buf ( n387352 , n36073 );
buf ( n387353 , n383072 );
nand ( n39848 , n387352 , n387353 );
buf ( n387355 , n39848 );
buf ( n387356 , n387355 );
nand ( n39851 , n39845 , n387356 );
buf ( n387358 , n39851 );
buf ( n387359 , n387358 );
not ( n39854 , n387359 );
or ( n39855 , n39840 , n39854 );
buf ( n387362 , n387293 );
not ( n39857 , n387362 );
buf ( n387364 , n383017 );
nand ( n39859 , n39857 , n387364 );
buf ( n387366 , n39859 );
buf ( n387367 , n387366 );
nand ( n39862 , n39855 , n387367 );
buf ( n387369 , n39862 );
xor ( n39864 , n39795 , n387369 );
buf ( n387371 , n383482 );
not ( n39866 , n387371 );
buf ( n387373 , n39826 );
not ( n39868 , n387373 );
or ( n39869 , n39866 , n39868 );
and ( n39870 , n383062 , n383429 );
not ( n39871 , n383062 );
and ( n39872 , n39871 , n383445 );
or ( n39873 , n39870 , n39872 );
buf ( n387380 , n39873 );
buf ( n387381 , n383409 );
nand ( n39876 , n387380 , n387381 );
buf ( n387383 , n39876 );
buf ( n387384 , n387383 );
nand ( n39879 , n39869 , n387384 );
buf ( n387386 , n39879 );
xor ( n39881 , n39864 , n387386 );
not ( n39882 , n39881 );
or ( n39883 , n39838 , n39882 );
or ( n39884 , n39881 , n39837 );
nand ( n39885 , n39883 , n39884 );
buf ( n387392 , n39885 );
not ( n39887 , n387392 );
and ( n39888 , n39779 , n39887 );
buf ( n387395 , n387283 );
buf ( n387396 , n39885 );
and ( n39891 , n387395 , n387396 );
nor ( n387398 , n39888 , n39891 );
buf ( n387399 , n387398 );
buf ( n387400 , n387399 );
xor ( n39895 , n387183 , n387400 );
buf ( n387402 , n39211 );
not ( n39897 , n387402 );
buf ( n387404 , n386776 );
not ( n39899 , n387404 );
or ( n39900 , n39897 , n39899 );
buf ( n387407 , n386753 );
nand ( n39902 , n39900 , n387407 );
buf ( n387409 , n39902 );
buf ( n387410 , n387409 );
buf ( n387411 , n39211 );
not ( n39906 , n387411 );
buf ( n387413 , n386779 );
nand ( n39908 , n39906 , n387413 );
buf ( n387415 , n39908 );
buf ( n387416 , n387415 );
and ( n39911 , n387410 , n387416 );
buf ( n387418 , n39911 );
not ( n39913 , n387418 );
xor ( n39914 , n387222 , n387201 );
xnor ( n39915 , n39914 , n387215 );
not ( n39916 , n39915 );
and ( n39917 , n39913 , n39916 );
buf ( n387424 , n39915 );
buf ( n387425 , n387418 );
nand ( n39920 , n387424 , n387425 );
buf ( n387427 , n39920 );
xor ( n39922 , n387238 , n387262 );
xor ( n39923 , n39922 , n387273 );
buf ( n387430 , n39923 );
and ( n39925 , n387427 , n387430 );
nor ( n39926 , n39917 , n39925 );
buf ( n387433 , n39926 );
not ( n39928 , n387433 );
buf ( n387435 , n39928 );
buf ( n387436 , n387313 );
not ( n39931 , n387436 );
buf ( n387438 , n385227 );
not ( n39933 , n387438 );
and ( n39934 , n39931 , n39933 );
buf ( n387441 , n386936 );
buf ( n387442 , n384627 );
and ( n39937 , n387441 , n387442 );
nor ( n39938 , n39934 , n39937 );
buf ( n387445 , n39938 );
buf ( n387446 , n387445 );
not ( n39941 , n387446 );
buf ( n387448 , n383409 );
not ( n39943 , n387448 );
buf ( n387450 , n39819 );
not ( n39945 , n387450 );
or ( n39946 , n39943 , n39945 );
buf ( n387453 , n386743 );
buf ( n387454 , n383482 );
nand ( n39949 , n387453 , n387454 );
buf ( n387456 , n39949 );
buf ( n387457 , n387456 );
nand ( n39952 , n39946 , n387457 );
buf ( n387459 , n39952 );
buf ( n387460 , n387459 );
not ( n39955 , n387460 );
buf ( n387462 , n39955 );
buf ( n387463 , n387462 );
not ( n39958 , n387463 );
or ( n39959 , n39941 , n39958 );
buf ( n387466 , n386839 );
buf ( n387467 , n386845 );
nand ( n39962 , n387466 , n387467 );
buf ( n387469 , n39962 );
not ( n39964 , n387469 );
not ( n39965 , n386873 );
or ( n39966 , n39964 , n39965 );
or ( n39967 , n386839 , n386845 );
nand ( n39968 , n39966 , n39967 );
buf ( n387475 , n39968 );
nand ( n39970 , n39959 , n387475 );
buf ( n387477 , n39970 );
buf ( n387478 , n387445 );
not ( n39973 , n387478 );
buf ( n387480 , n387459 );
nand ( n39975 , n39973 , n387480 );
buf ( n387482 , n39975 );
nand ( n39977 , n387477 , n387482 );
xor ( n39978 , n39795 , n39834 );
xnor ( n39979 , n39978 , n39810 );
or ( n39980 , n39977 , n39979 );
and ( n39981 , n387435 , n39980 );
and ( n39982 , n39979 , n39977 );
nor ( n39983 , n39981 , n39982 );
buf ( n387490 , n39983 );
xor ( n39985 , n39895 , n387490 );
buf ( n387492 , n39985 );
not ( n39987 , n39726 );
and ( n39988 , n387277 , n39723 );
not ( n39989 , n387277 );
and ( n39990 , n39989 , n387231 );
or ( n39991 , n39988 , n39990 );
not ( n39992 , n39991 );
or ( n39993 , n39987 , n39992 );
or ( n39994 , n39991 , n39726 );
nand ( n39995 , n39993 , n39994 );
not ( n39996 , n39995 );
not ( n39997 , n39926 );
xor ( n39998 , n39979 , n39977 );
not ( n39999 , n39998 );
or ( n40000 , n39997 , n39999 );
or ( n40001 , n39926 , n39998 );
nand ( n40002 , n40000 , n40001 );
not ( n40003 , n40002 );
and ( n40004 , n39996 , n40003 );
buf ( n387511 , n386891 );
buf ( n387512 , n386876 );
or ( n40007 , n387511 , n387512 );
buf ( n387514 , n39266 );
nand ( n40009 , n40007 , n387514 );
buf ( n387516 , n40009 );
buf ( n387517 , n387516 );
buf ( n387518 , n386891 );
buf ( n387519 , n386876 );
nand ( n40014 , n387518 , n387519 );
buf ( n387521 , n40014 );
buf ( n387522 , n387521 );
nand ( n40017 , n387517 , n387522 );
buf ( n387524 , n40017 );
not ( n40019 , n387524 );
xor ( n40020 , n387445 , n387459 );
xor ( n40021 , n40020 , n39968 );
nand ( n40022 , n40019 , n40021 );
buf ( n387529 , n40022 );
xor ( n40024 , n386922 , n386947 );
and ( n40025 , n40024 , n386954 );
and ( n40026 , n386922 , n386947 );
or ( n40027 , n40025 , n40026 );
buf ( n387534 , n40027 );
buf ( n40029 , n387534 );
buf ( n387536 , n40029 );
and ( n40031 , n387529 , n387536 );
not ( n40032 , n387524 );
nor ( n40033 , n40032 , n40021 );
buf ( n387540 , n40033 );
nor ( n40035 , n40031 , n387540 );
buf ( n387542 , n40035 );
nor ( n40037 , n40004 , n387542 );
and ( n40038 , n39995 , n40002 );
nor ( n40039 , n40037 , n40038 );
nand ( n40040 , n387492 , n40039 );
buf ( n387547 , n40040 );
not ( n40042 , n39837 );
nand ( n40043 , n40042 , n39881 );
buf ( n387550 , n40043 );
not ( n40045 , n387550 );
buf ( n387552 , n387283 );
not ( n40047 , n387552 );
buf ( n387554 , n40047 );
buf ( n387555 , n387554 );
not ( n40050 , n387555 );
or ( n40051 , n40045 , n40050 );
not ( n40052 , n39881 );
nand ( n40053 , n40052 , n39837 );
buf ( n387560 , n40053 );
nand ( n40055 , n40051 , n387560 );
buf ( n387562 , n40055 );
buf ( n387563 , n387562 );
buf ( n387564 , n387029 );
not ( n40059 , n387564 );
buf ( n387566 , n39670 );
not ( n40061 , n387566 );
or ( n40062 , n40059 , n40061 );
buf ( n387569 , n387029 );
buf ( n387570 , n39670 );
or ( n40065 , n387569 , n387570 );
buf ( n387572 , n387120 );
nand ( n40067 , n40065 , n387572 );
buf ( n387574 , n40067 );
buf ( n387575 , n387574 );
nand ( n40070 , n40062 , n387575 );
buf ( n387577 , n40070 );
buf ( n387578 , n387577 );
not ( n40073 , n387578 );
buf ( n387580 , n39795 );
not ( n40075 , n387580 );
buf ( n387582 , n387369 );
not ( n40077 , n387582 );
buf ( n387584 , n40077 );
buf ( n387585 , n387584 );
not ( n40080 , n387585 );
or ( n40081 , n40075 , n40080 );
buf ( n387588 , n387386 );
nand ( n40083 , n40081 , n387588 );
buf ( n387590 , n40083 );
buf ( n387591 , n387590 );
buf ( n387592 , n39795 );
not ( n40087 , n387592 );
buf ( n387594 , n387369 );
nand ( n40089 , n40087 , n387594 );
buf ( n387596 , n40089 );
buf ( n387597 , n387596 );
nand ( n40092 , n387591 , n387597 );
buf ( n387599 , n40092 );
buf ( n387600 , n387599 );
buf ( n387601 , n384627 );
not ( n40096 , n387601 );
buf ( n387603 , n387095 );
not ( n40098 , n387603 );
or ( n40099 , n40096 , n40098 );
buf ( n387606 , n384568 );
not ( n40101 , n387606 );
buf ( n387608 , n34863 );
not ( n40103 , n387608 );
or ( n40104 , n40101 , n40103 );
buf ( n387611 , n382473 );
buf ( n387612 , n384577 );
nand ( n40107 , n387611 , n387612 );
buf ( n387614 , n40107 );
buf ( n387615 , n387614 );
nand ( n40110 , n40104 , n387615 );
buf ( n387617 , n40110 );
buf ( n387618 , n387617 );
buf ( n387619 , n384557 );
nand ( n40114 , n387618 , n387619 );
buf ( n387621 , n40114 );
buf ( n387622 , n387621 );
nand ( n40117 , n40099 , n387622 );
buf ( n387624 , n40117 );
buf ( n387625 , n387624 );
and ( n40125 , n385774 , n382857 );
not ( n40126 , n385774 );
and ( n40127 , n40126 , n382903 );
or ( n40128 , n40125 , n40127 );
buf ( n387630 , n40128 );
buf ( n387631 , n382950 );
nand ( n40131 , n387630 , n387631 );
buf ( n387633 , n40131 );
buf ( n387634 , n387633 );
nand ( n40134 , C1 , n387634 );
buf ( n387636 , n40134 );
buf ( n387637 , n387636 );
not ( n40137 , n387637 );
buf ( n387639 , n40137 );
buf ( n387640 , n387639 );
xor ( n40140 , n387625 , n387640 );
buf ( n387642 , n383482 );
not ( n40142 , n387642 );
buf ( n387644 , n39873 );
not ( n40144 , n387644 );
or ( n40145 , n40142 , n40144 );
buf ( n387647 , n383429 );
not ( n40147 , n387647 );
buf ( n387649 , n383117 );
not ( n40149 , n387649 );
or ( n40150 , n40147 , n40149 );
buf ( n387652 , n383123 );
buf ( n387653 , n383445 );
nand ( n40153 , n387652 , n387653 );
buf ( n387655 , n40153 );
buf ( n387656 , n387655 );
nand ( n40156 , n40150 , n387656 );
buf ( n387658 , n40156 );
buf ( n387659 , n387658 );
buf ( n387660 , n383409 );
nand ( n40160 , n387659 , n387660 );
buf ( n387662 , n40160 );
buf ( n387663 , n387662 );
nand ( n40163 , n40145 , n387663 );
buf ( n387665 , n40163 );
buf ( n387666 , n387665 );
xor ( n40166 , n40140 , n387666 );
buf ( n387668 , n40166 );
buf ( n387669 , n387668 );
xor ( n40169 , n387600 , n387669 );
buf ( n387671 , n383137 );
not ( n40171 , n387671 );
buf ( n387673 , n383027 );
not ( n40173 , n387673 );
buf ( n387675 , n383578 );
not ( n40175 , n387675 );
or ( n40176 , n40173 , n40175 );
buf ( n387678 , n383584 );
buf ( n387679 , n383072 );
nand ( n40179 , n387678 , n387679 );
buf ( n387681 , n40179 );
buf ( n387682 , n387681 );
nand ( n40182 , n40176 , n387682 );
buf ( n387684 , n40182 );
buf ( n387685 , n387684 );
not ( n40185 , n387685 );
or ( n40186 , n40171 , n40185 );
buf ( n387688 , n387358 );
buf ( n387689 , n383017 );
nand ( n40189 , n387688 , n387689 );
buf ( n387691 , n40189 );
buf ( n387692 , n387691 );
nand ( n40192 , n40186 , n387692 );
buf ( n387694 , n40192 );
buf ( n387695 , n387694 );
xor ( n40195 , n387054 , n387080 );
and ( n40196 , n40195 , n387118 );
and ( n40197 , n387054 , n387080 );
or ( n40198 , n40196 , n40197 );
buf ( n387700 , n40198 );
buf ( n387701 , n387700 );
xor ( n40201 , n387695 , n387701 );
buf ( n387703 , n382607 );
not ( n40203 , n387703 );
buf ( n387705 , n387007 );
not ( n40205 , n387705 );
or ( n40206 , n40203 , n40205 );
and ( n40207 , n382924 , n379577 );
not ( n40208 , n382924 );
and ( n40209 , n40208 , n379574 );
or ( n40210 , n40207 , n40209 );
buf ( n387712 , n40210 );
buf ( n387713 , n379466 );
nand ( n40213 , n387712 , n387713 );
buf ( n387715 , n40213 );
buf ( n387716 , n387715 );
nand ( n40216 , n40206 , n387716 );
buf ( n387718 , n40216 );
buf ( n387719 , n387718 );
xor ( n40219 , n40201 , n387719 );
buf ( n387721 , n40219 );
buf ( n387722 , n387721 );
xor ( n40222 , n40169 , n387722 );
buf ( n387724 , n40222 );
buf ( n387725 , n387724 );
not ( n40225 , n387725 );
buf ( n387727 , n40225 );
buf ( n387728 , n387727 );
not ( n40228 , n387728 );
or ( n40229 , n40073 , n40228 );
buf ( n387731 , n387724 );
buf ( n387732 , n387577 );
not ( n40232 , n387732 );
buf ( n387734 , n40232 );
buf ( n387735 , n387734 );
nand ( n40235 , n387731 , n387735 );
buf ( n387737 , n40235 );
buf ( n387738 , n387737 );
nand ( n40238 , n40229 , n387738 );
buf ( n387740 , n40238 );
buf ( n387741 , n387740 );
not ( n40241 , n387741 );
xor ( n40242 , n387563 , n40241 );
buf ( n387744 , n40242 );
buf ( n387745 , n387744 );
xor ( n40245 , n387183 , n387400 );
and ( n40246 , n40245 , n387490 );
and ( n40247 , n387183 , n387400 );
or ( n40248 , n40246 , n40247 );
buf ( n387750 , n40248 );
buf ( n387751 , n387750 );
nand ( n40251 , n387745 , n387751 );
buf ( n387753 , n40251 );
buf ( n387754 , n387753 );
nand ( n40254 , n387547 , n387754 );
buf ( n387756 , n40254 );
buf ( n387757 , n387756 );
xor ( n40257 , n39995 , n40002 );
xnor ( n40258 , n40257 , n387542 );
buf ( n387760 , n40258 );
xor ( n40260 , n387418 , n39915 );
xor ( n40261 , n40260 , n387430 );
buf ( n387763 , n40261 );
and ( n40263 , n40021 , n387534 );
not ( n40264 , n40021 );
not ( n40265 , n387534 );
and ( n40266 , n40264 , n40265 );
nor ( n40267 , n40263 , n40266 );
xnor ( n40268 , n387524 , n40267 );
buf ( n387770 , n40268 );
xor ( n40270 , n387763 , n387770 );
buf ( n387772 , n39450 );
buf ( n387773 , n386964 );
nand ( n40273 , n387772 , n387773 );
buf ( n387775 , n40273 );
buf ( n387776 , n387775 );
not ( n40276 , n387776 );
buf ( n387778 , n386916 );
not ( n40278 , n387778 );
or ( n40279 , n40276 , n40278 );
buf ( n387781 , n386956 );
buf ( n387782 , n39444 );
nand ( n40282 , n387781 , n387782 );
buf ( n387784 , n40282 );
buf ( n387785 , n387784 );
nand ( n40285 , n40279 , n387785 );
buf ( n387787 , n40285 );
buf ( n387788 , n387787 );
and ( n40288 , n40270 , n387788 );
and ( n40289 , n387763 , n387770 );
or ( n40290 , n40288 , n40289 );
buf ( n387792 , n40290 );
buf ( n387793 , n387792 );
nor ( n40293 , n387760 , n387793 );
buf ( n387795 , n40293 );
not ( n40295 , n387795 );
not ( n40296 , n386895 );
not ( n40297 , n386976 );
or ( n40298 , n40296 , n40297 );
buf ( n387800 , n39375 );
not ( n40300 , n387800 );
buf ( n387802 , n39453 );
not ( n40302 , n387802 );
or ( n40303 , n40300 , n40302 );
buf ( n387805 , n386718 );
nand ( n40305 , n40303 , n387805 );
buf ( n387807 , n40305 );
nand ( n40307 , n40298 , n387807 );
xor ( n40308 , n387763 , n387770 );
xor ( n40309 , n40308 , n387788 );
buf ( n387811 , n40309 );
or ( n40311 , n40307 , n387811 );
nand ( n40312 , n40295 , n40311 );
buf ( n387814 , n40312 );
nor ( n40314 , n387757 , n387814 );
buf ( n387816 , n40314 );
buf ( n387817 , n387816 );
and ( n40317 , n386993 , n387817 );
buf ( n387819 , n40317 );
buf ( n387820 , n387734 );
not ( n40320 , n387820 );
buf ( n387822 , n387727 );
not ( n40322 , n387822 );
or ( n40323 , n40320 , n40322 );
buf ( n387825 , n387562 );
nand ( n40325 , n40323 , n387825 );
buf ( n387827 , n40325 );
buf ( n387828 , n387827 );
buf ( n387829 , n387724 );
buf ( n387830 , n387577 );
nand ( n40330 , n387829 , n387830 );
buf ( n387832 , n40330 );
buf ( n387833 , n387832 );
nand ( n40333 , n387828 , n387833 );
buf ( n387835 , n40333 );
buf ( n387836 , n387835 );
buf ( n387837 , n382950 );
not ( n40337 , n387837 );
buf ( n387839 , n383654 );
not ( n40339 , n387839 );
or ( n40340 , n40337 , n40339 );
buf ( n387842 , C1 );
buf ( n387843 , n387842 );
nand ( n40346 , n40340 , n387843 );
buf ( n387845 , n40346 );
buf ( n387846 , n387845 );
buf ( n387847 , n382607 );
not ( n40350 , n387847 );
buf ( n387849 , n40210 );
not ( n40352 , n387849 );
or ( n40353 , n40350 , n40352 );
buf ( n387852 , n383612 );
buf ( n387853 , n379466 );
nand ( n40356 , n387852 , n387853 );
buf ( n387855 , n40356 );
buf ( n387856 , n387855 );
nand ( n40359 , n40353 , n387856 );
buf ( n387858 , n40359 );
buf ( n387859 , n387858 );
xor ( n40362 , n387846 , n387859 );
buf ( n387861 , n383137 );
not ( n40364 , n387861 );
buf ( n387863 , n383683 );
not ( n40366 , n387863 );
or ( n40367 , n40364 , n40366 );
buf ( n387866 , n387684 );
buf ( n387867 , n383017 );
nand ( n40370 , n387866 , n387867 );
buf ( n387869 , n40370 );
buf ( n387870 , n387869 );
nand ( n40373 , n40367 , n387870 );
buf ( n387872 , n40373 );
buf ( n387873 , n387872 );
xor ( n40376 , n40362 , n387873 );
buf ( n387875 , n40376 );
buf ( n387876 , n387875 );
xor ( n40379 , n387625 , n387640 );
and ( n40380 , n40379 , n387666 );
and ( n40381 , n387625 , n387640 );
or ( n40382 , n40380 , n40381 );
buf ( n387881 , n40382 );
buf ( n387882 , n387881 );
buf ( n387883 , n385227 );
not ( n40386 , n387883 );
buf ( n387885 , n386127 );
not ( n40388 , n387885 );
or ( n40389 , n40386 , n40388 );
buf ( n387888 , n387617 );
nand ( n40391 , n40389 , n387888 );
buf ( n387890 , n40391 );
buf ( n387891 , n387890 );
buf ( n387892 , n383409 );
not ( n40395 , n387892 );
buf ( n387894 , n383451 );
not ( n40397 , n387894 );
or ( n40398 , n40395 , n40397 );
buf ( n387897 , n387658 );
buf ( n387898 , n383482 );
nand ( n40401 , n387897 , n387898 );
buf ( n387900 , n40401 );
buf ( n387901 , n387900 );
nand ( n40404 , n40398 , n387901 );
buf ( n387903 , n40404 );
buf ( n387904 , n387903 );
xor ( n40407 , n387891 , n387904 );
buf ( n387906 , n387636 );
xor ( n40409 , n40407 , n387906 );
buf ( n387908 , n40409 );
buf ( n387909 , n387908 );
xor ( n40412 , n387882 , n387909 );
xor ( n40413 , n387695 , n387701 );
and ( n40414 , n40413 , n387719 );
and ( n40415 , n387695 , n387701 );
or ( n40416 , n40414 , n40415 );
buf ( n387915 , n40416 );
buf ( n387916 , n387915 );
xor ( n40419 , n40412 , n387916 );
buf ( n387918 , n40419 );
buf ( n387919 , n387918 );
xor ( n40422 , n387876 , n387919 );
xor ( n40423 , n387600 , n387669 );
and ( n40424 , n40423 , n387722 );
and ( n40425 , n387600 , n387669 );
or ( n40426 , n40424 , n40425 );
buf ( n387925 , n40426 );
buf ( n387926 , n387925 );
xor ( n40429 , n40422 , n387926 );
buf ( n387928 , n40429 );
buf ( n387929 , n387928 );
or ( n40432 , n387836 , n387929 );
buf ( n387931 , n40432 );
buf ( n387932 , n387931 );
xor ( n40435 , n387846 , n387859 );
and ( n40436 , n40435 , n387873 );
and ( n40437 , n387846 , n387859 );
or ( n40438 , n40436 , n40437 );
buf ( n387937 , n40438 );
buf ( n387938 , n387937 );
xor ( n40441 , n387882 , n387909 );
and ( n40442 , n40441 , n387916 );
and ( n40443 , n387882 , n387909 );
or ( n40444 , n40442 , n40443 );
buf ( n387943 , n40444 );
buf ( n387944 , n387943 );
xor ( n40447 , n387938 , n387944 );
xor ( n40448 , n387891 , n387904 );
and ( n40449 , n40448 , n387906 );
and ( n40450 , n387891 , n387904 );
or ( n40451 , n40449 , n40450 );
buf ( n387950 , n40451 );
xor ( n40453 , n387950 , n383488 );
buf ( n387952 , n383617 );
not ( n40455 , n387952 );
buf ( n387954 , n383664 );
not ( n40457 , n387954 );
or ( n40458 , n40455 , n40457 );
buf ( n387957 , n383658 );
buf ( n387958 , n36040 );
nand ( n40461 , n387957 , n387958 );
buf ( n387960 , n40461 );
buf ( n387961 , n387960 );
nand ( n40464 , n40458 , n387961 );
buf ( n387963 , n40464 );
buf ( n387964 , n387963 );
buf ( n387965 , n383693 );
xnor ( n40468 , n387964 , n387965 );
buf ( n387967 , n40468 );
xor ( n40470 , n40453 , n387967 );
buf ( n387969 , n40470 );
xor ( n40472 , n40447 , n387969 );
buf ( n387971 , n40472 );
buf ( n387972 , n387971 );
xor ( n40475 , n387876 , n387919 );
and ( n40476 , n40475 , n387926 );
and ( n40477 , n387876 , n387919 );
or ( n40478 , n40476 , n40477 );
buf ( n387977 , n40478 );
buf ( n387978 , n387977 );
nor ( n40481 , n387972 , n387978 );
buf ( n387980 , n40481 );
buf ( n387981 , n387980 );
not ( n40484 , n387981 );
buf ( n387983 , n40484 );
buf ( n387984 , n387983 );
nand ( n40487 , n387932 , n387984 );
buf ( n387986 , n40487 );
xor ( n40489 , n387938 , n387944 );
and ( n40490 , n40489 , n387969 );
and ( n40491 , n387938 , n387944 );
or ( n40492 , n40490 , n40491 );
buf ( n387991 , n40492 );
buf ( n387992 , n387991 );
not ( n40495 , n387992 );
buf ( n387994 , n383505 );
not ( n40497 , n387994 );
buf ( n387996 , n383359 );
not ( n40499 , n387996 );
or ( n40500 , n40497 , n40499 );
buf ( n387999 , n383359 );
buf ( n388000 , n383505 );
or ( n40503 , n387999 , n388000 );
nand ( n40504 , n40500 , n40503 );
buf ( n388003 , n40504 );
xnor ( n40506 , n388003 , n383488 );
buf ( n388005 , n40506 );
buf ( n388006 , n36018 );
not ( n40509 , n388006 );
buf ( n388008 , n383555 );
not ( n40511 , n388008 );
and ( n40512 , n40509 , n40511 );
buf ( n388011 , n383555 );
buf ( n388012 , n36018 );
and ( n40515 , n388011 , n388012 );
nor ( n40516 , n40512 , n40515 );
buf ( n388015 , n40516 );
xor ( n40518 , n388015 , n383699 );
buf ( n388017 , n40518 );
xor ( n40520 , n388005 , n388017 );
buf ( n388019 , n387967 );
buf ( n388020 , n383488 );
nand ( n40523 , n388019 , n388020 );
buf ( n388022 , n40523 );
buf ( n388023 , n388022 );
buf ( n388024 , n387950 );
and ( n40527 , n388023 , n388024 );
buf ( n388026 , n387967 );
buf ( n388027 , n383488 );
nor ( n40530 , n388026 , n388027 );
buf ( n388029 , n40530 );
buf ( n388030 , n388029 );
nor ( n40533 , n40527 , n388030 );
buf ( n388032 , n40533 );
buf ( n388033 , n388032 );
xor ( n40536 , n40520 , n388033 );
buf ( n388035 , n40536 );
buf ( n388036 , n388035 );
nand ( n40539 , n40495 , n388036 );
buf ( n388038 , n40539 );
buf ( n388039 , n388038 );
xor ( n40542 , n383515 , n383530 );
xor ( n40543 , n40542 , n383711 );
buf ( n388042 , n40543 );
buf ( n388043 , n388042 );
not ( n40546 , n388043 );
xor ( n40547 , n388005 , n388017 );
and ( n40548 , n40547 , n388033 );
and ( n40549 , n388005 , n388017 );
or ( n40550 , n40548 , n40549 );
buf ( n388049 , n40550 );
buf ( n388050 , n388049 );
nand ( n40553 , n40546 , n388050 );
buf ( n388052 , n40553 );
buf ( n388053 , n388052 );
nand ( n40556 , n388039 , n388053 );
buf ( n388055 , n40556 );
nor ( n40558 , n387986 , n388055 );
nand ( n40559 , n387819 , n40558 );
buf ( n388058 , n40559 );
not ( n40561 , n388058 );
buf ( n388060 , n40561 );
not ( n40563 , n388060 );
buf ( n388062 , n24269 );
buf ( n40565 , n388062 );
buf ( n388064 , n40565 );
xnor ( n40567 , n388064 , n23868 );
buf ( n388066 , n40567 );
not ( n40569 , n388066 );
buf ( n388068 , n40569 );
buf ( n388069 , n388068 );
not ( n40572 , n388069 );
buf ( n388071 , n40572 );
buf ( n388072 , n388071 );
not ( n40575 , n388072 );
buf ( n388074 , n23868 );
not ( n40577 , n388074 );
buf ( n388076 , n40577 );
buf ( n388077 , n388076 );
buf ( n388078 , n24226 );
not ( n40581 , n388078 );
buf ( n388080 , n40581 );
buf ( n388081 , n388080 );
and ( n40584 , n388077 , n388081 );
not ( n40585 , n388077 );
buf ( n388084 , n24226 );
and ( n40587 , n40585 , n388084 );
nor ( n40588 , n40584 , n40587 );
buf ( n388087 , n40588 );
nand ( n40590 , n388087 , n40567 );
buf ( n40591 , n40590 );
not ( n40592 , n40591 );
buf ( n388091 , n40592 );
not ( n40594 , n388091 );
buf ( n388093 , n40594 );
buf ( n388094 , n388093 );
not ( n40597 , n388094 );
or ( n40598 , n40575 , n40597 );
nand ( n40599 , n24219 , n24222 );
and ( n40600 , n40599 , n24225 );
not ( n40601 , n40600 );
buf ( n388100 , n40601 );
buf ( n40603 , n388100 );
buf ( n388102 , n40603 );
buf ( n388103 , n388102 );
not ( n40606 , n388103 );
buf ( n388105 , n40606 );
buf ( n388106 , n388105 );
not ( n40609 , n388106 );
buf ( n388108 , n385499 );
not ( n40611 , n388108 );
or ( n40612 , n40609 , n40611 );
buf ( n388111 , n385499 );
not ( n40614 , n388111 );
buf ( n388113 , n40614 );
buf ( n388114 , n388113 );
buf ( n388115 , n388102 );
nand ( n40618 , n388114 , n388115 );
buf ( n388117 , n40618 );
buf ( n388118 , n388117 );
nand ( n40621 , n40612 , n388118 );
buf ( n388120 , n40621 );
buf ( n388121 , n388120 );
nand ( n40624 , n40598 , n388121 );
buf ( n388123 , n40624 );
buf ( n388124 , n388123 );
not ( n40627 , n23841 );
buf ( n388126 , n23899 );
not ( n40629 , n388126 );
buf ( n388128 , n40629 );
not ( n40631 , n388128 );
or ( n40632 , n40627 , n40631 );
not ( n40633 , n23898 );
nand ( n40634 , n371498 , n23884 );
not ( n40635 , n40634 );
or ( n40636 , n40633 , n40635 );
nand ( n40637 , n40636 , n23840 );
nand ( n40638 , n40632 , n40637 );
buf ( n40639 , n40638 );
not ( n40640 , n40639 );
buf ( n388139 , n40640 );
not ( n40642 , n388139 );
buf ( n388141 , n40642 );
buf ( n388142 , n388141 );
not ( n40645 , n388142 );
not ( n40646 , n371343 );
not ( n40647 , n371348 );
or ( n40648 , n40646 , n40647 );
not ( n40649 , n371343 );
nand ( n40650 , n40649 , n23745 );
nand ( n40651 , n40648 , n40650 );
not ( n40652 , n40651 );
buf ( n40653 , n40652 );
buf ( n388152 , n40653 );
buf ( n40655 , n388152 );
buf ( n388154 , n40655 );
buf ( n388155 , n388154 );
buf ( n40658 , n388155 );
buf ( n388157 , n40658 );
buf ( n388158 , n388157 );
not ( n40661 , n388158 );
buf ( n388160 , n40661 );
buf ( n388161 , n388160 );
not ( n40664 , n388161 );
buf ( n388163 , n36067 );
not ( n40666 , n388163 );
or ( n40667 , n40664 , n40666 );
buf ( n388166 , n36068 );
buf ( n388167 , n388157 );
nand ( n40670 , n388166 , n388167 );
buf ( n388169 , n40670 );
buf ( n388170 , n388169 );
nand ( n40673 , n40667 , n388170 );
buf ( n388172 , n40673 );
buf ( n388173 , n388172 );
not ( n40676 , n388173 );
or ( n40677 , n40645 , n40676 );
buf ( n388176 , n388160 );
not ( n40679 , n388176 );
buf ( n388178 , n36900 );
not ( n40681 , n388178 );
or ( n40682 , n40679 , n40681 );
buf ( n388181 , n38227 );
buf ( n388182 , n388157 );
nand ( n40685 , n388181 , n388182 );
buf ( n388184 , n40685 );
buf ( n388185 , n388184 );
nand ( n40688 , n40682 , n388185 );
buf ( n388187 , n40688 );
buf ( n388188 , n388187 );
not ( n40691 , n40638 );
buf ( n388190 , n40651 );
buf ( n40693 , n388190 );
buf ( n388192 , n40693 );
nand ( n40695 , n23900 , n388192 );
not ( n40696 , n371356 );
buf ( n40697 , n388128 );
nand ( n40698 , n40696 , n40697 );
nand ( n40699 , n40691 , n40695 , n40698 );
buf ( n40700 , n40699 );
not ( n40701 , n40700 );
buf ( n388200 , n40701 );
nand ( n40703 , n388188 , n388200 );
buf ( n388202 , n40703 );
buf ( n388203 , n388202 );
nand ( n40706 , n40677 , n388203 );
buf ( n388205 , n40706 );
buf ( n388206 , n388205 );
xor ( n40709 , n388124 , n388206 );
not ( n40710 , n12480 );
not ( n40711 , n38685 );
not ( n40712 , n40711 );
or ( n40713 , n40710 , n40712 );
not ( n40714 , n35435 );
buf ( n388213 , n12480 );
not ( n40716 , n388213 );
buf ( n388215 , n40716 );
nand ( n40718 , n40714 , n388215 );
nand ( n40719 , n40713 , n40718 );
not ( n40720 , n40719 );
buf ( n388219 , n40720 );
not ( n40722 , n388219 );
buf ( n388221 , n386300 );
not ( n40724 , n388221 );
or ( n40725 , n40722 , n40724 );
buf ( n388224 , n383137 );
buf ( n388225 , n27234 );
not ( n40728 , n388225 );
buf ( n388227 , n40728 );
buf ( n388228 , n388227 );
not ( n40731 , n388228 );
buf ( n388230 , n40731 );
buf ( n388231 , n388230 );
not ( n40734 , n388231 );
buf ( n388233 , n40711 );
not ( n40736 , n388233 );
buf ( n388235 , n40736 );
buf ( n388236 , n388235 );
not ( n40739 , n388236 );
or ( n40740 , n40734 , n40739 );
buf ( n388239 , n384965 );
buf ( n388240 , n388230 );
not ( n40743 , n388240 );
buf ( n388242 , n40743 );
buf ( n388243 , n388242 );
nand ( n40746 , n388239 , n388243 );
buf ( n388245 , n40746 );
buf ( n388246 , n388245 );
nand ( n40749 , n40740 , n388246 );
buf ( n388248 , n40749 );
buf ( n388249 , n388248 );
nand ( n40752 , n388224 , n388249 );
buf ( n388251 , n40752 );
buf ( n388252 , n388251 );
nand ( n40755 , n40725 , n388252 );
buf ( n388254 , n40755 );
buf ( n388255 , n388254 );
buf ( n40758 , n27610 );
not ( n40759 , n40758 );
not ( n40760 , n40759 );
buf ( n388259 , n40760 );
not ( n40762 , n388259 );
buf ( n388261 , n36259 );
buf ( n40764 , n388261 );
buf ( n388263 , n40764 );
buf ( n388264 , n388263 );
not ( n40767 , n388264 );
buf ( n388266 , n40767 );
buf ( n388267 , n388266 );
not ( n40770 , n388267 );
or ( n40771 , n40762 , n40770 );
buf ( n388270 , n36250 );
not ( n40773 , n388270 );
buf ( n388272 , n40773 );
not ( n40775 , n388272 );
buf ( n388274 , n40775 );
not ( n40777 , n27611 );
not ( n40778 , n40777 );
not ( n40779 , n40778 );
buf ( n388278 , n40779 );
nand ( n40781 , n388274 , n388278 );
buf ( n388280 , n40781 );
buf ( n388281 , n388280 );
nand ( n40784 , n40771 , n388281 );
buf ( n388283 , n40784 );
buf ( n388284 , n388283 );
not ( n40787 , n388284 );
buf ( n388286 , n383891 );
not ( n40789 , n388286 );
or ( n40790 , n40787 , n40789 );
not ( n40791 , n36252 );
not ( n40792 , n40791 );
buf ( n388291 , n375781 );
not ( n40794 , n388291 );
buf ( n388293 , n40794 );
not ( n40796 , n388293 );
or ( n40797 , n40792 , n40796 );
buf ( n388296 , n386147 );
buf ( n388297 , n388263 );
not ( n40800 , n388297 );
buf ( n388299 , n40800 );
buf ( n388300 , n388299 );
nand ( n40803 , n388296 , n388300 );
buf ( n388302 , n40803 );
nand ( n40805 , n40797 , n388302 );
nand ( n40806 , n40805 , n383907 );
buf ( n388305 , n40806 );
nand ( n40808 , n40790 , n388305 );
buf ( n388307 , n40808 );
buf ( n388308 , n388307 );
buf ( n388309 , n384008 );
not ( n40812 , n28213 );
not ( n40813 , n28209 );
not ( n40814 , n40813 );
or ( n40815 , n40812 , n40814 );
nand ( n40816 , n28209 , n28203 );
nand ( n40817 , n40815 , n40816 );
buf ( n40818 , n40817 );
buf ( n40819 , n40818 );
buf ( n388318 , n40819 );
buf ( n388319 , n36395 );
and ( n40822 , n388318 , n388319 );
not ( n40823 , n388318 );
not ( n40824 , n36395 );
buf ( n388323 , n40824 );
and ( n40826 , n40823 , n388323 );
nor ( n40827 , n40822 , n40826 );
buf ( n388326 , n40827 );
buf ( n388327 , n388326 );
or ( n40830 , n388309 , n388327 );
not ( n40831 , n27195 );
not ( n40832 , n40831 );
buf ( n40833 , n40832 );
buf ( n388332 , n40833 );
not ( n40835 , n40824 );
buf ( n388334 , n40835 );
and ( n40837 , n388332 , n388334 );
not ( n40838 , n388332 );
buf ( n40839 , n36424 );
buf ( n40840 , n40839 );
buf ( n388339 , n40840 );
and ( n40842 , n40838 , n388339 );
nor ( n40843 , n40837 , n40842 );
buf ( n388342 , n40843 );
buf ( n388343 , n388342 );
buf ( n388344 , n36363 );
buf ( n40847 , n388344 );
buf ( n388346 , n40847 );
buf ( n388347 , n388346 );
not ( n40850 , n388347 );
buf ( n388349 , n40850 );
buf ( n388350 , n388349 );
or ( n40853 , n388343 , n388350 );
nand ( n40854 , n40830 , n40853 );
buf ( n388353 , n40854 );
buf ( n388354 , n388353 );
xor ( n40857 , n388308 , n388354 );
buf ( n40858 , n36800 );
buf ( n388357 , n40858 );
not ( n40860 , n388357 );
buf ( n388359 , n40860 );
buf ( n388360 , n388359 );
and ( n40863 , n28261 , n28266 );
not ( n40864 , n28261 );
and ( n40865 , n40864 , n28265 );
nor ( n40866 , n40863 , n40865 );
buf ( n388365 , n40866 );
not ( n40868 , n388365 );
buf ( n388367 , n40868 );
buf ( n388368 , n388367 );
not ( n40871 , n388368 );
buf ( n388370 , n40871 );
buf ( n388371 , n388370 );
not ( n40874 , n388371 );
buf ( n388373 , n40874 );
buf ( n388374 , n388373 );
not ( n40877 , n388374 );
buf ( n388376 , n40877 );
buf ( n388377 , n388376 );
not ( n40880 , n388377 );
not ( n40881 , n36769 );
not ( n40882 , n36780 );
or ( n40883 , n40881 , n40882 );
nand ( n40884 , n40883 , n384351 );
buf ( n40885 , n40884 );
not ( n40886 , n40885 );
buf ( n388385 , n40886 );
not ( n40888 , n388385 );
or ( n40889 , n40880 , n40888 );
not ( n40890 , n40884 );
not ( n40891 , n40890 );
nand ( n40892 , n40891 , n388373 );
buf ( n388391 , n40892 );
nand ( n40894 , n40889 , n388391 );
buf ( n388393 , n40894 );
buf ( n388394 , n388393 );
not ( n40897 , n388394 );
buf ( n388396 , n40897 );
buf ( n388397 , n388396 );
or ( n40900 , n388360 , n388397 );
not ( n40901 , n36845 );
buf ( n388400 , n40901 );
not ( n40903 , n388400 );
buf ( n388402 , n40903 );
buf ( n388403 , n388402 );
buf ( n388404 , n28248 );
buf ( n40907 , n388404 );
buf ( n388406 , n40907 );
buf ( n388407 , n388406 );
not ( n40910 , n388407 );
buf ( n388409 , n40910 );
buf ( n388410 , n388409 );
buf ( n40913 , n388410 );
buf ( n388412 , n40913 );
buf ( n388413 , n388412 );
buf ( n388414 , n36810 );
and ( n40917 , n388413 , n388414 );
not ( n40918 , n388413 );
buf ( n388417 , n40885 );
not ( n40920 , n388417 );
buf ( n388419 , n40920 );
buf ( n388420 , n388419 );
and ( n40923 , n40918 , n388420 );
nor ( n40924 , n40917 , n40923 );
buf ( n388423 , n40924 );
buf ( n388424 , n388423 );
or ( n40927 , n388403 , n388424 );
nand ( n40928 , n40900 , n40927 );
buf ( n388427 , n40928 );
buf ( n388428 , n388427 );
and ( n40931 , n40857 , n388428 );
and ( n40932 , n388308 , n388354 );
or ( n40933 , n40931 , n40932 );
buf ( n388432 , n40933 );
buf ( n388433 , n388432 );
xor ( n40936 , n388255 , n388433 );
not ( n40937 , n384413 );
buf ( n388436 , n40819 );
not ( n40939 , n388436 );
buf ( n388438 , n388419 );
not ( n40941 , n388438 );
or ( n40942 , n40939 , n40941 );
buf ( n40943 , n40885 );
buf ( n388442 , n40943 );
buf ( n388443 , n40817 );
not ( n40946 , n388443 );
buf ( n388445 , n40946 );
buf ( n388446 , n388445 );
nand ( n40949 , n388442 , n388446 );
buf ( n388448 , n40949 );
buf ( n388449 , n388448 );
nand ( n40952 , n40942 , n388449 );
buf ( n388451 , n40952 );
not ( n40954 , n388451 );
or ( n40955 , n40937 , n40954 );
not ( n40956 , n388423 );
nand ( n40957 , n40956 , n36801 );
nand ( n40958 , n40955 , n40957 );
buf ( n388457 , n40958 );
buf ( n388458 , n36434 );
not ( n40961 , n388458 );
buf ( n388460 , n40961 );
buf ( n388461 , n388460 );
not ( n40964 , n388461 );
buf ( n388463 , n40964 );
buf ( n388464 , n388463 );
buf ( n388465 , n388342 );
or ( n40968 , n388464 , n388465 );
not ( n40969 , n36363 );
buf ( n388468 , n40969 );
not ( n40971 , n40758 );
not ( n40972 , n36395 );
not ( n40973 , n40972 );
not ( n40974 , n40973 );
and ( n40975 , n40971 , n40974 );
not ( n40976 , n40971 );
not ( n40977 , n36395 );
not ( n40978 , n40977 );
and ( n40979 , n40976 , n40978 );
nor ( n40980 , n40975 , n40979 );
buf ( n388479 , n40980 );
or ( n40982 , n388468 , n388479 );
nand ( n40983 , n40968 , n40982 );
buf ( n388482 , n40983 );
buf ( n388483 , n388482 );
xor ( n40986 , n388457 , n388483 );
buf ( n388485 , n40986 );
buf ( n388486 , n388485 );
buf ( n40990 , n27320 );
buf ( n388488 , n40990 );
buf ( n388489 , n384143 );
and ( n40993 , n388488 , n388489 );
not ( n40994 , n388488 );
buf ( n388492 , n385292 );
and ( n40996 , n40994 , n388492 );
nor ( n40997 , n40993 , n40996 );
buf ( n388495 , n40997 );
buf ( n388496 , n382938 );
not ( n41002 , n388496 );
buf ( n388498 , n41002 );
buf ( n388499 , n388498 );
buf ( n388500 , n28353 );
buf ( n41006 , n388500 );
buf ( n388502 , n41006 );
buf ( n388503 , n388502 );
not ( n41009 , n388503 );
buf ( n388505 , n384096 );
not ( n41011 , n388505 );
or ( n41012 , n41009 , n41011 );
buf ( n388508 , n382854 );
buf ( n388509 , n388502 );
not ( n41015 , n388509 );
buf ( n388511 , n41015 );
buf ( n388512 , n388511 );
nand ( n41018 , n388508 , n388512 );
buf ( n388514 , n41018 );
buf ( n388515 , n388514 );
nand ( n41021 , n41012 , n388515 );
buf ( n388517 , n41021 );
buf ( n388518 , n388517 );
not ( n41024 , n388518 );
buf ( n388520 , n41024 );
buf ( n388521 , n388520 );
or ( n41027 , n388499 , n388521 );
nand ( n41028 , C1 , n41027 );
buf ( n388524 , n41028 );
buf ( n388525 , n388524 );
xor ( n41031 , n388486 , n388525 );
buf ( n388527 , n41031 );
buf ( n388528 , n388527 );
and ( n41034 , n40936 , n388528 );
and ( n41035 , n388255 , n388433 );
or ( n41036 , n41034 , n41035 );
buf ( n388532 , n41036 );
buf ( n388533 , n388532 );
xor ( n41039 , n40709 , n388533 );
buf ( n388535 , n41039 );
buf ( n388536 , n388535 );
buf ( n388537 , n383467 );
buf ( n41043 , n388537 );
buf ( n388539 , n41043 );
buf ( n388540 , n388539 );
buf ( n388541 , n28644 );
buf ( n41047 , n388541 );
buf ( n388543 , n41047 );
buf ( n388544 , n388543 );
not ( n41050 , n388544 );
buf ( n388546 , n41050 );
buf ( n388547 , n388546 );
not ( n41053 , n388547 );
buf ( n388549 , n41053 );
buf ( n388550 , n388549 );
buf ( n388551 , n385633 );
and ( n41057 , n388550 , n388551 );
not ( n41058 , n388550 );
buf ( n388554 , n383414 );
buf ( n41060 , n388554 );
buf ( n388556 , n41060 );
buf ( n388557 , n388556 );
and ( n41063 , n41058 , n388557 );
nor ( n41064 , n41057 , n41063 );
buf ( n388560 , n41064 );
buf ( n388561 , n388560 );
or ( n41067 , n388540 , n388561 );
buf ( n388563 , n383403 );
buf ( n388564 , n27258 );
not ( n41070 , n388564 );
buf ( n388566 , n41070 );
buf ( n388567 , n388566 );
buf ( n41073 , n388567 );
buf ( n388569 , n41073 );
buf ( n388570 , n388569 );
buf ( n388571 , n388556 );
and ( n41077 , n388570 , n388571 );
not ( n41078 , n388570 );
buf ( n388574 , n383417 );
buf ( n41080 , n388574 );
buf ( n388576 , n41080 );
buf ( n388577 , n388576 );
and ( n41083 , n41078 , n388577 );
nor ( n41084 , n41077 , n41083 );
buf ( n388580 , n41084 );
buf ( n388581 , n388580 );
or ( n41087 , n388563 , n388581 );
nand ( n41088 , n41067 , n41087 );
buf ( n388584 , n41088 );
not ( n41090 , n388584 );
buf ( n388586 , n38765 );
not ( n41092 , n388586 );
buf ( n388588 , n41092 );
buf ( n388589 , n35435 );
not ( n41095 , n388589 );
buf ( n388591 , n388511 );
not ( n41097 , n388591 );
and ( n41098 , n41095 , n41097 );
buf ( n388594 , n35435 );
buf ( n388595 , n388511 );
and ( n41101 , n388594 , n388595 );
nor ( n41102 , n41098 , n41101 );
buf ( n388598 , n41102 );
or ( n41104 , n388588 , n388598 );
not ( n41105 , n383134 );
nand ( n41106 , n41105 , n40720 );
nand ( n41107 , n41104 , n41106 );
not ( n41108 , n41107 );
nand ( n41109 , n41090 , n41108 );
not ( n41110 , n41109 );
buf ( n388606 , n388299 );
not ( n41112 , n388606 );
buf ( n388608 , n41112 );
buf ( n388609 , n388608 );
buf ( n388610 , n27196 );
and ( n41116 , n388609 , n388610 );
not ( n41117 , n388609 );
not ( n41118 , n27195 );
buf ( n388614 , n41118 );
and ( n41120 , n41117 , n388614 );
nor ( n41121 , n41116 , n41120 );
buf ( n388617 , n41121 );
buf ( n388618 , n388617 );
not ( n41124 , n388618 );
buf ( n388620 , n383891 );
not ( n41126 , n388620 );
or ( n41127 , n41124 , n41126 );
buf ( n388623 , n388283 );
buf ( n388624 , n383904 );
not ( n41130 , n388624 );
buf ( n388626 , n41130 );
buf ( n388627 , n388626 );
not ( n41133 , n388627 );
buf ( n388629 , n41133 );
buf ( n388630 , n388629 );
nand ( n41136 , n388623 , n388630 );
buf ( n388632 , n41136 );
buf ( n388633 , n388632 );
nand ( n41139 , n41127 , n388633 );
buf ( n388635 , n41139 );
buf ( n388636 , n388635 );
and ( n41142 , n27280 , n374897 );
not ( n41143 , n27280 );
and ( n41144 , n41143 , n374902 );
nor ( n41145 , n41142 , n41144 );
buf ( n388641 , n41145 );
buf ( n41147 , n388641 );
buf ( n388643 , n41147 );
buf ( n388644 , n388643 );
buf ( n41150 , n388644 );
buf ( n388646 , n41150 );
buf ( n388647 , n388646 );
not ( n41153 , n388647 );
buf ( n388649 , n388419 );
not ( n41155 , n388649 );
or ( n41156 , n41153 , n41155 );
buf ( n388652 , n388646 );
not ( n41158 , n388652 );
buf ( n388654 , n41158 );
buf ( n388655 , n388654 );
buf ( n388656 , n40943 );
nand ( n41162 , n388655 , n388656 );
buf ( n388658 , n41162 );
buf ( n388659 , n388658 );
nand ( n41165 , n41156 , n388659 );
buf ( n388661 , n41165 );
buf ( n388662 , n388661 );
not ( n41168 , n388662 );
buf ( n388664 , n36801 );
not ( n41170 , n388664 );
or ( n41171 , n41168 , n41170 );
buf ( n388667 , n36845 );
not ( n41173 , n388667 );
buf ( n388669 , n41173 );
buf ( n388670 , n388669 );
buf ( n388671 , n388393 );
nand ( n41177 , n388670 , n388671 );
buf ( n388673 , n41177 );
buf ( n388674 , n388673 );
nand ( n41180 , n41171 , n388674 );
buf ( n388676 , n41180 );
buf ( n388677 , n388676 );
xor ( n41183 , n388636 , n388677 );
buf ( n388679 , n384008 );
buf ( n388680 , n388412 );
not ( n41186 , n388680 );
buf ( n388682 , n41186 );
buf ( n388683 , n388682 );
not ( n41189 , n388683 );
buf ( n388685 , n36395 );
not ( n41191 , n388685 );
or ( n41192 , n41189 , n41191 );
buf ( n388688 , n40977 );
buf ( n41194 , n28249 );
buf ( n41195 , n41194 );
buf ( n388691 , n41195 );
nand ( n41197 , n388688 , n388691 );
buf ( n388693 , n41197 );
buf ( n388694 , n388693 );
nand ( n41200 , n41192 , n388694 );
buf ( n388696 , n41200 );
buf ( n388697 , n388696 );
not ( n41203 , n388697 );
buf ( n388699 , n41203 );
buf ( n388700 , n388699 );
or ( n41206 , n388679 , n388700 );
buf ( n388702 , n383940 );
not ( n41208 , n388702 );
buf ( n388704 , n41208 );
buf ( n388705 , n388704 );
buf ( n388706 , n388326 );
or ( n41212 , n388705 , n388706 );
nand ( n41213 , n41206 , n41212 );
buf ( n388709 , n41213 );
buf ( n388710 , n388709 );
and ( n41216 , n41183 , n388710 );
and ( n41217 , n388636 , n388677 );
or ( n41218 , n41216 , n41217 );
buf ( n388714 , n41218 );
not ( n41220 , n388714 );
or ( n41221 , n41110 , n41220 );
nand ( n388717 , n41107 , n388584 );
nand ( n41223 , n41221 , n388717 );
buf ( n388719 , n41223 );
buf ( n388720 , n24226 );
buf ( n41226 , n388720 );
buf ( n388722 , n41226 );
xnor ( n41228 , n23773 , n388722 );
buf ( n388724 , n41228 );
buf ( n388725 , n371781 );
buf ( n388726 , n23773 );
nand ( n41232 , n388725 , n388726 );
buf ( n388728 , n41232 );
buf ( n388729 , n388728 );
buf ( n388730 , n371781 );
not ( n41236 , n388730 );
buf ( n388732 , n23774 );
nand ( n41238 , n41236 , n388732 );
buf ( n388734 , n41238 );
buf ( n388735 , n388734 );
nand ( n41241 , n388724 , n388729 , n388735 );
buf ( n388737 , n41241 );
buf ( n388738 , n388737 );
not ( n41244 , n388738 );
buf ( n388740 , n41244 );
buf ( n388741 , n388740 );
not ( n41247 , n388741 );
buf ( n388743 , n41247 );
buf ( n388744 , n388743 );
not ( n41250 , n388744 );
buf ( n388746 , n41250 );
buf ( n388747 , n388746 );
not ( n41253 , n388747 );
buf ( n388749 , n371781 );
not ( n41255 , n388749 );
buf ( n388751 , n41255 );
buf ( n388752 , n388751 );
buf ( n41258 , n388752 );
buf ( n388754 , n41258 );
buf ( n388755 , n388754 );
buf ( n41261 , n388755 );
buf ( n388757 , n41261 );
buf ( n388758 , n388757 );
not ( n41264 , n388758 );
buf ( n388760 , n41264 );
buf ( n388761 , n388760 );
not ( n41267 , n388761 );
buf ( n388763 , n383053 );
not ( n41269 , n388763 );
buf ( n388765 , n41269 );
buf ( n388766 , n388765 );
not ( n41272 , n388766 );
or ( n41273 , n41267 , n41272 );
buf ( n388769 , n383053 );
not ( n41275 , n388769 );
buf ( n388771 , n41275 );
buf ( n388772 , n388771 );
not ( n41278 , n388772 );
buf ( n388774 , n41278 );
buf ( n388775 , n388774 );
buf ( n388776 , n388757 );
nand ( n41282 , n388775 , n388776 );
buf ( n388778 , n41282 );
buf ( n388779 , n388778 );
nand ( n41285 , n41273 , n388779 );
buf ( n388781 , n41285 );
buf ( n388782 , n388781 );
not ( n41288 , n388782 );
or ( n41289 , n41253 , n41288 );
buf ( n388785 , n388760 );
not ( n41291 , n388785 );
buf ( n388787 , n38532 );
not ( n41293 , n388787 );
or ( n41294 , n41291 , n41293 );
buf ( n388790 , n35519 );
buf ( n388791 , n388757 );
nand ( n41297 , n388790 , n388791 );
buf ( n388793 , n41297 );
buf ( n388794 , n388793 );
nand ( n41300 , n41294 , n388794 );
buf ( n388796 , n41300 );
buf ( n388797 , n388796 );
buf ( n388798 , n41228 );
buf ( n41304 , n388798 );
buf ( n388800 , n41304 );
buf ( n388801 , n388800 );
not ( n41307 , n388801 );
buf ( n388803 , n41307 );
buf ( n388804 , n388803 );
not ( n41310 , n388804 );
buf ( n388806 , n41310 );
buf ( n388807 , n388806 );
not ( n41313 , n388807 );
buf ( n388809 , n41313 );
buf ( n388810 , n388809 );
nand ( n41316 , n388797 , n388810 );
buf ( n388812 , n41316 );
buf ( n388813 , n388812 );
nand ( n41319 , n41289 , n388813 );
buf ( n388815 , n41319 );
buf ( n388816 , n388815 );
xor ( n41322 , n388719 , n388816 );
not ( n41323 , n371719 );
not ( n41324 , n41323 );
not ( n41325 , n41324 );
not ( n41326 , n23813 );
not ( n41327 , n41326 );
or ( n41328 , n41325 , n41327 );
nand ( n41329 , n41323 , n23813 );
nand ( n41330 , n41328 , n41329 );
not ( n41331 , n41330 );
not ( n41332 , n41331 );
buf ( n388828 , n41332 );
not ( n41334 , n388828 );
buf ( n388830 , n41334 );
buf ( n388831 , n388830 );
buf ( n41337 , n388831 );
buf ( n388833 , n41337 );
buf ( n388834 , n388833 );
not ( n41340 , n388834 );
buf ( n41341 , n23840 );
not ( n41342 , n41341 );
buf ( n388838 , n41342 );
not ( n41344 , n388838 );
buf ( n388840 , n37027 );
not ( n41346 , n388840 );
or ( n41347 , n41344 , n41346 );
buf ( n388843 , n385834 );
not ( n41349 , n41342 );
buf ( n388845 , n41349 );
nand ( n41351 , n388843 , n388845 );
buf ( n388847 , n41351 );
buf ( n388848 , n388847 );
nand ( n41354 , n41347 , n388848 );
buf ( n388850 , n41354 );
buf ( n388851 , n388850 );
not ( n41357 , n388851 );
or ( n41358 , n41340 , n41357 );
not ( n41359 , n36066 );
and ( n41360 , n41342 , n41359 );
not ( n41361 , n41342 );
and ( n41362 , n41361 , n38822 );
or ( n41363 , n41360 , n41362 );
buf ( n388859 , n41363 );
not ( n41365 , n23840 );
nand ( n41366 , n41365 , n371420 );
buf ( n388862 , n23813 );
buf ( n388863 , n23840 );
nand ( n41369 , n388862 , n388863 );
buf ( n388865 , n41369 );
nand ( n41371 , n41330 , n41366 , n388865 );
buf ( n41372 , n41371 );
not ( n41373 , n41372 );
not ( n41374 , n41373 );
buf ( n388870 , n41374 );
not ( n41376 , n388870 );
buf ( n388872 , n41376 );
buf ( n388873 , n388872 );
nand ( n41379 , n388859 , n388873 );
buf ( n388875 , n41379 );
buf ( n388876 , n388875 );
nand ( n41382 , n41358 , n388876 );
buf ( n388878 , n41382 );
buf ( n388879 , n388878 );
and ( n41385 , n41322 , n388879 );
and ( n41386 , n388719 , n388816 );
or ( n41387 , n41385 , n41386 );
buf ( n388883 , n41387 );
buf ( n388884 , n388883 );
xor ( n41390 , n388536 , n388884 );
xor ( n41391 , n388255 , n388433 );
xor ( n41392 , n41391 , n388528 );
buf ( n388888 , n41392 );
buf ( n388889 , n388888 );
buf ( n388890 , n388293 );
not ( n41396 , n388890 );
buf ( n388892 , n41396 );
buf ( n388893 , n388892 );
not ( n41399 , n388893 );
buf ( n388895 , n384887 );
not ( n41401 , n388895 );
buf ( n388897 , n41401 );
buf ( n388898 , n388897 );
not ( n41404 , n388898 );
and ( n41405 , n41399 , n41404 );
buf ( n388901 , n386147 );
buf ( n41407 , n36304 );
buf ( n388903 , n41407 );
buf ( n41409 , n388903 );
buf ( n388905 , n41409 );
buf ( n388906 , n388905 );
not ( n41412 , n388906 );
buf ( n388908 , n41412 );
buf ( n388909 , n388908 );
and ( n41415 , n388901 , n388909 );
nor ( n41416 , n41405 , n41415 );
buf ( n388912 , n41416 );
not ( n41418 , n388912 );
not ( n41419 , n384901 );
and ( n41420 , n41418 , n41419 );
buf ( n388916 , n388908 );
buf ( n388917 , n28159 );
not ( n41423 , n388917 );
buf ( n388919 , n41423 );
buf ( n388920 , n388919 );
not ( n41426 , n388920 );
buf ( n388922 , n41426 );
buf ( n388923 , n388922 );
and ( n41429 , n388916 , n388923 );
not ( n41430 , n388916 );
buf ( n388926 , n28159 );
buf ( n41432 , n388926 );
buf ( n388928 , n41432 );
buf ( n388929 , n388928 );
not ( n41435 , n388929 );
buf ( n388931 , n41435 );
buf ( n388932 , n388931 );
and ( n41438 , n41430 , n388932 );
nor ( n41439 , n41429 , n41438 );
buf ( n388935 , n41439 );
buf ( n388936 , n388935 );
buf ( n388937 , n37317 );
nor ( n41443 , n388936 , n388937 );
buf ( n388939 , n41443 );
nor ( n41445 , n41420 , n388939 );
buf ( n388941 , n41445 );
not ( n41447 , n37923 );
buf ( n388943 , n41447 );
not ( n41449 , n388943 );
buf ( n388945 , n385473 );
not ( n41451 , n388945 );
buf ( n388947 , n37762 );
not ( n41453 , n388947 );
buf ( n388949 , n41453 );
buf ( n388950 , n388949 );
not ( n41456 , n388950 );
buf ( n388952 , n41456 );
buf ( n388953 , n388952 );
not ( n41459 , n388953 );
buf ( n388955 , n41459 );
buf ( n388956 , n388955 );
not ( n41462 , n388956 );
or ( n41463 , n41451 , n41462 );
buf ( n388959 , n37763 );
buf ( n388960 , n23528 );
buf ( n41466 , n388960 );
buf ( n388962 , n41466 );
buf ( n388963 , n388962 );
not ( n41469 , n388963 );
buf ( n388965 , n41469 );
buf ( n388966 , n388965 );
nand ( n41472 , n388959 , n388966 );
buf ( n388968 , n41472 );
buf ( n388969 , n388968 );
nand ( n41475 , n41463 , n388969 );
buf ( n388971 , n41475 );
buf ( n388972 , n388971 );
not ( n41478 , n388972 );
or ( n41479 , n41449 , n41478 );
buf ( n388975 , n385473 );
not ( n41481 , n388975 );
buf ( n388977 , n29077 );
not ( n41483 , n388977 );
buf ( n388979 , n41483 );
buf ( n388980 , n388979 );
not ( n41486 , n388980 );
or ( n41487 , n41481 , n41486 );
nand ( n41488 , n29077 , n388965 );
buf ( n388984 , n41488 );
nand ( n41490 , n41487 , n388984 );
buf ( n388986 , n41490 );
buf ( n388987 , n388986 );
buf ( n388988 , n385479 );
nand ( n41494 , n388987 , n388988 );
buf ( n388990 , n41494 );
buf ( n388991 , n388990 );
nand ( n41497 , n41479 , n388991 );
buf ( n388993 , n41497 );
buf ( n388994 , n388993 );
xor ( n41500 , n388941 , n388994 );
buf ( n388996 , n388215 );
not ( n41502 , n388996 );
buf ( n388998 , n41502 );
buf ( n388999 , n388998 );
not ( n41505 , n388999 );
buf ( n389001 , n385972 );
not ( n41507 , n389001 );
or ( n41508 , n41505 , n41507 );
buf ( n389004 , n31964 );
buf ( n389005 , n388215 );
nand ( n41511 , n389004 , n389005 );
buf ( n389007 , n41511 );
buf ( n389008 , n389007 );
nand ( n41514 , n41508 , n389008 );
buf ( n389010 , n41514 );
buf ( n389011 , n389010 );
not ( n41517 , n389011 );
buf ( n389013 , n382592 );
not ( n41519 , n389013 );
buf ( n389015 , n41519 );
buf ( n389016 , n389015 );
not ( n41522 , n389016 );
or ( n41523 , n41517 , n41522 );
buf ( n389019 , n31850 );
not ( n41525 , n389019 );
buf ( n389021 , n41525 );
buf ( n389022 , n389021 );
buf ( n41528 , n389022 );
buf ( n389024 , n41528 );
buf ( n389025 , n389024 );
buf ( n389026 , n388230 );
not ( n41532 , n389026 );
buf ( n389028 , n385972 );
not ( n41534 , n389028 );
or ( n41535 , n41532 , n41534 );
buf ( n389031 , n31964 );
buf ( n389032 , n388242 );
nand ( n41538 , n389031 , n389032 );
buf ( n389034 , n41538 );
buf ( n389035 , n389034 );
nand ( n41541 , n41535 , n389035 );
buf ( n389037 , n41541 );
buf ( n389038 , n389037 );
nand ( n41544 , n389025 , n389038 );
buf ( n389040 , n41544 );
buf ( n389041 , n389040 );
nand ( n41547 , n41523 , n389041 );
buf ( n389043 , n41547 );
buf ( n389044 , n389043 );
and ( n41550 , n41500 , n389044 );
and ( n41551 , n388941 , n388994 );
or ( n41552 , n41550 , n41551 );
buf ( n389048 , n41552 );
buf ( n389049 , n389048 );
not ( n41555 , n24069 );
and ( n41556 , n23960 , n41555 );
not ( n41557 , n23960 );
not ( n41558 , n24069 );
not ( n41559 , n41558 );
and ( n41560 , n41557 , n41559 );
nor ( n41561 , n41556 , n41560 );
buf ( n41562 , n41561 );
not ( n41563 , n41562 );
not ( n41564 , n41563 );
not ( n41565 , n41564 );
buf ( n389061 , n41565 );
not ( n41567 , n389061 );
buf ( n389063 , n24050 );
not ( n41569 , n389063 );
buf ( n389065 , n384199 );
not ( n41571 , n389065 );
buf ( n389067 , n41571 );
buf ( n389068 , n389067 );
not ( n41574 , n389068 );
or ( n41575 , n41569 , n41574 );
buf ( n389071 , n384186 );
buf ( n41577 , n24049 );
buf ( n389073 , n41577 );
not ( n41579 , n389073 );
buf ( n389075 , n41579 );
buf ( n389076 , n389075 );
nand ( n41582 , n389071 , n389076 );
buf ( n389078 , n41582 );
buf ( n389079 , n389078 );
nand ( n41585 , n41575 , n389079 );
buf ( n389081 , n41585 );
buf ( n389082 , n389081 );
not ( n41588 , n389082 );
or ( n41589 , n41567 , n41588 );
buf ( n389085 , n24050 );
not ( n41591 , n389085 );
not ( n41592 , n36655 );
not ( n41593 , n36663 );
or ( n41594 , n41592 , n41593 );
nand ( n41595 , n41594 , n36667 );
not ( n41596 , n41595 );
buf ( n389092 , n41596 );
not ( n41598 , n389092 );
or ( n41599 , n41591 , n41598 );
buf ( n389095 , n38472 );
buf ( n389096 , n389075 );
nand ( n41602 , n389095 , n389096 );
buf ( n389098 , n41602 );
buf ( n389099 , n389098 );
nand ( n41605 , n41599 , n389099 );
buf ( n389101 , n41605 );
buf ( n389102 , n389101 );
buf ( n389103 , n38935 );
not ( n41609 , n389103 );
buf ( n389105 , n23960 );
not ( n41611 , n389105 );
buf ( n389107 , n41611 );
buf ( n389108 , n389107 );
nand ( n41614 , n41609 , n389108 );
buf ( n389110 , n41614 );
buf ( n389111 , n389110 );
buf ( n389112 , n41561 );
nand ( n41618 , n23960 , n38935 );
buf ( n389114 , n41618 );
nand ( n41620 , n389111 , n389112 , n389114 );
buf ( n389116 , n41620 );
buf ( n389117 , n389116 );
buf ( n41623 , n389117 );
buf ( n389119 , n41623 );
buf ( n389120 , n389119 );
not ( n41626 , n389120 );
buf ( n389122 , n41626 );
buf ( n389123 , n389122 );
buf ( n41629 , n389123 );
buf ( n389125 , n41629 );
buf ( n389126 , n389125 );
nand ( n41632 , n389102 , n389126 );
buf ( n389128 , n41632 );
buf ( n389129 , n389128 );
nand ( n41635 , n41589 , n389129 );
buf ( n389131 , n41635 );
buf ( n389132 , n389131 );
xor ( n41638 , n389049 , n389132 );
xor ( n41639 , n388308 , n388354 );
xor ( n41640 , n41639 , n388428 );
buf ( n389136 , n41640 );
buf ( n389137 , n389136 );
and ( n41643 , n41638 , n389137 );
and ( n41644 , n389049 , n389132 );
or ( n41645 , n41643 , n41644 );
buf ( n389141 , n41645 );
buf ( n389142 , n389141 );
xor ( n41648 , n388889 , n389142 );
not ( n41649 , n388751 );
buf ( n389145 , n371736 );
buf ( n389146 , n371744 );
and ( n41652 , n389145 , n389146 );
not ( n41653 , n389145 );
buf ( n389149 , n371741 );
and ( n41655 , n41653 , n389149 );
nor ( n41656 , n41652 , n41655 );
buf ( n389152 , n41656 );
not ( n41658 , n389152 );
not ( n41659 , n41658 );
or ( n41660 , n41649 , n41659 );
not ( n41661 , n371797 );
nand ( n41662 , n389152 , n41661 );
nand ( n41663 , n41660 , n41662 );
not ( n41664 , n41663 );
buf ( n389160 , n41664 );
buf ( n41666 , n389160 );
buf ( n389162 , n41666 );
buf ( n389163 , n389162 );
not ( n41669 , n389163 );
buf ( n41670 , n24117 );
not ( n41671 , n41670 );
buf ( n389167 , n41671 );
not ( n41673 , n389167 );
buf ( n389169 , n386561 );
not ( n41675 , n389169 );
or ( n41676 , n41673 , n41675 );
buf ( n389172 , n382921 );
not ( n41678 , n41671 );
buf ( n389174 , n41678 );
nand ( n41680 , n389172 , n389174 );
buf ( n389176 , n41680 );
buf ( n389177 , n389176 );
nand ( n41683 , n41676 , n389177 );
buf ( n389179 , n41683 );
buf ( n389180 , n389179 );
not ( n41686 , n389180 );
or ( n41687 , n41669 , n41686 );
buf ( n389183 , n24118 );
not ( n41689 , n389183 );
buf ( n389185 , n386391 );
not ( n41691 , n389185 );
or ( n41692 , n41689 , n41691 );
buf ( n389188 , n35301 );
buf ( n389189 , n41678 );
nand ( n41695 , n389188 , n389189 );
buf ( n389191 , n41695 );
buf ( n389192 , n389191 );
nand ( n41698 , n41692 , n389192 );
buf ( n389194 , n41698 );
buf ( n389195 , n389194 );
buf ( n389196 , n371751 );
buf ( n389197 , n371719 );
nand ( n41703 , n389196 , n389197 );
buf ( n389199 , n41703 );
not ( n41705 , n371751 );
nand ( n41706 , n41705 , n41323 );
nand ( n41707 , n389199 , n41663 , n41706 );
not ( n41708 , n41707 );
not ( n41709 , n41708 );
buf ( n41710 , n41709 );
not ( n41711 , n41710 );
buf ( n389207 , n41711 );
nand ( n41713 , n389195 , n389207 );
buf ( n389209 , n41713 );
buf ( n389210 , n389209 );
nand ( n41716 , n41687 , n389210 );
buf ( n389212 , n41716 );
buf ( n389213 , n389212 );
and ( n41719 , n41648 , n389213 );
and ( n41720 , n388889 , n389142 );
or ( n41721 , n41719 , n41720 );
buf ( n389217 , n41721 );
buf ( n389218 , n389217 );
xor ( n41724 , n41390 , n389218 );
buf ( n389220 , n41724 );
buf ( n389221 , n388760 );
not ( n41727 , n389221 );
buf ( n389223 , n382924 );
not ( n41729 , n389223 );
or ( n41730 , n41727 , n41729 );
buf ( n389226 , n386561 );
not ( n41732 , n389226 );
buf ( n389228 , n388757 );
nand ( n41734 , n41732 , n389228 );
buf ( n389230 , n41734 );
buf ( n389231 , n389230 );
nand ( n41737 , n41730 , n389231 );
buf ( n389233 , n41737 );
buf ( n389234 , n389233 );
buf ( n389235 , n388746 );
and ( n41741 , n389234 , n389235 );
buf ( n389237 , n388781 );
not ( n41743 , n389237 );
buf ( n389239 , n388806 );
nor ( n41745 , n41743 , n389239 );
buf ( n389241 , n41745 );
buf ( n389242 , n389241 );
nor ( n41748 , n41741 , n389242 );
buf ( n389244 , n41748 );
buf ( n389245 , n389244 );
not ( n41751 , n389245 );
buf ( n389247 , n41751 );
buf ( n389248 , n389247 );
not ( n41754 , n389248 );
buf ( n389250 , n389162 );
not ( n41756 , n389250 );
buf ( n389252 , n389194 );
not ( n41758 , n389252 );
or ( n41759 , n41756 , n41758 );
buf ( n389255 , n41671 );
not ( n41761 , n389255 );
buf ( n389257 , n37027 );
not ( n41763 , n389257 );
or ( n41764 , n41761 , n41763 );
buf ( n389260 , n385834 );
buf ( n389261 , n41678 );
nand ( n41767 , n389260 , n389261 );
buf ( n389263 , n41767 );
buf ( n389264 , n389263 );
nand ( n41770 , n41764 , n389264 );
buf ( n389266 , n41770 );
buf ( n389267 , n389266 );
buf ( n389268 , n41711 );
nand ( n41774 , n389267 , n389268 );
buf ( n389270 , n41774 );
buf ( n389271 , n389270 );
nand ( n41777 , n41759 , n389271 );
buf ( n389273 , n41777 );
buf ( n389274 , n389273 );
not ( n41780 , n389274 );
or ( n41781 , n41754 , n41780 );
buf ( n389277 , n389273 );
buf ( n389278 , n389247 );
or ( n41784 , n389277 , n389278 );
buf ( n389280 , n41565 );
not ( n41786 , n389280 );
buf ( n389282 , n389101 );
not ( n41788 , n389282 );
or ( n41789 , n41786 , n41788 );
buf ( n389285 , n24050 );
not ( n41791 , n389285 );
buf ( n389287 , n37411 );
not ( n41793 , n389287 );
buf ( n389289 , n41793 );
buf ( n389290 , n389289 );
not ( n41796 , n389290 );
or ( n41797 , n41791 , n41796 );
buf ( n389293 , n36709 );
buf ( n389294 , n389075 );
nand ( n41800 , n389293 , n389294 );
buf ( n389296 , n41800 );
buf ( n389297 , n389296 );
nand ( n41803 , n41797 , n389297 );
buf ( n389299 , n41803 );
buf ( n389300 , n389299 );
buf ( n389301 , n389125 );
nand ( n41807 , n389300 , n389301 );
buf ( n389303 , n41807 );
buf ( n389304 , n389303 );
nand ( n41810 , n41789 , n389304 );
buf ( n389306 , n41810 );
buf ( n389307 , n389306 );
buf ( n389308 , n388502 );
not ( n41814 , n389308 );
buf ( n389310 , n385972 );
not ( n41816 , n389310 );
or ( n41817 , n41814 , n41816 );
buf ( n389313 , n31963 );
buf ( n389314 , n388511 );
nand ( n41820 , n389313 , n389314 );
buf ( n389316 , n41820 );
buf ( n389317 , n389316 );
nand ( n41823 , n41817 , n389317 );
buf ( n389319 , n41823 );
buf ( n389320 , n389319 );
not ( n41826 , n389320 );
buf ( n389322 , n382595 );
not ( n41828 , n389322 );
or ( n41829 , n41826 , n41828 );
buf ( n389325 , n389010 );
buf ( n389326 , n379460 );
not ( n41832 , n389326 );
buf ( n389328 , n41832 );
buf ( n389329 , n389328 );
nand ( n41835 , n389325 , n389329 );
buf ( n389331 , n41835 );
buf ( n389332 , n389331 );
nand ( n41838 , n41829 , n389332 );
buf ( n389334 , n41838 );
buf ( n389335 , n389334 );
buf ( n389336 , n372527 );
buf ( n41842 , n389336 );
buf ( n389338 , n41842 );
buf ( n389339 , n389338 );
buf ( n41845 , n389339 );
buf ( n389341 , n41845 );
and ( n41847 , n389341 , n384096 );
not ( n41848 , n389341 );
and ( n41849 , n41848 , n385328 );
or ( n41850 , n41847 , n41849 );
buf ( n389346 , n382938 );
not ( n41858 , n389346 );
buf ( n389348 , n41858 );
buf ( n389349 , n389348 );
buf ( n41861 , n376029 );
buf ( n389351 , n41861 );
not ( n41863 , n389351 );
buf ( n389353 , n41863 );
buf ( n389354 , n389353 );
buf ( n41866 , n389354 );
buf ( n389356 , n41866 );
buf ( n389357 , n389356 );
not ( n41869 , n389357 );
buf ( n389359 , n41869 );
buf ( n389360 , n389359 );
not ( n41872 , n389360 );
buf ( n389362 , n384096 );
not ( n41874 , n389362 );
or ( n41875 , n41872 , n41874 );
buf ( n389365 , n385292 );
buf ( n389366 , n389356 );
nand ( n389367 , n389365 , n389366 );
buf ( n389368 , n389367 );
buf ( n389369 , n389368 );
nand ( n41881 , n41875 , n389369 );
buf ( n389371 , n41881 );
not ( n41883 , n389371 );
buf ( n389373 , n41883 );
or ( n41885 , n389349 , n389373 );
nand ( n41886 , C1 , n41885 );
buf ( n389376 , n41886 );
buf ( n389377 , n389376 );
xor ( n41889 , n389335 , n389377 );
buf ( n389379 , n386480 );
not ( n41891 , n389379 );
buf ( n389381 , n38155 );
buf ( n389382 , n38971 );
nand ( n41894 , n389381 , n389382 );
buf ( n389384 , n41894 );
not ( n41896 , n38155 );
nand ( n41897 , n22982 , n41896 );
nand ( n41898 , n389384 , n41897 );
buf ( n389388 , n41898 );
not ( n41900 , n389388 );
or ( n41901 , n41891 , n41900 );
buf ( n389391 , n22982 );
not ( n41903 , n389391 );
not ( n41904 , n37763 );
buf ( n389394 , n41904 );
not ( n41906 , n389394 );
or ( n41907 , n41903 , n41906 );
not ( n41908 , n38972 );
nand ( n41909 , n41908 , n385324 );
buf ( n389399 , n41909 );
nand ( n41911 , n41907 , n389399 );
buf ( n389401 , n41911 );
buf ( n389402 , n389401 );
buf ( n389403 , n386496 );
nand ( n41915 , n389402 , n389403 );
buf ( n389405 , n41915 );
buf ( n389406 , n389405 );
nand ( n41918 , n41901 , n389406 );
buf ( n389408 , n41918 );
buf ( n389409 , n389408 );
and ( n41921 , n41889 , n389409 );
and ( n41922 , n389335 , n389377 );
or ( n41923 , n41921 , n41922 );
buf ( n389413 , n41923 );
buf ( n389414 , n389413 );
xor ( n41926 , n389307 , n389414 );
buf ( n389416 , n388833 );
not ( n41928 , n389416 );
buf ( n389418 , n36897 );
not ( n41930 , n389418 );
buf ( n389420 , n41930 );
buf ( n389421 , n389420 );
not ( n41933 , n389421 );
buf ( n389423 , n41933 );
xnor ( n41935 , n389423 , n41349 );
buf ( n389425 , n41935 );
not ( n41937 , n389425 );
or ( n41938 , n41928 , n41937 );
buf ( n389428 , n41342 );
not ( n41940 , n389428 );
buf ( n389430 , n37147 );
not ( n41942 , n389430 );
or ( n41943 , n41940 , n41942 );
buf ( n389433 , n38356 );
not ( n41945 , n389433 );
buf ( n389435 , n41945 );
buf ( n389436 , n389435 );
buf ( n389437 , n41349 );
nand ( n41949 , n389436 , n389437 );
buf ( n389439 , n41949 );
buf ( n389440 , n389439 );
nand ( n41952 , n41943 , n389440 );
buf ( n389442 , n41952 );
buf ( n389443 , n389442 );
buf ( n389444 , n388872 );
nand ( n41956 , n389443 , n389444 );
buf ( n389446 , n41956 );
buf ( n389447 , n389446 );
nand ( n41959 , n41938 , n389447 );
buf ( n389449 , n41959 );
buf ( n389450 , n389449 );
and ( n41962 , n41926 , n389450 );
and ( n41963 , n389307 , n389414 );
or ( n41964 , n41962 , n41963 );
buf ( n389454 , n41964 );
buf ( n389455 , n389454 );
nand ( n41967 , n41784 , n389455 );
buf ( n389457 , n41967 );
buf ( n389458 , n389457 );
nand ( n41970 , n41781 , n389458 );
buf ( n389460 , n41970 );
buf ( n389461 , n386480 );
not ( n41973 , n389461 );
buf ( n389463 , n22982 );
not ( n41975 , n389463 );
buf ( n389465 , n37411 );
not ( n41977 , n389465 );
buf ( n389467 , n41977 );
buf ( n389468 , n389467 );
not ( n41980 , n389468 );
or ( n41981 , n41975 , n41980 );
buf ( n389471 , n36709 );
buf ( n389472 , n38971 );
nand ( n41984 , n389471 , n389472 );
buf ( n389474 , n41984 );
buf ( n389475 , n389474 );
nand ( n41987 , n41981 , n389475 );
buf ( n389477 , n41987 );
buf ( n389478 , n389477 );
not ( n41990 , n389478 );
or ( n41991 , n41973 , n41990 );
buf ( n389481 , n38972 );
not ( n41993 , n389481 );
buf ( n389483 , n384092 );
not ( n41995 , n389483 );
buf ( n389485 , n41995 );
buf ( n389486 , n389485 );
not ( n41998 , n389486 );
or ( n41999 , n41993 , n41998 );
buf ( n389489 , n385983 );
buf ( n389490 , n38971 );
nand ( n42002 , n389489 , n389490 );
buf ( n389492 , n42002 );
buf ( n389493 , n389492 );
nand ( n42005 , n41999 , n389493 );
buf ( n389495 , n42005 );
buf ( n389496 , n389495 );
buf ( n389497 , n386496 );
nand ( n42009 , n389496 , n389497 );
buf ( n389499 , n42009 );
buf ( n389500 , n389499 );
nand ( n42012 , n41991 , n389500 );
buf ( n389502 , n42012 );
buf ( n389503 , n389502 );
buf ( n389504 , n388141 );
not ( n42016 , n389504 );
buf ( n389506 , n388160 );
not ( n42018 , n389506 );
buf ( n389508 , n38357 );
not ( n42020 , n389508 );
or ( n42021 , n42018 , n42020 );
buf ( n389511 , n389435 );
buf ( n389512 , n388157 );
nand ( n42024 , n389511 , n389512 );
buf ( n389514 , n42024 );
buf ( n389515 , n389514 );
nand ( n42027 , n42021 , n389515 );
buf ( n389517 , n42027 );
buf ( n389518 , n389517 );
not ( n42030 , n389518 );
or ( n42031 , n42016 , n42030 );
buf ( n389521 , n388160 );
not ( n42033 , n389521 );
buf ( n389523 , n37173 );
not ( n42035 , n389523 );
buf ( n389525 , n42035 );
buf ( n389526 , n389525 );
not ( n42038 , n389526 );
or ( n42039 , n42033 , n42038 );
buf ( n389529 , n37173 );
buf ( n389530 , n388157 );
nand ( n42042 , n389529 , n389530 );
buf ( n389532 , n42042 );
buf ( n389533 , n389532 );
nand ( n42045 , n42039 , n389533 );
buf ( n389535 , n42045 );
buf ( n389536 , n389535 );
buf ( n389537 , n40701 );
nand ( n42049 , n389536 , n389537 );
buf ( n389539 , n42049 );
buf ( n389540 , n389539 );
nand ( n42052 , n42031 , n389540 );
buf ( n389542 , n42052 );
buf ( n389543 , n389542 );
xor ( n42055 , n389503 , n389543 );
buf ( n389545 , n382938 );
buf ( n42062 , n389545 );
buf ( n389547 , n42062 );
buf ( n389548 , n389547 );
not ( n42065 , n375993 );
not ( n42066 , n42065 );
buf ( n389551 , n42066 );
not ( n42068 , n389551 );
buf ( n389553 , n384143 );
not ( n42070 , n389553 );
or ( n42071 , n42068 , n42070 );
buf ( n389556 , n382854 );
buf ( n42073 , n28390 );
not ( n42074 , n42073 );
buf ( n389559 , n42074 );
nand ( n42076 , n389556 , n389559 );
buf ( n389561 , n42076 );
buf ( n389562 , n389561 );
nand ( n42079 , n42071 , n389562 );
buf ( n389564 , n42079 );
buf ( n389565 , n389564 );
nand ( n42082 , n389548 , n389565 );
buf ( n389567 , n42082 );
buf ( n389568 , n389567 );
nand ( n42085 , C1 , n389568 );
buf ( n389570 , n42085 );
buf ( n389571 , n389570 );
buf ( n389572 , n386480 );
not ( n42089 , n389572 );
buf ( n389574 , n389495 );
not ( n42091 , n389574 );
or ( n42092 , n42089 , n42091 );
not ( n42093 , n41897 );
not ( n42094 , n389384 );
or ( n42095 , n42093 , n42094 );
nand ( n42096 , n42095 , n386496 );
buf ( n389581 , n42096 );
nand ( n42098 , n42092 , n389581 );
buf ( n389583 , n42098 );
buf ( n389584 , n389583 );
xor ( n42101 , n389571 , n389584 );
buf ( n389586 , n383476 );
buf ( n389587 , n388576 );
not ( n42104 , n389587 );
buf ( n389589 , n42104 );
buf ( n389590 , n389589 );
buf ( n389591 , n12471 );
not ( n42108 , n389591 );
buf ( n389593 , n42108 );
buf ( n389594 , n389593 );
and ( n42111 , n389590 , n389594 );
buf ( n389596 , n388556 );
not ( n42113 , n389596 );
buf ( n389598 , n42113 );
buf ( n389599 , n389598 );
buf ( n389600 , n389593 );
not ( n42117 , n389600 );
buf ( n389602 , n42117 );
buf ( n389603 , n389602 );
and ( n42120 , n389599 , n389603 );
nor ( n42121 , n42111 , n42120 );
buf ( n389606 , n42121 );
buf ( n389607 , n389606 );
or ( n42124 , n389586 , n389607 );
buf ( n389609 , n388560 );
buf ( n389610 , n383403 );
or ( n42127 , n389609 , n389610 );
nand ( n42128 , n42124 , n42127 );
buf ( n389613 , n42128 );
buf ( n389614 , n389613 );
and ( n42131 , n42101 , n389614 );
and ( n42132 , n389571 , n389584 );
or ( n42133 , n42131 , n42132 );
buf ( n389618 , n42133 );
buf ( n389619 , n389618 );
xor ( n42136 , n42055 , n389619 );
buf ( n389621 , n42136 );
not ( n42138 , n389621 );
xor ( n42139 , n389049 , n389132 );
xor ( n42140 , n42139 , n389137 );
buf ( n389625 , n42140 );
not ( n42142 , n389625 );
or ( n42143 , n42138 , n42142 );
or ( n42144 , n389621 , n389625 );
xor ( n42145 , n388941 , n388994 );
xor ( n42146 , n42145 , n389044 );
buf ( n389631 , n42146 );
buf ( n389632 , n389631 );
buf ( n389633 , n40701 );
not ( n42150 , n389633 );
not ( n42151 , n388160 );
buf ( n42152 , n36187 );
not ( n42153 , n42152 );
not ( n42154 , n42153 );
or ( n42155 , n42151 , n42154 );
buf ( n389640 , n36188 );
buf ( n389641 , n388157 );
nand ( n42158 , n389640 , n389641 );
buf ( n389643 , n42158 );
nand ( n42160 , n42155 , n389643 );
buf ( n389645 , n42160 );
not ( n42162 , n389645 );
or ( n42163 , n42150 , n42162 );
buf ( n389648 , n389535 );
buf ( n389649 , n388141 );
nand ( n42166 , n389648 , n389649 );
buf ( n389651 , n42166 );
buf ( n389652 , n389651 );
nand ( n42169 , n42163 , n389652 );
buf ( n389654 , n42169 );
buf ( n389655 , n389654 );
or ( n42172 , n389632 , n389655 );
xor ( n42173 , n389571 , n389584 );
xor ( n42174 , n42173 , n389614 );
buf ( n389659 , n42174 );
buf ( n389660 , n389659 );
nand ( n42177 , n42172 , n389660 );
buf ( n389662 , n42177 );
buf ( n389663 , n389662 );
buf ( n389664 , n389654 );
buf ( n389665 , n389631 );
nand ( n42182 , n389664 , n389665 );
buf ( n389667 , n42182 );
buf ( n389668 , n389667 );
nand ( n42185 , n389663 , n389668 );
buf ( n389670 , n42185 );
nand ( n42187 , n42144 , n389670 );
nand ( n42188 , n42143 , n42187 );
xor ( n42189 , n389460 , n42188 );
xor ( n42190 , n389503 , n389543 );
and ( n42191 , n42190 , n389619 );
and ( n42192 , n389503 , n389543 );
or ( n42193 , n42191 , n42192 );
buf ( n389678 , n42193 );
buf ( n389679 , n389678 );
buf ( n389680 , n386496 );
not ( n42197 , n389680 );
buf ( n389682 , n389477 );
not ( n42199 , n389682 );
or ( n42200 , n42197 , n42199 );
buf ( n389685 , n22982 );
not ( n42202 , n389685 );
buf ( n389687 , n384239 );
not ( n42204 , n389687 );
or ( n42205 , n42202 , n42204 );
buf ( n389690 , n36668 );
buf ( n42207 , n389690 );
buf ( n389692 , n42207 );
buf ( n389693 , n389692 );
buf ( n389694 , n38971 );
nand ( n42211 , n389693 , n389694 );
buf ( n389696 , n42211 );
buf ( n389697 , n389696 );
nand ( n42214 , n42205 , n389697 );
buf ( n389699 , n42214 );
buf ( n389700 , n389699 );
buf ( n389701 , n386480 );
nand ( n42218 , n389700 , n389701 );
buf ( n389703 , n42218 );
buf ( n389704 , n389703 );
nand ( n42221 , n42200 , n389704 );
buf ( n389706 , n42221 );
buf ( n389707 , n389706 );
buf ( n389708 , n389125 );
not ( n42225 , n389708 );
buf ( n389710 , n389081 );
not ( n42227 , n389710 );
or ( n42228 , n42225 , n42227 );
buf ( n389713 , n24050 );
not ( n42230 , n389713 );
buf ( n389715 , n36218 );
not ( n42232 , n389715 );
or ( n42233 , n42230 , n42232 );
not ( n42234 , n36216 );
buf ( n389719 , n42234 );
not ( n42236 , n389719 );
buf ( n389721 , n389075 );
nand ( n42238 , n42236 , n389721 );
buf ( n389723 , n42238 );
buf ( n389724 , n389723 );
nand ( n42241 , n42233 , n389724 );
buf ( n389726 , n42241 );
buf ( n389727 , n389726 );
buf ( n389728 , n41565 );
nand ( n42245 , n389727 , n389728 );
buf ( n389730 , n42245 );
buf ( n389731 , n389730 );
nand ( n42248 , n42228 , n389731 );
buf ( n389733 , n42248 );
buf ( n389734 , n389733 );
xor ( n42251 , n389707 , n389734 );
buf ( n389736 , n41445 );
not ( n42253 , n389736 );
buf ( n389738 , n42253 );
buf ( n389739 , n389738 );
buf ( n389740 , n389037 );
not ( n42257 , n389740 );
buf ( n389742 , n382589 );
not ( n42259 , n389742 );
buf ( n389744 , n42259 );
buf ( n389745 , n389744 );
not ( n42262 , n389745 );
or ( n42263 , n42257 , n42262 );
buf ( n389748 , n379463 );
buf ( n389749 , n389602 );
not ( n42266 , n389749 );
buf ( n389751 , n31963 );
not ( n42268 , n389751 );
buf ( n389753 , n42268 );
buf ( n389754 , n389753 );
not ( n42271 , n389754 );
or ( n42272 , n42266 , n42271 );
buf ( n389757 , n382994 );
not ( n42274 , n389757 );
buf ( n389759 , n42274 );
buf ( n389760 , n389759 );
buf ( n389761 , n389593 );
nand ( n42278 , n389760 , n389761 );
buf ( n389763 , n42278 );
buf ( n389764 , n389763 );
nand ( n42281 , n42272 , n389764 );
buf ( n389766 , n42281 );
buf ( n389767 , n389766 );
nand ( n42284 , n389748 , n389767 );
buf ( n389769 , n42284 );
buf ( n389770 , n389769 );
nand ( n42287 , n42263 , n389770 );
buf ( n389772 , n42287 );
buf ( n389773 , n389772 );
xor ( n42290 , n389739 , n389773 );
buf ( n389775 , n389547 );
not ( n42301 , n389775 );
buf ( n389777 , n42301 );
buf ( n389778 , n389777 );
buf ( n389779 , n388495 );
or ( n42305 , n389778 , n389779 );
nand ( n42306 , C1 , n42305 );
buf ( n389782 , n42306 );
buf ( n389783 , n389782 );
and ( n42309 , n42290 , n389783 );
and ( n42310 , n389739 , n389773 );
or ( n42311 , n42309 , n42310 );
buf ( n389787 , n42311 );
buf ( n389788 , n389787 );
xor ( n42314 , n42251 , n389788 );
buf ( n389790 , n42314 );
buf ( n389791 , n389790 );
xor ( n42317 , n389679 , n389791 );
buf ( n389793 , n37316 );
not ( n42319 , n389793 );
buf ( n389795 , n37347 );
not ( n42321 , n389795 );
buf ( n389797 , n385345 );
not ( n42323 , n389797 );
or ( n42324 , n42321 , n42323 );
buf ( n389800 , n29077 );
not ( n42326 , n389800 );
buf ( n389802 , n42326 );
buf ( n389803 , n389802 );
buf ( n42329 , n389803 );
buf ( n389805 , n42329 );
buf ( n389806 , n389805 );
not ( n42332 , n389806 );
buf ( n389808 , n42332 );
buf ( n389809 , n389808 );
buf ( n389810 , n37346 );
nand ( n42336 , n389809 , n389810 );
buf ( n389812 , n42336 );
buf ( n389813 , n389812 );
nand ( n42339 , n42324 , n389813 );
buf ( n389815 , n42339 );
buf ( n389816 , n389815 );
not ( n42342 , n389816 );
or ( n42343 , n42319 , n42342 );
buf ( n389819 , n388935 );
not ( n42345 , n389819 );
buf ( n389821 , n385269 );
nand ( n42347 , n42345 , n389821 );
buf ( n389823 , n42347 );
buf ( n389824 , n389823 );
nand ( n42350 , n42343 , n389824 );
buf ( n389826 , n42350 );
buf ( n389827 , n389826 );
buf ( n389828 , n41447 );
not ( n42354 , n389828 );
buf ( n389830 , n385494 );
not ( n42356 , n389830 );
buf ( n389832 , n36565 );
not ( n42358 , n389832 );
or ( n42359 , n42356 , n42358 );
buf ( n389835 , n38155 );
buf ( n389836 , n385491 );
nand ( n42362 , n389835 , n389836 );
buf ( n389838 , n42362 );
buf ( n389839 , n389838 );
nand ( n42365 , n42359 , n389839 );
buf ( n389841 , n42365 );
buf ( n389842 , n389841 );
not ( n42368 , n389842 );
or ( n42369 , n42354 , n42368 );
buf ( n389845 , n388971 );
buf ( n389846 , n385479 );
nand ( n42372 , n389845 , n389846 );
buf ( n389848 , n42372 );
buf ( n389849 , n389848 );
nand ( n42375 , n42369 , n389849 );
buf ( n389851 , n42375 );
buf ( n389852 , n389851 );
xor ( n42378 , n389827 , n389852 );
buf ( n389854 , n28297 );
not ( n42380 , n389854 );
buf ( n389856 , n42380 );
buf ( n389857 , n389856 );
buf ( n42383 , n389857 );
buf ( n389859 , n42383 );
buf ( n389860 , n389859 );
not ( n42386 , n389860 );
buf ( n389862 , n42386 );
buf ( n389863 , n389862 );
not ( n42389 , n389863 );
buf ( n42390 , n35797 );
buf ( n389866 , n42390 );
not ( n42392 , n389866 );
or ( n42393 , n42389 , n42392 );
buf ( n389869 , n37037 );
buf ( n389870 , n389859 );
nand ( n42396 , n389869 , n389870 );
buf ( n389872 , n42396 );
buf ( n389873 , n389872 );
nand ( n42399 , n42393 , n389873 );
buf ( n389875 , n42399 );
buf ( n389876 , n389875 );
not ( n42402 , n389876 );
buf ( n389878 , n384618 );
not ( n42404 , n389878 );
buf ( n389880 , n42404 );
buf ( n389881 , n389880 );
buf ( n42407 , n389881 );
buf ( n389883 , n42407 );
buf ( n389884 , n389883 );
not ( n42410 , n389884 );
or ( n42411 , n42402 , n42410 );
buf ( n389887 , n388646 );
not ( n42413 , n389887 );
buf ( n389889 , n384562 );
not ( n42415 , n389889 );
or ( n42416 , n42413 , n42415 );
buf ( n389892 , n35797 );
not ( n42418 , n389892 );
buf ( n389894 , n42418 );
buf ( n389895 , n389894 );
buf ( n42421 , n389895 );
buf ( n389897 , n42421 );
buf ( n389898 , n389897 );
buf ( n389899 , n388654 );
nand ( n42425 , n389898 , n389899 );
buf ( n389901 , n42425 );
buf ( n389902 , n389901 );
nand ( n42428 , n42416 , n389902 );
buf ( n389904 , n42428 );
buf ( n389905 , n389904 );
buf ( n389906 , n384551 );
not ( n42432 , n389906 );
buf ( n389908 , n42432 );
buf ( n389909 , n389908 );
nand ( n42435 , n389905 , n389909 );
buf ( n389911 , n42435 );
buf ( n389912 , n389911 );
nand ( n42438 , n42411 , n389912 );
buf ( n389914 , n42438 );
buf ( n389915 , n389914 );
and ( n42441 , n42378 , n389915 );
and ( n42442 , n389827 , n389852 );
or ( n42443 , n42441 , n42442 );
buf ( n389919 , n42443 );
buf ( n389920 , n389919 );
buf ( n389921 , n40805 );
not ( n42447 , n389921 );
buf ( n389923 , n383894 );
not ( n42449 , n389923 );
or ( n42450 , n42447 , n42449 );
buf ( n389926 , n36251 );
not ( n42452 , n389926 );
buf ( n389928 , n42452 );
buf ( n389929 , n389928 );
not ( n42455 , n389929 );
buf ( n389931 , n388919 );
not ( n42457 , n389931 );
or ( n42458 , n42455 , n42457 );
buf ( n389934 , n388263 );
not ( n42460 , n389934 );
buf ( n389936 , n42460 );
buf ( n389937 , n389936 );
buf ( n389938 , n386176 );
not ( n42464 , n389938 );
buf ( n389940 , n42464 );
buf ( n389941 , n389940 );
nand ( n42467 , n389937 , n389941 );
buf ( n389943 , n42467 );
buf ( n389944 , n389943 );
nand ( n42470 , n42458 , n389944 );
buf ( n389946 , n42470 );
buf ( n389947 , n389946 );
buf ( n389948 , n383907 );
nand ( n42474 , n389947 , n389948 );
buf ( n389950 , n42474 );
buf ( n389951 , n389950 );
nand ( n42477 , n42450 , n389951 );
buf ( n389953 , n42477 );
buf ( n389954 , n389953 );
buf ( n42480 , n389954 );
buf ( n389956 , n42480 );
buf ( n389957 , n389956 );
buf ( n389958 , n37346 );
buf ( n389959 , n385324 );
and ( n42485 , n389958 , n389959 );
not ( n42486 , n389958 );
buf ( n389962 , n388952 );
not ( n42488 , n389962 );
buf ( n389964 , n42488 );
buf ( n389965 , n389964 );
and ( n42491 , n42486 , n389965 );
nor ( n42492 , n42485 , n42491 );
buf ( n389968 , n42492 );
buf ( n389969 , n389968 );
not ( n42495 , n389969 );
buf ( n389971 , n37317 );
not ( n42497 , n389971 );
and ( n42498 , n42495 , n42497 );
buf ( n389974 , n389815 );
buf ( n389975 , n385269 );
and ( n42501 , n389974 , n389975 );
nor ( n42502 , n42498 , n42501 );
buf ( n389978 , n42502 );
buf ( n389979 , n389978 );
not ( n42505 , n389979 );
buf ( n389981 , n42505 );
buf ( n389982 , n389981 );
xor ( n42508 , n389957 , n389982 );
buf ( n389984 , n389766 );
not ( n42510 , n389984 );
buf ( n389986 , n382598 );
not ( n42512 , n389986 );
or ( n42513 , n42510 , n42512 );
buf ( n389989 , n386212 );
buf ( n389990 , n388549 );
not ( n42516 , n389990 );
buf ( n389992 , n385972 );
not ( n42518 , n389992 );
or ( n42519 , n42516 , n42518 );
buf ( n389995 , n385987 );
not ( n42521 , n389995 );
buf ( n389997 , n42521 );
buf ( n389998 , n389997 );
buf ( n389999 , n388546 );
nand ( n42525 , n389998 , n389999 );
buf ( n390001 , n42525 );
buf ( n390002 , n390001 );
nand ( n390003 , n42519 , n390002 );
buf ( n390004 , n390003 );
buf ( n390005 , n390004 );
nand ( n42531 , n389989 , n390005 );
buf ( n390007 , n42531 );
buf ( n390008 , n390007 );
nand ( n42534 , n42513 , n390008 );
buf ( n390010 , n42534 );
buf ( n390011 , n390010 );
xnor ( n42537 , n42508 , n390011 );
buf ( n390013 , n42537 );
buf ( n390014 , n390013 );
xor ( n42540 , n389920 , n390014 );
buf ( n390016 , n40701 );
not ( n42542 , n390016 );
buf ( n390018 , n389517 );
not ( n42544 , n390018 );
or ( n42545 , n42542 , n42544 );
buf ( n390021 , n388141 );
buf ( n390022 , n388187 );
nand ( n42548 , n390021 , n390022 );
buf ( n390024 , n42548 );
buf ( n390025 , n390024 );
nand ( n42551 , n42545 , n390025 );
buf ( n390027 , n42551 );
buf ( n390028 , n390027 );
xor ( n42554 , n42540 , n390028 );
buf ( n390030 , n42554 );
buf ( n390031 , n390030 );
xor ( n42557 , n42317 , n390031 );
buf ( n390033 , n42557 );
and ( n42559 , n42189 , n390033 );
and ( n42560 , n389460 , n42188 );
or ( n42561 , n42559 , n42560 );
xor ( n42562 , n389220 , n42561 );
buf ( n390038 , n389678 );
not ( n42564 , n390038 );
buf ( n390040 , n389790 );
not ( n42566 , n390040 );
or ( n42567 , n42564 , n42566 );
or ( n42568 , n389790 , n389678 );
nand ( n42569 , n42568 , n390030 );
buf ( n390045 , n42569 );
nand ( n42571 , n42567 , n390045 );
buf ( n390047 , n42571 );
buf ( n390048 , n390047 );
xor ( n42574 , n389707 , n389734 );
and ( n42575 , n42574 , n389788 );
and ( n42576 , n389707 , n389734 );
or ( n42577 , n42575 , n42576 );
buf ( n390053 , n42577 );
buf ( n390054 , n390053 );
buf ( n390055 , n41711 );
not ( n42581 , n390055 );
buf ( n390057 , n389179 );
not ( n42583 , n390057 );
or ( n42584 , n42581 , n42583 );
buf ( n390060 , n41671 );
not ( n42586 , n390060 );
buf ( n390062 , n386421 );
not ( n42588 , n390062 );
or ( n42589 , n42586 , n42588 );
buf ( n390065 , n386418 );
buf ( n390066 , n41670 );
nand ( n42592 , n390065 , n390066 );
buf ( n390068 , n42592 );
buf ( n390069 , n390068 );
nand ( n42595 , n42589 , n390069 );
buf ( n390071 , n42595 );
buf ( n390072 , n390071 );
buf ( n390073 , n389162 );
nand ( n42599 , n390072 , n390073 );
buf ( n390075 , n42599 );
buf ( n390076 , n390075 );
nand ( n42602 , n42584 , n390076 );
buf ( n390078 , n42602 );
buf ( n390079 , n390078 );
xor ( n42605 , n390054 , n390079 );
xor ( n42606 , n389920 , n390014 );
and ( n42607 , n42606 , n390028 );
and ( n42608 , n389920 , n390014 );
or ( n42609 , n42607 , n42608 );
buf ( n390085 , n42609 );
buf ( n390086 , n390085 );
xor ( n42612 , n42605 , n390086 );
buf ( n390088 , n42612 );
buf ( n390089 , n390088 );
xor ( n42615 , n390048 , n390089 );
not ( n42616 , n35300 );
xnor ( n42617 , n41342 , n42616 );
buf ( n390093 , n42617 );
buf ( n390094 , n388833 );
and ( n42620 , n390093 , n390094 );
buf ( n390096 , n388850 );
not ( n42622 , n390096 );
buf ( n390098 , n41374 );
nor ( n42624 , n42622 , n390098 );
buf ( n390100 , n42624 );
buf ( n390101 , n390100 );
nor ( n42627 , n42620 , n390101 );
buf ( n390103 , n42627 );
or ( n42629 , n40958 , n388482 );
nand ( n42630 , n388524 , n42629 );
and ( n42631 , n388457 , n388483 );
buf ( n390107 , n42631 );
not ( n42633 , n390107 );
nand ( n42634 , n42630 , n42633 );
buf ( n390110 , n42634 );
not ( n42636 , n390110 );
buf ( n390112 , n38972 );
not ( n42638 , n390112 );
buf ( n390114 , n389067 );
not ( n42640 , n390114 );
or ( n42641 , n42638 , n42640 );
buf ( n390117 , n384202 );
not ( n42643 , n390117 );
buf ( n390119 , n42643 );
buf ( n390120 , n390119 );
buf ( n390121 , n38971 );
nand ( n42647 , n390120 , n390121 );
buf ( n390123 , n42647 );
buf ( n390124 , n390123 );
nand ( n42650 , n42641 , n390124 );
buf ( n390126 , n42650 );
buf ( n390127 , n390126 );
buf ( n390128 , n386480 );
and ( n42654 , n390127 , n390128 );
buf ( n390130 , n389699 );
not ( n42656 , n390130 );
buf ( n390132 , n386499 );
nor ( n42658 , n42656 , n390132 );
buf ( n390134 , n42658 );
buf ( n390135 , n390134 );
nor ( n42661 , n42654 , n390135 );
buf ( n390137 , n42661 );
buf ( n390138 , n390137 );
buf ( n390139 , n389956 );
not ( n42665 , n390139 );
buf ( n390141 , n389978 );
not ( n42667 , n390141 );
or ( n42668 , n42665 , n42667 );
buf ( n390144 , n390010 );
nand ( n42670 , n42668 , n390144 );
buf ( n390146 , n42670 );
buf ( n390147 , n390146 );
buf ( n390148 , n389956 );
not ( n42674 , n390148 );
buf ( n390150 , n389981 );
nand ( n42676 , n42674 , n390150 );
buf ( n390152 , n42676 );
buf ( n390153 , n390152 );
nand ( n42679 , n390147 , n390153 );
buf ( n390155 , n42679 );
buf ( n390156 , n390155 );
xor ( n42682 , n390138 , n390156 );
buf ( n390158 , n42682 );
buf ( n390159 , n390158 );
not ( n42685 , n390159 );
or ( n42686 , n42636 , n42685 );
buf ( n390162 , n390158 );
buf ( n390163 , n42634 );
or ( n42689 , n390162 , n390163 );
nand ( n42690 , n42686 , n42689 );
buf ( n390166 , n42690 );
xor ( n42692 , n390103 , n390166 );
buf ( n390168 , n385494 );
not ( n42694 , n390168 );
buf ( n390170 , n37411 );
not ( n42696 , n390170 );
buf ( n390172 , n42696 );
buf ( n390173 , n390172 );
not ( n42699 , n390173 );
or ( n42700 , n42694 , n42699 );
buf ( n390176 , n389289 );
not ( n42702 , n390176 );
buf ( n390178 , n42702 );
buf ( n390179 , n390178 );
buf ( n390180 , n385491 );
nand ( n42706 , n390179 , n390180 );
buf ( n390182 , n42706 );
buf ( n390183 , n390182 );
nand ( n42709 , n42700 , n390183 );
buf ( n390185 , n42709 );
buf ( n390186 , n390185 );
buf ( n390187 , n38324 );
and ( n42713 , n390186 , n390187 );
buf ( n390189 , n385494 );
not ( n42715 , n390189 );
buf ( n390191 , n384089 );
not ( n42717 , n390191 );
or ( n42718 , n42715 , n42717 );
buf ( n390194 , n36509 );
buf ( n390195 , n385491 );
nand ( n42721 , n390194 , n390195 );
buf ( n390197 , n42721 );
buf ( n390198 , n390197 );
nand ( n42724 , n42718 , n390198 );
buf ( n390200 , n42724 );
buf ( n390201 , n390200 );
not ( n42727 , n390201 );
buf ( n390203 , n385482 );
nor ( n42729 , n42727 , n390203 );
buf ( n390205 , n42729 );
buf ( n390206 , n390205 );
nor ( n42732 , n42713 , n390206 );
buf ( n390208 , n42732 );
buf ( n390209 , n390208 );
not ( n42735 , n390209 );
buf ( n390211 , n386300 );
not ( n42737 , n390211 );
buf ( n390213 , n42737 );
buf ( n390214 , n390213 );
not ( n42740 , n390214 );
buf ( n390216 , n388248 );
not ( n42742 , n390216 );
buf ( n390218 , n42742 );
buf ( n390219 , n390218 );
not ( n42745 , n390219 );
and ( n42746 , n42740 , n42745 );
buf ( n390222 , n383134 );
buf ( n390223 , n389593 );
buf ( n390224 , n386223 );
and ( n42750 , n390223 , n390224 );
not ( n42751 , n390223 );
buf ( n390227 , n388235 );
and ( n42753 , n42751 , n390227 );
nor ( n42754 , n42750 , n42753 );
buf ( n390230 , n42754 );
buf ( n390231 , n390230 );
nor ( n42757 , n390222 , n390231 );
buf ( n390233 , n42757 );
buf ( n390234 , n390233 );
nor ( n42760 , n42746 , n390234 );
buf ( n390236 , n42760 );
buf ( n390237 , n390236 );
not ( n42763 , n390237 );
buf ( n390239 , n42763 );
buf ( n390240 , n390239 );
not ( n42766 , n390240 );
or ( n42767 , n42735 , n42766 );
buf ( n390243 , n390208 );
not ( n42769 , n390243 );
buf ( n390245 , n42769 );
buf ( n390246 , n390245 );
buf ( n390247 , n390236 );
nand ( n42773 , n390246 , n390247 );
buf ( n390249 , n42773 );
buf ( n390250 , n390249 );
nand ( n42776 , n42767 , n390250 );
buf ( n390252 , n42776 );
buf ( n390253 , n390252 );
buf ( n390254 , n389953 );
not ( n42780 , n40980 );
buf ( n390256 , n42780 );
not ( n42782 , n390256 );
buf ( n390258 , n384008 );
not ( n42784 , n390258 );
buf ( n390260 , n42784 );
buf ( n390261 , n390260 );
not ( n42787 , n390261 );
or ( n42788 , n42782 , n42787 );
buf ( n390264 , n40840 );
not ( n42790 , n390264 );
buf ( n390266 , n386150 );
not ( n42792 , n390266 );
or ( n42793 , n42790 , n42792 );
buf ( n390269 , n386150 );
buf ( n42795 , n390269 );
buf ( n390271 , n42795 );
buf ( n390272 , n390271 );
not ( n42798 , n390272 );
not ( n42799 , n40840 );
buf ( n390275 , n42799 );
nand ( n42801 , n42798 , n390275 );
buf ( n390277 , n42801 );
buf ( n390278 , n390277 );
nand ( n42804 , n42793 , n390278 );
buf ( n390280 , n42804 );
buf ( n390281 , n390280 );
buf ( n390282 , n388346 );
nand ( n42808 , n390281 , n390282 );
buf ( n390284 , n42808 );
buf ( n390285 , n390284 );
nand ( n42811 , n42788 , n390285 );
buf ( n390287 , n42811 );
buf ( n390288 , n390287 );
xor ( n42814 , n390254 , n390288 );
buf ( n390290 , n40858 );
not ( n42816 , n390290 );
buf ( n390292 , n42816 );
buf ( n390293 , n390292 );
buf ( n390294 , n388451 );
not ( n42820 , n390294 );
buf ( n390296 , n42820 );
buf ( n390297 , n390296 );
or ( n42823 , n390293 , n390297 );
buf ( n390299 , n388402 );
not ( n42825 , n40831 );
buf ( n390301 , n42825 );
buf ( n390302 , n388419 );
and ( n42828 , n390301 , n390302 );
not ( n42829 , n390301 );
buf ( n390305 , n388419 );
not ( n42831 , n390305 );
buf ( n390307 , n42831 );
buf ( n390308 , n390307 );
and ( n42834 , n42829 , n390308 );
nor ( n42835 , n42828 , n42834 );
buf ( n390311 , n42835 );
buf ( n390312 , n390311 );
or ( n42838 , n390299 , n390312 );
nand ( n42839 , n42823 , n42838 );
buf ( n390315 , n42839 );
buf ( n390316 , n390315 );
xor ( n42842 , n42814 , n390316 );
buf ( n390318 , n42842 );
buf ( n390319 , n390318 );
xnor ( n42845 , n390253 , n390319 );
buf ( n390321 , n42845 );
xor ( n42847 , n42692 , n390321 );
buf ( n390323 , n42847 );
xor ( n42849 , n42615 , n390323 );
buf ( n390325 , n42849 );
xor ( n42851 , n42562 , n390325 );
not ( n42852 , n42851 );
buf ( n390328 , n388105 );
buf ( n390329 , n35519 );
and ( n42855 , n390328 , n390329 );
not ( n42856 , n390328 );
buf ( n390332 , n383108 );
and ( n42858 , n42856 , n390332 );
nor ( n42859 , n42855 , n42858 );
buf ( n390335 , n42859 );
buf ( n390336 , n390335 );
not ( n42862 , n390336 );
buf ( n390338 , n388093 );
not ( n42864 , n390338 );
and ( n42865 , n42862 , n42864 );
buf ( n390341 , n388105 );
not ( n42867 , n390341 );
buf ( n390343 , n382526 );
not ( n42869 , n390343 );
buf ( n390345 , n42869 );
buf ( n390346 , n390345 );
not ( n42872 , n390346 );
or ( n42873 , n42867 , n42872 );
buf ( n390349 , n390345 );
not ( n42875 , n390349 );
buf ( n390351 , n42875 );
buf ( n390352 , n390351 );
buf ( n390353 , n388102 );
nand ( n42879 , n390352 , n390353 );
buf ( n390355 , n42879 );
buf ( n390356 , n390355 );
nand ( n42882 , n42873 , n390356 );
buf ( n390358 , n42882 );
buf ( n390359 , n390358 );
buf ( n390360 , n388071 );
not ( n42886 , n390360 );
buf ( n390362 , n42886 );
buf ( n390363 , n390362 );
and ( n42889 , n390359 , n390363 );
nor ( n42890 , n42865 , n42889 );
buf ( n390366 , n42890 );
buf ( n390367 , n390366 );
not ( n42893 , n390367 );
buf ( n390369 , n24074 );
not ( n42895 , n390369 );
buf ( n390371 , n36187 );
not ( n42897 , n390371 );
buf ( n390373 , n42897 );
buf ( n390374 , n390373 );
not ( n42900 , n390374 );
or ( n42901 , n42895 , n42900 );
buf ( n390377 , n390373 );
not ( n42903 , n390377 );
buf ( n390379 , n42903 );
buf ( n390380 , n390379 );
buf ( n390381 , n24073 );
nand ( n42907 , n390380 , n390381 );
buf ( n390383 , n42907 );
buf ( n390384 , n390383 );
nand ( n42910 , n42901 , n390384 );
buf ( n390386 , n42910 );
buf ( n390387 , n371522 );
not ( n42913 , n390387 );
buf ( n390389 , n42913 );
and ( n42915 , n388192 , n390389 );
not ( n42916 , n388192 );
buf ( n390392 , n23912 );
buf ( n390393 , n23915 );
xnor ( n42919 , n390392 , n390393 );
buf ( n390395 , n42919 );
and ( n42921 , n42916 , n390395 );
nor ( n42922 , n42915 , n42921 );
buf ( n42923 , n42922 );
not ( n42924 , n42923 );
not ( n42925 , n42924 );
buf ( n390401 , n42925 );
not ( n42927 , n390401 );
buf ( n390403 , n42927 );
and ( n42929 , n390386 , n390403 );
buf ( n390405 , n24074 );
not ( n42931 , n390405 );
buf ( n390407 , n37215 );
not ( n42933 , n390407 );
or ( n42934 , n42931 , n42933 );
buf ( n390410 , n36216 );
buf ( n390411 , n24073 );
nand ( n42937 , n390410 , n390411 );
buf ( n390413 , n42937 );
buf ( n390414 , n390413 );
nand ( n42940 , n42934 , n390414 );
buf ( n390416 , n42940 );
not ( n42942 , n390416 );
and ( n42943 , n24069 , n390395 );
not ( n42944 , n24069 );
buf ( n390420 , n390395 );
not ( n42946 , n390420 );
buf ( n390422 , n42946 );
and ( n42948 , n42944 , n390422 );
nor ( n42949 , n42943 , n42948 );
nand ( n42950 , n42949 , n42922 );
buf ( n42951 , n42950 );
buf ( n390427 , n42951 );
not ( n42953 , n390427 );
buf ( n390429 , n42953 );
buf ( n390430 , n390429 );
buf ( n42956 , n390430 );
buf ( n390432 , n42956 );
buf ( n390433 , n390432 );
not ( n42959 , n390433 );
buf ( n390435 , n42959 );
nor ( n42961 , n42942 , n390435 );
nor ( n42962 , n42929 , n42961 );
buf ( n390438 , n42962 );
not ( n42964 , n390438 );
buf ( n390440 , n42964 );
buf ( n390441 , n390440 );
not ( n42967 , n390441 );
or ( n42968 , n42893 , n42967 );
buf ( n390444 , n390440 );
buf ( n390445 , n390366 );
or ( n42971 , n390444 , n390445 );
nand ( n42972 , n42968 , n42971 );
buf ( n390448 , n42972 );
buf ( n390449 , n40990 );
not ( n42975 , n390449 );
buf ( n390451 , n35435 );
not ( n42977 , n390451 );
buf ( n390453 , n42977 );
buf ( n390454 , n390453 );
not ( n42980 , n390454 );
or ( n42981 , n42975 , n42980 );
buf ( n390457 , n35435 );
buf ( n390458 , n40990 );
not ( n42984 , n390458 );
buf ( n390460 , n42984 );
buf ( n390461 , n390460 );
nand ( n42987 , n390457 , n390461 );
buf ( n390463 , n42987 );
buf ( n390464 , n390463 );
nand ( n42990 , n42981 , n390464 );
buf ( n390466 , n42990 );
buf ( n390467 , n390466 );
not ( n42993 , n390467 );
buf ( n390469 , n383017 );
not ( n42995 , n390469 );
or ( n42996 , n42993 , n42995 );
buf ( n390472 , n388598 );
not ( n42998 , n390472 );
buf ( n390474 , n383134 );
not ( n43000 , n390474 );
buf ( n390476 , n43000 );
buf ( n390477 , n390476 );
nand ( n43003 , n42998 , n390477 );
buf ( n390479 , n43003 );
buf ( n390480 , n390479 );
nand ( n43006 , n42996 , n390480 );
buf ( n390482 , n43006 );
buf ( n390483 , n384621 );
not ( n43009 , n390483 );
buf ( n390485 , n43009 );
buf ( n390486 , n390485 );
not ( n43012 , n390486 );
buf ( n390488 , n388569 );
not ( n43014 , n390488 );
buf ( n390490 , n43014 );
buf ( n390491 , n390490 );
not ( n43017 , n390491 );
buf ( n390493 , n384562 );
not ( n43019 , n390493 );
or ( n43020 , n43017 , n43019 );
buf ( n390496 , n384562 );
not ( n43022 , n390496 );
buf ( n390498 , n43022 );
buf ( n390499 , n390498 );
buf ( n390500 , n388569 );
nand ( n43026 , n390499 , n390500 );
buf ( n390502 , n43026 );
buf ( n390503 , n390502 );
nand ( n43029 , n43020 , n390503 );
buf ( n390505 , n43029 );
buf ( n390506 , n390505 );
not ( n43032 , n390506 );
or ( n43033 , n43012 , n43032 );
buf ( n390509 , n389875 );
buf ( n390510 , n384554 );
nand ( n43036 , n390509 , n390510 );
buf ( n390512 , n43036 );
buf ( n390513 , n390512 );
nand ( n43039 , n43033 , n390513 );
buf ( n390515 , n43039 );
or ( n43041 , n390482 , n390515 );
buf ( n390517 , n388905 );
not ( n43043 , n390517 );
not ( n43044 , n27195 );
buf ( n390520 , n43044 );
not ( n43046 , n390520 );
or ( n43047 , n43043 , n43046 );
buf ( n390523 , n41118 );
not ( n43049 , n390523 );
buf ( n390525 , n388908 );
nand ( n43051 , n43049 , n390525 );
buf ( n390527 , n43051 );
buf ( n390528 , n390527 );
nand ( n43054 , n43047 , n390528 );
buf ( n390530 , n43054 );
buf ( n390531 , n390530 );
not ( n43057 , n390531 );
buf ( n43058 , n37337 );
buf ( n390534 , n43058 );
not ( n43060 , n390534 );
buf ( n390536 , n43060 );
buf ( n390537 , n390536 );
not ( n43063 , n390537 );
or ( n43064 , n43057 , n43063 );
buf ( n390540 , n388905 );
not ( n43066 , n390540 );
buf ( n390542 , n40779 );
not ( n43068 , n390542 );
or ( n43069 , n43066 , n43068 );
buf ( n390545 , n40760 );
buf ( n390546 , n388897 );
buf ( n43072 , n390546 );
buf ( n390548 , n43072 );
buf ( n390549 , n390548 );
nand ( n43075 , n390545 , n390549 );
buf ( n390551 , n43075 );
buf ( n390552 , n390551 );
nand ( n43078 , n43069 , n390552 );
buf ( n390554 , n43078 );
buf ( n390555 , n390554 );
buf ( n390556 , n37314 );
nand ( n43082 , n390555 , n390556 );
buf ( n390558 , n43082 );
buf ( n390559 , n390558 );
nand ( n43085 , n43064 , n390559 );
buf ( n390561 , n43085 );
buf ( n390562 , n390561 );
buf ( n390563 , n37316 );
not ( n43089 , n390563 );
buf ( n390565 , n388912 );
not ( n43091 , n390565 );
buf ( n390567 , n43091 );
buf ( n390568 , n390567 );
not ( n43094 , n390568 );
or ( n43095 , n43089 , n43094 );
buf ( n390571 , n384901 );
not ( n43097 , n390571 );
buf ( n390573 , n390554 );
nand ( n43099 , n43097 , n390573 );
buf ( n390575 , n43099 );
buf ( n390576 , n390575 );
nand ( n43102 , n43095 , n390576 );
buf ( n390578 , n43102 );
buf ( n390579 , n390578 );
xor ( n43105 , n390562 , n390579 );
buf ( n390581 , n40819 );
not ( n43107 , n390581 );
buf ( n390583 , n36251 );
not ( n43109 , n390583 );
or ( n43110 , n43107 , n43109 );
buf ( n390586 , n388263 );
buf ( n390587 , n388445 );
nand ( n43113 , n390586 , n390587 );
buf ( n390589 , n43113 );
buf ( n390590 , n390589 );
nand ( n43116 , n43110 , n390590 );
buf ( n390592 , n43116 );
buf ( n390593 , n390592 );
not ( n43119 , n390593 );
buf ( n390595 , n383894 );
not ( n43121 , n390595 );
or ( n43122 , n43119 , n43121 );
buf ( n390598 , n388617 );
buf ( n390599 , n383907 );
nand ( n43125 , n390598 , n390599 );
buf ( n390601 , n43125 );
buf ( n390602 , n390601 );
nand ( n43128 , n43122 , n390602 );
buf ( n390604 , n43128 );
buf ( n390605 , n390604 );
and ( n43131 , n43105 , n390605 );
and ( n43132 , n390562 , n390579 );
or ( n43133 , n43131 , n43132 );
buf ( n390609 , n43133 );
nand ( n43135 , n43041 , n390609 );
nand ( n43136 , n390515 , n390482 );
nand ( n43137 , n43135 , n43136 );
xor ( n43138 , n390448 , n43137 );
not ( n43139 , n43138 );
not ( n43140 , n42073 );
not ( n43141 , n40714 );
or ( n43142 , n43140 , n43141 );
buf ( n390618 , n35435 );
not ( n43144 , n42066 );
buf ( n390620 , n43144 );
nand ( n43146 , n390618 , n390620 );
buf ( n390622 , n43146 );
nand ( n43148 , n43142 , n390622 );
buf ( n390624 , n43148 );
not ( n43150 , n390624 );
buf ( n390626 , n383010 );
buf ( n390627 , n35405 );
and ( n43153 , n390626 , n390627 );
buf ( n390629 , n43153 );
buf ( n390630 , n390629 );
not ( n43156 , n390630 );
or ( n43157 , n43150 , n43156 );
buf ( n390633 , n383134 );
not ( n43159 , n390633 );
buf ( n390635 , n43159 );
buf ( n390636 , n390635 );
buf ( n390637 , n390466 );
nand ( n43163 , n390636 , n390637 );
buf ( n390639 , n43163 );
buf ( n390640 , n390639 );
nand ( n43166 , n43157 , n390640 );
buf ( n390642 , n43166 );
buf ( n390643 , n390642 );
not ( n43169 , n41565 );
not ( n43170 , n389299 );
or ( n43171 , n43169 , n43170 );
buf ( n390647 , n24050 );
not ( n43173 , n390647 );
buf ( n390649 , n36509 );
not ( n43175 , n390649 );
buf ( n390651 , n43175 );
buf ( n390652 , n390651 );
not ( n43178 , n390652 );
or ( n43179 , n43173 , n43178 );
buf ( n390655 , n384089 );
not ( n43181 , n390655 );
buf ( n390657 , n43181 );
buf ( n390658 , n390657 );
buf ( n390659 , n389075 );
nand ( n43185 , n390658 , n390659 );
buf ( n390661 , n43185 );
buf ( n390662 , n390661 );
nand ( n43188 , n43179 , n390662 );
buf ( n390664 , n43188 );
nand ( n43190 , n390664 , n389125 );
nand ( n43191 , n43171 , n43190 );
buf ( n390667 , n43191 );
xor ( n43193 , n390643 , n390667 );
not ( n43194 , n383891 );
not ( n43195 , n389936 );
buf ( n390671 , n41194 );
not ( n43197 , n390671 );
buf ( n390673 , n43197 );
not ( n43199 , n390673 );
or ( n43200 , n43195 , n43199 );
nand ( n43201 , n40775 , n41195 );
nand ( n43202 , n43200 , n43201 );
not ( n43203 , n43202 );
or ( n43204 , n43194 , n43203 );
buf ( n390680 , n390592 );
buf ( n390681 , n383907 );
nand ( n43207 , n390680 , n390681 );
buf ( n390683 , n43207 );
nand ( n43209 , n43204 , n390683 );
not ( n43210 , n41447 );
buf ( n390686 , n388962 );
not ( n43212 , n390686 );
buf ( n390688 , n388931 );
not ( n43214 , n390688 );
or ( n43215 , n43212 , n43214 );
buf ( n390691 , n28160 );
buf ( n390692 , n385488 );
nand ( n43218 , n390691 , n390692 );
buf ( n390694 , n43218 );
buf ( n390695 , n390694 );
nand ( n43221 , n43215 , n390695 );
buf ( n390697 , n43221 );
not ( n43223 , n390697 );
or ( n43224 , n43210 , n43223 );
buf ( n390700 , n388962 );
not ( n43226 , n390700 );
buf ( n390702 , n375781 );
not ( n43228 , n390702 );
buf ( n390704 , n43228 );
buf ( n390705 , n390704 );
not ( n43231 , n390705 );
or ( n43232 , n43226 , n43231 );
buf ( n390708 , n386147 );
buf ( n390709 , n388965 );
nand ( n43235 , n390708 , n390709 );
buf ( n390711 , n43235 );
buf ( n390712 , n390711 );
nand ( n43238 , n43232 , n390712 );
buf ( n390714 , n43238 );
not ( n43240 , n37932 );
nand ( n43241 , n390714 , n43240 );
nand ( n43242 , n43224 , n43241 );
xor ( n43243 , n43209 , n43242 );
buf ( n390719 , n388646 );
not ( n43245 , n390719 );
buf ( n390721 , n36395 );
not ( n43247 , n390721 );
or ( n43248 , n43245 , n43247 );
buf ( n390724 , n40839 );
buf ( n390725 , n388654 );
nand ( n43251 , n390724 , n390725 );
buf ( n390727 , n43251 );
buf ( n390728 , n390727 );
nand ( n43254 , n43248 , n390728 );
buf ( n390730 , n43254 );
not ( n43256 , n390730 );
not ( n43257 , n388460 );
or ( n43258 , n43256 , n43257 );
buf ( n390734 , n388370 );
not ( n43260 , n390734 );
buf ( n390736 , n40973 );
not ( n43262 , n390736 );
or ( n43263 , n43260 , n43262 );
buf ( n390739 , n40977 );
buf ( n390740 , n388373 );
nand ( n43266 , n390739 , n390740 );
buf ( n390742 , n43266 );
buf ( n390743 , n390742 );
nand ( n43269 , n43263 , n390743 );
buf ( n390745 , n43269 );
buf ( n390746 , n390745 );
buf ( n43272 , n36363 );
buf ( n390748 , n43272 );
nand ( n43274 , n390746 , n390748 );
buf ( n390750 , n43274 );
nand ( n43276 , n43258 , n390750 );
and ( n43277 , n43243 , n43276 );
and ( n43278 , n43209 , n43242 );
or ( n43279 , n43277 , n43278 );
buf ( n390755 , n43279 );
and ( n43281 , n43193 , n390755 );
and ( n43282 , n390643 , n390667 );
or ( n43283 , n43281 , n43282 );
buf ( n390759 , n43283 );
not ( n43285 , n390759 );
not ( n43286 , n388093 );
buf ( n390762 , n43286 );
not ( n43288 , n390762 );
buf ( n390764 , n388102 );
not ( n43290 , n390764 );
buf ( n390766 , n388771 );
not ( n43292 , n390766 );
or ( n43293 , n43290 , n43292 );
buf ( n390769 , n383056 );
buf ( n390770 , n388105 );
nand ( n43296 , n390769 , n390770 );
buf ( n390772 , n43296 );
buf ( n390773 , n390772 );
nand ( n43299 , n43293 , n390773 );
buf ( n390775 , n43299 );
buf ( n390776 , n390775 );
not ( n43302 , n390776 );
or ( n43303 , n43288 , n43302 );
buf ( n390779 , n390335 );
not ( n43305 , n390779 );
buf ( n390781 , n390362 );
nand ( n43307 , n43305 , n390781 );
buf ( n390783 , n43307 );
buf ( n390784 , n390783 );
nand ( n43310 , n43303 , n390784 );
buf ( n390786 , n43310 );
not ( n43312 , n390786 );
nand ( n43313 , n43285 , n43312 );
not ( n43314 , n43313 );
buf ( n390790 , n24074 );
not ( n43316 , n390790 );
buf ( n390792 , n384180 );
not ( n43318 , n390792 );
buf ( n390794 , n43318 );
buf ( n390795 , n390794 );
not ( n43321 , n390795 );
or ( n43322 , n43316 , n43321 );
buf ( n390798 , n384180 );
buf ( n390799 , n24073 );
nand ( n43325 , n390798 , n390799 );
buf ( n390801 , n43325 );
buf ( n390802 , n390801 );
nand ( n43328 , n43322 , n390802 );
buf ( n390804 , n43328 );
and ( n43330 , n390804 , n390403 );
buf ( n390806 , n24074 );
not ( n43332 , n390806 );
buf ( n390808 , n389692 );
not ( n43334 , n390808 );
buf ( n390810 , n43334 );
buf ( n390811 , n390810 );
not ( n43337 , n390811 );
or ( n43338 , n43332 , n43337 );
buf ( n390814 , n389692 );
buf ( n390815 , n24073 );
nand ( n43341 , n390814 , n390815 );
buf ( n390817 , n43341 );
buf ( n390818 , n390817 );
nand ( n43344 , n43338 , n390818 );
buf ( n390820 , n43344 );
not ( n43346 , n390820 );
nor ( n43347 , n43346 , n390435 );
nor ( n43348 , n43330 , n43347 );
buf ( n390824 , n43348 );
not ( n43350 , n390824 );
buf ( n390826 , n43350 );
not ( n43352 , n390826 );
buf ( n390828 , n390745 );
not ( n43354 , n390828 );
buf ( n390830 , n36434 );
not ( n43356 , n390830 );
buf ( n390832 , n43356 );
buf ( n390833 , n390832 );
not ( n43359 , n390833 );
or ( n43360 , n43354 , n43359 );
buf ( n390836 , n388696 );
buf ( n390837 , n388346 );
nand ( n43363 , n390836 , n390837 );
buf ( n390839 , n43363 );
buf ( n390840 , n390839 );
nand ( n43366 , n43360 , n390840 );
buf ( n390842 , n43366 );
buf ( n390843 , n390842 );
or ( n43369 , n29077 , n385488 );
nand ( n43370 , n43369 , n41488 );
not ( n43371 , n43370 );
not ( n43372 , n41447 );
or ( n43373 , n43371 , n43372 );
buf ( n390849 , n390697 );
buf ( n390850 , n43240 );
nand ( n43376 , n390849 , n390850 );
buf ( n390852 , n43376 );
nand ( n43378 , n43373 , n390852 );
not ( n43379 , n43378 );
buf ( n390855 , n43379 );
and ( n43381 , n390843 , n390855 );
not ( n43382 , n390843 );
buf ( n390858 , n41447 );
not ( n43384 , n390858 );
buf ( n390860 , n388986 );
not ( n43386 , n390860 );
or ( n43387 , n43384 , n43386 );
buf ( n390863 , n390852 );
nand ( n43389 , n43387 , n390863 );
buf ( n390865 , n43389 );
buf ( n390866 , n390865 );
and ( n43392 , n43382 , n390866 );
or ( n43393 , n43381 , n43392 );
buf ( n390869 , n43393 );
buf ( n390870 , n390869 );
buf ( n390871 , n389862 );
not ( n43397 , n390871 );
buf ( n390873 , n40885 );
not ( n43399 , n390873 );
buf ( n390875 , n43399 );
buf ( n390876 , n390875 );
not ( n43402 , n390876 );
or ( n43403 , n43397 , n43402 );
buf ( n390879 , n40943 );
buf ( n390880 , n389859 );
nand ( n43406 , n390879 , n390880 );
buf ( n390882 , n43406 );
buf ( n390883 , n390882 );
nand ( n43409 , n43403 , n390883 );
buf ( n390885 , n43409 );
buf ( n390886 , n390885 );
not ( n43412 , n390886 );
buf ( n390888 , n36801 );
not ( n43414 , n390888 );
or ( n43415 , n43412 , n43414 );
buf ( n390891 , n388661 );
buf ( n390892 , n388669 );
nand ( n43418 , n390891 , n390892 );
buf ( n390894 , n43418 );
buf ( n390895 , n390894 );
nand ( n43421 , n43415 , n390895 );
buf ( n390897 , n43421 );
buf ( n390898 , n390897 );
not ( n43424 , n390898 );
buf ( n390900 , n43424 );
buf ( n390901 , n390900 );
and ( n43427 , n390870 , n390901 );
not ( n43428 , n390870 );
buf ( n390904 , n390897 );
and ( n43430 , n43428 , n390904 );
nor ( n43431 , n43427 , n43430 );
buf ( n390907 , n43431 );
buf ( n390908 , n390907 );
not ( n43434 , n390908 );
buf ( n390910 , n43434 );
not ( n43436 , n390910 );
or ( n43437 , n43352 , n43436 );
buf ( n390913 , n43348 );
not ( n43439 , n390913 );
buf ( n390915 , n390907 );
not ( n43441 , n390915 );
or ( n43442 , n43439 , n43441 );
buf ( n390918 , n390561 );
not ( n43444 , n390918 );
buf ( n390920 , n43444 );
buf ( n390921 , n390920 );
buf ( n390922 , n390490 );
not ( n43448 , n390922 );
buf ( n390924 , n40886 );
not ( n43450 , n390924 );
or ( n43451 , n43448 , n43450 );
buf ( n390927 , n390875 );
not ( n43453 , n390927 );
buf ( n390929 , n43453 );
buf ( n390930 , n390929 );
buf ( n390931 , n388569 );
nand ( n43457 , n390930 , n390931 );
buf ( n390933 , n43457 );
buf ( n390934 , n390933 );
nand ( n43460 , n43451 , n390934 );
buf ( n390936 , n43460 );
buf ( n390937 , n390936 );
not ( n43463 , n390937 );
buf ( n390939 , n36801 );
not ( n43465 , n390939 );
or ( n43466 , n43463 , n43465 );
buf ( n390942 , n384413 );
buf ( n390943 , n390885 );
nand ( n43469 , n390942 , n390943 );
buf ( n390945 , n43469 );
buf ( n390946 , n390945 );
nand ( n43472 , n43466 , n390946 );
buf ( n390948 , n43472 );
buf ( n390949 , n390948 );
xor ( n43475 , n390921 , n390949 );
and ( n43476 , n40990 , n385987 );
not ( n43477 , n40990 );
and ( n43478 , n43477 , n31964 );
or ( n43479 , n43476 , n43478 );
buf ( n390955 , n43479 );
not ( n43481 , n390955 );
buf ( n390957 , n389744 );
not ( n43483 , n390957 );
or ( n43484 , n43481 , n43483 );
buf ( n390960 , n389024 );
buf ( n390961 , n389319 );
nand ( n43487 , n390960 , n390961 );
buf ( n390963 , n43487 );
buf ( n390964 , n390963 );
nand ( n43490 , n43484 , n390964 );
buf ( n390966 , n43490 );
buf ( n390967 , n390966 );
and ( n43493 , n43475 , n390967 );
and ( n43494 , n390921 , n390949 );
or ( n43495 , n43493 , n43494 );
buf ( n390971 , n43495 );
buf ( n390972 , n390971 );
nand ( n43498 , n43442 , n390972 );
buf ( n390974 , n43498 );
nand ( n43500 , n43437 , n390974 );
not ( n43501 , n43500 );
or ( n43502 , n43314 , n43501 );
nand ( n43503 , n390786 , n390759 );
nand ( n43504 , n43502 , n43503 );
not ( n43505 , n43504 );
or ( n43506 , n43139 , n43505 );
or ( n43507 , n43504 , n43138 );
buf ( n390983 , n23701 );
not ( n43509 , n390983 );
buf ( n390985 , n43509 );
buf ( n390986 , n390985 );
not ( n43512 , n390986 );
buf ( n390988 , n43512 );
xnor ( n43514 , n390988 , n23723 );
not ( n43515 , n43514 );
not ( n43516 , n43515 );
buf ( n390992 , n43516 );
not ( n43518 , n390992 );
not ( n43519 , n23725 );
buf ( n390995 , n371876 );
not ( n43521 , n390995 );
buf ( n390997 , n43521 );
not ( n43523 , n390997 );
or ( n43524 , n43519 , n43523 );
not ( n43525 , n23724 );
not ( n43526 , n24258 );
not ( n43527 , n371869 );
or ( n43528 , n43526 , n43527 );
nand ( n43529 , n43528 , n24268 );
not ( n43530 , n43529 );
not ( n43531 , n43530 );
or ( n43532 , n43525 , n43531 );
nand ( n43533 , n43532 , n43514 );
not ( n43534 , n43533 );
nand ( n43535 , n43524 , n43534 );
not ( n43536 , n43535 );
not ( n43537 , n43536 );
buf ( n391013 , n43537 );
not ( n43539 , n391013 );
or ( n43540 , n43518 , n43539 );
buf ( n391016 , n390997 );
buf ( n43542 , n391016 );
buf ( n391018 , n43542 );
buf ( n391019 , n391018 );
not ( n43545 , n391019 );
buf ( n391021 , n43545 );
buf ( n391022 , n391021 );
buf ( n43548 , n391022 );
buf ( n391024 , n43548 );
buf ( n391025 , n391024 );
not ( n43551 , n391025 );
buf ( n391027 , n43551 );
buf ( n391028 , n391027 );
not ( n43554 , n391028 );
buf ( n391030 , n34859 );
buf ( n43556 , n391030 );
buf ( n391032 , n43556 );
buf ( n391033 , n391032 );
not ( n43559 , n391033 );
or ( n43560 , n43554 , n43559 );
buf ( n391036 , n385499 );
buf ( n391037 , n391024 );
nand ( n43563 , n391036 , n391037 );
buf ( n391039 , n43563 );
buf ( n391040 , n391039 );
nand ( n43566 , n43560 , n391040 );
buf ( n391042 , n43566 );
buf ( n391043 , n391042 );
nand ( n43569 , n43540 , n391043 );
buf ( n391045 , n43569 );
buf ( n391046 , n391045 );
xor ( n43572 , n389739 , n389773 );
xor ( n43573 , n43572 , n389783 );
buf ( n391049 , n43573 );
buf ( n391050 , n391049 );
xor ( n43576 , n391046 , n391050 );
xor ( n43577 , n389827 , n389852 );
xor ( n43578 , n43577 , n389915 );
buf ( n391054 , n43578 );
buf ( n391055 , n391054 );
xor ( n43581 , n43576 , n391055 );
buf ( n391057 , n43581 );
nand ( n43583 , n43507 , n391057 );
nand ( n43584 , n43506 , n43583 );
buf ( n391060 , n43584 );
not ( n43586 , n390440 );
buf ( n391062 , n390366 );
not ( n43588 , n391062 );
buf ( n391064 , n43588 );
not ( n43590 , n391064 );
or ( n43591 , n43586 , n43590 );
not ( n43592 , n390366 );
not ( n43593 , n42962 );
or ( n43594 , n43592 , n43593 );
nand ( n43595 , n43594 , n43137 );
nand ( n43596 , n43591 , n43595 );
xor ( n43597 , n391046 , n391050 );
and ( n43598 , n43597 , n391055 );
and ( n43599 , n391046 , n391050 );
or ( n43600 , n43598 , n43599 );
buf ( n391076 , n43600 );
xor ( n43602 , n43596 , n391076 );
buf ( n391078 , n390435 );
not ( n43604 , n391078 );
buf ( n391080 , n43604 );
buf ( n391081 , n391080 );
not ( n43607 , n391081 );
buf ( n391083 , n390386 );
not ( n43609 , n391083 );
or ( n43610 , n43607 , n43609 );
buf ( n391086 , n389525 );
not ( n43612 , n391086 );
buf ( n391088 , n24074 );
not ( n43614 , n391088 );
or ( n43615 , n43612 , n43614 );
buf ( n391091 , n37173 );
buf ( n391092 , n24073 );
nand ( n43618 , n391091 , n391092 );
buf ( n391094 , n43618 );
buf ( n391095 , n391094 );
nand ( n43621 , n43615 , n391095 );
buf ( n391097 , n43621 );
buf ( n391098 , n391097 );
buf ( n391099 , n390403 );
nand ( n43625 , n391098 , n391099 );
buf ( n391101 , n43625 );
buf ( n391102 , n391101 );
nand ( n43628 , n43610 , n391102 );
buf ( n391104 , n43628 );
buf ( n391105 , n391104 );
buf ( n391106 , n43286 );
not ( n43632 , n391106 );
buf ( n391108 , n390358 );
not ( n43634 , n391108 );
or ( n43635 , n43632 , n43634 );
buf ( n391111 , n388120 );
buf ( n391112 , n390362 );
nand ( n43638 , n391111 , n391112 );
buf ( n391114 , n43638 );
buf ( n391115 , n391114 );
nand ( n43641 , n43635 , n391115 );
buf ( n391117 , n43641 );
buf ( n391118 , n391117 );
xor ( n43644 , n391105 , n391118 );
buf ( n391120 , n389904 );
not ( n43646 , n391120 );
buf ( n391122 , n384624 );
not ( n43648 , n391122 );
or ( n43649 , n43646 , n43648 );
buf ( n391125 , n388376 );
not ( n43651 , n391125 );
buf ( n391127 , n37037 );
not ( n43653 , n391127 );
buf ( n391129 , n43653 );
buf ( n391130 , n391129 );
not ( n43656 , n391130 );
or ( n43657 , n43651 , n43656 );
buf ( n391133 , n37037 );
buf ( n391134 , n388373 );
nand ( n43660 , n391133 , n391134 );
buf ( n391136 , n43660 );
buf ( n391137 , n391136 );
nand ( n43663 , n43657 , n391137 );
buf ( n391139 , n43663 );
buf ( n391140 , n391139 );
buf ( n391141 , n389908 );
nand ( n43667 , n391140 , n391141 );
buf ( n391143 , n43667 );
buf ( n391144 , n391143 );
nand ( n43670 , n43649 , n391144 );
buf ( n391146 , n43670 );
buf ( n391147 , n391146 );
buf ( n391148 , n41447 );
not ( n43674 , n391148 );
buf ( n391150 , n390200 );
not ( n43676 , n391150 );
or ( n43677 , n43674 , n43676 );
buf ( n391153 , n389841 );
buf ( n391154 , n385479 );
nand ( n43680 , n391153 , n391154 );
buf ( n391156 , n43680 );
buf ( n391157 , n391156 );
nand ( n43683 , n43677 , n391157 );
buf ( n391159 , n43683 );
buf ( n391160 , n391159 );
xor ( n43686 , n391147 , n391160 );
buf ( n391162 , n388539 );
buf ( n43688 , n391162 );
buf ( n391164 , n43688 );
buf ( n391165 , n391164 );
buf ( n391166 , n388580 );
or ( n43692 , n391165 , n391166 );
buf ( n391168 , n35825 );
not ( n43694 , n391168 );
buf ( n391170 , n43694 );
buf ( n391171 , n391170 );
buf ( n43697 , n391171 );
buf ( n391173 , n43697 );
buf ( n391174 , n391173 );
not ( n43700 , n391174 );
buf ( n391176 , n43700 );
buf ( n391177 , n391176 );
buf ( n391178 , n388556 );
buf ( n391179 , n389859 );
and ( n43705 , n391178 , n391179 );
buf ( n391181 , n389589 );
not ( n43707 , n391181 );
buf ( n391183 , n43707 );
buf ( n391184 , n391183 );
buf ( n391185 , n389862 );
and ( n43711 , n391184 , n391185 );
nor ( n43712 , n43705 , n43711 );
buf ( n391188 , n43712 );
buf ( n391189 , n391188 );
or ( n43715 , n391177 , n391189 );
nand ( n43716 , n43692 , n43715 );
buf ( n391192 , n43716 );
buf ( n391193 , n391192 );
xor ( n43719 , n43686 , n391193 );
buf ( n391195 , n43719 );
buf ( n391196 , n391195 );
xor ( n43722 , n43644 , n391196 );
buf ( n391198 , n43722 );
xor ( n43724 , n43602 , n391198 );
buf ( n391200 , n43724 );
xor ( n43726 , n391060 , n391200 );
not ( n43727 , n43537 );
buf ( n391203 , n43727 );
not ( n43729 , n391203 );
buf ( n391205 , n391027 );
not ( n43731 , n391205 );
buf ( n391207 , n382548 );
not ( n43733 , n391207 );
or ( n43734 , n43731 , n43733 );
buf ( n391210 , n382548 );
not ( n43736 , n391210 );
buf ( n391212 , n43736 );
buf ( n391213 , n391212 );
buf ( n391214 , n391024 );
nand ( n43740 , n391213 , n391214 );
buf ( n391216 , n43740 );
buf ( n391217 , n391216 );
nand ( n43743 , n43734 , n391217 );
buf ( n391219 , n43743 );
buf ( n391220 , n391219 );
not ( n43746 , n391220 );
or ( n43747 , n43729 , n43746 );
buf ( n391223 , n391042 );
buf ( n391224 , n43515 );
nand ( n43750 , n391223 , n391224 );
buf ( n391226 , n43750 );
buf ( n391227 , n391226 );
nand ( n43753 , n43747 , n391227 );
buf ( n391229 , n43753 );
buf ( n391230 , n388549 );
not ( n43756 , n391230 );
buf ( n391232 , n42390 );
not ( n43758 , n391232 );
or ( n43759 , n43756 , n43758 );
buf ( n391235 , n389897 );
buf ( n391236 , n388546 );
nand ( n43762 , n391235 , n391236 );
buf ( n391238 , n43762 );
buf ( n391239 , n391238 );
nand ( n43765 , n43759 , n391239 );
buf ( n391241 , n43765 );
buf ( n391242 , n391241 );
not ( n43768 , n391242 );
buf ( n391244 , n384624 );
not ( n43770 , n391244 );
or ( n43771 , n43768 , n43770 );
buf ( n391247 , n389908 );
buf ( n391248 , n390505 );
nand ( n43774 , n391247 , n391248 );
buf ( n391250 , n43774 );
buf ( n391251 , n391250 );
nand ( n43777 , n43771 , n391251 );
buf ( n391253 , n43777 );
buf ( n391254 , n391253 );
buf ( n391255 , n388242 );
buf ( n391256 , n383423 );
and ( n43782 , n391255 , n391256 );
not ( n43783 , n391255 );
buf ( n391259 , n388576 );
and ( n43785 , n43783 , n391259 );
nor ( n43786 , n43782 , n43785 );
buf ( n391262 , n43786 );
buf ( n391263 , n391262 );
not ( n43789 , n391263 );
buf ( n391265 , n43789 );
buf ( n391266 , n391265 );
not ( n43792 , n391266 );
buf ( n391268 , n388539 );
not ( n43794 , n391268 );
buf ( n391270 , n43794 );
buf ( n391271 , n391270 );
not ( n43797 , n391271 );
or ( n43798 , n43792 , n43797 );
buf ( n391274 , n389606 );
not ( n43800 , n391274 );
buf ( n391276 , n383406 );
nand ( n43802 , n43800 , n391276 );
buf ( n391278 , n43802 );
buf ( n391279 , n391278 );
nand ( n43805 , n43798 , n391279 );
buf ( n391281 , n43805 );
buf ( n391282 , n391281 );
xor ( n43808 , n391254 , n391282 );
xor ( n43809 , n390562 , n390579 );
xor ( n391285 , n43809 , n390605 );
buf ( n391286 , n391285 );
buf ( n391287 , n391286 );
and ( n43813 , n43808 , n391287 );
and ( n43814 , n391254 , n391282 );
or ( n43815 , n43813 , n43814 );
buf ( n391291 , n43815 );
xor ( n43817 , n391229 , n391291 );
buf ( n391293 , n41711 );
not ( n43819 , n391293 );
buf ( n391295 , n41671 );
not ( n43821 , n391295 );
buf ( n391297 , n37369 );
not ( n43823 , n391297 );
or ( n43824 , n43821 , n43823 );
buf ( n391300 , n36066 );
buf ( n391301 , n41678 );
nand ( n43827 , n391300 , n391301 );
buf ( n391303 , n43827 );
buf ( n391304 , n391303 );
nand ( n43830 , n43824 , n391304 );
buf ( n391306 , n43830 );
buf ( n391307 , n391306 );
not ( n43833 , n391307 );
or ( n43834 , n43819 , n43833 );
buf ( n391310 , n389266 );
buf ( n391311 , n389162 );
nand ( n43837 , n391310 , n391311 );
buf ( n391313 , n43837 );
buf ( n391314 , n391313 );
nand ( n43840 , n43834 , n391314 );
buf ( n391316 , n43840 );
and ( n43842 , n43817 , n391316 );
and ( n43843 , n391229 , n391291 );
or ( n43844 , n43842 , n43843 );
buf ( n391320 , n43844 );
xor ( n43846 , n388584 , n41107 );
xnor ( n43847 , n43846 , n388714 );
buf ( n391323 , n43847 );
buf ( n43849 , n391323 );
buf ( n391325 , n43849 );
buf ( n391326 , n391325 );
not ( n43852 , n391326 );
not ( n43853 , n388833 );
not ( n43854 , n41363 );
or ( n43855 , n43853 , n43854 );
nand ( n43856 , n41935 , n41373 );
nand ( n43857 , n43855 , n43856 );
not ( n43858 , n43857 );
buf ( n391334 , n390403 );
not ( n43860 , n391334 );
buf ( n391336 , n390416 );
not ( n43862 , n391336 );
or ( n43863 , n43860 , n43862 );
buf ( n391339 , n390804 );
buf ( n391340 , n391080 );
nand ( n43866 , n391339 , n391340 );
buf ( n391342 , n43866 );
buf ( n391343 , n391342 );
nand ( n43869 , n43863 , n391343 );
buf ( n391345 , n43869 );
buf ( n391346 , n391345 );
not ( n43872 , n391346 );
buf ( n391348 , n43872 );
buf ( n391349 , n391348 );
buf ( n391350 , n390897 );
not ( n43876 , n391350 );
buf ( n391352 , n390842 );
not ( n43878 , n391352 );
buf ( n391354 , n43379 );
nand ( n43880 , n43878 , n391354 );
buf ( n391356 , n43880 );
buf ( n391357 , n391356 );
not ( n43883 , n391357 );
or ( n43884 , n43876 , n43883 );
buf ( n391360 , n390865 );
buf ( n391361 , n390842 );
nand ( n43887 , n391360 , n391361 );
buf ( n391363 , n43887 );
buf ( n391364 , n391363 );
nand ( n43890 , n43884 , n391364 );
buf ( n391366 , n43890 );
buf ( n391367 , n391366 );
not ( n43893 , n391367 );
buf ( n391369 , n43893 );
buf ( n391370 , n391369 );
nand ( n43896 , n391349 , n391370 );
buf ( n391372 , n43896 );
buf ( n391373 , n391372 );
xor ( n43899 , n388636 , n388677 );
xor ( n43900 , n43899 , n388710 );
buf ( n391376 , n43900 );
buf ( n391377 , n391376 );
and ( n43903 , n391373 , n391377 );
and ( n43904 , n391345 , n391366 );
buf ( n391380 , n43904 );
nor ( n43906 , n43903 , n391380 );
buf ( n391382 , n43906 );
not ( n43908 , n391382 );
or ( n43909 , n43858 , n43908 );
or ( n43910 , n391382 , n43857 );
nand ( n43911 , n43909 , n43910 );
buf ( n391387 , n43911 );
not ( n43913 , n391387 );
or ( n43914 , n43852 , n43913 );
buf ( n391390 , n43911 );
buf ( n391391 , n391325 );
or ( n43917 , n391390 , n391391 );
nand ( n43918 , n43914 , n43917 );
buf ( n391394 , n43918 );
buf ( n391395 , n391394 );
xor ( n43921 , n391320 , n391395 );
buf ( n391397 , n390609 );
not ( n43923 , n391397 );
buf ( n391399 , n43923 );
and ( n43925 , n390515 , n391399 );
not ( n43926 , n390515 );
and ( n43927 , n43926 , n390609 );
or ( n43928 , n43925 , n43927 );
buf ( n391404 , n43928 );
buf ( n391405 , n390482 );
and ( n43931 , n391404 , n391405 );
not ( n43932 , n391404 );
buf ( n391408 , n390482 );
not ( n43934 , n391408 );
buf ( n391410 , n43934 );
buf ( n391411 , n391410 );
and ( n43937 , n43932 , n391411 );
nor ( n43938 , n43931 , n43937 );
buf ( n391414 , n43938 );
buf ( n391415 , n391414 );
buf ( n391416 , n388809 );
not ( n43942 , n391416 );
buf ( n391418 , n389233 );
not ( n43944 , n391418 );
or ( n43945 , n43942 , n43944 );
buf ( n391421 , n388760 );
buf ( n391422 , n35301 );
and ( n43948 , n391421 , n391422 );
not ( n43949 , n391421 );
buf ( n391425 , n42616 );
and ( n43951 , n43949 , n391425 );
nor ( n43952 , n43948 , n43951 );
buf ( n391428 , n43952 );
buf ( n391429 , n391428 );
buf ( n391430 , n388746 );
nand ( n43956 , n391429 , n391430 );
buf ( n391432 , n43956 );
buf ( n391433 , n391432 );
nand ( n43959 , n43945 , n391433 );
buf ( n391435 , n43959 );
buf ( n391436 , n391435 );
xor ( n43962 , n391415 , n391436 );
buf ( n391438 , n24887 );
not ( n43964 , n391438 );
buf ( n391440 , n43964 );
buf ( n391441 , n391440 );
buf ( n43967 , n391441 );
buf ( n391443 , n43967 );
buf ( n391444 , n391443 );
not ( n43970 , n391444 );
buf ( n391446 , n43970 );
buf ( n391447 , n391446 );
not ( n43973 , n391447 );
buf ( n391449 , n384143 );
not ( n43975 , n391449 );
or ( n43976 , n43973 , n43975 );
buf ( n391452 , n382854 );
buf ( n391453 , n391446 );
not ( n43979 , n391453 );
buf ( n391455 , n43979 );
buf ( n391456 , n391455 );
nand ( n43982 , n391452 , n391456 );
buf ( n391458 , n43982 );
buf ( n391459 , n391458 );
nand ( n43985 , n43976 , n391459 );
buf ( n391461 , n43985 );
buf ( n391462 , n389547 );
buf ( n391463 , n41850 );
nand ( n43994 , n391462 , n391463 );
buf ( n391465 , n43994 );
buf ( n391466 , n391465 );
nand ( n43997 , C1 , n391466 );
buf ( n391468 , n43997 );
buf ( n391469 , n391468 );
buf ( n391470 , n386480 );
not ( n44001 , n391470 );
buf ( n391472 , n389401 );
not ( n44003 , n391472 );
or ( n44004 , n44001 , n44003 );
buf ( n391475 , n22982 );
not ( n44006 , n391475 );
not ( n44007 , n29077 );
buf ( n391478 , n44007 );
not ( n44009 , n391478 );
or ( n44010 , n44006 , n44009 );
buf ( n391481 , n29077 );
not ( n44012 , n391481 );
buf ( n391483 , n44012 );
buf ( n391484 , n391483 );
not ( n44015 , n391484 );
buf ( n391486 , n44015 );
buf ( n391487 , n391486 );
buf ( n391488 , n38971 );
nand ( n44019 , n391487 , n391488 );
buf ( n391490 , n44019 );
buf ( n391491 , n391490 );
nand ( n44022 , n44010 , n391491 );
buf ( n391493 , n44022 );
buf ( n391494 , n391493 );
buf ( n391495 , n386496 );
nand ( n44026 , n391494 , n391495 );
buf ( n391497 , n44026 );
buf ( n391498 , n391497 );
nand ( n44029 , n44004 , n391498 );
buf ( n391500 , n44029 );
buf ( n391501 , n391500 );
or ( n44032 , n391469 , n391501 );
buf ( n391503 , n389125 );
not ( n44034 , n391503 );
buf ( n391505 , n24050 );
not ( n44036 , n391505 );
buf ( n391507 , n36565 );
not ( n44038 , n391507 );
or ( n44039 , n44036 , n44038 );
buf ( n391510 , n38155 );
buf ( n391511 , n389075 );
nand ( n44042 , n391510 , n391511 );
buf ( n391513 , n44042 );
buf ( n391514 , n391513 );
nand ( n44045 , n44039 , n391514 );
buf ( n391516 , n44045 );
buf ( n391517 , n391516 );
not ( n44048 , n391517 );
or ( n44049 , n44034 , n44048 );
buf ( n391520 , n390664 );
buf ( n391521 , n41565 );
nand ( n44052 , n391520 , n391521 );
buf ( n391523 , n44052 );
buf ( n391524 , n391523 );
nand ( n44055 , n44049 , n391524 );
buf ( n391526 , n44055 );
buf ( n391527 , n391526 );
nand ( n44058 , n44032 , n391527 );
buf ( n391529 , n44058 );
buf ( n391530 , n391529 );
buf ( n391531 , n391500 );
buf ( n391532 , n391468 );
nand ( n44063 , n391531 , n391532 );
buf ( n391534 , n44063 );
buf ( n391535 , n391534 );
nand ( n44066 , n391530 , n391535 );
buf ( n391537 , n44066 );
buf ( n391538 , n391537 );
xor ( n44069 , n389335 , n389377 );
xor ( n44070 , n44069 , n389409 );
buf ( n391541 , n44070 );
buf ( n391542 , n391541 );
xor ( n44073 , n391538 , n391542 );
not ( n44074 , n41447 );
not ( n44075 , n390714 );
or ( n44076 , n44074 , n44075 );
nand ( n44077 , n37922 , n37930 , n37931 );
buf ( n391548 , n44077 );
buf ( n44079 , n391548 );
buf ( n391550 , n44079 );
buf ( n391551 , n391550 );
not ( n44082 , n391551 );
buf ( n391553 , n44082 );
and ( n44084 , n385488 , n40758 );
not ( n44085 , n385488 );
and ( n44086 , n44085 , n27612 );
or ( n44087 , n44084 , n44086 );
nand ( n44088 , n391553 , n44087 );
nand ( n44089 , n44076 , n44088 );
buf ( n391560 , n44089 );
buf ( n391561 , n41407 );
not ( n44092 , n391561 );
buf ( n391563 , n44092 );
not ( n44094 , n391563 );
not ( n44095 , n40818 );
or ( n44096 , n44094 , n44095 );
buf ( n391567 , n28215 );
buf ( n44098 , n391567 );
buf ( n391569 , n44098 );
nand ( n44100 , n388905 , n391569 );
nand ( n44101 , n44096 , n44100 );
not ( n44102 , n44101 );
not ( n44103 , n37338 );
or ( n44104 , n44102 , n44103 );
buf ( n391575 , n390530 );
buf ( n391576 , n37314 );
nand ( n44107 , n391575 , n391576 );
buf ( n391578 , n44107 );
nand ( n44109 , n44104 , n391578 );
buf ( n391580 , n44109 );
xor ( n44111 , n391560 , n391580 );
buf ( n391582 , n389936 );
not ( n44113 , n391582 );
buf ( n391584 , n388370 );
not ( n44115 , n391584 );
or ( n44116 , n44113 , n44115 );
buf ( n391587 , n40775 );
buf ( n391588 , n388367 );
nand ( n44119 , n391587 , n391588 );
buf ( n391590 , n44119 );
buf ( n391591 , n391590 );
nand ( n44122 , n44116 , n391591 );
buf ( n391593 , n44122 );
buf ( n391594 , n391593 );
not ( n44125 , n391594 );
buf ( n391596 , n383891 );
not ( n44127 , n391596 );
or ( n44128 , n44125 , n44127 );
buf ( n391599 , n43202 );
buf ( n391600 , n383904 );
buf ( n44131 , n391600 );
buf ( n391602 , n44131 );
buf ( n391603 , n391602 );
nand ( n44134 , n391599 , n391603 );
buf ( n391605 , n44134 );
buf ( n391606 , n391605 );
nand ( n44137 , n44128 , n391606 );
buf ( n391608 , n44137 );
buf ( n391609 , n391608 );
and ( n44140 , n44111 , n391609 );
and ( n44141 , n391560 , n391580 );
or ( n44142 , n44140 , n44141 );
buf ( n391613 , n44142 );
buf ( n391614 , n391613 );
buf ( n391615 , n389602 );
not ( n44146 , n391615 );
buf ( n391617 , n391129 );
not ( n44148 , n391617 );
or ( n44149 , n44146 , n44148 );
buf ( n391620 , n389894 );
buf ( n391621 , n389593 );
nand ( n44152 , n391620 , n391621 );
buf ( n391623 , n44152 );
buf ( n391624 , n391623 );
nand ( n44155 , n44149 , n391624 );
buf ( n391626 , n44155 );
buf ( n391627 , n391626 );
not ( n44158 , n391627 );
buf ( n391629 , n389883 );
not ( n44160 , n391629 );
or ( n44161 , n44158 , n44160 );
buf ( n391632 , n391241 );
buf ( n391633 , n384548 );
not ( n44164 , n391633 );
buf ( n391635 , n44164 );
buf ( n391636 , n391635 );
not ( n44167 , n391636 );
buf ( n391638 , n44167 );
buf ( n391639 , n391638 );
nand ( n44170 , n391632 , n391639 );
buf ( n391641 , n44170 );
buf ( n391642 , n391641 );
nand ( n44173 , n44161 , n391642 );
buf ( n391644 , n44173 );
buf ( n391645 , n391644 );
xor ( n44176 , n391614 , n391645 );
buf ( n391647 , n383467 );
not ( n44178 , n391647 );
buf ( n391649 , n44178 );
buf ( n391650 , n391649 );
buf ( n44181 , n391650 );
buf ( n391652 , n44181 );
buf ( n391653 , n391652 );
not ( n44184 , n391653 );
buf ( n391655 , n44184 );
buf ( n391656 , n391655 );
buf ( n391657 , n388998 );
buf ( n391658 , n385633 );
and ( n44189 , n391657 , n391658 );
not ( n44190 , n391657 );
buf ( n391661 , n388556 );
and ( n44192 , n44190 , n391661 );
nor ( n44193 , n44189 , n44192 );
buf ( n391664 , n44193 );
buf ( n391665 , n391664 );
or ( n44196 , n391656 , n391665 );
buf ( n391667 , n391176 );
buf ( n391668 , n391262 );
or ( n44199 , n391667 , n391668 );
nand ( n44200 , n44196 , n44199 );
buf ( n391671 , n44200 );
buf ( n391672 , n391671 );
and ( n44203 , n44176 , n391672 );
and ( n44204 , n391614 , n391645 );
or ( n44205 , n44203 , n44204 );
buf ( n391676 , n44205 );
buf ( n391677 , n391676 );
and ( n44208 , n44073 , n391677 );
and ( n44209 , n391538 , n391542 );
or ( n44210 , n44208 , n44209 );
buf ( n391681 , n44210 );
buf ( n391682 , n391681 );
and ( n44213 , n43962 , n391682 );
and ( n44214 , n391415 , n391436 );
or ( n44215 , n44213 , n44214 );
buf ( n391686 , n44215 );
buf ( n391687 , n391686 );
and ( n44218 , n43921 , n391687 );
and ( n44219 , n391320 , n391395 );
or ( n44220 , n44218 , n44219 );
buf ( n391691 , n44220 );
buf ( n391692 , n391691 );
and ( n44223 , n43726 , n391692 );
and ( n44224 , n391060 , n391200 );
or ( n44225 , n44223 , n44224 );
buf ( n391696 , n44225 );
buf ( n391697 , n391696 );
not ( n44228 , n391697 );
buf ( n391699 , n44228 );
buf ( n391700 , n391699 );
not ( n44231 , n391700 );
xor ( n44232 , n43596 , n391076 );
and ( n44233 , n44232 , n391198 );
and ( n44234 , n43596 , n391076 );
or ( n44235 , n44233 , n44234 );
xor ( n44236 , n391105 , n391118 );
and ( n44237 , n44236 , n391196 );
and ( n44238 , n391105 , n391118 );
or ( n44239 , n44237 , n44238 );
buf ( n391710 , n44239 );
buf ( n391711 , n391710 );
buf ( n391712 , n390403 );
not ( n44243 , n391712 );
buf ( n391714 , n24074 );
not ( n44245 , n391714 );
buf ( n391716 , n38357 );
not ( n44247 , n391716 );
or ( n44248 , n44245 , n44247 );
buf ( n391719 , n37147 );
not ( n44250 , n391719 );
buf ( n391721 , n44250 );
buf ( n391722 , n391721 );
buf ( n391723 , n24073 );
nand ( n44254 , n391722 , n391723 );
buf ( n391725 , n44254 );
buf ( n391726 , n391725 );
nand ( n44257 , n44248 , n391726 );
buf ( n391728 , n44257 );
buf ( n391729 , n391728 );
not ( n44260 , n391729 );
or ( n44261 , n44243 , n44260 );
buf ( n391732 , n391080 );
buf ( n391733 , n391097 );
nand ( n44264 , n391732 , n391733 );
buf ( n391735 , n44264 );
buf ( n391736 , n391735 );
nand ( n44267 , n44261 , n391736 );
buf ( n391738 , n44267 );
buf ( n391739 , n391738 );
buf ( n391740 , n389547 );
buf ( n391741 , n388998 );
not ( n44277 , n391741 );
buf ( n391743 , n384096 );
not ( n44279 , n391743 );
or ( n44280 , n44277 , n44279 );
buf ( n391746 , n382854 );
buf ( n391747 , n388215 );
nand ( n44283 , n391746 , n391747 );
buf ( n391749 , n44283 );
buf ( n391750 , n391749 );
nand ( n44286 , n44280 , n391750 );
buf ( n391752 , n44286 );
buf ( n391753 , n391752 );
nand ( n44289 , n391740 , n391753 );
buf ( n391755 , n44289 );
buf ( n391756 , n391755 );
nand ( n44292 , C1 , n391756 );
buf ( n391758 , n44292 );
buf ( n391759 , n391758 );
buf ( n391760 , n384644 );
not ( n44296 , n391760 );
buf ( n391762 , n40775 );
not ( n44298 , n391762 );
buf ( n391764 , n44298 );
xor ( n44300 , n391764 , n389805 );
buf ( n391766 , n44300 );
not ( n44302 , n391766 );
or ( n44303 , n44296 , n44302 );
buf ( n391769 , n383894 );
buf ( n391770 , n389946 );
nand ( n44306 , n391769 , n391770 );
buf ( n391772 , n44306 );
buf ( n391773 , n391772 );
nand ( n44309 , n44303 , n391773 );
buf ( n391775 , n44309 );
buf ( n391776 , n391775 );
xor ( n44312 , n391759 , n391776 );
buf ( n391778 , n390004 );
not ( n44314 , n391778 );
buf ( n391780 , n382592 );
not ( n44316 , n391780 );
buf ( n391782 , n44316 );
buf ( n391783 , n391782 );
not ( n44319 , n391783 );
or ( n44320 , n44314 , n44319 );
buf ( n391786 , n389024 );
buf ( n391787 , n390490 );
not ( n44323 , n391787 );
buf ( n391789 , n385972 );
not ( n44325 , n391789 );
or ( n44326 , n44323 , n44325 );
buf ( n391792 , n385975 );
buf ( n391793 , n388569 );
nand ( n44329 , n391792 , n391793 );
buf ( n391795 , n44329 );
buf ( n391796 , n391795 );
nand ( n44332 , n44326 , n391796 );
buf ( n391798 , n44332 );
buf ( n391799 , n391798 );
nand ( n44335 , n391786 , n391799 );
buf ( n391801 , n44335 );
buf ( n391802 , n391801 );
nand ( n44338 , n44320 , n391802 );
buf ( n391804 , n44338 );
buf ( n391805 , n391804 );
xor ( n44341 , n44312 , n391805 );
buf ( n391807 , n44341 );
buf ( n391808 , n391807 );
xor ( n44344 , n391739 , n391808 );
xor ( n44345 , n391147 , n391160 );
and ( n44346 , n44345 , n391193 );
and ( n44347 , n391147 , n391160 );
or ( n44348 , n44346 , n44347 );
buf ( n391814 , n44348 );
buf ( n391815 , n391814 );
xor ( n44351 , n44344 , n391815 );
buf ( n391817 , n44351 );
buf ( n391818 , n391817 );
xor ( n44354 , n391711 , n391818 );
buf ( n391820 , n388809 );
not ( n44356 , n391820 );
buf ( n391822 , n388760 );
not ( n44358 , n391822 );
buf ( n391824 , n382548 );
not ( n44360 , n391824 );
or ( n44361 , n44358 , n44360 );
buf ( n391827 , n391212 );
buf ( n391828 , n388757 );
nand ( n44364 , n391827 , n391828 );
buf ( n391830 , n44364 );
buf ( n391831 , n391830 );
nand ( n44367 , n44361 , n391831 );
buf ( n391833 , n44367 );
buf ( n391834 , n391833 );
not ( n44370 , n391834 );
or ( n44371 , n44356 , n44370 );
buf ( n391837 , n388796 );
buf ( n391838 , n388746 );
nand ( n44374 , n391837 , n391838 );
buf ( n391840 , n44374 );
buf ( n391841 , n391840 );
nand ( n44377 , n44371 , n391841 );
buf ( n391843 , n44377 );
buf ( n391844 , n391843 );
not ( n44380 , n41565 );
and ( n44381 , n42152 , n389075 );
not ( n44382 , n42152 );
and ( n44383 , n44382 , n24050 );
or ( n44384 , n44381 , n44383 );
not ( n44385 , n44384 );
or ( n44386 , n44380 , n44385 );
buf ( n391852 , n389726 );
buf ( n391853 , n389125 );
nand ( n44389 , n391852 , n391853 );
buf ( n391855 , n44389 );
nand ( n44391 , n44386 , n391855 );
buf ( n391857 , n44391 );
xor ( n44393 , n391844 , n391857 );
buf ( n391859 , n391139 );
not ( n44395 , n391859 );
buf ( n391861 , n389883 );
not ( n44397 , n391861 );
or ( n44398 , n44395 , n44397 );
not ( n44399 , n41195 );
not ( n44400 , n44399 );
not ( n44401 , n384562 );
or ( n44402 , n44400 , n44401 );
buf ( n391868 , n384562 );
not ( n44404 , n391868 );
buf ( n391870 , n44404 );
buf ( n391871 , n391870 );
buf ( n391872 , n41195 );
nand ( n44408 , n391871 , n391872 );
buf ( n391874 , n44408 );
nand ( n44410 , n44402 , n391874 );
buf ( n391876 , n44410 );
buf ( n391877 , n389908 );
nand ( n44413 , n391876 , n391877 );
buf ( n391879 , n44413 );
buf ( n391880 , n391879 );
nand ( n44416 , n44398 , n391880 );
buf ( n391882 , n44416 );
buf ( n391883 , n391882 );
buf ( n391884 , n37695 );
not ( n44420 , n391884 );
buf ( n391886 , n37347 );
not ( n44422 , n391886 );
not ( n44423 , n36564 );
buf ( n391889 , n44423 );
not ( n44425 , n391889 );
or ( n44426 , n44422 , n44425 );
buf ( n391892 , n38155 );
buf ( n391893 , n37346 );
buf ( n44429 , n391893 );
buf ( n391895 , n44429 );
buf ( n391896 , n391895 );
nand ( n44432 , n391892 , n391896 );
buf ( n391898 , n44432 );
buf ( n391899 , n391898 );
nand ( n44435 , n44426 , n391899 );
buf ( n391901 , n44435 );
buf ( n391902 , n391901 );
not ( n44438 , n391902 );
or ( n44439 , n44420 , n44438 );
buf ( n391905 , n389968 );
not ( n44441 , n391905 );
buf ( n391907 , n385269 );
nand ( n44443 , n44441 , n391907 );
buf ( n391909 , n44443 );
buf ( n391910 , n391909 );
nand ( n44446 , n44439 , n391910 );
buf ( n391912 , n44446 );
buf ( n391913 , n391912 );
xor ( n44449 , n391883 , n391913 );
buf ( n391915 , n388539 );
not ( n44451 , n391915 );
buf ( n391917 , n44451 );
buf ( n391918 , n391917 );
not ( n44454 , n391918 );
buf ( n391920 , n44454 );
buf ( n391921 , n391920 );
buf ( n391922 , n391188 );
or ( n44458 , n391921 , n391922 );
buf ( n391924 , n391176 );
buf ( n391925 , n389589 );
buf ( n391926 , n388654 );
and ( n44462 , n391925 , n391926 );
buf ( n391928 , n391183 );
buf ( n391929 , n388646 );
and ( n44465 , n391928 , n391929 );
nor ( n44466 , n44462 , n44465 );
buf ( n391932 , n44466 );
buf ( n391933 , n391932 );
or ( n44469 , n391924 , n391933 );
nand ( n44470 , n44458 , n44469 );
buf ( n391936 , n44470 );
buf ( n391937 , n391936 );
xor ( n44473 , n44449 , n391937 );
buf ( n391939 , n44473 );
buf ( n391940 , n391939 );
xor ( n44476 , n44393 , n391940 );
buf ( n391942 , n44476 );
buf ( n391943 , n391942 );
xor ( n44479 , n44354 , n391943 );
buf ( n391945 , n44479 );
xor ( n44481 , n44235 , n391945 );
not ( n44482 , n43857 );
not ( n44483 , n44482 );
not ( n44484 , n43847 );
or ( n44485 , n44483 , n44484 );
buf ( n391951 , n391382 );
not ( n44487 , n391951 );
buf ( n391953 , n44487 );
nand ( n44489 , n44485 , n391953 );
buf ( n391955 , n44489 );
not ( n44491 , n43847 );
nand ( n44492 , n44491 , n43857 );
buf ( n391958 , n44492 );
nand ( n44494 , n391955 , n391958 );
buf ( n391960 , n44494 );
buf ( n391961 , n391960 );
xor ( n44497 , n388719 , n388816 );
xor ( n44498 , n44497 , n388879 );
buf ( n391964 , n44498 );
buf ( n391965 , n391964 );
xor ( n44501 , n391961 , n391965 );
xor ( n44502 , n388889 , n389142 );
xor ( n44503 , n44502 , n389213 );
buf ( n391969 , n44503 );
buf ( n391970 , n391969 );
and ( n44506 , n44501 , n391970 );
and ( n44507 , n391961 , n391965 );
or ( n44508 , n44506 , n44507 );
buf ( n391974 , n44508 );
xor ( n44510 , n44481 , n391974 );
buf ( n391976 , n44510 );
not ( n44512 , n391976 );
or ( n44513 , n44231 , n44512 );
xor ( n44514 , n44235 , n391945 );
xnor ( n44515 , n44514 , n391974 );
nand ( n44516 , n44515 , n391696 );
buf ( n391982 , n44516 );
nand ( n44518 , n44513 , n391982 );
buf ( n391984 , n44518 );
xor ( n44520 , n389244 , n389273 );
xor ( n44521 , n44520 , n389454 );
buf ( n391987 , n44521 );
not ( n44523 , n391987 );
buf ( n391989 , n389625 );
buf ( n391990 , n389670 );
xor ( n44526 , n391989 , n391990 );
buf ( n391992 , n389621 );
xnor ( n44528 , n44526 , n391992 );
buf ( n391994 , n44528 );
buf ( n391995 , n391994 );
not ( n44531 , n391995 );
or ( n44532 , n44523 , n44531 );
buf ( n391998 , n391366 );
buf ( n391999 , n391345 );
xor ( n44535 , n391998 , n391999 );
buf ( n392001 , n391376 );
xor ( n44537 , n44535 , n392001 );
buf ( n392003 , n44537 );
buf ( n392004 , n392003 );
xor ( n44540 , n389307 , n389414 );
xor ( n44541 , n44540 , n389450 );
buf ( n392007 , n44541 );
buf ( n392008 , n392007 );
xor ( n44544 , n392004 , n392008 );
buf ( n392010 , n388141 );
not ( n44546 , n392010 );
buf ( n392012 , n42160 );
not ( n44548 , n392012 );
or ( n44549 , n44546 , n44548 );
and ( n44550 , n36216 , n388157 );
not ( n44551 , n36216 );
and ( n44552 , n44551 , n388160 );
or ( n44553 , n44550 , n44552 );
buf ( n392019 , n44553 );
buf ( n392020 , n40701 );
nand ( n44556 , n392019 , n392020 );
buf ( n392022 , n44556 );
buf ( n392023 , n392022 );
nand ( n44559 , n44549 , n392023 );
buf ( n392025 , n44559 );
buf ( n392026 , n392025 );
buf ( n392027 , n389359 );
not ( n44563 , n392027 );
buf ( n392029 , n38685 );
not ( n44565 , n392029 );
or ( n44566 , n44563 , n44565 );
buf ( n392032 , n35435 );
buf ( n392033 , n389356 );
nand ( n44569 , n392032 , n392033 );
buf ( n392035 , n44569 );
buf ( n392036 , n392035 );
nand ( n44572 , n44566 , n392036 );
buf ( n392038 , n44572 );
buf ( n392039 , n392038 );
not ( n44575 , n392039 );
buf ( n392041 , n38765 );
not ( n44577 , n392041 );
or ( n44578 , n44575 , n44577 );
buf ( n392044 , n390635 );
buf ( n392045 , n43148 );
nand ( n44581 , n392044 , n392045 );
buf ( n392047 , n44581 );
buf ( n392048 , n392047 );
nand ( n44584 , n44578 , n392048 );
buf ( n392050 , n44584 );
buf ( n392051 , n392050 );
not ( n44587 , n388962 );
not ( n44588 , n43044 );
or ( n44589 , n44587 , n44588 );
buf ( n392055 , n27195 );
buf ( n392056 , n385488 );
nand ( n44592 , n392055 , n392056 );
buf ( n392058 , n44592 );
nand ( n44594 , n44589 , n392058 );
not ( n44595 , n44594 );
not ( n44596 , n43240 );
or ( n44597 , n44595 , n44596 );
nand ( n44598 , n41447 , n44087 );
nand ( n44599 , n44597 , n44598 );
buf ( n392065 , n44599 );
buf ( n392066 , n389862 );
not ( n44602 , n392066 );
buf ( n392068 , n40973 );
not ( n44604 , n392068 );
or ( n44605 , n44602 , n44604 );
buf ( n392071 , n40839 );
buf ( n392072 , n389859 );
nand ( n44608 , n392071 , n392072 );
buf ( n392074 , n44608 );
buf ( n392075 , n392074 );
nand ( n44611 , n44605 , n392075 );
buf ( n392077 , n44611 );
buf ( n392078 , n392077 );
not ( n44614 , n392078 );
buf ( n392080 , n390832 );
not ( n44616 , n392080 );
or ( n44617 , n44614 , n44616 );
buf ( n392083 , n388346 );
buf ( n392084 , n390730 );
nand ( n44620 , n392083 , n392084 );
buf ( n392086 , n44620 );
buf ( n392087 , n392086 );
nand ( n44623 , n44617 , n392087 );
buf ( n392089 , n44623 );
buf ( n392090 , n392089 );
xor ( n44626 , n392065 , n392090 );
buf ( n392092 , n388543 );
not ( n44628 , n392092 );
buf ( n392094 , n40886 );
not ( n44630 , n392094 );
or ( n44631 , n44628 , n44630 );
buf ( n392097 , n388546 );
buf ( n392098 , n40885 );
nand ( n44634 , n392097 , n392098 );
buf ( n392100 , n44634 );
buf ( n392101 , n392100 );
nand ( n44637 , n44631 , n392101 );
buf ( n392103 , n44637 );
buf ( n392104 , n392103 );
not ( n44640 , n392104 );
buf ( n392106 , n40858 );
not ( n44642 , n392106 );
or ( n44643 , n44640 , n44642 );
buf ( n392109 , n36845 );
not ( n44645 , n392109 );
buf ( n392111 , n44645 );
buf ( n392112 , n392111 );
buf ( n392113 , n390936 );
nand ( n44649 , n392112 , n392113 );
buf ( n392115 , n44649 );
buf ( n392116 , n392115 );
nand ( n44652 , n44643 , n392116 );
buf ( n392118 , n44652 );
buf ( n392119 , n392118 );
and ( n44655 , n44626 , n392119 );
and ( n44656 , n392065 , n392090 );
or ( n44657 , n44655 , n44656 );
buf ( n392123 , n44657 );
buf ( n392124 , n392123 );
xor ( n44660 , n392051 , n392124 );
xor ( n44661 , n43209 , n43242 );
xor ( n44662 , n44661 , n43276 );
buf ( n392128 , n44662 );
and ( n44664 , n44660 , n392128 );
and ( n44665 , n392051 , n392124 );
or ( n44666 , n44664 , n44665 );
buf ( n392132 , n44666 );
buf ( n392133 , n392132 );
xor ( n44669 , n392026 , n392133 );
buf ( n392135 , n43515 );
not ( n44671 , n392135 );
buf ( n392137 , n391219 );
not ( n44673 , n392137 );
or ( n44674 , n44671 , n44673 );
buf ( n392140 , n391027 );
not ( n44676 , n392140 );
buf ( n392142 , n35519 );
not ( n44678 , n392142 );
buf ( n392144 , n44678 );
buf ( n392145 , n392144 );
not ( n44681 , n392145 );
or ( n44682 , n44676 , n44681 );
buf ( n392148 , n35519 );
buf ( n392149 , n391024 );
nand ( n44685 , n392148 , n392149 );
buf ( n392151 , n44685 );
buf ( n392152 , n392151 );
nand ( n44688 , n44682 , n392152 );
buf ( n392154 , n44688 );
buf ( n392155 , n392154 );
buf ( n392156 , n43727 );
nand ( n44692 , n392155 , n392156 );
buf ( n392158 , n44692 );
buf ( n392159 , n392158 );
nand ( n44695 , n44674 , n392159 );
buf ( n392161 , n44695 );
buf ( n392162 , n392161 );
and ( n44698 , n44669 , n392162 );
and ( n44699 , n392026 , n392133 );
or ( n44700 , n44698 , n44699 );
buf ( n392166 , n44700 );
buf ( n392167 , n392166 );
and ( n44703 , n44544 , n392167 );
and ( n44704 , n392004 , n392008 );
or ( n44705 , n44703 , n44704 );
buf ( n392171 , n44705 );
buf ( n392172 , n392171 );
nand ( n44708 , n44532 , n392172 );
buf ( n392174 , n44708 );
buf ( n392175 , n392174 );
buf ( n392176 , n391994 );
not ( n44712 , n392176 );
buf ( n392178 , n44712 );
buf ( n392179 , n392178 );
buf ( n392180 , n44521 );
not ( n44716 , n392180 );
buf ( n392182 , n44716 );
buf ( n392183 , n392182 );
nand ( n44719 , n392179 , n392183 );
buf ( n392185 , n44719 );
buf ( n392186 , n392185 );
nand ( n44722 , n392175 , n392186 );
buf ( n392188 , n44722 );
xor ( n44724 , n391961 , n391965 );
xor ( n44725 , n44724 , n391970 );
buf ( n392191 , n44725 );
or ( n44727 , n392188 , n392191 );
xor ( n44728 , n389460 , n42188 );
xor ( n44729 , n44728 , n390033 );
nand ( n44730 , n44727 , n44729 );
nand ( n44731 , n392188 , n392191 );
nand ( n44732 , n44730 , n44731 );
and ( n44733 , n391984 , n44732 );
not ( n44734 , n391984 );
not ( n44735 , n44732 );
and ( n44736 , n44734 , n44735 );
nor ( n44737 , n44733 , n44736 );
not ( n44738 , n44737 );
xor ( n44739 , n42852 , n44738 );
not ( n44740 , n388833 );
not ( n44741 , n389442 );
or ( n44742 , n44740 , n44741 );
buf ( n392208 , n388872 );
xor ( n44744 , n41342 , n37173 );
buf ( n392210 , n44744 );
nand ( n44746 , n392208 , n392210 );
buf ( n392212 , n44746 );
nand ( n44748 , n44742 , n392212 );
buf ( n392214 , n44748 );
buf ( n392215 , n371925 );
buf ( n44751 , n392215 );
buf ( n392217 , n44751 );
buf ( n392218 , n392217 );
buf ( n392219 , n371278 );
xor ( n44755 , n392218 , n392219 );
buf ( n392221 , n44755 );
buf ( n392222 , n392221 );
not ( n44758 , n392222 );
buf ( n392224 , n44758 );
buf ( n392225 , n392224 );
not ( n44761 , n392225 );
and ( n44762 , n23701 , n371278 );
not ( n44763 , n23701 );
buf ( n392229 , n371278 );
not ( n44765 , n392229 );
buf ( n392231 , n44765 );
and ( n44767 , n44763 , n392231 );
nor ( n44768 , n44762 , n44767 );
nand ( n44769 , n44768 , n392224 );
not ( n44770 , n44769 );
not ( n44771 , n44770 );
buf ( n392237 , n44771 );
not ( n44773 , n392237 );
or ( n44774 , n44761 , n44773 );
buf ( n44775 , n23701 );
not ( n44776 , n44775 );
buf ( n392242 , n44776 );
buf ( n44778 , n392242 );
buf ( n392244 , n44778 );
buf ( n392245 , n392244 );
not ( n44781 , n392245 );
buf ( n392247 , n44781 );
buf ( n392248 , n392247 );
not ( n44784 , n392248 );
buf ( n392250 , n388113 );
not ( n44786 , n392250 );
or ( n44787 , n44784 , n44786 );
buf ( n392253 , n385499 );
buf ( n392254 , n392244 );
nand ( n44790 , n392253 , n392254 );
buf ( n392256 , n44790 );
buf ( n392257 , n392256 );
nand ( n44793 , n44787 , n392257 );
buf ( n392259 , n44793 );
buf ( n392260 , n392259 );
nand ( n44796 , n44774 , n392260 );
buf ( n392262 , n44796 );
buf ( n392263 , n392262 );
nor ( n44799 , n392214 , n392263 );
buf ( n392265 , n44799 );
buf ( n392266 , n392265 );
not ( n44802 , n392266 );
buf ( n392268 , n44802 );
buf ( n392269 , n392268 );
not ( n44805 , n392269 );
xor ( n44806 , n391254 , n391282 );
xor ( n44807 , n44806 , n391287 );
buf ( n392273 , n44807 );
buf ( n392274 , n392273 );
not ( n44810 , n392274 );
or ( n44811 , n44805 , n44810 );
nand ( n44812 , n44748 , n392262 );
buf ( n392278 , n44812 );
nand ( n44814 , n44811 , n392278 );
buf ( n392280 , n44814 );
not ( n44816 , n392280 );
buf ( n392282 , n389631 );
buf ( n392283 , n389654 );
xor ( n44819 , n392282 , n392283 );
buf ( n392285 , n389659 );
xnor ( n44821 , n44819 , n392285 );
buf ( n392287 , n44821 );
nand ( n44823 , n44816 , n392287 );
xor ( n44824 , n391229 , n391291 );
xor ( n44825 , n44824 , n391316 );
and ( n44826 , n44823 , n44825 );
nor ( n44827 , n392287 , n44816 );
nor ( n44828 , n44826 , n44827 );
buf ( n392294 , n44828 );
not ( n44830 , n392294 );
buf ( n392296 , n44830 );
buf ( n392297 , n392296 );
not ( n44833 , n392297 );
buf ( n392299 , n388102 );
not ( n44835 , n392299 );
buf ( n392301 , n386561 );
not ( n44837 , n392301 );
or ( n44838 , n44835 , n44837 );
buf ( n392304 , n382921 );
buf ( n392305 , n388105 );
nand ( n44841 , n392304 , n392305 );
buf ( n392307 , n44841 );
buf ( n392308 , n392307 );
nand ( n44844 , n44838 , n392308 );
buf ( n392310 , n44844 );
buf ( n392311 , n392310 );
buf ( n392312 , n43286 );
and ( n44848 , n392311 , n392312 );
not ( n44849 , n390775 );
nor ( n44850 , n44849 , n388071 );
buf ( n392316 , n44850 );
nor ( n44852 , n44848 , n392316 );
buf ( n392318 , n44852 );
buf ( n392319 , n392318 );
not ( n44855 , n392319 );
buf ( n392321 , n44855 );
buf ( n392322 , n392321 );
not ( n44858 , n392322 );
buf ( n392324 , n388809 );
not ( n44860 , n392324 );
buf ( n392326 , n391428 );
not ( n44862 , n392326 );
or ( n44863 , n44860 , n44862 );
buf ( n392329 , n388760 );
not ( n44865 , n392329 );
buf ( n392331 , n35997 );
not ( n44867 , n392331 );
buf ( n392333 , n44867 );
buf ( n392334 , n392333 );
not ( n44870 , n392334 );
or ( n44871 , n44865 , n44870 );
buf ( n392337 , n35997 );
buf ( n392338 , n388757 );
nand ( n44874 , n392337 , n392338 );
buf ( n392340 , n44874 );
buf ( n392341 , n392340 );
nand ( n44877 , n44871 , n392341 );
buf ( n392343 , n44877 );
buf ( n392344 , n392343 );
buf ( n392345 , n388746 );
nand ( n44881 , n392344 , n392345 );
buf ( n392347 , n44881 );
buf ( n392348 , n392347 );
nand ( n44884 , n44863 , n392348 );
buf ( n392350 , n44884 );
buf ( n392351 , n392350 );
not ( n44887 , n392351 );
or ( n44888 , n44858 , n44887 );
buf ( n392354 , n392321 );
buf ( n392355 , n392350 );
or ( n44891 , n392354 , n392355 );
xor ( n44892 , n43348 , n390971 );
xor ( n44893 , n44892 , n390907 );
buf ( n392359 , n44893 );
nand ( n44895 , n44891 , n392359 );
buf ( n392361 , n44895 );
buf ( n392362 , n392361 );
nand ( n44898 , n44888 , n392362 );
buf ( n392364 , n44898 );
buf ( n392365 , n392364 );
not ( n44901 , n392365 );
xor ( n44902 , n390759 , n43312 );
xnor ( n44903 , n44902 , n43500 );
buf ( n392369 , n44903 );
not ( n44905 , n392369 );
or ( n44906 , n44901 , n44905 );
buf ( n392372 , n44903 );
buf ( n392373 , n392364 );
or ( n44909 , n392372 , n392373 );
xor ( n44910 , n390643 , n390667 );
xor ( n44911 , n44910 , n390755 );
buf ( n392377 , n44911 );
buf ( n392378 , n392377 );
xor ( n44914 , n390921 , n390949 );
xor ( n44915 , n44914 , n390967 );
buf ( n392381 , n44915 );
not ( n44917 , n392381 );
buf ( n392383 , n40701 );
not ( n44919 , n392383 );
buf ( n392385 , n388157 );
buf ( n392386 , n389067 );
and ( n44922 , n392385 , n392386 );
not ( n44923 , n392385 );
buf ( n392389 , n384180 );
and ( n44925 , n44923 , n392389 );
nor ( n44926 , n44922 , n44925 );
buf ( n392392 , n44926 );
buf ( n392393 , n392392 );
not ( n44929 , n392393 );
or ( n44930 , n44919 , n44929 );
buf ( n392396 , n44553 );
buf ( n392397 , n388141 );
nand ( n44933 , n392396 , n392397 );
buf ( n392399 , n44933 );
buf ( n392400 , n392399 );
nand ( n44936 , n44930 , n392400 );
buf ( n392402 , n44936 );
buf ( n392403 , n391080 );
not ( n44939 , n392403 );
buf ( n392405 , n24074 );
not ( n44941 , n392405 );
buf ( n392407 , n389467 );
not ( n44943 , n392407 );
or ( n44944 , n44941 , n44943 );
not ( n44945 , n36708 );
buf ( n392411 , n44945 );
buf ( n392412 , n24073 );
nand ( n44948 , n392411 , n392412 );
buf ( n392414 , n44948 );
buf ( n392415 , n392414 );
nand ( n44951 , n44944 , n392415 );
buf ( n392417 , n44951 );
buf ( n392418 , n392417 );
not ( n44954 , n392418 );
or ( n44955 , n44939 , n44954 );
buf ( n392421 , n390820 );
buf ( n392422 , n390403 );
nand ( n44958 , n392421 , n392422 );
buf ( n392424 , n44958 );
buf ( n392425 , n392424 );
nand ( n44961 , n44955 , n392425 );
buf ( n392427 , n44961 );
or ( n44963 , n392402 , n392427 );
not ( n44964 , n44963 );
or ( n44965 , n44917 , n44964 );
nand ( n44966 , n392402 , n392427 );
nand ( n44967 , n44965 , n44966 );
buf ( n392433 , n44967 );
xor ( n44969 , n392378 , n392433 );
buf ( n392435 , n389162 );
not ( n44971 , n392435 );
buf ( n392437 , n391306 );
not ( n44973 , n392437 );
or ( n44974 , n44971 , n44973 );
buf ( n392440 , n41671 );
not ( n44976 , n392440 );
buf ( n392442 , n385774 );
not ( n44978 , n392442 );
or ( n44979 , n44976 , n44978 );
buf ( n392445 , n38227 );
buf ( n392446 , n41678 );
nand ( n44982 , n392445 , n392446 );
buf ( n392448 , n44982 );
buf ( n392449 , n392448 );
nand ( n44985 , n44979 , n392449 );
buf ( n392451 , n44985 );
buf ( n392452 , n392451 );
buf ( n392453 , n41711 );
nand ( n44989 , n392452 , n392453 );
buf ( n392455 , n44989 );
buf ( n392456 , n392455 );
nand ( n44992 , n44974 , n392456 );
buf ( n392458 , n44992 );
buf ( n392459 , n392458 );
and ( n44995 , n44969 , n392459 );
and ( n44996 , n392378 , n392433 );
or ( n44997 , n44995 , n44996 );
buf ( n392463 , n44997 );
buf ( n392464 , n392463 );
nand ( n45000 , n44909 , n392464 );
buf ( n392466 , n45000 );
buf ( n392467 , n392466 );
nand ( n45003 , n44906 , n392467 );
buf ( n392469 , n45003 );
buf ( n392470 , n392469 );
not ( n45006 , n392470 );
or ( n45007 , n44833 , n45006 );
buf ( n392473 , n392469 );
not ( n45009 , n392473 );
buf ( n392475 , n45009 );
buf ( n392476 , n392475 );
not ( n45012 , n392476 );
buf ( n392478 , n44828 );
not ( n45014 , n392478 );
or ( n45015 , n45012 , n45014 );
xor ( n45016 , n43504 , n391057 );
xor ( n45017 , n45016 , n43138 );
buf ( n392483 , n45017 );
nand ( n45019 , n45015 , n392483 );
buf ( n392485 , n45019 );
buf ( n392486 , n392485 );
nand ( n45022 , n45007 , n392486 );
buf ( n392488 , n45022 );
buf ( n392489 , n392488 );
not ( n45025 , n392489 );
xor ( n45026 , n391060 , n391200 );
xor ( n45027 , n45026 , n391692 );
buf ( n392493 , n45027 );
buf ( n392494 , n392493 );
not ( n45030 , n392494 );
buf ( n392496 , n45030 );
buf ( n392497 , n392496 );
nand ( n45033 , n45025 , n392497 );
buf ( n392499 , n45033 );
not ( n45035 , n392499 );
xor ( n45036 , n391320 , n391395 );
xor ( n45037 , n45036 , n391687 );
buf ( n392503 , n45037 );
buf ( n392504 , n392503 );
not ( n45040 , n392504 );
buf ( n392506 , n392171 );
buf ( n392507 , n392182 );
xor ( n45043 , n392506 , n392507 );
buf ( n392509 , n392178 );
xnor ( n45045 , n45043 , n392509 );
buf ( n392511 , n45045 );
buf ( n392512 , n392511 );
not ( n45048 , n392512 );
buf ( n392514 , n45048 );
buf ( n392515 , n392514 );
not ( n45051 , n392515 );
or ( n45052 , n45040 , n45051 );
buf ( n392518 , n392503 );
not ( n45054 , n392518 );
buf ( n392520 , n45054 );
buf ( n392521 , n392520 );
not ( n45057 , n392521 );
buf ( n392523 , n392511 );
not ( n45059 , n392523 );
or ( n45060 , n45057 , n45059 );
xor ( n45061 , n391415 , n391436 );
xor ( n45062 , n45061 , n391682 );
buf ( n392528 , n45062 );
buf ( n392529 , n392528 );
not ( n45065 , n389162 );
not ( n45066 , n392451 );
or ( n45067 , n45065 , n45066 );
not ( n392533 , n41671 );
not ( n45069 , n37147 );
or ( n45070 , n392533 , n45069 );
buf ( n392536 , n391721 );
buf ( n392537 , n41678 );
nand ( n45073 , n392536 , n392537 );
buf ( n392539 , n45073 );
nand ( n45075 , n45070 , n392539 );
not ( n45076 , n41709 );
nand ( n45077 , n45075 , n45076 );
nand ( n45078 , n45067 , n45077 );
not ( n45079 , n45078 );
buf ( n392545 , n391500 );
buf ( n392546 , n391468 );
xor ( n45082 , n392545 , n392546 );
buf ( n392548 , n391526 );
xnor ( n45084 , n45082 , n392548 );
buf ( n392550 , n45084 );
buf ( n392551 , n392550 );
not ( n45087 , n392551 );
buf ( n392553 , n45087 );
not ( n45089 , n392553 );
or ( n45090 , n45079 , n45089 );
not ( n45091 , n392550 );
buf ( n392557 , n45078 );
not ( n45093 , n392557 );
buf ( n392559 , n45093 );
not ( n45095 , n392559 );
or ( n45096 , n45091 , n45095 );
buf ( n392562 , n386480 );
not ( n45098 , n392562 );
buf ( n392564 , n391493 );
not ( n45100 , n392564 );
or ( n45101 , n45098 , n45100 );
not ( n45102 , n22982 );
and ( n45103 , n28159 , n45102 );
not ( n45104 , n28159 );
and ( n45105 , n45104 , n22982 );
or ( n45106 , n45103 , n45105 );
buf ( n392572 , n45106 );
buf ( n392573 , n386496 );
nand ( n45109 , n392572 , n392573 );
buf ( n392575 , n45109 );
buf ( n392576 , n392575 );
nand ( n45112 , n45101 , n392576 );
buf ( n392578 , n45112 );
buf ( n392579 , n392578 );
buf ( n392580 , n42073 );
not ( n45116 , n392580 );
buf ( n392582 , n385972 );
not ( n45118 , n392582 );
or ( n45119 , n45116 , n45118 );
buf ( n392585 , n389759 );
buf ( n392586 , n42074 );
nand ( n45122 , n392585 , n392586 );
buf ( n392588 , n45122 );
buf ( n392589 , n392588 );
nand ( n45125 , n45119 , n392589 );
buf ( n392591 , n45125 );
buf ( n392592 , n392591 );
not ( n45128 , n392592 );
buf ( n392594 , n389015 );
not ( n45130 , n392594 );
or ( n45131 , n45128 , n45130 );
buf ( n392597 , n386209 );
buf ( n392598 , n43479 );
nand ( n45134 , n392597 , n392598 );
buf ( n392600 , n45134 );
buf ( n392601 , n392600 );
nand ( n45137 , n45131 , n392601 );
buf ( n392603 , n45137 );
buf ( n392604 , n392603 );
xor ( n45140 , n392579 , n392604 );
buf ( n392606 , n372471 );
buf ( n45143 , n392606 );
buf ( n392608 , n45143 );
buf ( n392609 , n392608 );
buf ( n45146 , n392609 );
buf ( n392611 , n45146 );
buf ( n392612 , n392611 );
not ( n45149 , n392612 );
buf ( n392614 , n384096 );
not ( n45151 , n392614 );
or ( n45152 , n45149 , n45151 );
buf ( n392617 , n385292 );
buf ( n392618 , n392611 );
not ( n45155 , n392618 );
buf ( n392620 , n45155 );
buf ( n392621 , n392620 );
nand ( n45158 , n392617 , n392621 );
buf ( n392623 , n45158 );
buf ( n392624 , n392623 );
nand ( n45161 , n45152 , n392624 );
buf ( n392626 , n45161 );
buf ( n392627 , n386161 );
buf ( n392628 , n391461 );
not ( n45170 , n392628 );
buf ( n392630 , n45170 );
buf ( n392631 , n392630 );
or ( n45173 , n392627 , n392631 );
nand ( n45174 , C1 , n45173 );
buf ( n392634 , n45174 );
buf ( n392635 , n392634 );
and ( n45177 , n45140 , n392635 );
and ( n45178 , n392579 , n392604 );
or ( n45179 , n45177 , n45178 );
buf ( n392639 , n45179 );
nand ( n45181 , n45096 , n392639 );
nand ( n45182 , n45090 , n45181 );
buf ( n392642 , n45182 );
buf ( n392643 , n388230 );
not ( n45185 , n392643 );
buf ( n392645 , n391129 );
not ( n45187 , n392645 );
or ( n45188 , n45185 , n45187 );
buf ( n392648 , n389894 );
buf ( n392649 , n388242 );
nand ( n45191 , n392648 , n392649 );
buf ( n392651 , n45191 );
buf ( n392652 , n392651 );
nand ( n45194 , n45188 , n392652 );
buf ( n392654 , n45194 );
buf ( n392655 , n392654 );
not ( n45197 , n392655 );
buf ( n392657 , n384621 );
not ( n45199 , n392657 );
buf ( n392659 , n45199 );
buf ( n392660 , n392659 );
not ( n45202 , n392660 );
or ( n45203 , n45197 , n45202 );
buf ( n392663 , n391626 );
buf ( n392664 , n384548 );
buf ( n45206 , n392664 );
buf ( n392666 , n45206 );
buf ( n392667 , n392666 );
nand ( n45209 , n392663 , n392667 );
buf ( n392669 , n45209 );
buf ( n392670 , n392669 );
nand ( n45212 , n45203 , n392670 );
buf ( n392672 , n45212 );
buf ( n392673 , n392672 );
not ( n45215 , n392673 );
buf ( n392675 , n45215 );
buf ( n392676 , n392675 );
not ( n45218 , n392676 );
and ( n45219 , n391516 , n41565 );
and ( n45220 , n24050 , n388949 );
not ( n45221 , n24050 );
and ( n45222 , n45221 , n37763 );
or ( n45223 , n45220 , n45222 );
and ( n45224 , n45223 , n389125 );
nor ( n45225 , n45219 , n45224 );
buf ( n392685 , n45225 );
not ( n45227 , n392685 );
or ( n45228 , n45218 , n45227 );
buf ( n392688 , n383476 );
buf ( n392689 , n388502 );
buf ( n392690 , n383420 );
and ( n45232 , n392689 , n392690 );
not ( n45233 , n392689 );
buf ( n392693 , n388556 );
and ( n45235 , n45233 , n392693 );
nor ( n45236 , n45232 , n45235 );
buf ( n392696 , n45236 );
buf ( n392697 , n392696 );
or ( n45239 , n392688 , n392697 );
buf ( n392699 , n383403 );
buf ( n392700 , n391664 );
or ( n45242 , n392699 , n392700 );
nand ( n45243 , n45239 , n45242 );
buf ( n392703 , n45243 );
buf ( n392704 , n392703 );
nand ( n45246 , n45228 , n392704 );
buf ( n392706 , n45246 );
buf ( n392707 , n392706 );
buf ( n392708 , n45225 );
not ( n45250 , n392708 );
buf ( n392710 , n45250 );
buf ( n392711 , n392710 );
buf ( n392712 , n392672 );
nand ( n45254 , n392711 , n392712 );
buf ( n392714 , n45254 );
buf ( n392715 , n392714 );
nand ( n45257 , n392707 , n392715 );
buf ( n392717 , n45257 );
buf ( n392718 , n392717 );
buf ( n45260 , n44770 );
buf ( n392720 , n45260 );
not ( n45262 , n392720 );
buf ( n392722 , n392247 );
not ( n45264 , n392722 );
buf ( n392724 , n382548 );
not ( n45266 , n392724 );
or ( n45267 , n45264 , n45266 );
buf ( n392727 , n390345 );
buf ( n392728 , n392244 );
nand ( n45270 , n392727 , n392728 );
buf ( n392730 , n45270 );
buf ( n392731 , n392730 );
nand ( n45273 , n45267 , n392731 );
buf ( n392733 , n45273 );
buf ( n392734 , n392733 );
not ( n45276 , n392734 );
or ( n45277 , n45262 , n45276 );
buf ( n392737 , n392259 );
buf ( n392738 , n392224 );
not ( n45280 , n392738 );
buf ( n392740 , n45280 );
buf ( n392741 , n392740 );
nand ( n45283 , n392737 , n392741 );
buf ( n392743 , n45283 );
buf ( n392744 , n392743 );
nand ( n45286 , n45277 , n392744 );
buf ( n392746 , n45286 );
buf ( n392747 , n392746 );
xor ( n45289 , n392718 , n392747 );
xor ( n45290 , n391614 , n391645 );
xor ( n45291 , n45290 , n391672 );
buf ( n392751 , n45291 );
buf ( n392752 , n392751 );
and ( n45294 , n45289 , n392752 );
and ( n45295 , n392718 , n392747 );
or ( n45296 , n45294 , n45295 );
buf ( n392756 , n45296 );
buf ( n392757 , n392756 );
xor ( n45299 , n392642 , n392757 );
xor ( n45300 , n391538 , n391542 );
xor ( n45301 , n45300 , n391677 );
buf ( n392761 , n45301 );
buf ( n392762 , n392761 );
and ( n45304 , n45299 , n392762 );
and ( n45305 , n392642 , n392757 );
or ( n45306 , n45304 , n45305 );
buf ( n392766 , n45306 );
buf ( n392767 , n392766 );
xor ( n45309 , n392529 , n392767 );
buf ( n392769 , n388746 );
not ( n45311 , n392769 );
and ( n45312 , n36066 , n388757 );
not ( n45313 , n36066 );
and ( n45314 , n45313 , n388760 );
or ( n45315 , n45312 , n45314 );
buf ( n392775 , n45315 );
not ( n45317 , n392775 );
or ( n45318 , n45311 , n45317 );
buf ( n392778 , n392343 );
buf ( n392779 , n388809 );
nand ( n45321 , n392778 , n392779 );
buf ( n392781 , n45321 );
buf ( n392782 , n392781 );
nand ( n45324 , n45318 , n392782 );
buf ( n392784 , n45324 );
buf ( n392785 , n392784 );
buf ( n392786 , n42925 );
not ( n45328 , n392786 );
buf ( n392788 , n45328 );
buf ( n392789 , n392788 );
not ( n45331 , n392789 );
buf ( n392791 , n392417 );
not ( n45333 , n392791 );
or ( n45334 , n45331 , n45333 );
buf ( n392794 , n24074 );
not ( n45336 , n392794 );
buf ( n392796 , n384083 );
not ( n45338 , n392796 );
or ( n45339 , n45336 , n45338 );
buf ( n392799 , n384092 );
buf ( n392800 , n24073 );
nand ( n45342 , n392799 , n392800 );
buf ( n392802 , n45342 );
buf ( n392803 , n392802 );
nand ( n45345 , n45339 , n392803 );
buf ( n392805 , n45345 );
buf ( n392806 , n392805 );
buf ( n392807 , n391080 );
nand ( n45349 , n392806 , n392807 );
buf ( n392809 , n45349 );
buf ( n392810 , n392809 );
nand ( n45352 , n45334 , n392810 );
buf ( n392812 , n45352 );
buf ( n392813 , n392812 );
not ( n45355 , n392813 );
buf ( n392815 , n45355 );
not ( n45357 , n392815 );
buf ( n392817 , n389359 );
not ( n45359 , n392817 );
buf ( n392819 , n382994 );
not ( n45361 , n392819 );
or ( n45362 , n45359 , n45361 );
buf ( n392822 , n389759 );
buf ( n392823 , n389356 );
nand ( n45365 , n392822 , n392823 );
buf ( n392825 , n45365 );
buf ( n392826 , n392825 );
nand ( n45368 , n45362 , n392826 );
buf ( n392828 , n45368 );
buf ( n392829 , n392828 );
not ( n45371 , n392829 );
buf ( n392831 , n31850 );
buf ( n392832 , n382586 );
and ( n45374 , n392831 , n392832 );
buf ( n392834 , n45374 );
buf ( n392835 , n392834 );
not ( n45377 , n392835 );
or ( n45378 , n45371 , n45377 );
buf ( n392838 , n31850 );
not ( n45380 , n392838 );
buf ( n392840 , n392591 );
nand ( n45382 , n45380 , n392840 );
buf ( n392842 , n45382 );
buf ( n392843 , n392842 );
nand ( n45385 , n45378 , n392843 );
buf ( n392845 , n45385 );
buf ( n392846 , n392845 );
not ( n45388 , n392846 );
buf ( n392848 , n389125 );
not ( n45390 , n392848 );
not ( n45391 , n24049 );
buf ( n392851 , n45391 );
buf ( n392852 , n388979 );
and ( n45394 , n392851 , n392852 );
not ( n45395 , n392851 );
buf ( n392855 , n29077 );
and ( n45397 , n45395 , n392855 );
nor ( n45398 , n45394 , n45397 );
buf ( n392858 , n45398 );
buf ( n392859 , n392858 );
not ( n45401 , n392859 );
or ( n45402 , n45390 , n45401 );
buf ( n392862 , n45223 );
buf ( n392863 , n41565 );
nand ( n45405 , n392862 , n392863 );
buf ( n392865 , n45405 );
buf ( n392866 , n392865 );
nand ( n45408 , n45402 , n392866 );
buf ( n392868 , n45408 );
buf ( n392869 , n392868 );
not ( n45411 , n392869 );
buf ( n392871 , n45411 );
buf ( n392872 , n392871 );
nand ( n45414 , n45388 , n392872 );
buf ( n392874 , n45414 );
buf ( n392875 , n392874 );
buf ( n392876 , n24841 );
not ( n45418 , n392876 );
buf ( n392878 , n45418 );
buf ( n392879 , n392878 );
buf ( n45421 , n392879 );
buf ( n392881 , n45421 );
buf ( n392882 , n392881 );
not ( n45424 , n392882 );
buf ( n392884 , n45424 );
buf ( n392885 , n392884 );
not ( n45427 , n392885 );
buf ( n392887 , n45427 );
buf ( n392888 , n392887 );
buf ( n392889 , n385328 );
and ( n45431 , n392888 , n392889 );
not ( n45432 , n392888 );
buf ( n392892 , n384143 );
and ( n45434 , n45432 , n392892 );
nor ( n45435 , n45431 , n45434 );
buf ( n392895 , n45435 );
buf ( n392896 , n389547 );
buf ( n392897 , n392626 );
nand ( n45446 , n392896 , n392897 );
buf ( n392899 , n45446 );
buf ( n392900 , n392899 );
nand ( n45449 , C1 , n392900 );
buf ( n392902 , n45449 );
buf ( n392903 , n392902 );
and ( n45452 , n392875 , n392903 );
buf ( n392905 , n392845 );
buf ( n392906 , n392868 );
and ( n45455 , n392905 , n392906 );
buf ( n392908 , n45455 );
buf ( n392909 , n392908 );
nor ( n45458 , n45452 , n392909 );
buf ( n392911 , n45458 );
not ( n45460 , n392911 );
or ( n45461 , n45357 , n45460 );
buf ( n392914 , n44599 );
not ( n45463 , n392914 );
buf ( n392916 , n389602 );
not ( n45465 , n392916 );
buf ( n392918 , n390875 );
not ( n45467 , n392918 );
or ( n45468 , n45465 , n45467 );
buf ( n392921 , n36810 );
buf ( n392922 , n389593 );
nand ( n45471 , n392921 , n392922 );
buf ( n392924 , n45471 );
buf ( n392925 , n392924 );
nand ( n45474 , n45468 , n392925 );
buf ( n392927 , n45474 );
not ( n45476 , n392927 );
not ( n45477 , n40858 );
or ( n45478 , n45476 , n45477 );
nand ( n45479 , n392103 , n392111 );
nand ( n45480 , n45478 , n45479 );
buf ( n392933 , n45480 );
not ( n45482 , n392933 );
buf ( n392935 , n45482 );
buf ( n392936 , n392935 );
not ( n45485 , n392936 );
or ( n45486 , n45463 , n45485 );
buf ( n392939 , n388463 );
buf ( n392940 , n40977 );
not ( n45489 , n392940 );
buf ( n392942 , n388569 );
not ( n45491 , n392942 );
and ( n45492 , n45489 , n45491 );
buf ( n392945 , n40840 );
buf ( n392946 , n388569 );
and ( n45495 , n392945 , n392946 );
nor ( n45496 , n45492 , n45495 );
buf ( n392949 , n45496 );
buf ( n392950 , n392949 );
or ( n45499 , n392939 , n392950 );
buf ( n392952 , n392077 );
not ( n45501 , n392952 );
buf ( n392954 , n45501 );
buf ( n392955 , n392954 );
buf ( n392956 , n388704 );
or ( n45505 , n392955 , n392956 );
nand ( n45506 , n45499 , n45505 );
buf ( n392959 , n45506 );
buf ( n392960 , n392959 );
nand ( n45509 , n45486 , n392960 );
buf ( n392962 , n45509 );
buf ( n392963 , n392962 );
buf ( n392964 , n44599 );
not ( n45513 , n392964 );
buf ( n392966 , n45480 );
nand ( n45515 , n45513 , n392966 );
buf ( n392968 , n45515 );
buf ( n392969 , n392968 );
nand ( n45518 , n392963 , n392969 );
buf ( n392971 , n45518 );
not ( n45520 , n392971 );
not ( n45521 , n45520 );
nand ( n45522 , n45461 , n45521 );
buf ( n392975 , n392874 );
buf ( n392976 , n392902 );
and ( n45525 , n392975 , n392976 );
buf ( n392978 , n392908 );
nor ( n45527 , n45525 , n392978 );
buf ( n392980 , n45527 );
buf ( n392981 , n392980 );
not ( n45530 , n392981 );
buf ( n392983 , n392812 );
nand ( n45532 , n45530 , n392983 );
buf ( n392985 , n45532 );
nand ( n45534 , n45522 , n392985 );
buf ( n392987 , n45534 );
xor ( n45536 , n392785 , n392987 );
xor ( n45537 , n392051 , n392124 );
xor ( n45538 , n45537 , n392128 );
buf ( n392991 , n45538 );
buf ( n392992 , n392991 );
and ( n45541 , n45536 , n392992 );
and ( n45542 , n392785 , n392987 );
or ( n45543 , n45541 , n45542 );
buf ( n392996 , n45543 );
buf ( n392997 , n392996 );
buf ( n392998 , n392265 );
not ( n45547 , n392998 );
buf ( n393000 , n44812 );
nand ( n45549 , n45547 , n393000 );
buf ( n393002 , n45549 );
xnor ( n45551 , n393002 , n392273 );
buf ( n393004 , n45551 );
xor ( n45553 , n392997 , n393004 );
xor ( n45554 , n392026 , n392133 );
xor ( n45555 , n45554 , n392162 );
buf ( n393008 , n45555 );
buf ( n393009 , n393008 );
and ( n45558 , n45553 , n393009 );
and ( n45559 , n392997 , n393004 );
or ( n45560 , n45558 , n45559 );
buf ( n393013 , n45560 );
buf ( n393014 , n393013 );
and ( n45563 , n45309 , n393014 );
and ( n45564 , n392529 , n392767 );
or ( n45565 , n45563 , n45564 );
buf ( n393018 , n45565 );
buf ( n393019 , n393018 );
nand ( n45568 , n45060 , n393019 );
buf ( n393021 , n45568 );
buf ( n393022 , n393021 );
nand ( n45571 , n45052 , n393022 );
buf ( n393024 , n45571 );
not ( n45573 , n393024 );
or ( n45574 , n45035 , n45573 );
buf ( n393027 , n392493 );
buf ( n393028 , n392488 );
nand ( n45577 , n393027 , n393028 );
buf ( n393030 , n45577 );
nand ( n45579 , n45574 , n393030 );
xnor ( n45580 , n44739 , n45579 );
buf ( n393033 , n45580 );
buf ( n393034 , n392174 );
buf ( n393035 , n392185 );
nand ( n45584 , n393034 , n393035 );
buf ( n393037 , n45584 );
xor ( n45586 , n392191 , n393037 );
not ( n45587 , n44729 );
and ( n45588 , n45586 , n45587 );
not ( n45589 , n45586 );
and ( n45590 , n45589 , n44729 );
nor ( n45591 , n45588 , n45590 );
buf ( n393044 , n45591 );
buf ( n393045 , n44828 );
buf ( n393046 , n392475 );
and ( n45595 , n393045 , n393046 );
not ( n45596 , n393045 );
buf ( n393049 , n392469 );
and ( n45598 , n45596 , n393049 );
nor ( n45599 , n45595 , n45598 );
buf ( n393052 , n45599 );
buf ( n393053 , n45017 );
not ( n45602 , n393053 );
buf ( n393055 , n45602 );
and ( n45604 , n393052 , n393055 );
not ( n45605 , n393052 );
and ( n45606 , n45605 , n45017 );
nor ( n45607 , n45604 , n45606 );
xor ( n45608 , n392004 , n392008 );
xor ( n45609 , n45608 , n392167 );
buf ( n393062 , n45609 );
buf ( n393063 , n393062 );
buf ( n393064 , n392280 );
buf ( n393065 , n392287 );
xor ( n45614 , n393064 , n393065 );
buf ( n393067 , n44825 );
xnor ( n45616 , n45614 , n393067 );
buf ( n393069 , n45616 );
buf ( n393070 , n393069 );
xor ( n45619 , n393063 , n393070 );
buf ( n393072 , n388872 );
not ( n45621 , n393072 );
not ( n45622 , n41342 );
not ( n45623 , n37679 );
or ( n45624 , n45622 , n45623 );
or ( n45625 , n37679 , n41342 );
nand ( n45626 , n45624 , n45625 );
buf ( n393079 , n45626 );
not ( n45628 , n393079 );
or ( n45629 , n45621 , n45628 );
buf ( n393082 , n44744 );
buf ( n393083 , n388833 );
nand ( n45632 , n393082 , n393083 );
buf ( n393085 , n45632 );
buf ( n393086 , n393085 );
nand ( n45635 , n45629 , n393086 );
buf ( n393088 , n45635 );
buf ( n393089 , n393088 );
buf ( n393090 , n384868 );
buf ( n393091 , n23528 );
and ( n45640 , n393090 , n393091 );
not ( n45641 , n393090 );
buf ( n393094 , n37282 );
and ( n45643 , n45641 , n393094 );
nor ( n45644 , n45640 , n45643 );
buf ( n393097 , n45644 );
buf ( n393098 , n393097 );
not ( n45647 , n393098 );
buf ( n393100 , n45647 );
not ( n45649 , n393100 );
not ( n45650 , n44101 );
or ( n45651 , n45649 , n45650 );
nand ( n45652 , n393097 , n384891 );
not ( n45653 , n45652 );
buf ( n393106 , n388897 );
buf ( n393107 , n37305 );
not ( n45656 , n393107 );
buf ( n393109 , n45656 );
buf ( n393110 , n393109 );
nand ( n45659 , n393106 , n393110 );
buf ( n393112 , n45659 );
nand ( n45661 , n45653 , n393112 );
not ( n45662 , n45661 );
buf ( n393115 , n388897 );
not ( n45664 , n393115 );
buf ( n393117 , n45664 );
and ( n45666 , n393117 , n41194 );
not ( n45667 , n393117 );
and ( n45668 , n45667 , n28250 );
or ( n45669 , n45666 , n45668 );
nand ( n45670 , n45662 , n45669 );
nand ( n45671 , n45651 , n45670 );
not ( n45672 , n45671 );
buf ( n393125 , n386474 );
not ( n45674 , n393125 );
buf ( n393127 , n45674 );
not ( n45676 , n393127 );
not ( n45677 , n45106 );
or ( n45678 , n45676 , n45677 );
buf ( n393131 , n22982 );
not ( n45680 , n393131 );
buf ( n393133 , n375781 );
not ( n45682 , n393133 );
buf ( n393135 , n45682 );
buf ( n393136 , n393135 );
not ( n45685 , n393136 );
or ( n45686 , n45680 , n45685 );
buf ( n393139 , n386147 );
buf ( n393140 , n38971 );
nand ( n45689 , n393139 , n393140 );
buf ( n393142 , n45689 );
buf ( n393143 , n393142 );
nand ( n45692 , n45686 , n393143 );
buf ( n393145 , n45692 );
nand ( n45694 , n393145 , n386496 );
nand ( n45695 , n45678 , n45694 );
not ( n45696 , n45695 );
or ( n45697 , n45672 , n45696 );
or ( n45698 , n45695 , n45671 );
not ( n45699 , n27300 );
buf ( n393152 , n45699 );
not ( n45701 , n393152 );
buf ( n393154 , n45701 );
buf ( n393155 , n393154 );
not ( n45704 , n393155 );
buf ( n393157 , n388272 );
not ( n45706 , n393157 );
or ( n45707 , n45704 , n45706 );
not ( n45708 , n27301 );
nand ( n45709 , n45708 , n388263 );
buf ( n393162 , n45709 );
nand ( n45711 , n45707 , n393162 );
buf ( n393164 , n45711 );
not ( n45713 , n393164 );
not ( n45714 , n383891 );
or ( n45715 , n45713 , n45714 );
buf ( n393168 , n388626 );
not ( n45717 , n393168 );
buf ( n393170 , n391593 );
nand ( n45719 , n45717 , n393170 );
buf ( n393172 , n45719 );
nand ( n45721 , n45715 , n393172 );
nand ( n45722 , n45698 , n45721 );
nand ( n45723 , n45697 , n45722 );
not ( n45724 , n45723 );
buf ( n393177 , n389341 );
not ( n45726 , n393177 );
buf ( n393179 , n390453 );
not ( n45728 , n393179 );
or ( n45729 , n45726 , n45728 );
buf ( n393182 , n35435 );
buf ( n393183 , n389341 );
not ( n45732 , n393183 );
buf ( n393185 , n45732 );
buf ( n393186 , n393185 );
nand ( n45735 , n393182 , n393186 );
buf ( n393188 , n45735 );
buf ( n393189 , n393188 );
nand ( n45738 , n45729 , n393189 );
buf ( n393191 , n45738 );
not ( n45740 , n393191 );
not ( n45741 , n390629 );
or ( n45742 , n45740 , n45741 );
nand ( n45743 , n390476 , n392038 );
nand ( n45744 , n45742 , n45743 );
not ( n45745 , n45744 );
or ( n45746 , n45724 , n45745 );
buf ( n393199 , n45723 );
not ( n45748 , n393199 );
buf ( n393201 , n45748 );
buf ( n393202 , n393201 );
not ( n45751 , n393202 );
not ( n45752 , n45744 );
buf ( n393205 , n45752 );
not ( n45754 , n393205 );
or ( n45755 , n45751 , n45754 );
xor ( n45756 , n391560 , n391580 );
xor ( n45757 , n45756 , n391609 );
buf ( n393210 , n45757 );
buf ( n393211 , n393210 );
nand ( n45760 , n45755 , n393211 );
buf ( n393213 , n45760 );
nand ( n45762 , n45746 , n393213 );
buf ( n393215 , n45762 );
xor ( n45764 , n393089 , n393215 );
buf ( n393217 , n43727 );
not ( n45766 , n393217 );
buf ( n393219 , n391027 );
not ( n45768 , n393219 );
buf ( n393221 , n388765 );
not ( n45770 , n393221 );
or ( n45771 , n45768 , n45770 );
buf ( n393224 , n383053 );
buf ( n393225 , n391024 );
nand ( n45774 , n393224 , n393225 );
buf ( n393227 , n45774 );
buf ( n393228 , n393227 );
nand ( n45777 , n45771 , n393228 );
buf ( n393230 , n45777 );
buf ( n393231 , n393230 );
not ( n45780 , n393231 );
or ( n45781 , n45766 , n45780 );
buf ( n393234 , n392154 );
buf ( n393235 , n43515 );
nand ( n45784 , n393234 , n393235 );
buf ( n393237 , n45784 );
buf ( n393238 , n393237 );
nand ( n45787 , n45781 , n393238 );
buf ( n393240 , n45787 );
buf ( n393241 , n393240 );
and ( n45790 , n45764 , n393241 );
and ( n45791 , n393089 , n393215 );
or ( n45792 , n45790 , n45791 );
buf ( n393245 , n45792 );
buf ( n393246 , n393245 );
xor ( n45795 , n392378 , n392433 );
xor ( n45796 , n45795 , n392459 );
buf ( n393249 , n45796 );
buf ( n393250 , n393249 );
xor ( n45799 , n393246 , n393250 );
xor ( n45800 , n392065 , n392090 );
xor ( n45801 , n45800 , n392119 );
buf ( n393254 , n45801 );
not ( n45803 , n393254 );
buf ( n393256 , n388141 );
not ( n45805 , n393256 );
buf ( n393258 , n392392 );
not ( n45807 , n393258 );
or ( n45808 , n45805 , n45807 );
buf ( n393261 , n388160 );
not ( n45810 , n393261 );
buf ( n393263 , n390810 );
not ( n45812 , n393263 );
or ( n45813 , n45810 , n45812 );
buf ( n393266 , n389692 );
buf ( n393267 , n388157 );
nand ( n45816 , n393266 , n393267 );
buf ( n393269 , n45816 );
buf ( n393270 , n393269 );
nand ( n45819 , n45813 , n393270 );
buf ( n393272 , n45819 );
buf ( n393273 , n393272 );
buf ( n393274 , n40701 );
nand ( n45823 , n393273 , n393274 );
buf ( n393276 , n45823 );
buf ( n393277 , n393276 );
nand ( n45826 , n45808 , n393277 );
buf ( n393279 , n45826 );
not ( n45828 , n393279 );
nand ( n45829 , n45803 , n45828 );
not ( n45830 , n45829 );
xor ( n45831 , n392579 , n392604 );
xor ( n45832 , n45831 , n392635 );
buf ( n393285 , n45832 );
not ( n45834 , n393285 );
or ( n45835 , n45830 , n45834 );
nand ( n45836 , n393279 , n393254 );
nand ( n45837 , n45835 , n45836 );
xor ( n45838 , n392427 , n392402 );
xor ( n45839 , n45838 , n392381 );
xor ( n45840 , n45837 , n45839 );
not ( n45841 , n43286 );
buf ( n393294 , n388102 );
not ( n45843 , n393294 );
buf ( n393296 , n42616 );
not ( n45845 , n393296 );
or ( n45846 , n45843 , n45845 );
buf ( n393299 , n35301 );
buf ( n393300 , n388105 );
nand ( n45849 , n393299 , n393300 );
buf ( n393302 , n45849 );
buf ( n393303 , n393302 );
nand ( n45852 , n45846 , n393303 );
buf ( n393305 , n45852 );
not ( n45854 , n393305 );
or ( n45855 , n45841 , n45854 );
buf ( n393308 , n392310 );
buf ( n393309 , n390362 );
nand ( n45858 , n393308 , n393309 );
buf ( n393311 , n45858 );
nand ( n45860 , n45855 , n393311 );
and ( n45861 , n45840 , n45860 );
and ( n45862 , n45837 , n45839 );
or ( n45863 , n45861 , n45862 );
buf ( n393316 , n45863 );
and ( n45865 , n45799 , n393316 );
and ( n45866 , n393246 , n393250 );
or ( n45867 , n45865 , n45866 );
buf ( n393320 , n45867 );
buf ( n393321 , n393320 );
and ( n45870 , n45619 , n393321 );
and ( n45871 , n393063 , n393070 );
or ( n45872 , n45870 , n45871 );
buf ( n393325 , n45872 );
buf ( n393326 , n393325 );
not ( n45875 , n393326 );
buf ( n393328 , n45875 );
nand ( n45877 , n45607 , n393328 );
not ( n45878 , n45877 );
xor ( n45879 , n392529 , n392767 );
xor ( n45880 , n45879 , n393014 );
buf ( n393333 , n45880 );
not ( n45882 , n393333 );
xor ( n45883 , n392350 , n392318 );
xnor ( n45884 , n45883 , n44893 );
buf ( n393337 , n45884 );
buf ( n393338 , n388833 );
not ( n45887 , n393338 );
buf ( n393340 , n45626 );
not ( n45889 , n393340 );
or ( n45890 , n45887 , n45889 );
buf ( n393343 , n41342 );
not ( n45892 , n393343 );
not ( n45893 , n36216 );
buf ( n393346 , n45893 );
not ( n45895 , n393346 );
or ( n45896 , n45892 , n45895 );
buf ( n45897 , n41341 );
buf ( n393350 , n45897 );
buf ( n393351 , n36216 );
nand ( n45900 , n393350 , n393351 );
buf ( n393353 , n45900 );
buf ( n393354 , n393353 );
nand ( n45903 , n45896 , n393354 );
buf ( n393356 , n45903 );
buf ( n393357 , n393356 );
buf ( n393358 , n388872 );
nand ( n45907 , n393357 , n393358 );
buf ( n393360 , n45907 );
buf ( n393361 , n393360 );
nand ( n45910 , n45890 , n393361 );
buf ( n393363 , n45910 );
not ( n45912 , n393363 );
buf ( n393365 , n45912 );
not ( n45914 , n393365 );
buf ( n393367 , n392217 );
buf ( n45916 , n393367 );
buf ( n393369 , n45916 );
buf ( n393370 , n393369 );
not ( n45919 , n393370 );
buf ( n393372 , n34858 );
not ( n45921 , n393372 );
buf ( n393374 , n45921 );
buf ( n393375 , n393374 );
not ( n45924 , n393375 );
or ( n45925 , n45919 , n45924 );
buf ( n393378 , n34858 );
buf ( n393379 , n393369 );
not ( n45928 , n393379 );
buf ( n393381 , n45928 );
buf ( n393382 , n393381 );
buf ( n45931 , n393382 );
buf ( n393384 , n45931 );
buf ( n393385 , n393384 );
nand ( n45934 , n393378 , n393385 );
buf ( n393387 , n45934 );
buf ( n393388 , n393387 );
nand ( n45937 , n45925 , n393388 );
buf ( n393390 , n45937 );
buf ( n393391 , n393390 );
xor ( n45940 , n371244 , n371925 );
and ( n45941 , n371244 , n23604 );
not ( n45942 , n371244 );
buf ( n393395 , n23604 );
not ( n45944 , n393395 );
buf ( n393397 , n45944 );
and ( n45946 , n45942 , n393397 );
or ( n45947 , n45941 , n45946 );
nand ( n45948 , n45940 , n45947 );
not ( n45949 , n45948 );
buf ( n393402 , n45949 );
not ( n45951 , n393402 );
buf ( n393404 , n45951 );
buf ( n393405 , n393404 );
not ( n45954 , n45947 );
buf ( n393407 , n45954 );
not ( n45956 , n393407 );
buf ( n393409 , n45956 );
buf ( n393410 , n393409 );
nand ( n45959 , n393405 , n393410 );
buf ( n393412 , n45959 );
buf ( n393413 , n393412 );
nand ( n45962 , n393391 , n393413 );
buf ( n393415 , n45962 );
buf ( n393416 , n393415 );
not ( n45965 , n393416 );
buf ( n393418 , n45965 );
buf ( n393419 , n393418 );
not ( n45968 , n393419 );
or ( n45969 , n45914 , n45968 );
buf ( n393422 , n392740 );
not ( n45971 , n393422 );
buf ( n393424 , n392733 );
not ( n45973 , n393424 );
or ( n45974 , n45971 , n45973 );
buf ( n393427 , n392247 );
not ( n45976 , n393427 );
buf ( n393429 , n392144 );
not ( n45978 , n393429 );
or ( n45979 , n45976 , n45978 );
buf ( n393432 , n35519 );
buf ( n393433 , n392244 );
nand ( n45982 , n393432 , n393433 );
buf ( n393435 , n45982 );
buf ( n393436 , n393435 );
nand ( n45985 , n45979 , n393436 );
buf ( n393438 , n45985 );
buf ( n393439 , n393438 );
buf ( n393440 , n45260 );
nand ( n45989 , n393439 , n393440 );
buf ( n393442 , n45989 );
buf ( n393443 , n393442 );
nand ( n45992 , n45974 , n393443 );
buf ( n393445 , n45992 );
buf ( n393446 , n393445 );
nand ( n45995 , n45969 , n393446 );
buf ( n393448 , n45995 );
buf ( n393449 , n393448 );
buf ( n393450 , n393415 );
buf ( n393451 , n393363 );
nand ( n46000 , n393450 , n393451 );
buf ( n393453 , n46000 );
buf ( n393454 , n393453 );
nand ( n46003 , n393449 , n393454 );
buf ( n393456 , n46003 );
buf ( n393457 , n393456 );
not ( n46006 , n393457 );
buf ( n393459 , n392639 );
buf ( n393460 , n45078 );
xor ( n46009 , n393459 , n393460 );
buf ( n393462 , n392553 );
xnor ( n46011 , n46009 , n393462 );
buf ( n393464 , n46011 );
buf ( n393465 , n393464 );
not ( n46014 , n393465 );
buf ( n393467 , n46014 );
buf ( n393468 , n393467 );
not ( n46017 , n393468 );
or ( n46018 , n46006 , n46017 );
buf ( n393471 , n393456 );
not ( n46020 , n393471 );
buf ( n393473 , n46020 );
not ( n46022 , n393473 );
not ( n46023 , n393464 );
or ( n46024 , n46022 , n46023 );
not ( n46025 , n389162 );
not ( n46026 , n45075 );
or ( n46027 , n46025 , n46026 );
and ( n46028 , n37173 , n41678 );
not ( n46029 , n37173 );
and ( n46030 , n46029 , n41671 );
or ( n46031 , n46028 , n46030 );
buf ( n393484 , n46031 );
buf ( n393485 , n41711 );
nand ( n46034 , n393484 , n393485 );
buf ( n393487 , n46034 );
nand ( n46036 , n46027 , n393487 );
buf ( n393489 , n385473 );
not ( n46038 , n393489 );
not ( n46039 , n375838 );
not ( n46040 , n375845 );
or ( n46041 , n46039 , n46040 );
nand ( n46042 , n46041 , n375851 );
not ( n46043 , n46042 );
buf ( n393496 , n46043 );
not ( n46045 , n393496 );
or ( n46046 , n46038 , n46045 );
buf ( n393499 , n28250 );
buf ( n393500 , n388965 );
nand ( n46049 , n393499 , n393500 );
buf ( n393502 , n46049 );
buf ( n393503 , n393502 );
nand ( n46052 , n46046 , n393503 );
buf ( n393505 , n46052 );
buf ( n393506 , n393505 );
not ( n46055 , n393506 );
and ( n46056 , n37922 , n37930 , n37931 );
buf ( n393509 , n46056 );
not ( n46058 , n393509 );
or ( n46059 , n46055 , n46058 );
not ( n46060 , n37922 );
not ( n46061 , n46060 );
buf ( n46062 , n46061 );
buf ( n393515 , n46062 );
not ( n46064 , n393515 );
buf ( n393517 , n385473 );
not ( n46066 , n393517 );
buf ( n393519 , n388445 );
not ( n46068 , n393519 );
or ( n46069 , n46066 , n46068 );
buf ( n393522 , n40817 );
buf ( n393523 , n385473 );
not ( n46072 , n393523 );
buf ( n393525 , n46072 );
buf ( n393526 , n393525 );
nand ( n46075 , n393522 , n393526 );
buf ( n393528 , n46075 );
buf ( n393529 , n393528 );
nand ( n46078 , n46069 , n393529 );
buf ( n393531 , n46078 );
buf ( n393532 , n393531 );
nand ( n46081 , n46064 , n393532 );
buf ( n393534 , n46081 );
buf ( n393535 , n393534 );
nand ( n46084 , n46059 , n393535 );
buf ( n393537 , n46084 );
buf ( n393538 , n393537 );
not ( n46087 , n44594 );
not ( n46088 , n41447 );
or ( n46089 , n46087 , n46088 );
buf ( n393542 , n44077 );
not ( n46091 , n393542 );
buf ( n393544 , n46091 );
buf ( n393545 , n393544 );
buf ( n393546 , n393531 );
nand ( n46095 , n393545 , n393546 );
buf ( n393548 , n46095 );
nand ( n46097 , n46089 , n393548 );
buf ( n393550 , n46097 );
xor ( n46099 , n393538 , n393550 );
not ( n46100 , n45669 );
not ( n46101 , n37314 );
or ( n46102 , n46100 , n46101 );
buf ( n393555 , n388367 );
not ( n46104 , n393555 );
buf ( n393557 , n46104 );
buf ( n393558 , n393557 );
not ( n46107 , n393558 );
buf ( n393560 , n37345 );
not ( n46109 , n393560 );
buf ( n393562 , n46109 );
buf ( n393563 , n393562 );
nor ( n46112 , n46107 , n393563 );
buf ( n393565 , n46112 );
not ( n46114 , n28270 );
and ( n46115 , n393117 , n46114 );
nor ( n46116 , n393565 , n46115 );
or ( n46117 , n46116 , n43058 );
nand ( n46118 , n46102 , n46117 );
buf ( n393571 , n46118 );
and ( n46120 , n46099 , n393571 );
and ( n46121 , n393538 , n393550 );
or ( n46122 , n46120 , n46121 );
buf ( n393575 , n46122 );
buf ( n393576 , n388998 );
not ( n46125 , n393576 );
buf ( n393578 , n42390 );
not ( n46127 , n393578 );
or ( n46128 , n46125 , n46127 );
buf ( n393581 , n391870 );
buf ( n393582 , n388215 );
nand ( n46131 , n393581 , n393582 );
buf ( n393584 , n46131 );
buf ( n393585 , n393584 );
nand ( n46134 , n46128 , n393585 );
buf ( n393587 , n46134 );
buf ( n393588 , n393587 );
not ( n46137 , n393588 );
buf ( n393590 , n389880 );
not ( n46139 , n393590 );
buf ( n393592 , n46139 );
buf ( n393593 , n393592 );
not ( n46142 , n393593 );
buf ( n393595 , n46142 );
buf ( n393596 , n393595 );
not ( n46145 , n393596 );
or ( n46146 , n46137 , n46145 );
buf ( n393599 , n392654 );
buf ( n393600 , n391635 );
not ( n46149 , n393600 );
buf ( n393602 , n46149 );
buf ( n393603 , n393602 );
nand ( n46152 , n393599 , n393603 );
buf ( n393605 , n46152 );
buf ( n393606 , n393605 );
nand ( n46155 , n46146 , n393606 );
buf ( n393608 , n46155 );
xor ( n46157 , n393575 , n393608 );
not ( n46158 , n391080 );
buf ( n393611 , n24074 );
not ( n46160 , n393611 );
not ( n46161 , n36564 );
buf ( n393614 , n46161 );
not ( n46163 , n393614 );
or ( n46164 , n46160 , n46163 );
buf ( n393617 , n38155 );
buf ( n393618 , n24073 );
nand ( n46167 , n393617 , n393618 );
buf ( n393620 , n46167 );
buf ( n393621 , n393620 );
nand ( n46170 , n46164 , n393621 );
buf ( n393623 , n46170 );
not ( n46172 , n393623 );
or ( n46173 , n46158 , n46172 );
nand ( n46174 , n390403 , n392805 );
nand ( n46175 , n46173 , n46174 );
and ( n46176 , n46157 , n46175 );
and ( n46177 , n393575 , n393608 );
or ( n46178 , n46176 , n46177 );
xor ( n46179 , n46036 , n46178 );
buf ( n393632 , n392703 );
buf ( n393633 , n392672 );
not ( n46182 , n393633 );
buf ( n393635 , n45225 );
not ( n46184 , n393635 );
or ( n46185 , n46182 , n46184 );
buf ( n393638 , n392710 );
buf ( n393639 , n392675 );
nand ( n46188 , n393638 , n393639 );
buf ( n393641 , n46188 );
buf ( n393642 , n393641 );
nand ( n46191 , n46185 , n393642 );
buf ( n393644 , n46191 );
buf ( n393645 , n393644 );
xor ( n46194 , n393632 , n393645 );
buf ( n393647 , n46194 );
and ( n46196 , n46179 , n393647 );
and ( n46197 , n46036 , n46178 );
or ( n46198 , n46196 , n46197 );
buf ( n46199 , n46198 );
nand ( n46200 , n46024 , n46199 );
buf ( n393653 , n46200 );
nand ( n46202 , n46018 , n393653 );
buf ( n393655 , n46202 );
buf ( n393656 , n393655 );
xor ( n46205 , n393337 , n393656 );
xor ( n46206 , n392642 , n392757 );
xor ( n46207 , n46206 , n392762 );
buf ( n393660 , n46207 );
buf ( n393661 , n393660 );
and ( n46210 , n46205 , n393661 );
and ( n46211 , n393337 , n393656 );
or ( n46212 , n46210 , n46211 );
buf ( n393665 , n46212 );
buf ( n393666 , n393665 );
not ( n46215 , n393666 );
buf ( n393668 , n46215 );
buf ( n393669 , n393668 );
and ( n46218 , n392463 , n392364 );
not ( n46219 , n392463 );
buf ( n393672 , n392364 );
not ( n46221 , n393672 );
buf ( n393674 , n46221 );
and ( n46223 , n46219 , n393674 );
or ( n46224 , n46218 , n46223 );
buf ( n46225 , n44903 );
xor ( n46226 , n46224 , n46225 );
buf ( n393679 , n46226 );
nand ( n46228 , n393669 , n393679 );
buf ( n393681 , n46228 );
not ( n46230 , n393681 );
or ( n46231 , n45882 , n46230 );
buf ( n393684 , n393665 );
buf ( n393685 , n46226 );
not ( n46234 , n393685 );
buf ( n393687 , n46234 );
buf ( n393688 , n393687 );
nand ( n46237 , n393684 , n393688 );
buf ( n393690 , n46237 );
nand ( n46239 , n46231 , n393690 );
not ( n46240 , n46239 );
or ( n46241 , n45878 , n46240 );
not ( n46242 , n45607 );
nand ( n46243 , n46242 , n393325 );
nand ( n46244 , n46241 , n46243 );
buf ( n393697 , n46244 );
not ( n46246 , n393697 );
buf ( n393699 , n46246 );
buf ( n393700 , n393699 );
xor ( n46249 , n393044 , n393700 );
buf ( n393702 , n392488 );
buf ( n393703 , n392496 );
and ( n46252 , n393702 , n393703 );
not ( n46253 , n393702 );
buf ( n393706 , n392493 );
and ( n46255 , n46253 , n393706 );
nor ( n46256 , n46252 , n46255 );
buf ( n393709 , n46256 );
xor ( n46258 , n393709 , n393024 );
buf ( n393711 , n46258 );
and ( n46260 , n46249 , n393711 );
and ( n46261 , n393044 , n393700 );
or ( n46262 , n46260 , n46261 );
buf ( n393715 , n46262 );
buf ( n393716 , n393715 );
nand ( n46265 , n393033 , n393716 );
buf ( n393718 , n46265 );
buf ( n393719 , n393718 );
xor ( n46268 , n393044 , n393700 );
xor ( n46269 , n46268 , n393711 );
buf ( n393722 , n46269 );
buf ( n393723 , n393722 );
buf ( n393724 , n392503 );
buf ( n393725 , n393018 );
xor ( n46274 , n393724 , n393725 );
buf ( n393727 , n392514 );
xnor ( n46276 , n46274 , n393727 );
buf ( n393729 , n46276 );
xor ( n46278 , n393246 , n393250 );
xor ( n46279 , n46278 , n393316 );
buf ( n393732 , n46279 );
buf ( n393733 , n393732 );
not ( n46282 , n393733 );
xor ( n46283 , n393337 , n393656 );
xor ( n46284 , n46283 , n393661 );
buf ( n393737 , n46284 );
buf ( n393738 , n393737 );
not ( n46287 , n393738 );
or ( n46288 , n46282 , n46287 );
buf ( n393741 , n393737 );
buf ( n393742 , n393732 );
or ( n46291 , n393741 , n393742 );
xor ( n46292 , n45837 , n45839 );
xor ( n46293 , n46292 , n45860 );
buf ( n393746 , n46293 );
not ( n46295 , n393746 );
xor ( n46296 , n393456 , n46198 );
xnor ( n46297 , n46296 , n393464 );
buf ( n393750 , n46297 );
not ( n46299 , n393750 );
or ( n46300 , n46295 , n46299 );
not ( n46301 , n46293 );
not ( n393754 , n46301 );
or ( n46303 , n393754 , n46297 );
xor ( n46304 , n46036 , n46178 );
xor ( n46305 , n46304 , n393647 );
not ( n46306 , n46305 );
buf ( n393759 , n392902 );
buf ( n393760 , n392845 );
buf ( n393761 , n392868 );
and ( n46310 , n393760 , n393761 );
not ( n46311 , n393760 );
buf ( n393764 , n392871 );
and ( n46313 , n46311 , n393764 );
nor ( n46314 , n46310 , n46313 );
buf ( n393767 , n46314 );
buf ( n393768 , n393767 );
xor ( n46317 , n393759 , n393768 );
buf ( n393770 , n46317 );
buf ( n393771 , n393770 );
buf ( n393772 , n44599 );
buf ( n393773 , n45480 );
xor ( n46322 , n393772 , n393773 );
buf ( n393775 , n392959 );
xnor ( n46324 , n46322 , n393775 );
buf ( n393777 , n46324 );
buf ( n393778 , n393777 );
xor ( n46327 , n393771 , n393778 );
buf ( n393780 , n388833 );
not ( n46329 , n393780 );
buf ( n393782 , n393356 );
not ( n46331 , n393782 );
or ( n46332 , n46329 , n46331 );
buf ( n393785 , n41342 );
not ( n46334 , n393785 );
buf ( n393787 , n389067 );
not ( n46336 , n393787 );
or ( n46337 , n46334 , n46336 );
buf ( n393790 , n384177 );
buf ( n393791 , n45897 );
nand ( n46340 , n393790 , n393791 );
buf ( n393793 , n46340 );
buf ( n393794 , n393793 );
nand ( n46343 , n46337 , n393794 );
buf ( n393796 , n46343 );
buf ( n393797 , n393796 );
buf ( n393798 , n388872 );
nand ( n46347 , n393797 , n393798 );
buf ( n393800 , n46347 );
buf ( n393801 , n393800 );
nand ( n46350 , n46332 , n393801 );
buf ( n393803 , n46350 );
buf ( n393804 , n393803 );
and ( n46353 , n46327 , n393804 );
and ( n46354 , n393771 , n393778 );
or ( n46355 , n46353 , n46354 );
buf ( n393808 , n46355 );
not ( n46357 , n393808 );
or ( n46358 , n46306 , n46357 );
or ( n46359 , n46305 , n393808 );
not ( n46360 , n41671 );
not ( n46361 , n37680 );
not ( n46362 , n46361 );
or ( n46363 , n46360 , n46362 );
nand ( n46364 , n41678 , n37680 );
nand ( n46365 , n46363 , n46364 );
and ( n46366 , n46365 , n41711 );
and ( n46367 , n46031 , n389162 );
nor ( n46368 , n46366 , n46367 );
not ( n46369 , n46368 );
not ( n46370 , n46369 );
buf ( n393823 , n393404 );
not ( n46372 , n393823 );
buf ( n393825 , n46372 );
buf ( n393826 , n393825 );
not ( n46375 , n393826 );
buf ( n393828 , n393369 );
not ( n46377 , n393828 );
buf ( n393830 , n382526 );
not ( n46379 , n393830 );
or ( n46380 , n46377 , n46379 );
buf ( n393833 , n390345 );
buf ( n393834 , n393384 );
nand ( n46383 , n393833 , n393834 );
buf ( n393836 , n46383 );
buf ( n393837 , n393836 );
nand ( n46386 , n46380 , n393837 );
buf ( n393839 , n46386 );
buf ( n393840 , n393839 );
not ( n46389 , n393840 );
or ( n46390 , n46375 , n46389 );
buf ( n393843 , n393390 );
buf ( n393844 , n45954 );
nand ( n46393 , n393843 , n393844 );
buf ( n393846 , n46393 );
buf ( n393847 , n393846 );
nand ( n46396 , n46390 , n393847 );
buf ( n393849 , n46396 );
not ( n46398 , n393849 );
or ( n46399 , n46370 , n46398 );
or ( n46400 , n393849 , n46369 );
xor ( n46401 , n393575 , n393608 );
xor ( n46402 , n46401 , n46175 );
buf ( n46403 , n46402 );
nand ( n46404 , n46400 , n46403 );
nand ( n46405 , n46399 , n46404 );
nand ( n46406 , n46359 , n46405 );
nand ( n46407 , n46358 , n46406 );
buf ( n46408 , n46407 );
nand ( n46409 , n46303 , n46408 );
buf ( n393862 , n46409 );
nand ( n46411 , n46300 , n393862 );
buf ( n393864 , n46411 );
buf ( n393865 , n393864 );
nand ( n46414 , n46291 , n393865 );
buf ( n393867 , n46414 );
buf ( n393868 , n393867 );
nand ( n46417 , n46288 , n393868 );
buf ( n393870 , n46417 );
not ( n46419 , n393870 );
xor ( n46420 , n393063 , n393070 );
xor ( n46421 , n46420 , n393321 );
buf ( n393874 , n46421 );
buf ( n393875 , n393874 );
not ( n46424 , n393875 );
buf ( n393877 , n46424 );
buf ( n393878 , n393877 );
xor ( n46427 , n393089 , n393215 );
xor ( n46428 , n46427 , n393241 );
buf ( n393881 , n46428 );
buf ( n393882 , n393881 );
buf ( n393883 , n40990 );
buf ( n393884 , n383420 );
and ( n46433 , n393883 , n393884 );
not ( n46434 , n393883 );
buf ( n393887 , n388556 );
and ( n46436 , n46434 , n393887 );
nor ( n46437 , n46433 , n46436 );
buf ( n393890 , n46437 );
buf ( n393891 , n393890 );
not ( n46440 , n393891 );
buf ( n393893 , n46440 );
buf ( n393894 , n393893 );
not ( n46443 , n393894 );
buf ( n393896 , n391270 );
not ( n46445 , n393896 );
or ( n46446 , n46443 , n46445 );
buf ( n393899 , n392696 );
not ( n46448 , n393899 );
buf ( n393901 , n383403 );
not ( n46450 , n393901 );
buf ( n393903 , n46450 );
buf ( n393904 , n393903 );
nand ( n46453 , n46448 , n393904 );
buf ( n393906 , n46453 );
buf ( n393907 , n393906 );
nand ( n46456 , n46446 , n393907 );
buf ( n393909 , n46456 );
buf ( n393910 , n393909 );
xor ( n46459 , n45671 , n45695 );
and ( n46460 , n46459 , n45721 );
not ( n46461 , n46459 );
not ( n46462 , n45721 );
and ( n46463 , n46461 , n46462 );
nor ( n46464 , n46460 , n46463 );
buf ( n393917 , n46464 );
or ( n46466 , n393910 , n393917 );
buf ( n393919 , n46466 );
buf ( n393920 , n393919 );
buf ( n393921 , n388272 );
not ( n46470 , n393921 );
buf ( n393923 , n46470 );
not ( n46472 , n393923 );
not ( n46473 , n28289 );
nand ( n46474 , n46473 , n28284 );
not ( n46475 , n28284 );
nand ( n46476 , n46475 , n28289 );
nand ( n46477 , n46474 , n46476 );
not ( n46478 , n46477 );
not ( n46479 , n46478 );
or ( n46480 , n46472 , n46479 );
buf ( n46481 , n28297 );
nand ( n46482 , n46481 , n36251 );
nand ( n46483 , n46480 , n46482 );
buf ( n393936 , n46483 );
not ( n46485 , n393936 );
buf ( n393938 , n36317 );
not ( n46487 , n393938 );
or ( n46488 , n46485 , n46487 );
buf ( n393941 , n393164 );
buf ( n393942 , n383904 );
nand ( n46491 , n393941 , n393942 );
buf ( n393944 , n46491 );
buf ( n393945 , n393944 );
nand ( n46494 , n46488 , n393945 );
buf ( n393947 , n46494 );
buf ( n393948 , n393947 );
not ( n46497 , n393948 );
buf ( n393950 , n46497 );
not ( n46499 , n393950 );
buf ( n393952 , n386477 );
not ( n46501 , n393952 );
buf ( n393954 , n393145 );
not ( n46503 , n393954 );
or ( n46504 , n46501 , n46503 );
buf ( n393957 , n27611 );
not ( n46506 , n393957 );
buf ( n393959 , n38971 );
not ( n46508 , n393959 );
and ( n46509 , n46506 , n46508 );
buf ( n393962 , n40778 );
not ( n46511 , n22982 );
buf ( n393964 , n46511 );
and ( n46513 , n393962 , n393964 );
nor ( n46514 , n46509 , n46513 );
buf ( n393967 , n46514 );
buf ( n393968 , n393967 );
not ( n46517 , n393968 );
buf ( n393970 , n386496 );
nand ( n46519 , n46517 , n393970 );
buf ( n393972 , n46519 );
buf ( n393973 , n393972 );
nand ( n46522 , n46504 , n393973 );
buf ( n393975 , n46522 );
buf ( n393976 , n393975 );
buf ( n46525 , n393976 );
buf ( n393978 , n46525 );
nor ( n46527 , n46499 , n393978 );
not ( n46528 , n36422 );
not ( n46529 , n36425 );
or ( n46530 , n46528 , n46529 );
nand ( n46531 , n46530 , n36428 );
nand ( n46532 , n46531 , n384003 );
buf ( n393985 , n46532 );
not ( n46534 , n393985 );
buf ( n393987 , n388546 );
buf ( n393988 , n40977 );
and ( n46537 , n393987 , n393988 );
not ( n46538 , n393987 );
buf ( n393991 , n40973 );
and ( n46540 , n46538 , n393991 );
nor ( n46541 , n46537 , n46540 );
buf ( n393994 , n46541 );
buf ( n393995 , n393994 );
not ( n46544 , n393995 );
and ( n46545 , n46534 , n46544 );
buf ( n393998 , n392949 );
buf ( n393999 , n383937 );
nor ( n46548 , n393998 , n393999 );
buf ( n394001 , n46548 );
buf ( n394002 , n394001 );
nor ( n46551 , n46545 , n394002 );
buf ( n394004 , n46551 );
or ( n46553 , n46527 , n394004 );
buf ( n394006 , n393947 );
buf ( n394007 , n393978 );
nand ( n46556 , n394006 , n394007 );
buf ( n394009 , n46556 );
nand ( n46558 , n46553 , n394009 );
buf ( n394011 , n46558 );
and ( n46560 , n393920 , n394011 );
buf ( n394013 , n46464 );
buf ( n394014 , n393909 );
and ( n46563 , n394013 , n394014 );
buf ( n394016 , n46563 );
buf ( n394017 , n394016 );
nor ( n46566 , n46560 , n394017 );
buf ( n394019 , n46566 );
buf ( n394020 , n394019 );
not ( n46569 , n394020 );
buf ( n394022 , n388809 );
not ( n46571 , n394022 );
buf ( n394024 , n45315 );
not ( n46573 , n394024 );
or ( n46574 , n46571 , n46573 );
buf ( n394027 , n388760 );
not ( n46576 , n394027 );
buf ( n394029 , n389420 );
not ( n46578 , n394029 );
or ( n46579 , n46576 , n46578 );
buf ( n394032 , n38227 );
buf ( n394033 , n388757 );
nand ( n46582 , n394032 , n394033 );
buf ( n394035 , n46582 );
buf ( n394036 , n394035 );
nand ( n46585 , n46579 , n394036 );
buf ( n394038 , n46585 );
buf ( n394039 , n394038 );
buf ( n394040 , n388746 );
nand ( n46589 , n394039 , n394040 );
buf ( n394042 , n46589 );
buf ( n394043 , n394042 );
nand ( n46592 , n46574 , n394043 );
buf ( n394045 , n46592 );
buf ( n394046 , n394045 );
not ( n46595 , n394046 );
buf ( n394048 , n46595 );
buf ( n394049 , n394048 );
not ( n46598 , n394049 );
or ( n46599 , n46569 , n46598 );
not ( n46600 , n45744 );
not ( n46601 , n45723 );
or ( n46602 , n46600 , n46601 );
nand ( n46603 , n393201 , n45752 );
nand ( n46604 , n46602 , n46603 );
not ( n46605 , n393210 );
and ( n46606 , n46604 , n46605 );
not ( n46607 , n46604 );
and ( n46608 , n46607 , n393210 );
nor ( n46609 , n46606 , n46608 );
buf ( n394062 , n46609 );
nand ( n46611 , n46599 , n394062 );
buf ( n394064 , n46611 );
buf ( n394065 , n394064 );
buf ( n394066 , n394019 );
not ( n46615 , n394066 );
buf ( n394068 , n394045 );
nand ( n46617 , n46615 , n394068 );
buf ( n394070 , n46617 );
buf ( n394071 , n394070 );
nand ( n46620 , n394065 , n394071 );
buf ( n394073 , n46620 );
buf ( n394074 , n394073 );
xor ( n46623 , n393882 , n394074 );
xor ( n46624 , n392718 , n392747 );
xor ( n46625 , n46624 , n392752 );
buf ( n394078 , n46625 );
buf ( n394079 , n394078 );
and ( n46628 , n46623 , n394079 );
and ( n46629 , n393882 , n394074 );
or ( n46630 , n46628 , n46629 );
buf ( n394083 , n46630 );
not ( n46632 , n394083 );
xor ( n46633 , n392997 , n393004 );
xor ( n46634 , n46633 , n393009 );
buf ( n394087 , n46634 );
not ( n46636 , n394087 );
xor ( n46637 , n392785 , n392987 );
xor ( n46638 , n46637 , n392992 );
buf ( n394091 , n46638 );
buf ( n394092 , n394091 );
buf ( n394093 , n391446 );
not ( n46642 , n394093 );
buf ( n394095 , n40714 );
not ( n46644 , n394095 );
or ( n46645 , n46642 , n46644 );
buf ( n394098 , n38685 );
not ( n46647 , n394098 );
buf ( n394100 , n391455 );
nand ( n46649 , n46647 , n394100 );
buf ( n394102 , n46649 );
buf ( n394103 , n394102 );
nand ( n46652 , n46645 , n394103 );
buf ( n394105 , n46652 );
not ( n46654 , n394105 );
not ( n46655 , n38765 );
or ( n46656 , n46654 , n46655 );
buf ( n394109 , n390476 );
buf ( n394110 , n393191 );
nand ( n46659 , n394109 , n394110 );
buf ( n394112 , n46659 );
nand ( n46661 , n46656 , n394112 );
buf ( n394114 , n46661 );
buf ( n394115 , n40701 );
not ( n46664 , n394115 );
buf ( n394117 , n388154 );
buf ( n394118 , n37411 );
not ( n46667 , n394118 );
buf ( n394120 , n46667 );
buf ( n394121 , n394120 );
and ( n46670 , n394117 , n394121 );
not ( n46671 , n394117 );
buf ( n394124 , n44945 );
and ( n46673 , n46671 , n394124 );
nor ( n46674 , n46670 , n46673 );
buf ( n394127 , n46674 );
buf ( n394128 , n394127 );
not ( n46677 , n394128 );
or ( n46678 , n46664 , n46677 );
buf ( n394131 , n393272 );
buf ( n394132 , n40640 );
not ( n46681 , n394132 );
buf ( n394134 , n46681 );
buf ( n394135 , n394134 );
nand ( n46684 , n394131 , n394135 );
buf ( n394137 , n46684 );
buf ( n394138 , n394137 );
nand ( n46687 , n46678 , n394138 );
buf ( n394140 , n46687 );
buf ( n394141 , n394140 );
xor ( n46690 , n394114 , n394141 );
buf ( n394143 , n41565 );
not ( n46692 , n394143 );
buf ( n394145 , n392858 );
not ( n46694 , n394145 );
or ( n46695 , n46692 , n46694 );
not ( n46696 , n24049 );
and ( n46697 , n28153 , n46696 );
not ( n46698 , n28153 );
not ( n46699 , n45391 );
and ( n46700 , n46698 , n46699 );
or ( n46701 , n46697 , n46700 );
and ( n46702 , n27908 , n46701 );
not ( n46703 , n27908 );
not ( n46704 , n24049 );
and ( n46705 , n28156 , n46704 );
not ( n46706 , n28156 );
not ( n46707 , n45391 );
and ( n46708 , n46706 , n46707 );
or ( n46709 , n46705 , n46708 );
and ( n46710 , n46703 , n46709 );
or ( n46711 , n46702 , n46710 );
buf ( n394164 , n46711 );
not ( n46713 , n394164 );
buf ( n394166 , n389125 );
nand ( n46715 , n46713 , n394166 );
buf ( n394168 , n46715 );
buf ( n394169 , n394168 );
nand ( n46718 , n46695 , n394169 );
buf ( n394171 , n46718 );
buf ( n394172 , n394171 );
not ( n46721 , n394172 );
buf ( n394174 , n388230 );
not ( n46723 , n394174 );
buf ( n394176 , n40886 );
not ( n46725 , n394176 );
or ( n46726 , n46723 , n46725 );
buf ( n394179 , n40885 );
buf ( n394180 , n388242 );
nand ( n46729 , n394179 , n394180 );
buf ( n394182 , n46729 );
buf ( n394183 , n394182 );
nand ( n46732 , n46726 , n394183 );
buf ( n394185 , n46732 );
buf ( n394186 , n394185 );
not ( n46735 , n394186 );
buf ( n394188 , n40858 );
not ( n46737 , n394188 );
or ( n46738 , n46735 , n46737 );
buf ( n394191 , n384413 );
buf ( n394192 , n392927 );
nand ( n46741 , n394191 , n394192 );
buf ( n394194 , n46741 );
buf ( n394195 , n394194 );
nand ( n46744 , n46738 , n394195 );
buf ( n394197 , n46744 );
buf ( n394198 , n394197 );
not ( n46747 , n394198 );
buf ( n394200 , n46747 );
buf ( n394201 , n394200 );
nand ( n46750 , n46721 , n394201 );
buf ( n394203 , n46750 );
not ( n46752 , n394203 );
buf ( n394205 , n24828 );
not ( n46754 , n394205 );
buf ( n394207 , n46754 );
buf ( n394208 , n394207 );
not ( n46757 , n394208 );
buf ( n394210 , n46757 );
buf ( n394211 , n394210 );
not ( n46760 , n394211 );
buf ( n394213 , n384143 );
not ( n46762 , n394213 );
or ( n46763 , n46760 , n46762 );
buf ( n394216 , n385328 );
buf ( n394217 , n394210 );
not ( n46766 , n394217 );
buf ( n394219 , n46766 );
buf ( n394220 , n394219 );
nand ( n46769 , n394216 , n394220 );
buf ( n394222 , n46769 );
buf ( n394223 , n394222 );
nand ( n46772 , n46763 , n394223 );
buf ( n394225 , n46772 );
or ( n46781 , n382941 , n392895 );
nand ( n46782 , C1 , n46781 );
not ( n46783 , n46782 );
or ( n46784 , n46752 , n46783 );
buf ( n394230 , n394197 );
buf ( n394231 , n394171 );
nand ( n46787 , n394230 , n394231 );
buf ( n394233 , n46787 );
nand ( n46789 , n46784 , n394233 );
buf ( n394235 , n46789 );
and ( n46791 , n46690 , n394235 );
and ( n46792 , n394114 , n394141 );
or ( n46793 , n46791 , n46792 );
buf ( n394239 , n46793 );
buf ( n394240 , n394239 );
not ( n46796 , n392911 );
not ( n46797 , n46796 );
and ( n46798 , n392812 , n45520 );
not ( n46799 , n392812 );
and ( n46800 , n46799 , n392971 );
nor ( n46801 , n46798 , n46800 );
not ( n46802 , n46801 );
or ( n46803 , n46797 , n46802 );
or ( n46804 , n46801 , n46796 );
nand ( n46805 , n46803 , n46804 );
buf ( n394251 , n46805 );
xor ( n46807 , n394240 , n394251 );
not ( n46808 , n393279 );
not ( n46809 , n45803 );
or ( n46810 , n46808 , n46809 );
nand ( n46811 , n393254 , n45828 );
nand ( n46812 , n46810 , n46811 );
and ( n46813 , n46812 , n393285 );
not ( n46814 , n46812 );
not ( n46815 , n393285 );
and ( n46816 , n46814 , n46815 );
nor ( n46817 , n46813 , n46816 );
buf ( n394263 , n46817 );
and ( n46819 , n46807 , n394263 );
and ( n46820 , n394240 , n394251 );
or ( n46821 , n46819 , n46820 );
buf ( n394267 , n46821 );
buf ( n394268 , n394267 );
xor ( n46824 , n394092 , n394268 );
buf ( n394270 , n43727 );
not ( n46826 , n394270 );
buf ( n394272 , n391027 );
not ( n46828 , n394272 );
buf ( n394274 , n386561 );
not ( n46830 , n394274 );
or ( n46831 , n46828 , n46830 );
buf ( n394277 , n382921 );
buf ( n394278 , n391024 );
nand ( n46834 , n394277 , n394278 );
buf ( n394280 , n46834 );
buf ( n394281 , n394280 );
nand ( n46837 , n46831 , n394281 );
buf ( n394283 , n46837 );
buf ( n394284 , n394283 );
not ( n46840 , n394284 );
or ( n46841 , n46826 , n46840 );
buf ( n394287 , n393230 );
buf ( n394288 , n43515 );
nand ( n46844 , n394287 , n394288 );
buf ( n394290 , n46844 );
buf ( n394291 , n394290 );
nand ( n46847 , n46841 , n394291 );
buf ( n394293 , n46847 );
buf ( n394294 , n394293 );
buf ( n394295 , n390362 );
not ( n46851 , n394295 );
buf ( n394297 , n393305 );
not ( n46853 , n394297 );
or ( n46854 , n46851 , n46853 );
buf ( n394300 , n388102 );
not ( n46856 , n394300 );
buf ( n394302 , n37027 );
not ( n46858 , n394302 );
or ( n46859 , n46856 , n46858 );
buf ( n394305 , n35997 );
not ( n46861 , n394305 );
buf ( n394307 , n46861 );
buf ( n394308 , n394307 );
not ( n46864 , n394308 );
buf ( n394310 , n388105 );
nand ( n46866 , n46864 , n394310 );
buf ( n394312 , n46866 );
buf ( n394313 , n394312 );
nand ( n46869 , n46859 , n394313 );
buf ( n394315 , n46869 );
buf ( n394316 , n394315 );
buf ( n394317 , n43286 );
nand ( n46873 , n394316 , n394317 );
buf ( n394319 , n46873 );
buf ( n394320 , n394319 );
nand ( n46876 , n46854 , n394320 );
buf ( n394322 , n46876 );
buf ( n394323 , n394322 );
xor ( n46879 , n394294 , n394323 );
not ( n46880 , n46116 );
not ( n46881 , n37313 );
and ( n46882 , n46880 , n46881 );
buf ( n394328 , n393154 );
not ( n46884 , n394328 );
buf ( n394330 , n46884 );
buf ( n394331 , n394330 );
buf ( n394332 , n390548 );
and ( n46888 , n394331 , n394332 );
not ( n46889 , n394331 );
buf ( n394335 , n393117 );
and ( n46891 , n46889 , n394335 );
or ( n46892 , n46888 , n46891 );
buf ( n394338 , n46892 );
not ( n46894 , n394338 );
and ( n46895 , n390536 , n46894 );
nor ( n46896 , n46882 , n46895 );
not ( n46897 , n46896 );
not ( n46898 , n46897 );
or ( n46899 , n393967 , n386474 );
buf ( n394345 , n22982 );
not ( n46901 , n394345 );
buf ( n394347 , n43044 );
not ( n46903 , n394347 );
or ( n46904 , n46901 , n46903 );
buf ( n394350 , n27195 );
not ( n46906 , n22982 );
buf ( n394352 , n46906 );
nand ( n46908 , n394350 , n394352 );
buf ( n394354 , n46908 );
buf ( n394355 , n394354 );
nand ( n46911 , n46904 , n394355 );
buf ( n394357 , n46911 );
nand ( n46913 , n394357 , n38961 );
nand ( n46914 , n46899 , n46913 );
not ( n46915 , n46914 );
or ( n46916 , n46898 , n46915 );
not ( n46917 , n46914 );
not ( n46918 , n46917 );
not ( n46919 , n46896 );
or ( n46920 , n46918 , n46919 );
not ( n46921 , n41562 );
not ( n46922 , n46921 );
not ( n46923 , n46711 );
not ( n46924 , n46923 );
or ( n46925 , n46922 , n46924 );
buf ( n394371 , n24050 );
not ( n46927 , n394371 );
buf ( n394373 , n393135 );
not ( n46929 , n394373 );
or ( n46930 , n46927 , n46929 );
buf ( n394376 , n375781 );
buf ( n394377 , n45391 );
nand ( n46933 , n394376 , n394377 );
buf ( n394379 , n46933 );
buf ( n394380 , n394379 );
nand ( n46936 , n46930 , n394380 );
buf ( n394382 , n46936 );
nand ( n46938 , n394382 , n389122 );
nand ( n46939 , n46925 , n46938 );
nand ( n46940 , n46920 , n46939 );
nand ( n46941 , n46916 , n46940 );
buf ( n394387 , n46941 );
buf ( n394388 , n388502 );
not ( n46944 , n394388 );
buf ( n394390 , n389894 );
not ( n46946 , n394390 );
buf ( n394392 , n46946 );
buf ( n394393 , n394392 );
not ( n46949 , n394393 );
or ( n46950 , n46944 , n46949 );
buf ( n394396 , n391870 );
buf ( n394397 , n388511 );
nand ( n46953 , n394396 , n394397 );
buf ( n394399 , n46953 );
buf ( n394400 , n394399 );
nand ( n46956 , n46950 , n394400 );
buf ( n394402 , n46956 );
buf ( n394403 , n394402 );
not ( n46959 , n394403 );
buf ( n394405 , n389880 );
not ( n46961 , n394405 );
or ( n46962 , n46959 , n46961 );
buf ( n394408 , n391638 );
buf ( n394409 , n393587 );
nand ( n46965 , n394408 , n394409 );
buf ( n394411 , n46965 );
buf ( n394412 , n394411 );
nand ( n46968 , n46962 , n394412 );
buf ( n394414 , n46968 );
buf ( n394415 , n394414 );
xor ( n46971 , n394387 , n394415 );
buf ( n394417 , n392788 );
not ( n46973 , n394417 );
buf ( n394419 , n393623 );
not ( n46975 , n394419 );
or ( n46976 , n46973 , n46975 );
buf ( n394422 , n24072 );
not ( n46978 , n394422 );
buf ( n394424 , n37763 );
not ( n46980 , n394424 );
buf ( n394426 , n46980 );
buf ( n394427 , n394426 );
not ( n46983 , n394427 );
or ( n46984 , n46978 , n46983 );
buf ( n394430 , n388952 );
buf ( n394431 , n24071 );
nand ( n46987 , n394430 , n394431 );
buf ( n394433 , n46987 );
buf ( n394434 , n394433 );
nand ( n46990 , n46984 , n394434 );
buf ( n394436 , n46990 );
buf ( n394437 , n394436 );
buf ( n394438 , n391080 );
nand ( n46994 , n394437 , n394438 );
buf ( n394440 , n46994 );
buf ( n394441 , n394440 );
nand ( n46997 , n46976 , n394441 );
buf ( n394443 , n46997 );
buf ( n394444 , n394443 );
and ( n47000 , n46971 , n394444 );
and ( n47001 , n394387 , n394415 );
or ( n47002 , n47000 , n47001 );
buf ( n394448 , n47002 );
buf ( n394449 , n394448 );
buf ( n47005 , n394449 );
buf ( n394451 , n47005 );
buf ( n394452 , n394451 );
not ( n47008 , n394452 );
buf ( n394454 , n388746 );
not ( n47010 , n394454 );
buf ( n394456 , n388760 );
not ( n47012 , n394456 );
buf ( n394458 , n37147 );
not ( n47014 , n394458 );
or ( n47015 , n47012 , n47014 );
buf ( n394461 , n38356 );
not ( n47017 , n394461 );
buf ( n394463 , n47017 );
buf ( n394464 , n394463 );
buf ( n394465 , n388757 );
nand ( n47021 , n394464 , n394465 );
buf ( n394467 , n47021 );
buf ( n394468 , n394467 );
nand ( n47024 , n47015 , n394468 );
buf ( n394470 , n47024 );
buf ( n394471 , n394470 );
not ( n47027 , n394471 );
or ( n47028 , n47010 , n47027 );
buf ( n394474 , n394038 );
buf ( n394475 , n388809 );
nand ( n47031 , n394474 , n394475 );
buf ( n394477 , n47031 );
buf ( n394478 , n394477 );
nand ( n47034 , n47028 , n394478 );
buf ( n394480 , n47034 );
buf ( n394481 , n394480 );
not ( n47037 , n394481 );
or ( n47038 , n47008 , n47037 );
buf ( n394484 , n394451 );
buf ( n394485 , n394480 );
or ( n47041 , n394484 , n394485 );
buf ( n394487 , n389341 );
not ( n47043 , n394487 );
buf ( n394489 , n389753 );
not ( n47045 , n394489 );
or ( n47046 , n47043 , n47045 );
buf ( n394492 , n389997 );
buf ( n394493 , n393185 );
nand ( n47049 , n394492 , n394493 );
buf ( n394495 , n47049 );
buf ( n394496 , n394495 );
nand ( n47052 , n47046 , n394496 );
buf ( n394498 , n47052 );
buf ( n394499 , n394498 );
not ( n47055 , n394499 );
buf ( n394501 , n389015 );
not ( n47057 , n394501 );
or ( n47058 , n47055 , n47057 );
buf ( n394504 , n389024 );
buf ( n394505 , n392828 );
nand ( n47061 , n394504 , n394505 );
buf ( n394507 , n47061 );
buf ( n394508 , n394507 );
nand ( n47064 , n47058 , n394508 );
buf ( n394510 , n47064 );
buf ( n394511 , n394510 );
xor ( n47067 , n393538 , n393550 );
xor ( n47068 , n47067 , n393571 );
buf ( n394514 , n47068 );
buf ( n394515 , n394514 );
xor ( n47071 , n394511 , n394515 );
buf ( n394517 , n42073 );
not ( n47073 , n394517 );
buf ( n394519 , n388576 );
not ( n47075 , n394519 );
or ( n47076 , n47073 , n47075 );
buf ( n394522 , n388556 );
buf ( n394523 , n43144 );
nand ( n47079 , n394522 , n394523 );
buf ( n394525 , n47079 );
buf ( n394526 , n394525 );
nand ( n47082 , n47076 , n394526 );
buf ( n394528 , n47082 );
buf ( n394529 , n394528 );
not ( n47085 , n394529 );
buf ( n394531 , n391652 );
not ( n47087 , n394531 );
or ( n47088 , n47085 , n47087 );
buf ( n394534 , n393890 );
not ( n47090 , n394534 );
buf ( n394536 , n383406 );
nand ( n47092 , n47090 , n394536 );
buf ( n394538 , n47092 );
buf ( n394539 , n394538 );
nand ( n47095 , n47088 , n394539 );
buf ( n394541 , n47095 );
buf ( n394542 , n394541 );
and ( n47098 , n47071 , n394542 );
and ( n47099 , n394511 , n394515 );
or ( n47100 , n47098 , n47099 );
buf ( n394546 , n47100 );
buf ( n394547 , n394546 );
nand ( n47103 , n47041 , n394547 );
buf ( n394549 , n47103 );
buf ( n394550 , n394549 );
nand ( n47106 , n47038 , n394550 );
buf ( n394552 , n47106 );
buf ( n394553 , n394552 );
and ( n47109 , n46879 , n394553 );
and ( n47110 , n394294 , n394323 );
or ( n47111 , n47109 , n47110 );
buf ( n394557 , n47111 );
buf ( n394558 , n394557 );
and ( n47114 , n46824 , n394558 );
and ( n47115 , n394092 , n394268 );
or ( n47116 , n47114 , n47115 );
buf ( n394562 , n47116 );
buf ( n394563 , n394562 );
not ( n47119 , n394563 );
buf ( n394565 , n47119 );
nand ( n47121 , n46636 , n394565 );
not ( n47122 , n47121 );
or ( n47123 , n46632 , n47122 );
buf ( n394569 , n394562 );
buf ( n394570 , n394087 );
nand ( n47126 , n394569 , n394570 );
buf ( n394572 , n47126 );
nand ( n47128 , n47123 , n394572 );
buf ( n394574 , n47128 );
not ( n47130 , n394574 );
buf ( n394576 , n47130 );
buf ( n394577 , n394576 );
nand ( n47133 , n393878 , n394577 );
buf ( n394579 , n47133 );
not ( n47135 , n394579 );
or ( n47136 , n46419 , n47135 );
buf ( n394582 , n393877 );
buf ( n394583 , n394576 );
or ( n47139 , n394582 , n394583 );
buf ( n394585 , n47139 );
nand ( n47141 , n47136 , n394585 );
not ( n47142 , n47141 );
xor ( n47143 , n393729 , n47142 );
xor ( n47144 , n393325 , n45607 );
xor ( n47145 , n47144 , n46239 );
and ( n47146 , n47143 , n47145 );
and ( n47147 , n393729 , n47142 );
or ( n47148 , n47146 , n47147 );
buf ( n394594 , n47148 );
nand ( n47150 , n393723 , n394594 );
buf ( n394596 , n47150 );
buf ( n394597 , n394596 );
xor ( n47153 , n393729 , n47142 );
xor ( n47154 , n47153 , n47145 );
buf ( n394600 , n393665 );
buf ( n394601 , n393687 );
and ( n47157 , n394600 , n394601 );
not ( n47158 , n394600 );
buf ( n394604 , n46226 );
and ( n47160 , n47158 , n394604 );
nor ( n47161 , n47157 , n47160 );
buf ( n394607 , n47161 );
buf ( n394608 , n394607 );
buf ( n394609 , n393333 );
not ( n47165 , n394609 );
buf ( n394611 , n47165 );
buf ( n394612 , n394611 );
and ( n47168 , n394608 , n394612 );
not ( n47169 , n394608 );
buf ( n394615 , n393333 );
and ( n47171 , n47169 , n394615 );
nor ( n47172 , n47168 , n47171 );
buf ( n394618 , n47172 );
buf ( n394619 , n394618 );
and ( n47175 , n393874 , n47128 );
not ( n47176 , n393874 );
and ( n47177 , n47176 , n394576 );
nor ( n47178 , n47175 , n47177 );
not ( n47179 , n393870 );
and ( n47180 , n47178 , n47179 );
not ( n47181 , n47178 );
and ( n47182 , n47181 , n393870 );
nor ( n47183 , n47180 , n47182 );
buf ( n394629 , n47183 );
xor ( n47185 , n394619 , n394629 );
buf ( n394631 , n394083 );
buf ( n394632 , n394087 );
xor ( n47188 , n394631 , n394632 );
buf ( n394634 , n394562 );
xnor ( n47190 , n47188 , n394634 );
buf ( n394636 , n47190 );
buf ( n394637 , n394636 );
xor ( n47193 , n393882 , n394074 );
xor ( n47194 , n47193 , n394079 );
buf ( n394640 , n47194 );
buf ( n394641 , n394640 );
not ( n47197 , n394641 );
buf ( n394643 , n47197 );
buf ( n394644 , n394643 );
buf ( n47200 , n394644 );
buf ( n394646 , n47200 );
not ( n47202 , n394646 );
xor ( n47203 , n394092 , n394268 );
xor ( n47204 , n47203 , n394558 );
buf ( n394650 , n47204 );
buf ( n394651 , n394650 );
not ( n47207 , n394651 );
buf ( n394653 , n47207 );
not ( n47209 , n394653 );
or ( n47210 , n47202 , n47209 );
or ( n47211 , n394646 , n394653 );
buf ( n394657 , n36317 );
not ( n47213 , n394657 );
buf ( n394659 , n47213 );
not ( n47215 , n394659 );
buf ( n394661 , n27258 );
not ( n47217 , n394661 );
buf ( n394663 , n47217 );
buf ( n394664 , n394663 );
not ( n47220 , n394664 );
buf ( n394666 , n47220 );
buf ( n394667 , n394666 );
buf ( n394668 , n388272 );
and ( n47224 , n394667 , n394668 );
not ( n47225 , n394667 );
buf ( n394671 , n393923 );
and ( n47227 , n47225 , n394671 );
nor ( n47228 , n47224 , n47227 );
buf ( n394674 , n47228 );
not ( n47230 , n394674 );
and ( n47231 , n47215 , n47230 );
not ( n47232 , n388626 );
buf ( n394678 , n388263 );
not ( n47234 , n394678 );
buf ( n394680 , n389856 );
not ( n47236 , n394680 );
and ( n47237 , n47234 , n47236 );
buf ( n394683 , n393923 );
buf ( n394684 , n46478 );
and ( n47240 , n394683 , n394684 );
nor ( n47241 , n47237 , n47240 );
buf ( n394687 , n47241 );
not ( n47243 , n394687 );
and ( n47244 , n47232 , n47243 );
nor ( n47245 , n47231 , n47244 );
buf ( n394691 , n47245 );
not ( n47247 , n394691 );
buf ( n394693 , n393537 );
not ( n47249 , n394693 );
or ( n47250 , n47247 , n47249 );
buf ( n394696 , n46532 );
buf ( n394697 , n389593 );
buf ( n394698 , n40824 );
and ( n47254 , n394697 , n394698 );
not ( n47255 , n394697 );
not ( n47256 , n40839 );
buf ( n394702 , n47256 );
and ( n47258 , n47255 , n394702 );
nor ( n47259 , n47254 , n47258 );
buf ( n394705 , n47259 );
buf ( n394706 , n394705 );
or ( n47262 , n394696 , n394706 );
buf ( n394708 , n383937 );
buf ( n394709 , n393994 );
or ( n47265 , n394708 , n394709 );
nand ( n47266 , n47262 , n47265 );
buf ( n394712 , n47266 );
buf ( n394713 , n394712 );
nand ( n47269 , n47250 , n394713 );
buf ( n394715 , n47269 );
buf ( n394716 , n394715 );
buf ( n394717 , n393537 );
not ( n47273 , n394717 );
buf ( n394719 , n47245 );
not ( n47275 , n394719 );
buf ( n394721 , n47275 );
buf ( n394722 , n394721 );
nand ( n47278 , n47273 , n394722 );
buf ( n394724 , n47278 );
buf ( n394725 , n394724 );
nand ( n47281 , n394716 , n394725 );
buf ( n394727 , n47281 );
buf ( n394728 , n394727 );
buf ( n394729 , n392611 );
not ( n47285 , n394729 );
buf ( n394731 , n390453 );
not ( n47287 , n394731 );
or ( n47288 , n47285 , n47287 );
buf ( n394734 , n38685 );
not ( n47290 , n394734 );
buf ( n394736 , n392620 );
nand ( n47292 , n47290 , n394736 );
buf ( n394738 , n47292 );
buf ( n394739 , n394738 );
nand ( n47295 , n47288 , n394739 );
buf ( n394741 , n47295 );
buf ( n394742 , n394741 );
not ( n47298 , n394742 );
buf ( n394744 , n390629 );
not ( n47300 , n394744 );
or ( n47301 , n47298 , n47300 );
buf ( n394747 , n383134 );
not ( n47303 , n394747 );
buf ( n394749 , n394105 );
nand ( n47305 , n47303 , n394749 );
buf ( n394751 , n47305 );
buf ( n394752 , n394751 );
nand ( n47308 , n47301 , n394752 );
buf ( n394754 , n47308 );
buf ( n394755 , n394754 );
xor ( n47311 , n394728 , n394755 );
buf ( n394757 , n394004 );
not ( n47313 , n394757 );
buf ( n394759 , n393950 );
not ( n47315 , n394759 );
buf ( n394761 , n393975 );
not ( n47317 , n394761 );
or ( n47318 , n47315 , n47317 );
buf ( n394764 , n393950 );
buf ( n394765 , n393975 );
or ( n47321 , n394764 , n394765 );
nand ( n47322 , n47318 , n47321 );
buf ( n394768 , n47322 );
buf ( n394769 , n394768 );
not ( n47325 , n394769 );
or ( n47326 , n47313 , n47325 );
buf ( n394772 , n394004 );
buf ( n394773 , n394768 );
or ( n47329 , n394772 , n394773 );
nand ( n47330 , n47326 , n47329 );
buf ( n394776 , n47330 );
buf ( n394777 , n394776 );
and ( n47333 , n47311 , n394777 );
and ( n47334 , n394728 , n394755 );
or ( n47335 , n47333 , n47334 );
buf ( n394781 , n47335 );
buf ( n394782 , n394781 );
not ( n47338 , n394782 );
buf ( n394784 , n47338 );
buf ( n394785 , n394784 );
not ( n47341 , n394785 );
buf ( n394787 , n40858 );
not ( n47343 , n394787 );
buf ( n394789 , n388998 );
not ( n47345 , n394789 );
buf ( n394791 , n40886 );
not ( n47347 , n394791 );
or ( n47348 , n47345 , n47347 );
buf ( n394794 , n40943 );
buf ( n394795 , n388215 );
nand ( n47351 , n394794 , n394795 );
buf ( n394797 , n47351 );
buf ( n394798 , n394797 );
nand ( n47354 , n47348 , n394798 );
buf ( n394800 , n47354 );
buf ( n394801 , n394800 );
not ( n47357 , n394801 );
or ( n47358 , n47343 , n47357 );
buf ( n394804 , n392111 );
buf ( n394805 , n394185 );
nand ( n47361 , n394804 , n394805 );
buf ( n394807 , n47361 );
buf ( n394808 , n394807 );
nand ( n47364 , n47358 , n394808 );
buf ( n394810 , n47364 );
not ( n47366 , n394810 );
buf ( n394812 , n372419 );
not ( n47368 , n394812 );
buf ( n394814 , n47368 );
buf ( n394815 , n394814 );
not ( n47371 , n394815 );
buf ( n394817 , n47371 );
buf ( n394818 , n394817 );
not ( n47374 , n394818 );
buf ( n394820 , n384143 );
not ( n47376 , n394820 );
or ( n47377 , n47374 , n47376 );
buf ( n394823 , n385328 );
buf ( n394824 , n394814 );
nand ( n47380 , n394823 , n394824 );
buf ( n394826 , n47380 );
buf ( n394827 , n394826 );
nand ( n47383 , n47377 , n394827 );
buf ( n394829 , n47383 );
buf ( n394830 , n382938 );
buf ( n394831 , n394225 );
nand ( n47393 , n394830 , n394831 );
buf ( n394833 , n47393 );
buf ( n394834 , n394833 );
nand ( n47396 , C1 , n394834 );
buf ( n394836 , n47396 );
not ( n47398 , n394836 );
or ( n47399 , n47366 , n47398 );
buf ( n394839 , n394836 );
buf ( n394840 , n394810 );
nor ( n47402 , n394839 , n394840 );
buf ( n394842 , n47402 );
buf ( n394843 , n391080 );
not ( n47405 , n394843 );
buf ( n394845 , n24072 );
not ( n47407 , n394845 );
buf ( n394847 , n391483 );
not ( n47409 , n394847 );
or ( n47410 , n47407 , n47409 );
buf ( n47411 , n24070 );
buf ( n47412 , n47411 );
buf ( n394852 , n47412 );
not ( n47414 , n394852 );
buf ( n394854 , n29077 );
nand ( n47416 , n47414 , n394854 );
buf ( n394856 , n47416 );
buf ( n394857 , n394856 );
nand ( n47419 , n47410 , n394857 );
buf ( n394859 , n47419 );
buf ( n394860 , n394859 );
not ( n47422 , n394860 );
or ( n47423 , n47405 , n47422 );
buf ( n394863 , n394436 );
buf ( n394864 , n392788 );
nand ( n47426 , n394863 , n394864 );
buf ( n394866 , n47426 );
buf ( n394867 , n394866 );
nand ( n47429 , n47423 , n394867 );
buf ( n394869 , n47429 );
buf ( n394870 , n394869 );
not ( n47432 , n394870 );
buf ( n394872 , n47432 );
or ( n47434 , n394842 , n394872 );
nand ( n47435 , n47399 , n47434 );
buf ( n394875 , n47435 );
not ( n47437 , n394875 );
buf ( n394877 , n388141 );
not ( n47439 , n394877 );
buf ( n394879 , n394127 );
not ( n47441 , n394879 );
or ( n47442 , n47439 , n47441 );
buf ( n394882 , n388154 );
not ( n47444 , n394882 );
buf ( n394884 , n47444 );
buf ( n394885 , n394884 );
not ( n47447 , n394885 );
buf ( n394887 , n384089 );
not ( n47449 , n394887 );
or ( n47450 , n47447 , n47449 );
buf ( n394890 , n36509 );
buf ( n394891 , n388154 );
nand ( n47453 , n394890 , n394891 );
buf ( n394893 , n47453 );
buf ( n394894 , n394893 );
nand ( n47456 , n47450 , n394894 );
buf ( n394896 , n47456 );
buf ( n394897 , n394896 );
buf ( n394898 , n40701 );
nand ( n47460 , n394897 , n394898 );
buf ( n394900 , n47460 );
buf ( n394901 , n394900 );
nand ( n47463 , n47442 , n394901 );
buf ( n394903 , n47463 );
buf ( n394904 , n394903 );
not ( n47466 , n394904 );
buf ( n394906 , n41342 );
buf ( n394907 , n384239 );
and ( n47469 , n394906 , n394907 );
not ( n47470 , n394906 );
buf ( n394910 , n41595 );
and ( n47472 , n47470 , n394910 );
nor ( n47473 , n47469 , n47472 );
buf ( n394913 , n47473 );
buf ( n394914 , n394913 );
not ( n47476 , n394914 );
buf ( n394916 , n41374 );
not ( n47478 , n394916 );
and ( n47479 , n47476 , n47478 );
buf ( n394919 , n393796 );
buf ( n394920 , n388833 );
and ( n47482 , n394919 , n394920 );
nor ( n47483 , n47479 , n47482 );
buf ( n394923 , n47483 );
buf ( n394924 , n394923 );
nand ( n47486 , n47466 , n394924 );
buf ( n394926 , n47486 );
buf ( n394927 , n394926 );
not ( n47489 , n394927 );
or ( n47490 , n47437 , n47489 );
buf ( n394930 , n394923 );
not ( n47492 , n394930 );
buf ( n394932 , n394903 );
buf ( n47494 , n394932 );
buf ( n394934 , n47494 );
buf ( n394935 , n394934 );
nand ( n47497 , n47492 , n394935 );
buf ( n394937 , n47497 );
buf ( n394938 , n394937 );
nand ( n47500 , n47490 , n394938 );
buf ( n394940 , n47500 );
buf ( n394941 , n394940 );
not ( n47503 , n394941 );
buf ( n394943 , n47503 );
buf ( n394944 , n394943 );
not ( n47506 , n394944 );
or ( n47507 , n47341 , n47506 );
xor ( n47508 , n394013 , n394014 );
buf ( n394948 , n47508 );
xor ( n47510 , n46558 , n394948 );
buf ( n394950 , n47510 );
nand ( n394951 , n47507 , n394950 );
buf ( n394952 , n394951 );
buf ( n394953 , n394952 );
buf ( n394954 , n394940 );
buf ( n394955 , n394781 );
nand ( n47517 , n394954 , n394955 );
buf ( n394957 , n47517 );
buf ( n394958 , n394957 );
nand ( n47520 , n394953 , n394958 );
buf ( n394960 , n47520 );
buf ( n394961 , n394960 );
not ( n47523 , n394961 );
buf ( n394963 , n47523 );
buf ( n394964 , n394963 );
not ( n47526 , n394964 );
buf ( n394966 , n393415 );
buf ( n394967 , n393363 );
and ( n47529 , n394966 , n394967 );
not ( n47530 , n394966 );
buf ( n394970 , n45912 );
and ( n47532 , n47530 , n394970 );
nor ( n47533 , n47529 , n47532 );
buf ( n394973 , n47533 );
buf ( n394974 , n394973 );
buf ( n394975 , n393445 );
xnor ( n47537 , n394974 , n394975 );
buf ( n394977 , n47537 );
buf ( n394978 , n394977 );
not ( n47540 , n394978 );
or ( n47541 , n47526 , n47540 );
buf ( n394981 , n45260 );
not ( n47543 , n394981 );
buf ( n394983 , n392247 );
not ( n47545 , n394983 );
buf ( n394985 , n386421 );
not ( n47547 , n394985 );
or ( n47548 , n47545 , n47547 );
buf ( n394988 , n383056 );
buf ( n394989 , n392244 );
nand ( n47551 , n394988 , n394989 );
buf ( n394991 , n47551 );
buf ( n394992 , n394991 );
nand ( n47554 , n47548 , n394992 );
buf ( n394994 , n47554 );
buf ( n394995 , n394994 );
not ( n47557 , n394995 );
or ( n47558 , n47543 , n47557 );
buf ( n394998 , n393438 );
buf ( n394999 , n392740 );
nand ( n47561 , n394998 , n394999 );
buf ( n395001 , n47561 );
buf ( n395002 , n395001 );
nand ( n47564 , n47558 , n395002 );
buf ( n395004 , n47564 );
buf ( n395005 , n395004 );
not ( n47567 , n395005 );
buf ( n395007 , n36066 );
not ( n47569 , n395007 );
buf ( n395009 , n388105 );
not ( n47571 , n395009 );
and ( n47572 , n47569 , n47571 );
buf ( n395012 , n38822 );
buf ( n395013 , n388105 );
and ( n47575 , n395012 , n395013 );
nor ( n47576 , n47572 , n47575 );
buf ( n395016 , n47576 );
buf ( n395017 , n395016 );
not ( n47579 , n395017 );
buf ( n395019 , n388093 );
not ( n47581 , n395019 );
and ( n47582 , n47579 , n47581 );
buf ( n395022 , n394315 );
buf ( n395023 , n390362 );
and ( n47585 , n395022 , n395023 );
nor ( n47586 , n47582 , n47585 );
buf ( n395026 , n47586 );
buf ( n395027 , n395026 );
not ( n47589 , n395027 );
buf ( n395029 , n47589 );
buf ( n395030 , n395029 );
not ( n47592 , n395030 );
or ( n47593 , n47567 , n47592 );
buf ( n395033 , n395029 );
buf ( n395034 , n395004 );
or ( n47596 , n395033 , n395034 );
xor ( n47597 , n393771 , n393778 );
xor ( n47598 , n47597 , n393804 );
buf ( n395038 , n47598 );
buf ( n395039 , n395038 );
nand ( n47601 , n47596 , n395039 );
buf ( n395041 , n47601 );
buf ( n395042 , n395041 );
nand ( n47604 , n47593 , n395042 );
buf ( n395044 , n47604 );
buf ( n395045 , n395044 );
nand ( n47607 , n47541 , n395045 );
buf ( n395047 , n47607 );
buf ( n395048 , n395047 );
buf ( n395049 , n394977 );
not ( n47611 , n395049 );
buf ( n395051 , n394960 );
nand ( n47613 , n47611 , n395051 );
buf ( n395053 , n47613 );
buf ( n395054 , n395053 );
nand ( n47616 , n395048 , n395054 );
buf ( n395056 , n47616 );
not ( n47618 , n395056 );
nand ( n47619 , n47211 , n47618 );
nand ( n47620 , n47210 , n47619 );
buf ( n395060 , n47620 );
xor ( n47622 , n394637 , n395060 );
not ( n47623 , n46609 );
not ( n47624 , n394048 );
or ( n47625 , n47623 , n47624 );
not ( n47626 , n46609 );
nand ( n47627 , n47626 , n394045 );
nand ( n47628 , n47625 , n47627 );
buf ( n395068 , n47628 );
buf ( n395069 , n394019 );
buf ( n47631 , n395069 );
buf ( n395071 , n47631 );
buf ( n395072 , n395071 );
not ( n47634 , n395072 );
buf ( n395074 , n47634 );
buf ( n395075 , n395074 );
and ( n47637 , n395068 , n395075 );
not ( n47638 , n395068 );
buf ( n395078 , n395071 );
and ( n47640 , n47638 , n395078 );
nor ( n47641 , n47637 , n47640 );
buf ( n395081 , n47641 );
buf ( n395082 , n395081 );
xor ( n47644 , n394114 , n394141 );
xor ( n47645 , n47644 , n394235 );
buf ( n395085 , n47645 );
buf ( n395086 , n395085 );
not ( n47648 , n395086 );
buf ( n395088 , n43727 );
not ( n47650 , n395088 );
buf ( n395090 , n391027 );
not ( n47652 , n395090 );
buf ( n395092 , n42616 );
not ( n47654 , n395092 );
or ( n47655 , n47652 , n47654 );
buf ( n395095 , n35301 );
buf ( n395096 , n391024 );
nand ( n47658 , n395095 , n395096 );
buf ( n395098 , n47658 );
buf ( n395099 , n395098 );
nand ( n47661 , n47655 , n395099 );
buf ( n395101 , n47661 );
buf ( n395102 , n395101 );
not ( n47664 , n395102 );
or ( n47665 , n47650 , n47664 );
buf ( n395105 , n394283 );
buf ( n395106 , n43515 );
nand ( n47668 , n395105 , n395106 );
buf ( n395108 , n47668 );
buf ( n395109 , n395108 );
nand ( n47671 , n47665 , n395109 );
buf ( n395111 , n47671 );
buf ( n395112 , n395111 );
not ( n47674 , n395112 );
or ( n47675 , n47648 , n47674 );
buf ( n395115 , n395111 );
buf ( n395116 , n395085 );
or ( n47678 , n395115 , n395116 );
xor ( n47679 , n394171 , n394200 );
xnor ( n47680 , n47679 , n46782 );
buf ( n395120 , n47680 );
buf ( n395121 , n40990 );
not ( n47683 , n395121 );
buf ( n395123 , n394392 );
not ( n47685 , n395123 );
or ( n47686 , n47683 , n47685 );
buf ( n395126 , n390498 );
buf ( n395127 , n390460 );
nand ( n47689 , n395126 , n395127 );
buf ( n395129 , n47689 );
buf ( n395130 , n395129 );
nand ( n47692 , n47686 , n395130 );
buf ( n395132 , n47692 );
buf ( n395133 , n395132 );
not ( n47695 , n395133 );
buf ( n395135 , n389880 );
not ( n47697 , n395135 );
or ( n47698 , n47695 , n47697 );
buf ( n395138 , n394402 );
buf ( n395139 , n392666 );
nand ( n47701 , n395138 , n395139 );
buf ( n395141 , n47701 );
buf ( n395142 , n395141 );
nand ( n47704 , n47698 , n395142 );
buf ( n395144 , n47704 );
buf ( n395145 , n395144 );
not ( n47707 , n395145 );
buf ( n395147 , n40701 );
not ( n47709 , n395147 );
buf ( n395149 , n394884 );
not ( n47711 , n395149 );
buf ( n395151 , n38660 );
not ( n47713 , n395151 );
or ( n47714 , n47711 , n47713 );
buf ( n395154 , n36564 );
buf ( n395155 , n388154 );
nand ( n47717 , n395154 , n395155 );
buf ( n395157 , n47717 );
buf ( n395158 , n395157 );
nand ( n47720 , n47714 , n395158 );
buf ( n395160 , n47720 );
buf ( n395161 , n395160 );
not ( n47723 , n395161 );
or ( n47724 , n47709 , n47723 );
buf ( n395164 , n394896 );
buf ( n47726 , n40639 );
buf ( n395166 , n47726 );
nand ( n47728 , n395164 , n395166 );
buf ( n395168 , n47728 );
buf ( n395169 , n395168 );
nand ( n47731 , n47724 , n395169 );
buf ( n395171 , n47731 );
buf ( n395172 , n395171 );
not ( n47734 , n395172 );
or ( n47735 , n47707 , n47734 );
buf ( n395175 , n395171 );
buf ( n395176 , n395144 );
or ( n47738 , n395175 , n395176 );
not ( n47739 , n38961 );
buf ( n395179 , n22982 );
not ( n47741 , n395179 );
buf ( n395181 , n388409 );
not ( n47743 , n395181 );
or ( n47744 , n47741 , n47743 );
buf ( n395184 , n388406 );
buf ( n395185 , n46906 );
nand ( n47747 , n395184 , n395185 );
buf ( n395187 , n47747 );
buf ( n395188 , n395187 );
nand ( n47750 , n47744 , n395188 );
buf ( n395190 , n47750 );
not ( n47752 , n395190 );
or ( n47753 , n47739 , n47752 );
not ( n47754 , n22982 );
or ( n47755 , n391569 , n47754 );
not ( n47756 , n375822 );
nand ( n47757 , n47756 , n47754 );
buf ( n395197 , n386474 );
not ( n47759 , n395197 );
buf ( n395199 , n47759 );
nand ( n47761 , n47755 , n47757 , n395199 );
nand ( n47762 , n47753 , n47761 );
buf ( n395202 , n47762 );
buf ( n395203 , n41565 );
not ( n47765 , n395203 );
buf ( n395205 , n394382 );
not ( n47767 , n395205 );
or ( n47768 , n47765 , n47767 );
buf ( n395208 , n40758 );
not ( n47770 , n395208 );
buf ( n395210 , n45391 );
not ( n47772 , n395210 );
and ( n47773 , n47770 , n47772 );
buf ( n395213 , n27613 );
buf ( n395214 , n45391 );
and ( n47776 , n395213 , n395214 );
nor ( n47777 , n47773 , n47776 );
buf ( n395217 , n47777 );
buf ( n395218 , n395217 );
not ( n47780 , n395218 );
buf ( n395220 , n389125 );
nand ( n47782 , n47780 , n395220 );
buf ( n395222 , n47782 );
buf ( n395223 , n395222 );
nand ( n47785 , n47768 , n395223 );
buf ( n395225 , n47785 );
buf ( n395226 , n395225 );
xor ( n47788 , n395202 , n395226 );
not ( n47789 , n388546 );
not ( n47790 , n388608 );
or ( n47791 , n47789 , n47790 );
nand ( n47792 , n388266 , n388543 );
nand ( n47793 , n47791 , n47792 );
buf ( n395233 , n47793 );
not ( n47795 , n395233 );
buf ( n395235 , n383891 );
not ( n47797 , n395235 );
or ( n47798 , n47795 , n47797 );
buf ( n395238 , n394674 );
not ( n47800 , n395238 );
buf ( n395240 , n383907 );
nand ( n47802 , n47800 , n395240 );
buf ( n395242 , n47802 );
buf ( n395243 , n395242 );
nand ( n47805 , n47798 , n395243 );
buf ( n395245 , n47805 );
buf ( n395246 , n395245 );
and ( n47808 , n47788 , n395246 );
and ( n47809 , n395202 , n395226 );
or ( n47810 , n47808 , n47809 );
buf ( n395250 , n47810 );
buf ( n395251 , n395250 );
nand ( n47813 , n47738 , n395251 );
buf ( n395253 , n47813 );
buf ( n395254 , n395253 );
nand ( n47816 , n47735 , n395254 );
buf ( n395256 , n47816 );
buf ( n395257 , n395256 );
xor ( n47819 , n395120 , n395257 );
buf ( n395259 , n388809 );
not ( n47821 , n395259 );
buf ( n395261 , n394470 );
not ( n47823 , n395261 );
or ( n47824 , n47821 , n47823 );
buf ( n395264 , n388760 );
not ( n47826 , n395264 );
buf ( n395266 , n389525 );
not ( n47828 , n395266 );
or ( n47829 , n47826 , n47828 );
buf ( n395269 , n37173 );
buf ( n395270 , n388757 );
nand ( n47832 , n395269 , n395270 );
buf ( n395272 , n47832 );
buf ( n395273 , n395272 );
nand ( n47835 , n47829 , n395273 );
buf ( n395275 , n47835 );
buf ( n395276 , n395275 );
buf ( n395277 , n388746 );
nand ( n47839 , n395276 , n395277 );
buf ( n395279 , n47839 );
buf ( n395280 , n395279 );
nand ( n47842 , n47824 , n395280 );
buf ( n395282 , n47842 );
buf ( n395283 , n395282 );
and ( n47845 , n47819 , n395283 );
and ( n47846 , n395120 , n395257 );
or ( n47847 , n47845 , n47846 );
buf ( n395287 , n47847 );
buf ( n395288 , n395287 );
nand ( n47850 , n47678 , n395288 );
buf ( n395290 , n47850 );
buf ( n395291 , n395290 );
nand ( n47853 , n47675 , n395291 );
buf ( n395293 , n47853 );
buf ( n395294 , n395293 );
xor ( n47856 , n395082 , n395294 );
xor ( n47857 , n394448 , n394480 );
xnor ( n47858 , n47857 , n394546 );
buf ( n395298 , n47858 );
not ( n47860 , n395298 );
buf ( n395300 , n47860 );
not ( n47862 , n395300 );
not ( n47863 , n23603 );
buf ( n395303 , n47863 );
not ( n47865 , n395303 );
buf ( n395305 , n34859 );
not ( n47867 , n395305 );
or ( n47868 , n47865 , n47867 );
buf ( n395308 , n393374 );
not ( n47870 , n395308 );
buf ( n395310 , n47863 );
not ( n47872 , n395310 );
buf ( n395312 , n47872 );
buf ( n395313 , n395312 );
buf ( n47875 , n395313 );
buf ( n395315 , n47875 );
buf ( n395316 , n395315 );
nand ( n47878 , n47870 , n395316 );
buf ( n395318 , n47878 );
buf ( n395319 , n395318 );
nand ( n47881 , n47868 , n395319 );
buf ( n395321 , n47881 );
buf ( n395322 , n395321 );
buf ( n395323 , n371183 );
not ( n47885 , n395323 );
buf ( n395325 , n47885 );
buf ( n395326 , n395325 );
not ( n47888 , n395326 );
buf ( n395328 , n47888 );
nand ( n47890 , n23604 , n395328 );
buf ( n47891 , n23551 );
buf ( n395331 , n47891 );
not ( n47893 , n395331 );
buf ( n395333 , n47893 );
buf ( n395334 , n395333 );
buf ( n395335 , n371183 );
xor ( n47897 , n395334 , n395335 );
buf ( n395337 , n47897 );
buf ( n395338 , n23603 );
buf ( n395339 , n395325 );
nand ( n47901 , n395338 , n395339 );
buf ( n395341 , n47901 );
and ( n47903 , n47890 , n395337 , n395341 );
not ( n47904 , n47903 );
buf ( n395344 , n47904 );
not ( n47906 , n395344 );
buf ( n395346 , n47906 );
buf ( n395347 , n395346 );
buf ( n47909 , n395347 );
buf ( n395349 , n47909 );
buf ( n395350 , n395349 );
not ( n47912 , n395350 );
buf ( n395352 , n47912 );
buf ( n395353 , n395352 );
buf ( n395354 , n395337 );
not ( n47916 , n395354 );
buf ( n395356 , n47916 );
buf ( n395357 , n395356 );
buf ( n47919 , n395357 );
buf ( n395359 , n47919 );
buf ( n395360 , n395359 );
buf ( n47922 , n395360 );
buf ( n395362 , n47922 );
buf ( n395363 , n395362 );
not ( n47925 , n395363 );
buf ( n395365 , n47925 );
buf ( n395366 , n395365 );
nand ( n47928 , n395353 , n395366 );
buf ( n395368 , n47928 );
buf ( n395369 , n395368 );
nand ( n47931 , n395322 , n395369 );
buf ( n395371 , n47931 );
buf ( n395372 , n395371 );
buf ( n395373 , n45954 );
not ( n47935 , n395373 );
buf ( n395375 , n393839 );
not ( n47937 , n395375 );
or ( n47938 , n47935 , n47937 );
buf ( n395378 , n393369 );
not ( n47940 , n395378 );
buf ( n395380 , n392144 );
not ( n47942 , n395380 );
or ( n47943 , n47940 , n47942 );
buf ( n395383 , n35519 );
buf ( n395384 , n393381 );
nand ( n47946 , n395383 , n395384 );
buf ( n395386 , n47946 );
buf ( n395387 , n395386 );
nand ( n47949 , n47943 , n395387 );
buf ( n395389 , n47949 );
buf ( n395390 , n395389 );
buf ( n395391 , n393825 );
nand ( n47953 , n395390 , n395391 );
buf ( n395393 , n47953 );
buf ( n395394 , n395393 );
nand ( n47956 , n47938 , n395394 );
buf ( n395396 , n47956 );
buf ( n395397 , n395396 );
xor ( n47959 , n395372 , n395397 );
not ( n47960 , n389162 );
not ( n47961 , n46365 );
or ( n47962 , n47960 , n47961 );
buf ( n395402 , n41671 );
not ( n47964 , n395402 );
buf ( n395404 , n42234 );
not ( n47966 , n395404 );
or ( n47967 , n47964 , n47966 );
buf ( n395407 , n36217 );
buf ( n395408 , n41670 );
nand ( n47970 , n395407 , n395408 );
buf ( n395410 , n47970 );
buf ( n395411 , n395410 );
nand ( n47973 , n47967 , n395411 );
buf ( n395413 , n47973 );
buf ( n395414 , n395413 );
buf ( n395415 , n41711 );
nand ( n47977 , n395414 , n395415 );
buf ( n395417 , n47977 );
nand ( n47979 , n47962 , n395417 );
buf ( n395419 , n47979 );
and ( n47981 , n47959 , n395419 );
and ( n47982 , n395372 , n395397 );
or ( n47983 , n47981 , n47982 );
buf ( n395423 , n47983 );
not ( n47985 , n395423 );
or ( n47986 , n47862 , n47985 );
buf ( n395426 , n395423 );
not ( n47988 , n395426 );
buf ( n395428 , n47988 );
not ( n47990 , n395428 );
not ( n47991 , n47858 );
or ( n47992 , n47990 , n47991 );
buf ( n395432 , n41447 );
not ( n47994 , n395432 );
buf ( n395434 , n393505 );
not ( n47996 , n395434 );
or ( n47997 , n47994 , n47996 );
buf ( n395437 , n46056 );
buf ( n395438 , n393557 );
not ( n48000 , n395438 );
buf ( n395440 , n393525 );
not ( n48002 , n395440 );
or ( n48003 , n48000 , n48002 );
buf ( n395443 , n385473 );
buf ( n395444 , n388367 );
nand ( n48006 , n395443 , n395444 );
buf ( n395446 , n48006 );
buf ( n395447 , n395446 );
nand ( n48009 , n48003 , n395447 );
buf ( n395449 , n48009 );
buf ( n395450 , n395449 );
nand ( n48012 , n395437 , n395450 );
buf ( n395452 , n48012 );
buf ( n395453 , n395452 );
nand ( n48015 , n47997 , n395453 );
buf ( n395455 , n48015 );
buf ( n395456 , n395455 );
not ( n48018 , n395456 );
buf ( n395458 , n48018 );
buf ( n395459 , n395458 );
not ( n48021 , n395459 );
or ( n48022 , n391569 , n47754 );
nand ( n48023 , n48022 , n47757 );
not ( n48024 , n48023 );
buf ( n48025 , n38960 );
not ( n48026 , n48025 );
and ( n48027 , n48024 , n48026 );
buf ( n395467 , n386474 );
not ( n48029 , n395467 );
buf ( n395469 , n48029 );
and ( n48031 , n394357 , n395469 );
nor ( n48032 , n48027 , n48031 );
buf ( n395472 , n48032 );
not ( n48034 , n395472 );
or ( n48035 , n48021 , n48034 );
buf ( n395475 , n43058 );
buf ( n395476 , n391563 );
not ( n48038 , n395476 );
buf ( n395478 , n48038 );
buf ( n395479 , n395478 );
not ( n48041 , n395479 );
buf ( n395481 , n46478 );
not ( n48043 , n395481 );
and ( n48044 , n48041 , n48043 );
buf ( n395484 , n393562 );
buf ( n395485 , n46478 );
and ( n48047 , n395484 , n395485 );
nor ( n48048 , n48044 , n48047 );
buf ( n395488 , n48048 );
buf ( n395489 , n395488 );
or ( n48051 , n395475 , n395489 );
buf ( n395491 , n394338 );
buf ( n395492 , n37315 );
or ( n48054 , n395491 , n395492 );
nand ( n48055 , n48051 , n48054 );
buf ( n395495 , n48055 );
buf ( n395496 , n395495 );
nand ( n48058 , n48035 , n395496 );
buf ( n395498 , n48058 );
buf ( n395499 , n395498 );
buf ( n395500 , n48032 );
not ( n48062 , n395500 );
buf ( n395502 , n395455 );
nand ( n48064 , n48062 , n395502 );
buf ( n395504 , n48064 );
buf ( n395505 , n395504 );
nand ( n48067 , n395499 , n395505 );
buf ( n395507 , n48067 );
buf ( n395508 , n391446 );
not ( n48070 , n395508 );
buf ( n395510 , n389753 );
not ( n48072 , n395510 );
or ( n48073 , n48070 , n48072 );
buf ( n395513 , n389997 );
buf ( n395514 , n391455 );
nand ( n48076 , n395513 , n395514 );
buf ( n395516 , n48076 );
buf ( n395517 , n395516 );
nand ( n48079 , n48073 , n395517 );
buf ( n395519 , n48079 );
not ( n48081 , n395519 );
not ( n48082 , n389015 );
or ( n48083 , n48081 , n48082 );
buf ( n395523 , n394498 );
buf ( n395524 , n389328 );
nand ( n48086 , n395523 , n395524 );
buf ( n395526 , n48086 );
nand ( n48088 , n48083 , n395526 );
xor ( n48089 , n395507 , n48088 );
not ( n48090 , n46917 );
not ( n48091 , n46939 );
and ( n48092 , n48090 , n48091 );
and ( n48093 , n46917 , n46939 );
nor ( n48094 , n48092 , n48093 );
buf ( n48095 , n46896 );
and ( n48096 , n48094 , n48095 );
not ( n48097 , n48094 );
not ( n48098 , n48095 );
and ( n48099 , n48097 , n48098 );
nor ( n48100 , n48096 , n48099 );
and ( n48101 , n48089 , n48100 );
and ( n48102 , n395507 , n48088 );
or ( n48103 , n48101 , n48102 );
not ( n48104 , n48103 );
not ( n48105 , n48104 );
xor ( n48106 , n394387 , n394415 );
xor ( n48107 , n48106 , n394444 );
buf ( n395547 , n48107 );
not ( n48109 , n395547 );
not ( n48110 , n48109 );
or ( n48111 , n48105 , n48110 );
xor ( n48112 , n394511 , n394515 );
xor ( n48113 , n48112 , n394542 );
buf ( n395553 , n48113 );
nand ( n48115 , n48111 , n395553 );
not ( n48116 , n48109 );
nand ( n48117 , n48116 , n48103 );
nand ( n48118 , n48115 , n48117 );
nand ( n48119 , n47992 , n48118 );
nand ( n48120 , n47986 , n48119 );
buf ( n395560 , n48120 );
and ( n48122 , n47856 , n395560 );
and ( n48123 , n395082 , n395294 );
or ( n48124 , n48122 , n48123 );
buf ( n395564 , n48124 );
not ( n48126 , n395564 );
buf ( n395566 , n46407 );
buf ( n395567 , n46293 );
and ( n48129 , n395566 , n395567 );
not ( n48130 , n395566 );
buf ( n395570 , n46301 );
and ( n48132 , n48130 , n395570 );
nor ( n48133 , n48129 , n48132 );
buf ( n395573 , n48133 );
not ( n48135 , n46297 );
and ( n48136 , n395573 , n48135 );
not ( n48137 , n395573 );
and ( n48138 , n48137 , n46297 );
nor ( n48139 , n48136 , n48138 );
nand ( n48140 , n48126 , n48139 );
buf ( n395580 , n48140 );
xor ( n48142 , n394294 , n394323 );
xor ( n48143 , n48142 , n394553 );
buf ( n395583 , n48143 );
buf ( n48145 , n395583 );
not ( n48146 , n48145 );
xor ( n48147 , n394240 , n394251 );
xor ( n48148 , n48147 , n394263 );
buf ( n395588 , n48148 );
not ( n48150 , n395588 );
nand ( n48151 , n48146 , n48150 );
not ( n48152 , n48151 );
not ( n48153 , n46305 );
not ( n48154 , n48153 );
xor ( n48155 , n393808 , n46405 );
not ( n48156 , n48155 );
or ( n48157 , n48154 , n48156 );
or ( n48158 , n48155 , n48153 );
nand ( n48159 , n48157 , n48158 );
not ( n48160 , n48159 );
or ( n48161 , n48152 , n48160 );
nand ( n48162 , n48145 , n395588 );
nand ( n48163 , n48161 , n48162 );
buf ( n395603 , n48163 );
and ( n48165 , n395580 , n395603 );
buf ( n395605 , n395564 );
not ( n48167 , n395605 );
buf ( n395607 , n48139 );
nor ( n48169 , n48167 , n395607 );
buf ( n395609 , n48169 );
buf ( n395610 , n395609 );
nor ( n48172 , n48165 , n395610 );
buf ( n395612 , n48172 );
buf ( n395613 , n395612 );
and ( n48175 , n47622 , n395613 );
and ( n48176 , n394637 , n395060 );
or ( n48177 , n48175 , n48176 );
buf ( n395617 , n48177 );
buf ( n395618 , n395617 );
and ( n48180 , n47185 , n395618 );
and ( n48181 , n394619 , n394629 );
or ( n48182 , n48180 , n48181 );
buf ( n395622 , n48182 );
nand ( n48184 , n47154 , n395622 );
buf ( n395624 , n48184 );
nand ( n48186 , n42852 , n44738 );
not ( n48187 , n48186 );
not ( n48188 , n45579 );
or ( n48189 , n48187 , n48188 );
nand ( n48190 , n42851 , n44737 );
nand ( n48191 , n48189 , n48190 );
buf ( n395631 , n48191 );
not ( n48193 , n395631 );
xor ( n48194 , n389220 , n42561 );
and ( n48195 , n48194 , n390325 );
and ( n48196 , n389220 , n42561 );
or ( n48197 , n48195 , n48196 );
buf ( n395637 , n48197 );
not ( n48199 , n44510 );
not ( n48200 , n391696 );
or ( n48201 , n48199 , n48200 );
not ( n48202 , n44510 );
not ( n48203 , n48202 );
not ( n48204 , n391699 );
or ( n48205 , n48203 , n48204 );
nand ( n48206 , n48205 , n44732 );
nand ( n48207 , n48201 , n48206 );
buf ( n395647 , n48207 );
xor ( n48209 , n395637 , n395647 );
xor ( n48210 , n44235 , n391945 );
and ( n48211 , n48210 , n391974 );
and ( n48212 , n44235 , n391945 );
or ( n48213 , n48211 , n48212 );
xor ( n48214 , n391711 , n391818 );
and ( n48215 , n48214 , n391943 );
and ( n48216 , n391711 , n391818 );
or ( n48217 , n48215 , n48216 );
buf ( n395657 , n48217 );
buf ( n395658 , n395657 );
xor ( n48220 , n391844 , n391857 );
and ( n48221 , n48220 , n391940 );
and ( n48222 , n391844 , n391857 );
or ( n48223 , n48221 , n48222 );
buf ( n395663 , n48223 );
buf ( n395664 , n395663 );
buf ( n395665 , n386480 );
not ( n48227 , n395665 );
buf ( n395667 , n38972 );
not ( n48229 , n395667 );
buf ( n395669 , n37215 );
not ( n48231 , n395669 );
or ( n48232 , n48229 , n48231 );
not ( n48233 , n36216 );
not ( n48234 , n48233 );
buf ( n395674 , n48234 );
buf ( n395675 , n38971 );
nand ( n48237 , n395674 , n395675 );
buf ( n395677 , n48237 );
buf ( n395678 , n395677 );
nand ( n48240 , n48232 , n395678 );
buf ( n395680 , n48240 );
buf ( n395681 , n395680 );
not ( n48243 , n395681 );
or ( n48244 , n48227 , n48243 );
buf ( n395684 , n390126 );
buf ( n395685 , n386496 );
nand ( n48247 , n395684 , n395685 );
buf ( n395687 , n48247 );
buf ( n395688 , n395687 );
nand ( n48250 , n48244 , n395688 );
buf ( n395690 , n48250 );
buf ( n395691 , n395690 );
xor ( n48253 , n391883 , n391913 );
and ( n48254 , n48253 , n391937 );
and ( n48255 , n391883 , n391913 );
or ( n48256 , n48254 , n48255 );
buf ( n395696 , n48256 );
buf ( n395697 , n395696 );
xor ( n48259 , n395691 , n395697 );
not ( n48260 , n388498 );
buf ( n395700 , n385328 );
not ( n48262 , n395700 );
buf ( n395702 , n388242 );
not ( n48264 , n395702 );
and ( n48265 , n48262 , n48264 );
buf ( n395705 , n385292 );
buf ( n395706 , n388242 );
and ( n48268 , n395705 , n395706 );
nor ( n48269 , n48265 , n48268 );
buf ( n395709 , n48269 );
not ( n48271 , n395709 );
and ( n48272 , n48260 , n48271 );
nor ( n48275 , n48272 , C0 );
buf ( n395713 , n390292 );
not ( n48277 , n395713 );
buf ( n395715 , n390311 );
not ( n48279 , n395715 );
and ( n48280 , n48277 , n48279 );
buf ( n395718 , n36845 );
buf ( n395719 , n40971 );
buf ( n395720 , n36809 );
not ( n48284 , n395720 );
buf ( n395722 , n48284 );
buf ( n395723 , n395722 );
and ( n48287 , n395719 , n395723 );
not ( n48288 , n395719 );
buf ( n395726 , n40890 );
and ( n48290 , n48288 , n395726 );
nor ( n48291 , n48287 , n48290 );
buf ( n395729 , n48291 );
buf ( n395730 , n395729 );
nor ( n48294 , n395718 , n395730 );
buf ( n395732 , n48294 );
buf ( n395733 , n395732 );
nor ( n48297 , n48280 , n395733 );
buf ( n395735 , n48297 );
buf ( n395736 , n395735 );
not ( n48300 , n395736 );
buf ( n395738 , n48300 );
buf ( n395739 , n395738 );
buf ( n395740 , n391798 );
not ( n48304 , n395740 );
buf ( n395742 , n382598 );
not ( n48306 , n395742 );
or ( n48307 , n48304 , n48306 );
buf ( n395745 , n386212 );
buf ( n395746 , n389862 );
not ( n48310 , n395746 );
buf ( n395748 , n385987 );
not ( n48312 , n395748 );
or ( n48313 , n48310 , n48312 );
buf ( n395751 , n389997 );
buf ( n395752 , n389859 );
nand ( n48316 , n395751 , n395752 );
buf ( n395754 , n48316 );
buf ( n395755 , n395754 );
nand ( n48319 , n48313 , n395755 );
buf ( n395757 , n48319 );
buf ( n395758 , n395757 );
nand ( n48322 , n395745 , n395758 );
buf ( n395760 , n48322 );
buf ( n395761 , n395760 );
nand ( n48325 , n48307 , n395761 );
buf ( n395763 , n48325 );
buf ( n395764 , n395763 );
xor ( n48328 , n395739 , n395764 );
buf ( n395766 , n48328 );
not ( n48330 , n395766 );
xor ( n48331 , n48275 , n48330 );
buf ( n395769 , n48331 );
xor ( n48333 , n48259 , n395769 );
buf ( n395771 , n48333 );
buf ( n395772 , n395771 );
xor ( n48336 , n395664 , n395772 );
buf ( n395774 , n384644 );
not ( n48338 , n395774 );
buf ( n395776 , n389928 );
not ( n48340 , n395776 );
buf ( n395778 , n41904 );
not ( n48342 , n395778 );
or ( n48343 , n48340 , n48342 );
buf ( n395781 , n385324 );
buf ( n395782 , n36251 );
nand ( n48346 , n395781 , n395782 );
buf ( n395784 , n48346 );
buf ( n395785 , n395784 );
nand ( n48349 , n48343 , n395785 );
buf ( n395787 , n48349 );
buf ( n395788 , n395787 );
not ( n48352 , n395788 );
or ( n48353 , n48338 , n48352 );
buf ( n395791 , n383894 );
buf ( n395792 , n44300 );
nand ( n48356 , n395791 , n395792 );
buf ( n395794 , n48356 );
buf ( n395795 , n395794 );
nand ( n48359 , n48353 , n395795 );
buf ( n395797 , n48359 );
buf ( n395798 , n395797 );
buf ( n395799 , n390280 );
not ( n48363 , n395799 );
buf ( n395801 , n390260 );
not ( n48365 , n395801 );
or ( n48366 , n48363 , n48365 );
and ( n48367 , n388928 , n42799 );
not ( n48368 , n388928 );
and ( n48369 , n48368 , n40840 );
nor ( n48370 , n48367 , n48369 );
buf ( n395808 , n48370 );
not ( n48372 , n395808 );
buf ( n395810 , n43272 );
nand ( n48374 , n48372 , n395810 );
buf ( n395812 , n48374 );
buf ( n395813 , n395812 );
nand ( n48377 , n48366 , n395813 );
buf ( n395815 , n48377 );
buf ( n395816 , n395815 );
not ( n48380 , n395816 );
buf ( n395818 , n48380 );
buf ( n395819 , n395818 );
xor ( n48383 , n395798 , n395819 );
buf ( n395821 , n385269 );
not ( n48385 , n395821 );
buf ( n395823 , n391901 );
not ( n48387 , n395823 );
or ( n48388 , n48385 , n48387 );
buf ( n395826 , n37347 );
not ( n48390 , n395826 );
buf ( n395828 , n385983 );
not ( n48392 , n395828 );
buf ( n395830 , n48392 );
buf ( n395831 , n395830 );
not ( n48395 , n395831 );
or ( n48396 , n48390 , n48395 );
buf ( n395834 , n385983 );
buf ( n395835 , n391895 );
nand ( n48399 , n395834 , n395835 );
buf ( n395837 , n48399 );
buf ( n395838 , n395837 );
nand ( n48402 , n48396 , n395838 );
buf ( n395840 , n48402 );
buf ( n395841 , n395840 );
buf ( n395842 , n37695 );
nand ( n48406 , n395841 , n395842 );
buf ( n395844 , n48406 );
buf ( n395845 , n395844 );
nand ( n48409 , n48388 , n395845 );
buf ( n395847 , n48409 );
buf ( n395848 , n395847 );
xor ( n48412 , n48383 , n395848 );
buf ( n395850 , n48412 );
buf ( n395851 , n395850 );
buf ( n395852 , n41711 );
not ( n48416 , n395852 );
buf ( n395854 , n390071 );
not ( n48418 , n395854 );
or ( n48419 , n48416 , n48418 );
and ( n48420 , n38532 , n24118 );
not ( n48421 , n38532 );
and ( n48422 , n48421 , n41670 );
or ( n48423 , n48420 , n48422 );
buf ( n395861 , n48423 );
buf ( n395862 , n389162 );
nand ( n48426 , n395861 , n395862 );
buf ( n395864 , n48426 );
buf ( n395865 , n395864 );
nand ( n48429 , n48419 , n395865 );
buf ( n395867 , n48429 );
buf ( n395868 , n395867 );
xor ( n48432 , n395851 , n395868 );
buf ( n395870 , n384621 );
buf ( n395871 , n44410 );
not ( n48435 , n395871 );
buf ( n395873 , n48435 );
buf ( n395874 , n395873 );
or ( n48438 , n395870 , n395874 );
buf ( n395876 , n40819 );
buf ( n395877 , n389897 );
not ( n48441 , n395877 );
buf ( n395879 , n48441 );
buf ( n395880 , n395879 );
and ( n48444 , n395876 , n395880 );
not ( n48445 , n395876 );
buf ( n395883 , n42390 );
not ( n48447 , n395883 );
buf ( n395885 , n48447 );
buf ( n395886 , n395885 );
and ( n48450 , n48445 , n395886 );
nor ( n48451 , n48444 , n48450 );
buf ( n395889 , n48451 );
buf ( n395890 , n395889 );
buf ( n395891 , n384551 );
or ( n48455 , n395890 , n395891 );
nand ( n48456 , n48438 , n48455 );
buf ( n395894 , n48456 );
buf ( n395895 , n395894 );
buf ( n395896 , n390230 );
not ( n48460 , n395896 );
buf ( n395898 , n48460 );
not ( n48462 , n395898 );
not ( n48463 , n383017 );
or ( n48464 , n48462 , n48463 );
not ( n48465 , n383027 );
not ( n48466 , n388546 );
or ( n48467 , n48465 , n48466 );
nand ( n48468 , n383024 , n388549 );
nand ( n48469 , n48467 , n48468 );
nand ( n48470 , n48469 , n390635 );
nand ( n48471 , n48464 , n48470 );
buf ( n395909 , n48471 );
xor ( n48473 , n395895 , n395909 );
buf ( n395911 , n391164 );
buf ( n395912 , n391932 );
or ( n48476 , n395911 , n395912 );
buf ( n395914 , n383499 );
buf ( n395915 , n388376 );
not ( n48479 , n395915 );
buf ( n395917 , n385630 );
not ( n48481 , n395917 );
buf ( n395919 , n48481 );
buf ( n395920 , n395919 );
not ( n48484 , n395920 );
or ( n48485 , n48479 , n48484 );
buf ( n395923 , n389589 );
buf ( n395924 , n388373 );
nand ( n48488 , n395923 , n395924 );
buf ( n395926 , n48488 );
buf ( n395927 , n395926 );
nand ( n48491 , n48485 , n395927 );
buf ( n395929 , n48491 );
buf ( n395930 , n395929 );
not ( n48494 , n395930 );
buf ( n395932 , n48494 );
buf ( n395933 , n395932 );
or ( n48497 , n395914 , n395933 );
nand ( n48498 , n48476 , n48497 );
buf ( n395936 , n48498 );
buf ( n395937 , n395936 );
xor ( n48501 , n48473 , n395937 );
buf ( n395939 , n48501 );
buf ( n395940 , n395939 );
xor ( n48504 , n48432 , n395940 );
buf ( n395942 , n48504 );
buf ( n395943 , n395942 );
xor ( n48507 , n48336 , n395943 );
buf ( n395945 , n48507 );
buf ( n395946 , n395945 );
xor ( n48510 , n395658 , n395946 );
xor ( n48511 , n388124 , n388206 );
and ( n48512 , n48511 , n388533 );
and ( n48513 , n388124 , n388206 );
or ( n48514 , n48512 , n48513 );
buf ( n395952 , n48514 );
buf ( n395953 , n395952 );
not ( n48517 , n388809 );
buf ( n395955 , n385502 );
not ( n48519 , n395955 );
buf ( n395957 , n388757 );
nand ( n48521 , n48519 , n395957 );
buf ( n395959 , n48521 );
nand ( n48523 , n388760 , n388113 );
nand ( n48524 , n395959 , n48523 );
not ( n48525 , n48524 );
or ( n48526 , n48517 , n48525 );
buf ( n395964 , n391833 );
buf ( n395965 , n388746 );
nand ( n48529 , n395964 , n395965 );
buf ( n395967 , n48529 );
nand ( n48531 , n48526 , n395967 );
not ( n48532 , n44384 );
not ( n48533 , n389125 );
or ( n48534 , n48532 , n48533 );
buf ( n395972 , n24050 );
not ( n48536 , n395972 );
buf ( n395974 , n389525 );
not ( n48538 , n395974 );
or ( n48539 , n48536 , n48538 );
buf ( n395977 , n384741 );
buf ( n395978 , n389075 );
nand ( n48542 , n395977 , n395978 );
buf ( n395980 , n48542 );
buf ( n395981 , n395980 );
nand ( n48545 , n48539 , n395981 );
buf ( n395983 , n48545 );
buf ( n395984 , n395983 );
buf ( n395985 , n41565 );
nand ( n48549 , n395984 , n395985 );
buf ( n395987 , n48549 );
nand ( n48551 , n48534 , n395987 );
xor ( n48552 , n48531 , n48551 );
not ( n48553 , n391080 );
not ( n48554 , n391728 );
or ( n48555 , n48553 , n48554 );
not ( n48556 , n42925 );
buf ( n395994 , n24074 );
not ( n48558 , n395994 );
buf ( n395996 , n385774 );
not ( n48560 , n395996 );
or ( n48561 , n48558 , n48560 );
buf ( n395999 , n38227 );
buf ( n396000 , n24073 );
nand ( n48564 , n395999 , n396000 );
buf ( n396002 , n48564 );
buf ( n396003 , n396002 );
nand ( n48567 , n48561 , n396003 );
buf ( n396005 , n48567 );
nand ( n48569 , n48556 , n396005 );
nand ( n48570 , n48555 , n48569 );
xor ( n48571 , n48552 , n48570 );
buf ( n396009 , n48571 );
xor ( n48573 , n395953 , n396009 );
xor ( n48574 , n390054 , n390079 );
and ( n48575 , n48574 , n390086 );
and ( n48576 , n390054 , n390079 );
or ( n48577 , n48575 , n48576 );
buf ( n396015 , n48577 );
buf ( n396016 , n396015 );
xor ( n48580 , n48573 , n396016 );
buf ( n396018 , n48580 );
buf ( n396019 , n396018 );
xor ( n48583 , n48510 , n396019 );
buf ( n396021 , n48583 );
not ( n48585 , n396021 );
xor ( n48586 , n48213 , n48585 );
xor ( n48587 , n388536 , n388884 );
and ( n48588 , n48587 , n389218 );
and ( n48589 , n388536 , n388884 );
or ( n48590 , n48588 , n48589 );
buf ( n396028 , n48590 );
buf ( n396029 , n396028 );
xor ( n48593 , n390048 , n390089 );
and ( n48594 , n48593 , n390323 );
and ( n48595 , n390048 , n390089 );
or ( n48596 , n48594 , n48595 );
buf ( n396034 , n48596 );
buf ( n396035 , n396034 );
xor ( n48599 , n396029 , n396035 );
buf ( n396037 , n390239 );
not ( n48601 , n396037 );
buf ( n396039 , n390245 );
not ( n48603 , n396039 );
or ( n48604 , n48601 , n48603 );
buf ( n396042 , n390236 );
not ( n48606 , n396042 );
buf ( n396044 , n390208 );
not ( n48608 , n396044 );
or ( n48609 , n48606 , n48608 );
buf ( n396047 , n390318 );
nand ( n48611 , n48609 , n396047 );
buf ( n396049 , n48611 );
buf ( n396050 , n396049 );
nand ( n48614 , n48604 , n396050 );
buf ( n396052 , n48614 );
buf ( n396053 , n396052 );
nand ( n48617 , n390137 , n42630 , n42633 );
not ( n48618 , n48617 );
not ( n48619 , n390155 );
or ( n48620 , n48618 , n48619 );
not ( n48621 , n42633 );
not ( n48622 , n42630 );
or ( n48623 , n48621 , n48622 );
not ( n48624 , n390137 );
nand ( n48625 , n48623 , n48624 );
nand ( n48626 , n48620 , n48625 );
buf ( n396064 , n48626 );
xor ( n48628 , n396053 , n396064 );
buf ( n396066 , n388141 );
not ( n48630 , n396066 );
buf ( n396068 , n388160 );
not ( n48632 , n396068 );
buf ( n396070 , n383575 );
not ( n48634 , n396070 );
or ( n48635 , n48632 , n48634 );
nand ( n48636 , n39051 , n388157 );
buf ( n396074 , n48636 );
nand ( n48638 , n48635 , n396074 );
buf ( n396076 , n48638 );
buf ( n396077 , n396076 );
not ( n48641 , n396077 );
or ( n48642 , n48630 , n48641 );
buf ( n396080 , n388172 );
buf ( n396081 , n40701 );
nand ( n48645 , n396080 , n396081 );
buf ( n396083 , n48645 );
buf ( n396084 , n396083 );
nand ( n48648 , n48642 , n396084 );
buf ( n396086 , n48648 );
buf ( n396087 , n396086 );
xor ( n48651 , n48628 , n396087 );
buf ( n396089 , n48651 );
buf ( n396090 , n396089 );
buf ( n396091 , n390103 );
not ( n48655 , n396091 );
buf ( n396093 , n390321 );
not ( n48657 , n396093 );
or ( n48658 , n48655 , n48657 );
buf ( n396096 , n390166 );
nand ( n48660 , n48658 , n396096 );
buf ( n396098 , n48660 );
buf ( n396099 , n396098 );
buf ( n396100 , n390321 );
buf ( n396101 , n390103 );
or ( n48665 , n396100 , n396101 );
buf ( n396103 , n48665 );
buf ( n396104 , n396103 );
nand ( n48668 , n396099 , n396104 );
buf ( n396106 , n48668 );
buf ( n396107 , n396106 );
xor ( n48671 , n396090 , n396107 );
xor ( n48672 , n390254 , n390288 );
and ( n48673 , n48672 , n390316 );
and ( n48674 , n390254 , n390288 );
or ( n48675 , n48673 , n48674 );
buf ( n396113 , n48675 );
buf ( n396114 , n396113 );
buf ( n396115 , n385479 );
not ( n48679 , n396115 );
buf ( n396117 , n390185 );
not ( n48681 , n396117 );
or ( n48682 , n48679 , n48681 );
buf ( n396120 , n385494 );
not ( n48684 , n396120 );
buf ( n396122 , n386012 );
not ( n48686 , n396122 );
or ( n48687 , n48684 , n48686 );
buf ( n396125 , n38472 );
buf ( n396126 , n385491 );
nand ( n48690 , n396125 , n396126 );
buf ( n396128 , n48690 );
buf ( n396129 , n396128 );
nand ( n48693 , n48687 , n396129 );
buf ( n396131 , n48693 );
buf ( n396132 , n396131 );
buf ( n396133 , n41447 );
nand ( n48697 , n396132 , n396133 );
buf ( n396135 , n48697 );
buf ( n396136 , n396135 );
nand ( n48700 , n48682 , n396136 );
buf ( n396138 , n48700 );
buf ( n396139 , n396138 );
xor ( n48703 , n396114 , n396139 );
xor ( n48704 , n391759 , n391776 );
and ( n48705 , n48704 , n391805 );
and ( n48706 , n391759 , n391776 );
or ( n48707 , n48705 , n48706 );
buf ( n396145 , n48707 );
buf ( n396146 , n396145 );
xor ( n48710 , n48703 , n396146 );
buf ( n396148 , n48710 );
buf ( n396149 , n388833 );
not ( n48713 , n396149 );
and ( n48714 , n41342 , n382924 );
not ( n48715 , n41342 );
and ( n48716 , n48715 , n382921 );
or ( n48717 , n48714 , n48716 );
buf ( n396155 , n48717 );
not ( n48719 , n396155 );
or ( n48720 , n48713 , n48719 );
buf ( n396158 , n42617 );
buf ( n396159 , n388872 );
nand ( n48723 , n396158 , n396159 );
buf ( n396161 , n48723 );
buf ( n396162 , n396161 );
nand ( n48726 , n48720 , n396162 );
buf ( n396164 , n48726 );
xor ( n48728 , n396148 , n396164 );
xor ( n48729 , n391739 , n391808 );
and ( n48730 , n48729 , n391815 );
and ( n48731 , n391739 , n391808 );
or ( n48732 , n48730 , n48731 );
buf ( n396170 , n48732 );
xor ( n48734 , n48728 , n396170 );
buf ( n396172 , n48734 );
xor ( n48736 , n48671 , n396172 );
buf ( n396174 , n48736 );
buf ( n396175 , n396174 );
xor ( n48739 , n48599 , n396175 );
buf ( n396177 , n48739 );
xnor ( n48741 , n48586 , n396177 );
buf ( n396179 , n48741 );
xnor ( n48743 , n48209 , n396179 );
buf ( n396181 , n48743 );
buf ( n396182 , n396181 );
nand ( n48746 , n48193 , n396182 );
buf ( n396184 , n48746 );
buf ( n396185 , n396184 );
and ( n48749 , n393719 , n394597 , n395624 , n396185 );
buf ( n396187 , n48749 );
xor ( n48751 , n48126 , n48163 );
buf ( n48752 , n48139 );
xnor ( n48753 , n48751 , n48752 );
buf ( n396191 , n395056 );
not ( n48755 , n396191 );
buf ( n396193 , n394643 );
not ( n48757 , n396193 );
or ( n48758 , n48755 , n48757 );
buf ( n396196 , n394640 );
buf ( n396197 , n395056 );
not ( n48761 , n396197 );
buf ( n396199 , n48761 );
buf ( n396200 , n396199 );
nand ( n48764 , n396196 , n396200 );
buf ( n396202 , n48764 );
buf ( n396203 , n396202 );
nand ( n48767 , n48758 , n396203 );
buf ( n396205 , n48767 );
and ( n48769 , n396205 , n394650 );
not ( n48770 , n396205 );
and ( n48771 , n48770 , n394653 );
nor ( n48772 , n48769 , n48771 );
not ( n48773 , n46402 );
not ( n48774 , n393849 );
not ( n48775 , n46368 );
or ( n48776 , n48774 , n48775 );
not ( n48777 , n393849 );
nand ( n48778 , n48777 , n46369 );
nand ( n48779 , n48776 , n48778 );
xor ( n48780 , n48773 , n48779 );
buf ( n396218 , n48780 );
not ( n48782 , n396218 );
buf ( n396220 , n48782 );
not ( n48784 , n396220 );
buf ( n396222 , n392884 );
not ( n48786 , n396222 );
buf ( n396224 , n37402 );
not ( n48788 , n396224 );
or ( n48789 , n48786 , n48788 );
buf ( n396227 , n35435 );
buf ( n396228 , n392887 );
nand ( n48792 , n396227 , n396228 );
buf ( n396230 , n48792 );
buf ( n396231 , n396230 );
nand ( n48795 , n48789 , n396231 );
buf ( n396233 , n48795 );
buf ( n396234 , n396233 );
not ( n48798 , n396234 );
buf ( n396236 , n390629 );
not ( n48800 , n396236 );
or ( n48801 , n48798 , n48800 );
buf ( n396239 , n383134 );
not ( n48803 , n396239 );
buf ( n396241 , n394741 );
nand ( n48805 , n48803 , n396241 );
buf ( n396243 , n48805 );
buf ( n396244 , n396243 );
nand ( n48808 , n48801 , n396244 );
buf ( n396246 , n48808 );
buf ( n396247 , n396246 );
not ( n48811 , n396247 );
buf ( n396249 , n389359 );
not ( n48813 , n396249 );
buf ( n396251 , n388576 );
not ( n48815 , n396251 );
or ( n48816 , n48813 , n48815 );
buf ( n396254 , n388556 );
buf ( n396255 , n389356 );
nand ( n48819 , n396254 , n396255 );
buf ( n396257 , n48819 );
buf ( n396258 , n396257 );
nand ( n48822 , n48816 , n396258 );
buf ( n396260 , n48822 );
buf ( n396261 , n396260 );
not ( n48825 , n396261 );
buf ( n396263 , n391649 );
not ( n48827 , n396263 );
or ( n48828 , n48825 , n48827 );
not ( n48829 , n383403 );
nand ( n48830 , n48829 , n394528 );
buf ( n396268 , n48830 );
nand ( n48832 , n48828 , n396268 );
buf ( n396270 , n48832 );
buf ( n396271 , n396270 );
not ( n48835 , n396271 );
or ( n48836 , n48811 , n48835 );
buf ( n396274 , n396270 );
buf ( n396275 , n396246 );
or ( n48839 , n396274 , n396275 );
xor ( n48840 , n393537 , n394721 );
xnor ( n48841 , n48840 , n394712 );
buf ( n396279 , n48841 );
nand ( n48843 , n48839 , n396279 );
buf ( n396281 , n48843 );
buf ( n396282 , n396281 );
nand ( n48846 , n48836 , n396282 );
buf ( n396284 , n48846 );
buf ( n396285 , n396284 );
xor ( n48849 , n394728 , n394755 );
xor ( n48850 , n48849 , n394777 );
buf ( n396288 , n48850 );
buf ( n396289 , n396288 );
xor ( n48853 , n396285 , n396289 );
buf ( n396291 , n388102 );
not ( n48855 , n396291 );
buf ( n396293 , n389420 );
not ( n48857 , n396293 );
or ( n48858 , n48855 , n48857 );
buf ( n396296 , n36897 );
buf ( n48860 , n396296 );
buf ( n396298 , n48860 );
buf ( n396299 , n396298 );
buf ( n396300 , n388105 );
nand ( n48864 , n396299 , n396300 );
buf ( n396302 , n48864 );
buf ( n396303 , n396302 );
nand ( n48867 , n48858 , n396303 );
buf ( n396305 , n48867 );
not ( n48869 , n396305 );
not ( n48870 , n43286 );
or ( n48871 , n48869 , n48870 );
or ( n48872 , n395016 , n388071 );
nand ( n48873 , n48871 , n48872 );
buf ( n396311 , n48873 );
and ( n48875 , n48853 , n396311 );
and ( n48876 , n396285 , n396289 );
or ( n48877 , n48875 , n48876 );
buf ( n396315 , n48877 );
not ( n48879 , n396315 );
or ( n48880 , n48784 , n48879 );
buf ( n396318 , n48780 );
not ( n48882 , n396318 );
buf ( n396320 , n396315 );
not ( n48884 , n396320 );
buf ( n396322 , n48884 );
buf ( n396323 , n396322 );
not ( n48887 , n396323 );
or ( n48888 , n48882 , n48887 );
buf ( n396326 , n394903 );
buf ( n396327 , n394923 );
xor ( n48891 , n396326 , n396327 );
buf ( n396329 , n47435 );
xor ( n48893 , n48891 , n396329 );
buf ( n396331 , n48893 );
buf ( n396332 , n396331 );
not ( n48896 , n396332 );
buf ( n396334 , n48896 );
buf ( n396335 , n396334 );
not ( n48899 , n396335 );
buf ( n396337 , n388872 );
not ( n48901 , n396337 );
buf ( n396339 , n41342 );
not ( n48903 , n396339 );
buf ( n396341 , n389289 );
not ( n48905 , n396341 );
or ( n48906 , n48903 , n48905 );
buf ( n396344 , n36709 );
buf ( n396345 , n45897 );
nand ( n48909 , n396344 , n396345 );
buf ( n396347 , n48909 );
buf ( n396348 , n396347 );
nand ( n48912 , n48906 , n396348 );
buf ( n396350 , n48912 );
buf ( n396351 , n396350 );
not ( n48915 , n396351 );
or ( n48916 , n48901 , n48915 );
buf ( n396354 , n394913 );
not ( n48918 , n396354 );
buf ( n396356 , n388833 );
nand ( n48920 , n48918 , n396356 );
buf ( n396358 , n48920 );
buf ( n396359 , n396358 );
nand ( n48923 , n48916 , n396359 );
buf ( n396361 , n48923 );
buf ( n396362 , n396361 );
buf ( n396363 , n40901 );
buf ( n396364 , n394800 );
nand ( n48928 , n396363 , n396364 );
buf ( n396366 , n48928 );
buf ( n396367 , n388511 );
buf ( n396368 , n40885 );
and ( n48932 , n396367 , n396368 );
not ( n48933 , n396367 );
buf ( n396371 , n36810 );
not ( n48935 , n396371 );
buf ( n396373 , n48935 );
buf ( n396374 , n396373 );
and ( n48938 , n48933 , n396374 );
nor ( n48939 , n48932 , n48938 );
buf ( n396377 , n48939 );
not ( n48941 , n396377 );
nand ( n48942 , n48941 , n40858 );
nand ( n48943 , n396366 , n48942 );
buf ( n396381 , n48943 );
buf ( n396382 , n388230 );
not ( n48946 , n396382 );
buf ( n396384 , n47256 );
not ( n48948 , n396384 );
or ( n48949 , n48946 , n48948 );
buf ( n396387 , n388242 );
buf ( n396388 , n36396 );
nand ( n48952 , n396387 , n396388 );
buf ( n396390 , n48952 );
buf ( n396391 , n396390 );
nand ( n48955 , n48949 , n396391 );
buf ( n396393 , n48955 );
not ( n48957 , n396393 );
not ( n48958 , n390832 );
or ( n48959 , n48957 , n48958 );
buf ( n396397 , n394705 );
not ( n48961 , n396397 );
buf ( n396399 , n388346 );
nand ( n48963 , n48961 , n396399 );
buf ( n396401 , n48963 );
nand ( n48965 , n48959 , n396401 );
buf ( n396403 , n48965 );
or ( n48967 , n396381 , n396403 );
buf ( n396405 , n389744 );
not ( n48969 , n396405 );
buf ( n396407 , n392611 );
not ( n48971 , n396407 );
buf ( n396409 , n389753 );
not ( n48973 , n396409 );
or ( n48974 , n48971 , n48973 );
buf ( n396412 , n389997 );
buf ( n396413 , n392620 );
nand ( n48977 , n396412 , n396413 );
buf ( n396415 , n48977 );
buf ( n396416 , n396415 );
nand ( n48980 , n48974 , n396416 );
buf ( n396418 , n48980 );
buf ( n396419 , n396418 );
not ( n48983 , n396419 );
or ( n48984 , n48969 , n48983 );
buf ( n396422 , n389328 );
buf ( n396423 , n395519 );
nand ( n48987 , n396422 , n396423 );
buf ( n396425 , n48987 );
buf ( n396426 , n396425 );
nand ( n48990 , n48984 , n396426 );
buf ( n396428 , n48990 );
buf ( n396429 , n396428 );
nand ( n48993 , n48967 , n396429 );
buf ( n396431 , n48993 );
buf ( n396432 , n396431 );
not ( n48996 , n48942 );
not ( n48997 , n396366 );
or ( n48998 , n48996 , n48997 );
not ( n48999 , n396393 );
not ( n49000 , n390832 );
or ( n49001 , n48999 , n49000 );
nand ( n49002 , n49001 , n396401 );
nand ( n49003 , n48998 , n49002 );
buf ( n396441 , n49003 );
nand ( n49005 , n396432 , n396441 );
buf ( n396443 , n49005 );
buf ( n396444 , n396443 );
xor ( n49008 , n396362 , n396444 );
buf ( n396446 , n389162 );
not ( n49010 , n396446 );
buf ( n396448 , n395413 );
not ( n49012 , n396448 );
or ( n49013 , n49010 , n49012 );
buf ( n396451 , n41671 );
not ( n49015 , n396451 );
buf ( n396453 , n384208 );
not ( n49017 , n396453 );
or ( n49018 , n49015 , n49017 );
buf ( n396456 , n390119 );
buf ( n396457 , n41670 );
nand ( n49021 , n396456 , n396457 );
buf ( n396459 , n49021 );
buf ( n396460 , n396459 );
nand ( n49024 , n49018 , n396460 );
buf ( n396462 , n49024 );
buf ( n396463 , n396462 );
buf ( n396464 , n41711 );
nand ( n49028 , n396463 , n396464 );
buf ( n396466 , n49028 );
buf ( n396467 , n396466 );
nand ( n49031 , n49013 , n396467 );
buf ( n396469 , n49031 );
buf ( n396470 , n396469 );
and ( n49034 , n49008 , n396470 );
and ( n49035 , n396362 , n396444 );
or ( n49036 , n49034 , n49035 );
buf ( n396474 , n49036 );
buf ( n396475 , n396474 );
not ( n49039 , n396475 );
or ( n49040 , n48899 , n49039 );
buf ( n396478 , n396331 );
not ( n49042 , n396478 );
buf ( n396480 , n396474 );
not ( n49044 , n396480 );
buf ( n396482 , n49044 );
buf ( n396483 , n396482 );
not ( n49047 , n396483 );
or ( n49048 , n49042 , n49047 );
xor ( n49049 , n394869 , n394810 );
xor ( n49050 , n49049 , n394836 );
buf ( n396488 , n49050 );
not ( n49052 , n396488 );
buf ( n396490 , n43286 );
not ( n49054 , n396490 );
buf ( n396492 , n388105 );
not ( n49056 , n396492 );
buf ( n396494 , n389435 );
not ( n49058 , n396494 );
or ( n49059 , n49056 , n49058 );
buf ( n396497 , n394463 );
not ( n49061 , n396497 );
buf ( n396499 , n388102 );
nand ( n49063 , n49061 , n396499 );
buf ( n396501 , n49063 );
buf ( n396502 , n396501 );
nand ( n49066 , n49059 , n396502 );
buf ( n396504 , n49066 );
buf ( n396505 , n396504 );
not ( n49069 , n396505 );
or ( n49070 , n49054 , n49069 );
buf ( n396508 , n396305 );
buf ( n396509 , n390362 );
nand ( n49073 , n396508 , n396509 );
buf ( n396511 , n49073 );
buf ( n396512 , n396511 );
nand ( n49076 , n49070 , n396512 );
buf ( n396514 , n49076 );
buf ( n396515 , n396514 );
not ( n49079 , n396515 );
or ( n49080 , n49052 , n49079 );
buf ( n396518 , n396514 );
buf ( n396519 , n49050 );
or ( n49083 , n396518 , n396519 );
buf ( n396521 , n392788 );
not ( n49085 , n396521 );
buf ( n396523 , n394859 );
not ( n49087 , n396523 );
or ( n49088 , n49085 , n49087 );
buf ( n396526 , n390432 );
buf ( n396527 , n24072 );
not ( n49091 , n396527 );
buf ( n396529 , n38630 );
not ( n49093 , n396529 );
or ( n49094 , n49091 , n49093 );
buf ( n396532 , n28159 );
not ( n49096 , n396532 );
buf ( n396534 , n49096 );
buf ( n396535 , n396534 );
not ( n49099 , n396535 );
buf ( n396537 , n49099 );
buf ( n396538 , n396537 );
not ( n49102 , n47412 );
buf ( n396540 , n49102 );
nand ( n49104 , n396538 , n396540 );
buf ( n396542 , n49104 );
buf ( n396543 , n396542 );
nand ( n49107 , n49094 , n396543 );
buf ( n396545 , n49107 );
buf ( n396546 , n396545 );
nand ( n49110 , n396526 , n396546 );
buf ( n396548 , n49110 );
buf ( n396549 , n396548 );
nand ( n49113 , n49088 , n396549 );
buf ( n396551 , n49113 );
buf ( n396552 , n396551 );
and ( n49116 , n24783 , n24785 , n24788 , n24789 );
not ( n49117 , n49116 );
buf ( n396555 , n49117 );
not ( n49119 , n396555 );
buf ( n396557 , n384096 );
not ( n49121 , n396557 );
or ( n49122 , n49119 , n49121 );
buf ( n396560 , n385328 );
not ( n49124 , n49117 );
buf ( n396562 , n49124 );
nand ( n49126 , n396560 , n396562 );
buf ( n396564 , n49126 );
buf ( n396565 , n396564 );
nand ( n49129 , n49122 , n396565 );
buf ( n396567 , n49129 );
buf ( n396568 , n382938 );
buf ( n396569 , n394829 );
nand ( n49138 , n396568 , n396569 );
buf ( n396571 , n49138 );
buf ( n396572 , n396571 );
nand ( n49141 , C1 , n396572 );
buf ( n396574 , n49141 );
buf ( n396575 , n396574 );
xor ( n49144 , n396552 , n396575 );
buf ( n396577 , n388646 );
not ( n49146 , n396577 );
buf ( n396579 , n385488 );
not ( n49148 , n396579 );
or ( n49149 , n49146 , n49148 );
buf ( n396582 , n385473 );
buf ( n396583 , n388643 );
not ( n49152 , n396583 );
buf ( n396585 , n49152 );
buf ( n396586 , n396585 );
nand ( n49155 , n396582 , n396586 );
buf ( n396588 , n49155 );
buf ( n396589 , n396588 );
nand ( n49158 , n49149 , n396589 );
buf ( n396591 , n49158 );
buf ( n396592 , n396591 );
not ( n49161 , n396592 );
buf ( n396594 , n393544 );
not ( n49163 , n396594 );
or ( n49164 , n49161 , n49163 );
buf ( n396597 , n395449 );
not ( n49166 , n37923 );
buf ( n396599 , n49166 );
nand ( n49168 , n396597 , n396599 );
buf ( n396601 , n49168 );
buf ( n396602 , n396601 );
nand ( n49171 , n49164 , n396602 );
buf ( n396604 , n49171 );
buf ( n396605 , n396604 );
not ( n49174 , n396605 );
buf ( n396607 , n41577 );
not ( n49176 , n396607 );
buf ( n396609 , n40831 );
not ( n49178 , n396609 );
or ( n49179 , n49176 , n49178 );
buf ( n396612 , n27196 );
buf ( n396613 , n45391 );
nand ( n49182 , n396612 , n396613 );
buf ( n396615 , n49182 );
buf ( n396616 , n396615 );
nand ( n49185 , n49179 , n396616 );
buf ( n396618 , n49185 );
buf ( n396619 , n396618 );
buf ( n396620 , n389116 );
not ( n49189 , n396620 );
buf ( n396622 , n49189 );
buf ( n396623 , n396622 );
and ( n49192 , n396619 , n396623 );
buf ( n396625 , n395217 );
buf ( n396626 , n41564 );
nor ( n49195 , n396625 , n396626 );
buf ( n396628 , n49195 );
buf ( n396629 , n396628 );
nor ( n49198 , n49192 , n396629 );
buf ( n396631 , n49198 );
buf ( n396632 , n396631 );
not ( n49201 , n396632 );
buf ( n396634 , n49201 );
buf ( n396635 , n396634 );
not ( n49204 , n396635 );
or ( n49205 , n49174 , n49204 );
buf ( n396638 , n396604 );
not ( n49207 , n396638 );
buf ( n396640 , n49207 );
buf ( n396641 , n396640 );
not ( n49210 , n396641 );
buf ( n396643 , n396631 );
not ( n49212 , n396643 );
or ( n49213 , n49210 , n49212 );
not ( n49214 , n37338 );
buf ( n396647 , n388905 );
not ( n49216 , n396647 );
buf ( n396649 , n388566 );
not ( n49218 , n396649 );
and ( n49219 , n49216 , n49218 );
buf ( n396652 , n395478 );
buf ( n396653 , n388566 );
and ( n49222 , n396652 , n396653 );
nor ( n49223 , n49219 , n49222 );
buf ( n396656 , n49223 );
not ( n49225 , n396656 );
not ( n49226 , n49225 );
or ( n49227 , n49214 , n49226 );
buf ( n396660 , n395488 );
not ( n49229 , n396660 );
buf ( n396662 , n37316 );
nand ( n49231 , n49229 , n396662 );
buf ( n396664 , n49231 );
nand ( n49233 , n49227 , n396664 );
buf ( n396666 , n49233 );
nand ( n49235 , n49213 , n396666 );
buf ( n396668 , n49235 );
buf ( n396669 , n396668 );
nand ( n49238 , n49205 , n396669 );
buf ( n396671 , n49238 );
buf ( n396672 , n396671 );
and ( n49241 , n49144 , n396672 );
and ( n49242 , n396552 , n396575 );
or ( n49243 , n49241 , n49242 );
buf ( n396676 , n49243 );
buf ( n396677 , n396676 );
nand ( n49246 , n49083 , n396677 );
buf ( n396679 , n49246 );
buf ( n396680 , n396679 );
nand ( n49249 , n49080 , n396680 );
buf ( n396682 , n49249 );
buf ( n396683 , n396682 );
nand ( n49252 , n49048 , n396683 );
buf ( n396685 , n49252 );
buf ( n396686 , n396685 );
nand ( n49255 , n49040 , n396686 );
buf ( n396688 , n49255 );
buf ( n396689 , n396688 );
nand ( n49258 , n48888 , n396689 );
buf ( n396691 , n49258 );
nand ( n49260 , n48880 , n396691 );
not ( n49261 , n49260 );
not ( n49262 , n395044 );
not ( n49263 , n394977 );
not ( n49264 , n394960 );
or ( n49265 , n49263 , n49264 );
or ( n49266 , n394977 , n394960 );
nand ( n49267 , n49265 , n49266 );
not ( n49268 , n49267 );
or ( n49269 , n49262 , n49268 );
or ( n49270 , n395044 , n49267 );
nand ( n49271 , n49269 , n49270 );
nand ( n49272 , n49261 , n49271 );
not ( n49273 , n49272 );
xor ( n49274 , n395082 , n395294 );
xor ( n49275 , n49274 , n395560 );
buf ( n396708 , n49275 );
not ( n49277 , n396708 );
or ( n49278 , n49273 , n49277 );
not ( n49279 , n49271 );
nand ( n49280 , n49279 , n49260 );
nand ( n49281 , n49278 , n49280 );
and ( n396714 , n48772 , n49281 );
not ( n49283 , n48772 );
buf ( n396716 , n49281 );
not ( n49285 , n396716 );
buf ( n396718 , n49285 );
and ( n49287 , n49283 , n396718 );
nor ( n49288 , n396714 , n49287 );
xor ( n49289 , n395004 , n395026 );
xnor ( n49290 , n49289 , n395038 );
not ( n49291 , n49290 );
xor ( n49292 , n394781 , n394943 );
xnor ( n49293 , n49292 , n47510 );
buf ( n396726 , n49293 );
buf ( n49295 , n396726 );
buf ( n396728 , n49295 );
not ( n49297 , n396728 );
or ( n49298 , n49291 , n49297 );
buf ( n396731 , n396728 );
buf ( n396732 , n49290 );
or ( n49301 , n396731 , n396732 );
xor ( n49302 , n395120 , n395257 );
xor ( n49303 , n49302 , n395283 );
buf ( n396736 , n49303 );
not ( n49305 , n396736 );
buf ( n396738 , n45260 );
not ( n49307 , n396738 );
buf ( n396740 , n392247 );
not ( n49309 , n396740 );
buf ( n396742 , n386561 );
not ( n49311 , n396742 );
or ( n49312 , n49309 , n49311 );
buf ( n396745 , n382921 );
buf ( n396746 , n392244 );
nand ( n49315 , n396745 , n396746 );
buf ( n396748 , n49315 );
buf ( n396749 , n396748 );
nand ( n49318 , n49312 , n396749 );
buf ( n396751 , n49318 );
buf ( n396752 , n396751 );
not ( n49321 , n396752 );
or ( n49322 , n49307 , n49321 );
buf ( n396755 , n392224 );
not ( n49324 , n396755 );
buf ( n396757 , n394994 );
nand ( n49326 , n49324 , n396757 );
buf ( n396759 , n49326 );
buf ( n396760 , n396759 );
nand ( n49329 , n49322 , n396760 );
buf ( n396762 , n49329 );
buf ( n396763 , n43515 );
not ( n49332 , n396763 );
buf ( n396765 , n395101 );
not ( n49334 , n396765 );
or ( n49335 , n49332 , n49334 );
buf ( n396768 , n391027 );
not ( n49337 , n396768 );
buf ( n396770 , n37027 );
not ( n49339 , n396770 );
or ( n49340 , n49337 , n49339 );
buf ( n396773 , n383575 );
not ( n49342 , n396773 );
buf ( n396775 , n391024 );
nand ( n49344 , n49342 , n396775 );
buf ( n396777 , n49344 );
buf ( n396778 , n396777 );
nand ( n49347 , n49340 , n396778 );
buf ( n396780 , n49347 );
buf ( n396781 , n396780 );
buf ( n396782 , n43727 );
nand ( n49351 , n396781 , n396782 );
buf ( n396784 , n49351 );
buf ( n396785 , n396784 );
nand ( n49354 , n49335 , n396785 );
buf ( n396787 , n49354 );
or ( n49356 , n396762 , n396787 );
not ( n49357 , n49356 );
or ( n49358 , n49305 , n49357 );
buf ( n396791 , n396762 );
buf ( n396792 , n396787 );
nand ( n49361 , n396791 , n396792 );
buf ( n396794 , n49361 );
nand ( n49363 , n49358 , n396794 );
buf ( n396796 , n49363 );
nand ( n49365 , n49301 , n396796 );
buf ( n396798 , n49365 );
nand ( n49367 , n49298 , n396798 );
not ( n49368 , n49367 );
not ( n49369 , n395588 );
not ( n49370 , n395583 );
not ( n49371 , n49370 );
or ( n49372 , n49369 , n49371 );
nand ( n49373 , n395583 , n48150 );
nand ( n49374 , n49372 , n49373 );
xor ( n49375 , n48153 , n48155 );
and ( n49376 , n49374 , n49375 );
not ( n49377 , n49374 );
and ( n49378 , n49377 , n48159 );
nor ( n49379 , n49376 , n49378 );
not ( n49380 , n49379 );
not ( n49381 , n49380 );
or ( n49382 , n49368 , n49381 );
not ( n49383 , n49367 );
not ( n49384 , n49383 );
not ( n49385 , n49379 );
or ( n49386 , n49384 , n49385 );
buf ( n396819 , n395085 );
buf ( n396820 , n395111 );
xor ( n49389 , n396819 , n396820 );
buf ( n396822 , n395287 );
xor ( n49391 , n49389 , n396822 );
buf ( n396824 , n49391 );
buf ( n396825 , n396824 );
buf ( n396826 , n393825 );
not ( n49395 , n396826 );
buf ( n396828 , n393369 );
not ( n49397 , n396828 );
buf ( n396830 , n388771 );
not ( n49399 , n396830 );
or ( n49400 , n49397 , n49399 );
buf ( n396833 , n386418 );
buf ( n396834 , n393381 );
nand ( n49403 , n396833 , n396834 );
buf ( n396836 , n49403 );
buf ( n396837 , n396836 );
nand ( n49406 , n49400 , n396837 );
buf ( n396839 , n49406 );
buf ( n396840 , n396839 );
not ( n49409 , n396840 );
or ( n49410 , n49395 , n49409 );
buf ( n396843 , n395389 );
buf ( n396844 , n45954 );
nand ( n49413 , n396843 , n396844 );
buf ( n396846 , n49413 );
buf ( n396847 , n396846 );
nand ( n49416 , n49410 , n396847 );
buf ( n396849 , n49416 );
buf ( n396850 , n396849 );
not ( n49419 , n396850 );
xor ( n49420 , n395202 , n395226 );
xor ( n49421 , n49420 , n395246 );
buf ( n396854 , n49421 );
buf ( n396855 , n396854 );
not ( n49424 , n394210 );
not ( n49425 , n388235 );
or ( n49426 , n49424 , n49425 );
buf ( n396859 , n35435 );
buf ( n396860 , n394219 );
nand ( n49429 , n396859 , n396860 );
buf ( n396862 , n49429 );
nand ( n49431 , n49426 , n396862 );
buf ( n396864 , n49431 );
not ( n49433 , n396864 );
buf ( n396866 , n383014 );
not ( n49435 , n396866 );
buf ( n396868 , n49435 );
buf ( n396869 , n396868 );
not ( n49438 , n396869 );
or ( n49439 , n49433 , n49438 );
buf ( n396872 , n390476 );
buf ( n396873 , n396233 );
nand ( n49442 , n396872 , n396873 );
buf ( n396875 , n49442 );
buf ( n396876 , n396875 );
nand ( n49445 , n49439 , n396876 );
buf ( n396878 , n49445 );
buf ( n396879 , n396878 );
xor ( n49448 , n396855 , n396879 );
buf ( n396881 , n388833 );
not ( n49450 , n396881 );
buf ( n396883 , n396350 );
not ( n49452 , n396883 );
or ( n49453 , n49450 , n49452 );
buf ( n396886 , n41342 );
not ( n49455 , n396886 );
buf ( n396888 , n389485 );
not ( n49457 , n396888 );
or ( n49458 , n49455 , n49457 );
buf ( n396891 , n390657 );
buf ( n396892 , n45897 );
nand ( n49461 , n396891 , n396892 );
buf ( n396894 , n49461 );
buf ( n396895 , n396894 );
nand ( n49464 , n49458 , n396895 );
buf ( n396897 , n49464 );
buf ( n396898 , n396897 );
buf ( n396899 , n388872 );
nand ( n49468 , n396898 , n396899 );
buf ( n396901 , n49468 );
buf ( n396902 , n396901 );
nand ( n49471 , n49453 , n396902 );
buf ( n396904 , n49471 );
buf ( n396905 , n396904 );
and ( n49474 , n49448 , n396905 );
and ( n49475 , n396855 , n396879 );
or ( n49476 , n49474 , n49475 );
buf ( n396909 , n49476 );
buf ( n396910 , n396909 );
not ( n49479 , n396910 );
or ( n49480 , n49419 , n49479 );
buf ( n396913 , n396849 );
buf ( n396914 , n396909 );
or ( n49483 , n396913 , n396914 );
xor ( n49484 , n48841 , n396246 );
xor ( n49485 , n49484 , n396270 );
buf ( n396918 , n49485 );
nand ( n49487 , n49483 , n396918 );
buf ( n396920 , n49487 );
buf ( n396921 , n396920 );
nand ( n49490 , n49480 , n396921 );
buf ( n396923 , n49490 );
not ( n49492 , n396923 );
buf ( n396925 , n395362 );
not ( n49494 , n396925 );
buf ( n396927 , n395321 );
not ( n49496 , n396927 );
or ( n49497 , n49494 , n49496 );
buf ( n396930 , n47863 );
not ( n49499 , n396930 );
buf ( n396932 , n390351 );
not ( n49501 , n396932 );
or ( n49502 , n49499 , n49501 );
buf ( n396935 , n382545 );
buf ( n396936 , n395312 );
nand ( n49505 , n396935 , n396936 );
buf ( n396938 , n49505 );
buf ( n396939 , n396938 );
nand ( n49508 , n49502 , n396939 );
buf ( n396941 , n49508 );
buf ( n396942 , n396941 );
buf ( n396943 , n395349 );
nand ( n49512 , n396942 , n396943 );
buf ( n396945 , n49512 );
buf ( n396946 , n396945 );
nand ( n49515 , n49497 , n396946 );
buf ( n396948 , n49515 );
not ( n49517 , n396948 );
buf ( n396950 , n388746 );
not ( n49519 , n396950 );
buf ( n396952 , n388760 );
not ( n49521 , n396952 );
buf ( n396954 , n390373 );
not ( n49523 , n396954 );
or ( n49524 , n49521 , n49523 );
not ( n49525 , n37679 );
buf ( n396958 , n49525 );
buf ( n396959 , n388757 );
nand ( n49528 , n396958 , n396959 );
buf ( n396961 , n49528 );
buf ( n396962 , n396961 );
nand ( n49531 , n49524 , n396962 );
buf ( n396964 , n49531 );
buf ( n396965 , n396964 );
not ( n49534 , n396965 );
or ( n49535 , n49519 , n49534 );
buf ( n396968 , n395275 );
buf ( n396969 , n388809 );
nand ( n49538 , n396968 , n396969 );
buf ( n396971 , n49538 );
buf ( n396972 , n396971 );
nand ( n49541 , n49535 , n396972 );
buf ( n396974 , n49541 );
buf ( n396975 , n396974 );
not ( n49544 , n396975 );
buf ( n396977 , n49544 );
nand ( n49546 , n49517 , n396977 );
not ( n49547 , n49546 );
buf ( n396980 , n389341 );
buf ( n396981 , n388556 );
and ( n49550 , n396980 , n396981 );
not ( n49551 , n396980 );
buf ( n396984 , n388576 );
and ( n49553 , n49551 , n396984 );
nor ( n49554 , n49550 , n49553 );
buf ( n396987 , n49554 );
buf ( n396988 , n396987 );
not ( n49557 , n396988 );
buf ( n396990 , n391270 );
not ( n49559 , n396990 );
or ( n49560 , n49557 , n49559 );
buf ( n396993 , n391170 );
buf ( n396994 , n396260 );
nand ( n49563 , n396993 , n396994 );
buf ( n396996 , n49563 );
buf ( n396997 , n396996 );
nand ( n49566 , n49560 , n396997 );
buf ( n396999 , n49566 );
not ( n49568 , n396999 );
not ( n49569 , n49568 );
buf ( n397002 , n49569 );
not ( n49571 , n397002 );
buf ( n397004 , n42073 );
not ( n49573 , n397004 );
buf ( n397006 , n394392 );
not ( n49575 , n397006 );
or ( n49576 , n49573 , n49575 );
buf ( n397009 , n37037 );
buf ( n397010 , n42074 );
nand ( n49579 , n397009 , n397010 );
buf ( n397012 , n49579 );
buf ( n397013 , n397012 );
nand ( n49582 , n49576 , n397013 );
buf ( n397015 , n49582 );
buf ( n397016 , n397015 );
not ( n49585 , n397016 );
buf ( n397018 , n389880 );
not ( n49587 , n397018 );
or ( n49588 , n49585 , n49587 );
buf ( n397021 , n395132 );
buf ( n397022 , n391638 );
nand ( n49591 , n397021 , n397022 );
buf ( n397024 , n49591 );
buf ( n397025 , n397024 );
nand ( n49594 , n49588 , n397025 );
buf ( n397027 , n49594 );
buf ( n397028 , n397027 );
not ( n49597 , n397028 );
or ( n49598 , n49571 , n49597 );
buf ( n397031 , n397027 );
not ( n49600 , n397031 );
buf ( n397033 , n49600 );
buf ( n397034 , n397033 );
not ( n49603 , n397034 );
buf ( n397036 , n49568 );
not ( n49605 , n397036 );
or ( n49606 , n49603 , n49605 );
buf ( n397039 , n40990 );
not ( n49608 , n397039 );
buf ( n397041 , n40890 );
not ( n49610 , n397041 );
or ( n49611 , n49608 , n49610 );
buf ( n397044 , n40885 );
buf ( n397045 , n390460 );
nand ( n49614 , n397044 , n397045 );
buf ( n397047 , n49614 );
buf ( n397048 , n397047 );
nand ( n49617 , n49611 , n397048 );
buf ( n397050 , n49617 );
buf ( n397051 , n397050 );
not ( n49620 , n397051 );
buf ( n397053 , n36801 );
not ( n49622 , n397053 );
or ( n49623 , n49620 , n49622 );
buf ( n397056 , n396377 );
not ( n49625 , n397056 );
buf ( n397058 , n392111 );
nand ( n49627 , n49625 , n397058 );
buf ( n397060 , n49627 );
buf ( n397061 , n397060 );
nand ( n49630 , n49623 , n397061 );
buf ( n397063 , n49630 );
not ( n49632 , n397063 );
not ( n49633 , n395199 );
not ( n49634 , n22982 );
buf ( n397067 , n40866 );
buf ( n49636 , n397067 );
buf ( n397069 , n49636 );
buf ( n397070 , n397069 );
not ( n49639 , n397070 );
buf ( n397072 , n49639 );
not ( n49641 , n397072 );
or ( n49642 , n49634 , n49641 );
buf ( n397075 , n46114 );
not ( n49644 , n397075 );
buf ( n397077 , n49644 );
buf ( n397078 , n397077 );
buf ( n397079 , n45102 );
nand ( n49648 , n397078 , n397079 );
buf ( n397081 , n49648 );
nand ( n49650 , n49642 , n397081 );
not ( n49651 , n49650 );
or ( n49652 , n49633 , n49651 );
buf ( n49653 , n37913 );
buf ( n397086 , n49653 );
not ( n49655 , n397086 );
buf ( n397088 , n45699 );
not ( n49657 , n397088 );
or ( n49658 , n49655 , n49657 );
buf ( n397091 , n388643 );
buf ( n49660 , n37913 );
not ( n49661 , n49660 );
buf ( n397094 , n49661 );
nand ( n49663 , n397091 , n397094 );
buf ( n397096 , n49663 );
buf ( n397097 , n397096 );
nand ( n49666 , n49658 , n397097 );
buf ( n397099 , n49666 );
buf ( n397100 , n38960 );
not ( n49669 , n397100 );
buf ( n397102 , n49669 );
nand ( n49671 , n397099 , n397102 );
nand ( n49672 , n49652 , n49671 );
buf ( n397105 , n49672 );
buf ( n397106 , n386477 );
not ( n49675 , n397106 );
buf ( n397108 , n395190 );
not ( n49677 , n397108 );
or ( n49678 , n49675 , n49677 );
nand ( n49679 , n49650 , n38961 );
buf ( n397112 , n49679 );
nand ( n49681 , n49678 , n397112 );
buf ( n397114 , n49681 );
buf ( n397115 , n397114 );
xor ( n49684 , n397105 , n397115 );
buf ( n397117 , n391550 );
not ( n49686 , n28296 );
buf ( n397119 , n49686 );
not ( n49688 , n397119 );
buf ( n397121 , n393525 );
not ( n49690 , n397121 );
or ( n49691 , n49688 , n49690 );
buf ( n397124 , n388962 );
buf ( n397125 , n389856 );
nand ( n49694 , n397124 , n397125 );
buf ( n397127 , n49694 );
buf ( n397128 , n397127 );
nand ( n49697 , n49691 , n397128 );
buf ( n397130 , n49697 );
buf ( n397131 , n397130 );
not ( n49700 , n397131 );
buf ( n397133 , n49700 );
buf ( n397134 , n397133 );
or ( n49703 , n397117 , n397134 );
buf ( n397136 , n396591 );
not ( n49705 , n397136 );
buf ( n397138 , n49705 );
buf ( n397139 , n397138 );
buf ( n397140 , n46062 );
or ( n49709 , n397139 , n397140 );
nand ( n49710 , n49703 , n49709 );
buf ( n397143 , n49710 );
buf ( n397144 , n397143 );
and ( n49713 , n49684 , n397144 );
and ( n49714 , n397105 , n397115 );
or ( n49715 , n49713 , n49714 );
buf ( n397148 , n49715 );
buf ( n397149 , n388998 );
not ( n49718 , n397149 );
buf ( n397151 , n36395 );
not ( n49720 , n397151 );
or ( n49721 , n49718 , n49720 );
buf ( n397154 , n36396 );
buf ( n397155 , n388215 );
nand ( n49724 , n397154 , n397155 );
buf ( n397157 , n49724 );
buf ( n397158 , n397157 );
nand ( n49727 , n49721 , n397158 );
buf ( n397160 , n49727 );
buf ( n397161 , n397160 );
not ( n49730 , n397161 );
buf ( n397163 , n46532 );
not ( n49732 , n397163 );
buf ( n397165 , n49732 );
buf ( n397166 , n397165 );
not ( n49735 , n397166 );
or ( n49736 , n49730 , n49735 );
buf ( n397169 , n388346 );
buf ( n397170 , n396393 );
nand ( n49739 , n397169 , n397170 );
buf ( n397172 , n49739 );
buf ( n397173 , n397172 );
nand ( n49742 , n49736 , n397173 );
buf ( n397175 , n49742 );
or ( n49744 , n397148 , n397175 );
not ( n49745 , n49744 );
or ( n49746 , n49632 , n49745 );
nand ( n49747 , n397148 , n397175 );
nand ( n49748 , n49746 , n49747 );
buf ( n397181 , n49748 );
nand ( n49750 , n49606 , n397181 );
buf ( n397183 , n49750 );
buf ( n397184 , n397183 );
nand ( n49753 , n49598 , n397184 );
buf ( n397186 , n49753 );
not ( n49755 , n397186 );
or ( n49756 , n49547 , n49755 );
buf ( n397189 , n396948 );
buf ( n397190 , n396974 );
nand ( n49759 , n397189 , n397190 );
buf ( n397192 , n49759 );
nand ( n49761 , n49756 , n397192 );
not ( n49762 , n49761 );
buf ( n397195 , n395160 );
buf ( n397196 , n47726 );
and ( n49765 , n397195 , n397196 );
not ( n49766 , n394884 );
not ( n49767 , n394426 );
or ( n49768 , n49766 , n49767 );
buf ( n397201 , n37763 );
buf ( n397202 , n388154 );
nand ( n49771 , n397201 , n397202 );
buf ( n397204 , n49771 );
nand ( n49773 , n49768 , n397204 );
and ( n49774 , n49773 , n40701 );
buf ( n397207 , n49774 );
nor ( n49776 , n49765 , n397207 );
buf ( n397209 , n49776 );
buf ( n397210 , n397209 );
not ( n49779 , n397210 );
buf ( n397212 , n49779 );
not ( n49781 , n397212 );
buf ( n397214 , n48032 );
buf ( n397215 , n395458 );
and ( n49784 , n397214 , n397215 );
not ( n49785 , n397214 );
buf ( n397218 , n395455 );
and ( n49787 , n49785 , n397218 );
nor ( n49788 , n49784 , n49787 );
buf ( n397221 , n49788 );
buf ( n397222 , n397221 );
buf ( n397223 , n395495 );
not ( n49792 , n397223 );
buf ( n397225 , n49792 );
buf ( n397226 , n397225 );
and ( n49795 , n397222 , n397226 );
not ( n49796 , n397222 );
buf ( n397229 , n395495 );
and ( n49798 , n49796 , n397229 );
nor ( n49799 , n49795 , n49798 );
buf ( n397232 , n49799 );
buf ( n397233 , n397232 );
not ( n49802 , n397233 );
buf ( n397235 , n49802 );
not ( n49804 , n397235 );
or ( n49805 , n49781 , n49804 );
not ( n49806 , n397209 );
not ( n49807 , n397232 );
or ( n49808 , n49806 , n49807 );
buf ( n397241 , n47762 );
not ( n49810 , n397241 );
buf ( n397243 , n49810 );
buf ( n397244 , n397243 );
buf ( n397245 , n389602 );
not ( n49814 , n397245 );
buf ( n397247 , n36251 );
not ( n49816 , n397247 );
or ( n49817 , n49814 , n49816 );
buf ( n397250 , n40775 );
buf ( n397251 , n389593 );
nand ( n49820 , n397250 , n397251 );
buf ( n397253 , n49820 );
buf ( n397254 , n397253 );
nand ( n49823 , n49817 , n397254 );
buf ( n397256 , n49823 );
buf ( n397257 , n397256 );
not ( n49826 , n397257 );
buf ( n397259 , n383891 );
not ( n49828 , n397259 );
or ( n49829 , n49826 , n49828 );
nand ( n49830 , n391602 , n47793 );
buf ( n397263 , n49830 );
nand ( n49832 , n49829 , n397263 );
buf ( n397265 , n49832 );
buf ( n397266 , n397265 );
xor ( n49835 , n397244 , n397266 );
buf ( n397268 , n390432 );
not ( n49837 , n397268 );
buf ( n397270 , n47412 );
not ( n49839 , n397270 );
buf ( n397272 , n388293 );
not ( n49841 , n397272 );
or ( n49842 , n49839 , n49841 );
buf ( n397275 , n390704 );
not ( n49844 , n397275 );
buf ( n397277 , n49844 );
buf ( n397278 , n397277 );
buf ( n397279 , n49102 );
nand ( n49848 , n397278 , n397279 );
buf ( n397281 , n49848 );
buf ( n397282 , n397281 );
nand ( n49851 , n49842 , n397282 );
buf ( n397284 , n49851 );
buf ( n397285 , n397284 );
not ( n49854 , n397285 );
or ( n49855 , n49837 , n49854 );
buf ( n397288 , n396545 );
buf ( n397289 , n392788 );
nand ( n49858 , n397288 , n397289 );
buf ( n397291 , n49858 );
buf ( n397292 , n397291 );
nand ( n49861 , n49855 , n397292 );
buf ( n397294 , n49861 );
buf ( n397295 , n397294 );
and ( n49864 , n49835 , n397295 );
and ( n49865 , n397244 , n397266 );
or ( n49866 , n49864 , n49865 );
buf ( n397299 , n49866 );
nand ( n49868 , n49808 , n397299 );
nand ( n49869 , n49805 , n49868 );
buf ( n397302 , n49869 );
xor ( n49871 , n395507 , n48088 );
xor ( n49872 , n49871 , n48100 );
buf ( n397305 , n49872 );
xor ( n49874 , n397302 , n397305 );
xor ( n49875 , n395144 , n395171 );
xor ( n49876 , n49875 , n395250 );
buf ( n397309 , n49876 );
and ( n49878 , n49874 , n397309 );
and ( n49879 , n397302 , n397305 );
or ( n49880 , n49878 , n49879 );
buf ( n397313 , n49880 );
buf ( n397314 , n397313 );
not ( n49883 , n397314 );
buf ( n397316 , n49883 );
nand ( n49885 , n49762 , n397316 );
not ( n49886 , n49885 );
or ( n49887 , n49492 , n49886 );
not ( n49888 , n397316 );
nand ( n49889 , n49888 , n49761 );
nand ( n49890 , n49887 , n49889 );
buf ( n397323 , n49890 );
xor ( n49892 , n396825 , n397323 );
not ( n49893 , n395428 );
not ( n49894 , n48118 );
not ( n49895 , n49894 );
or ( n49896 , n49893 , n49895 );
or ( n49897 , n395428 , n49894 );
nand ( n49898 , n49896 , n49897 );
not ( n49899 , n49898 );
xor ( n49900 , n395300 , n49899 );
buf ( n397333 , n49900 );
and ( n49902 , n49892 , n397333 );
and ( n49903 , n396825 , n397323 );
or ( n49904 , n49902 , n49903 );
buf ( n397337 , n49904 );
nand ( n49906 , n49386 , n397337 );
nand ( n49907 , n49382 , n49906 );
not ( n49908 , n49907 );
and ( n49909 , n49288 , n49908 );
not ( n49910 , n49288 );
and ( n49911 , n49910 , n49907 );
nor ( n49912 , n49909 , n49911 );
xor ( n49913 , n48753 , n49912 );
buf ( n397346 , n49260 );
buf ( n397347 , n49279 );
xor ( n49916 , n397346 , n397347 );
buf ( n397349 , n396708 );
xnor ( n49918 , n49916 , n397349 );
buf ( n397351 , n49918 );
buf ( n397352 , n397351 );
xor ( n49921 , n395547 , n48104 );
xor ( n49922 , n49921 , n395553 );
xor ( n49923 , n395372 , n395397 );
xor ( n49924 , n49923 , n395419 );
buf ( n397357 , n49924 );
not ( n49926 , n397357 );
nand ( n49927 , n49922 , n49926 );
buf ( n397360 , n49927 );
not ( n49929 , n397360 );
buf ( n397362 , n43727 );
not ( n49931 , n397362 );
not ( n49932 , n391027 );
not ( n49933 , n36068 );
not ( n49934 , n49933 );
or ( n49935 , n49932 , n49934 );
buf ( n397368 , n391027 );
not ( n49937 , n397368 );
not ( n49938 , n41359 );
buf ( n397371 , n49938 );
nand ( n49940 , n49937 , n397371 );
buf ( n397373 , n49940 );
nand ( n49942 , n49935 , n397373 );
buf ( n397375 , n49942 );
not ( n49944 , n397375 );
or ( n49945 , n49931 , n49944 );
buf ( n397378 , n396780 );
buf ( n397379 , n43515 );
nand ( n49948 , n397378 , n397379 );
buf ( n397381 , n49948 );
buf ( n397382 , n397381 );
nand ( n49951 , n49945 , n397382 );
buf ( n397384 , n49951 );
buf ( n397385 , n397384 );
not ( n49954 , n397385 );
buf ( n397387 , n49954 );
buf ( n397388 , n397387 );
not ( n49957 , n397388 );
buf ( n397390 , n45260 );
not ( n49959 , n397390 );
and ( n49960 , n392247 , n386391 );
not ( n49961 , n392247 );
and ( n49962 , n49961 , n35301 );
or ( n49963 , n49960 , n49962 );
buf ( n397396 , n49963 );
not ( n49965 , n397396 );
or ( n49966 , n49959 , n49965 );
buf ( n397399 , n396751 );
buf ( n397400 , n392740 );
nand ( n49969 , n397399 , n397400 );
buf ( n397402 , n49969 );
buf ( n397403 , n397402 );
nand ( n49972 , n49966 , n397403 );
buf ( n397405 , n49972 );
not ( n49974 , n397405 );
buf ( n397407 , n49974 );
not ( n49976 , n397407 );
or ( n49977 , n49957 , n49976 );
buf ( n397410 , n389162 );
not ( n49979 , n397410 );
buf ( n397412 , n396462 );
not ( n49981 , n397412 );
or ( n49982 , n49979 , n49981 );
buf ( n397415 , n41671 );
not ( n49984 , n397415 );
buf ( n397417 , n389692 );
not ( n49986 , n397417 );
buf ( n397419 , n49986 );
buf ( n397420 , n397419 );
not ( n49989 , n397420 );
or ( n49990 , n49984 , n49989 );
buf ( n397423 , n389692 );
buf ( n397424 , n41670 );
nand ( n49993 , n397423 , n397424 );
buf ( n397426 , n49993 );
buf ( n397427 , n397426 );
nand ( n49996 , n49990 , n397427 );
buf ( n397429 , n49996 );
buf ( n397430 , n397429 );
buf ( n397431 , n41711 );
nand ( n50000 , n397430 , n397431 );
buf ( n397433 , n50000 );
buf ( n397434 , n397433 );
nand ( n50003 , n49982 , n397434 );
buf ( n397436 , n50003 );
not ( n50005 , n397436 );
buf ( n397438 , n48965 );
buf ( n397439 , n48943 );
xor ( n50008 , n397438 , n397439 );
buf ( n397441 , n396428 );
xnor ( n50010 , n50008 , n397441 );
buf ( n397443 , n50010 );
buf ( n397444 , n397443 );
not ( n50013 , n397444 );
buf ( n397446 , n50013 );
not ( n50015 , n397446 );
or ( n50016 , n50005 , n50015 );
buf ( n397449 , n397436 );
not ( n50018 , n397449 );
buf ( n397451 , n50018 );
not ( n50020 , n397451 );
not ( n50021 , n397443 );
or ( n50022 , n50020 , n50021 );
buf ( n397455 , n47726 );
not ( n50024 , n397455 );
buf ( n397457 , n49773 );
not ( n50026 , n397457 );
or ( n50027 , n50024 , n50026 );
buf ( n397460 , n394884 );
not ( n50029 , n397460 );
buf ( n397462 , n391483 );
not ( n50031 , n397462 );
or ( n50032 , n50029 , n50031 );
buf ( n397465 , n29077 );
buf ( n397466 , n388154 );
nand ( n50035 , n397465 , n397466 );
buf ( n397468 , n50035 );
buf ( n397469 , n397468 );
nand ( n50038 , n50032 , n397469 );
buf ( n397471 , n50038 );
buf ( n397472 , n397471 );
buf ( n50041 , n40699 );
buf ( n397474 , n50041 );
not ( n50043 , n397474 );
buf ( n397476 , n50043 );
buf ( n397477 , n397476 );
nand ( n50046 , n397472 , n397477 );
buf ( n397479 , n50046 );
buf ( n397480 , n397479 );
nand ( n50049 , n50027 , n397480 );
buf ( n397482 , n50049 );
buf ( n397483 , n397482 );
buf ( n397484 , n372373 );
not ( n50053 , n397484 );
buf ( n397486 , n50053 );
buf ( n397487 , n397486 );
not ( n50056 , n397487 );
buf ( n397489 , n50056 );
buf ( n397490 , n397489 );
not ( n50059 , n397490 );
buf ( n397492 , n50059 );
buf ( n397493 , n397492 );
buf ( n50062 , n397493 );
buf ( n397495 , n50062 );
buf ( n397496 , n397495 );
not ( n50065 , n397496 );
buf ( n397498 , n50065 );
buf ( n397499 , n397498 );
not ( n50068 , n397499 );
buf ( n397501 , n384143 );
not ( n50070 , n397501 );
or ( n50071 , n50068 , n50070 );
buf ( n397504 , n382854 );
buf ( n397505 , n397495 );
nand ( n50074 , n397504 , n397505 );
buf ( n397507 , n50074 );
buf ( n397508 , n397507 );
nand ( n50077 , n50071 , n397508 );
buf ( n397510 , n50077 );
buf ( n397511 , n389547 );
buf ( n397512 , n396567 );
nand ( n50086 , n397511 , n397512 );
buf ( n397514 , n50086 );
buf ( n397515 , n397514 );
nand ( n50089 , C1 , n397515 );
buf ( n397517 , n50089 );
buf ( n397518 , n397517 );
xor ( n50092 , n397483 , n397518 );
and ( n50093 , n392884 , n389753 );
not ( n50094 , n392884 );
buf ( n397522 , n385972 );
not ( n50096 , n397522 );
buf ( n397524 , n50096 );
and ( n50098 , n50094 , n397524 );
or ( n50099 , n50093 , n50098 );
buf ( n397527 , n50099 );
not ( n50101 , n397527 );
buf ( n397529 , n382595 );
not ( n50103 , n397529 );
or ( n50104 , n50101 , n50103 );
buf ( n397532 , n389024 );
buf ( n397533 , n396418 );
nand ( n50107 , n397532 , n397533 );
buf ( n397535 , n50107 );
buf ( n397536 , n397535 );
nand ( n50110 , n50104 , n397536 );
buf ( n397538 , n50110 );
buf ( n397539 , n397538 );
and ( n50113 , n50092 , n397539 );
and ( n50114 , n397483 , n397518 );
or ( n50115 , n50113 , n50114 );
buf ( n397543 , n50115 );
nand ( n50117 , n50022 , n397543 );
nand ( n50118 , n50016 , n50117 );
buf ( n397546 , n50118 );
buf ( n50120 , n397546 );
buf ( n397548 , n50120 );
buf ( n397549 , n397548 );
nand ( n50123 , n49977 , n397549 );
buf ( n397551 , n50123 );
buf ( n397552 , n397551 );
buf ( n397553 , n397384 );
buf ( n397554 , n397405 );
nand ( n50128 , n397553 , n397554 );
buf ( n397556 , n50128 );
buf ( n397557 , n397556 );
nand ( n50131 , n397552 , n397557 );
buf ( n397559 , n50131 );
buf ( n397560 , n397559 );
not ( n50134 , n397560 );
or ( n50135 , n49929 , n50134 );
not ( n50136 , n49922 );
nand ( n50137 , n50136 , n397357 );
buf ( n397565 , n50137 );
nand ( n50139 , n50135 , n397565 );
buf ( n397567 , n50139 );
not ( n50141 , n397567 );
buf ( n397569 , n49293 );
buf ( n397570 , n49363 );
xor ( n50144 , n397569 , n397570 );
buf ( n397572 , n49290 );
xnor ( n50146 , n50144 , n397572 );
buf ( n397574 , n50146 );
not ( n50148 , n397574 );
not ( n50149 , n50148 );
or ( n50150 , n50141 , n50149 );
buf ( n397578 , n397567 );
not ( n50152 , n397578 );
buf ( n397580 , n50152 );
buf ( n397581 , n397580 );
not ( n50155 , n397581 );
buf ( n397583 , n397574 );
not ( n50157 , n397583 );
or ( n50158 , n50155 , n50157 );
xor ( n50159 , n48780 , n396315 );
xor ( n50160 , n50159 , n396688 );
buf ( n397588 , n50160 );
not ( n50162 , n397588 );
buf ( n397590 , n50162 );
buf ( n397591 , n397590 );
nand ( n50165 , n50158 , n397591 );
buf ( n397593 , n50165 );
nand ( n50167 , n50150 , n397593 );
not ( n50168 , n50167 );
buf ( n397596 , n50168 );
xor ( n50170 , n397352 , n397596 );
xor ( n50171 , n396285 , n396289 );
xor ( n50172 , n50171 , n396311 );
buf ( n397600 , n50172 );
not ( n50174 , n397600 );
buf ( n397602 , n396787 );
buf ( n397603 , n396762 );
xor ( n50177 , n397602 , n397603 );
buf ( n397605 , n396736 );
xnor ( n50179 , n50177 , n397605 );
buf ( n397607 , n50179 );
nand ( n50181 , n50174 , n397607 );
not ( n50182 , n50181 );
xor ( n50183 , n396362 , n396444 );
xor ( n50184 , n50183 , n396470 );
buf ( n397612 , n50184 );
buf ( n397613 , n397612 );
not ( n50187 , n397613 );
xor ( n50188 , n396552 , n396575 );
xor ( n50189 , n50188 , n396672 );
buf ( n397617 , n50189 );
buf ( n397618 , n397617 );
not ( n50192 , n397618 );
buf ( n397620 , n50192 );
buf ( n397621 , n397620 );
not ( n50195 , n397621 );
buf ( n397623 , n396504 );
buf ( n397624 , n390362 );
and ( n50198 , n397623 , n397624 );
and ( n50199 , n37173 , n388105 );
not ( n50200 , n37173 );
and ( n50201 , n50200 , n388102 );
or ( n50202 , n50199 , n50201 );
buf ( n397630 , n50202 );
buf ( n397631 , n43286 );
and ( n50205 , n397630 , n397631 );
buf ( n397633 , n50205 );
buf ( n397634 , n397633 );
nor ( n50208 , n50198 , n397634 );
buf ( n397636 , n50208 );
buf ( n397637 , n397636 );
not ( n50211 , n397637 );
or ( n50212 , n50195 , n50211 );
buf ( n397640 , n393592 );
buf ( n397641 , n389356 );
buf ( n397642 , n37037 );
and ( n50216 , n397641 , n397642 );
not ( n50217 , n397641 );
buf ( n397645 , n395879 );
and ( n50219 , n50217 , n397645 );
nor ( n50220 , n50216 , n50219 );
buf ( n397648 , n50220 );
buf ( n397649 , n397648 );
or ( n50223 , n397640 , n397649 );
buf ( n397651 , n392666 );
not ( n50225 , n397651 );
buf ( n397653 , n50225 );
buf ( n397654 , n397653 );
buf ( n397655 , n397015 );
not ( n50229 , n397655 );
buf ( n397657 , n50229 );
buf ( n397658 , n397657 );
or ( n50232 , n397654 , n397658 );
nand ( n50233 , n50223 , n50232 );
buf ( n397661 , n50233 );
buf ( n397662 , n397661 );
buf ( n397663 , n396604 );
buf ( n397664 , n396634 );
xor ( n50238 , n397663 , n397664 );
buf ( n397666 , n49233 );
xor ( n50240 , n50238 , n397666 );
buf ( n397668 , n50240 );
buf ( n397669 , n397668 );
xor ( n50243 , n397662 , n397669 );
buf ( n397671 , n391164 );
and ( n50245 , n391446 , n391183 );
not ( n50246 , n391446 );
and ( n50247 , n50246 , n385729 );
nor ( n50248 , n50245 , n50247 );
buf ( n397676 , n50248 );
or ( n50250 , n397671 , n397676 );
buf ( n397678 , n391176 );
buf ( n397679 , n396987 );
not ( n50253 , n397679 );
buf ( n397681 , n50253 );
buf ( n397682 , n397681 );
or ( n50256 , n397678 , n397682 );
nand ( n50257 , n50250 , n50256 );
buf ( n397685 , n50257 );
buf ( n397686 , n397685 );
and ( n50260 , n50243 , n397686 );
and ( n50261 , n397662 , n397669 );
or ( n50262 , n50260 , n50261 );
buf ( n397690 , n50262 );
buf ( n397691 , n397690 );
nand ( n50265 , n50212 , n397691 );
buf ( n397693 , n50265 );
buf ( n397694 , n397693 );
buf ( n397695 , n397636 );
not ( n50269 , n397695 );
buf ( n397697 , n50269 );
buf ( n397698 , n397697 );
buf ( n397699 , n397617 );
nand ( n50273 , n397698 , n397699 );
buf ( n397701 , n50273 );
buf ( n397702 , n397701 );
nand ( n50276 , n397694 , n397702 );
buf ( n397704 , n50276 );
buf ( n397705 , n397704 );
not ( n50279 , n397705 );
or ( n50280 , n50187 , n50279 );
buf ( n397708 , n397612 );
not ( n50282 , n397708 );
buf ( n397710 , n50282 );
buf ( n397711 , n397710 );
not ( n50285 , n397711 );
not ( n50286 , n397704 );
buf ( n397714 , n50286 );
not ( n50288 , n397714 );
or ( n50289 , n50285 , n50288 );
buf ( n397717 , n397033 );
not ( n50291 , n397717 );
buf ( n397719 , n396999 );
not ( n50293 , n397719 );
or ( n50294 , n50291 , n50293 );
buf ( n397722 , n396999 );
buf ( n397723 , n397033 );
or ( n50297 , n397722 , n397723 );
nand ( n50298 , n50294 , n50297 );
buf ( n397726 , n50298 );
buf ( n397727 , n397726 );
buf ( n397728 , n49748 );
not ( n50302 , n397728 );
buf ( n397730 , n50302 );
buf ( n397731 , n397730 );
and ( n50305 , n397727 , n397731 );
not ( n50306 , n397727 );
buf ( n397734 , n49748 );
and ( n50308 , n50306 , n397734 );
nor ( n50309 , n50305 , n50308 );
buf ( n397737 , n50309 );
not ( n50311 , n397737 );
not ( n50312 , n46921 );
not ( n50313 , n396618 );
or ( n50314 , n50312 , n50313 );
buf ( n397742 , n24050 );
not ( n50316 , n397742 );
not ( n50317 , n40817 );
buf ( n397745 , n50317 );
not ( n50319 , n397745 );
or ( n50320 , n50316 , n50319 );
buf ( n397748 , n40818 );
buf ( n397749 , n45391 );
nand ( n50323 , n397748 , n397749 );
buf ( n397751 , n50323 );
buf ( n397752 , n397751 );
nand ( n50326 , n50320 , n397752 );
buf ( n397754 , n50326 );
buf ( n397755 , n397754 );
buf ( n397756 , n396622 );
nand ( n50330 , n397755 , n397756 );
buf ( n397758 , n50330 );
nand ( n50332 , n50314 , n397758 );
not ( n50333 , n50332 );
not ( n50334 , n50333 );
not ( n50335 , n37338 );
buf ( n397763 , n388543 );
not ( n50337 , n397763 );
buf ( n397765 , n388897 );
not ( n50339 , n397765 );
or ( n50340 , n50337 , n50339 );
buf ( n397768 , n395478 );
buf ( n397769 , n388546 );
nand ( n50343 , n397768 , n397769 );
buf ( n397771 , n50343 );
buf ( n397772 , n397771 );
nand ( n50346 , n50340 , n397772 );
buf ( n397774 , n50346 );
not ( n50348 , n397774 );
or ( n50349 , n50335 , n50348 );
nand ( n50350 , n49225 , n37314 );
nand ( n50351 , n50349 , n50350 );
buf ( n397779 , n50351 );
not ( n50353 , n397779 );
buf ( n397781 , n50353 );
not ( n50355 , n397781 );
or ( n50356 , n50334 , n50355 );
not ( n50357 , n383894 );
buf ( n397785 , n388230 );
not ( n50359 , n397785 );
buf ( n397787 , n389936 );
not ( n50361 , n397787 );
or ( n50362 , n50359 , n50361 );
buf ( n397790 , n388272 );
not ( n50364 , n397790 );
buf ( n397792 , n388242 );
nand ( n50366 , n50364 , n397792 );
buf ( n397794 , n50366 );
buf ( n397795 , n397794 );
nand ( n50369 , n50362 , n397795 );
buf ( n397797 , n50369 );
not ( n50371 , n397797 );
or ( n50372 , n50357 , n50371 );
buf ( n397800 , n397256 );
buf ( n397801 , n383907 );
nand ( n50375 , n397800 , n397801 );
buf ( n397803 , n50375 );
nand ( n50377 , n50372 , n397803 );
nand ( n50378 , n50356 , n50377 );
buf ( n397806 , n50332 );
buf ( n397807 , n50351 );
nand ( n50381 , n397806 , n397807 );
buf ( n397809 , n50381 );
and ( n50383 , n50378 , n397809 );
buf ( n397811 , n396897 );
buf ( n397812 , n388833 );
and ( n50386 , n397811 , n397812 );
not ( n50387 , n44423 );
not ( n50388 , n41342 );
or ( n50389 , n50387 , n50388 );
buf ( n397817 , n36564 );
buf ( n397818 , n45897 );
nand ( n50392 , n397817 , n397818 );
buf ( n397820 , n50392 );
nand ( n50394 , n50389 , n397820 );
not ( n50395 , n50394 );
nor ( n50396 , n50395 , n41374 );
buf ( n397824 , n50396 );
nor ( n50398 , n50386 , n397824 );
buf ( n397826 , n50398 );
xor ( n50400 , n50383 , n397826 );
buf ( n397828 , n394817 );
not ( n50402 , n397828 );
buf ( n397830 , n388235 );
not ( n50404 , n397830 );
or ( n50405 , n50402 , n50404 );
buf ( n397833 , n384965 );
buf ( n397834 , n394814 );
nand ( n50408 , n397833 , n397834 );
buf ( n397836 , n50408 );
buf ( n397837 , n397836 );
nand ( n50411 , n50405 , n397837 );
buf ( n397839 , n50411 );
buf ( n397840 , n397839 );
not ( n50414 , n397840 );
buf ( n397842 , n50414 );
buf ( n397843 , n397842 );
not ( n50417 , n397843 );
buf ( n397845 , n383014 );
not ( n50419 , n397845 );
and ( n50420 , n50417 , n50419 );
not ( n50421 , n49431 );
nor ( n50422 , n50421 , n386307 );
buf ( n397850 , n50422 );
nor ( n50424 , n50420 , n397850 );
buf ( n397852 , n50424 );
and ( n50426 , n50400 , n397852 );
and ( n50427 , n50383 , n397826 );
or ( n50428 , n50426 , n50427 );
not ( n50429 , n50428 );
and ( n50430 , n50311 , n50429 );
buf ( n397858 , n50428 );
buf ( n397859 , n397737 );
nand ( n50433 , n397858 , n397859 );
buf ( n397861 , n50433 );
not ( n50435 , n397209 );
not ( n50436 , n397235 );
or ( n50437 , n50435 , n50436 );
buf ( n397865 , n397212 );
buf ( n397866 , n397232 );
nand ( n50440 , n397865 , n397866 );
buf ( n397868 , n50440 );
nand ( n50442 , n50437 , n397868 );
xor ( n50443 , n50442 , n397299 );
and ( n50444 , n397861 , n50443 );
nor ( n50445 , n50430 , n50444 );
buf ( n397873 , n50445 );
not ( n50447 , n397873 );
buf ( n397875 , n50447 );
buf ( n397876 , n397875 );
nand ( n50450 , n50289 , n397876 );
buf ( n397878 , n50450 );
buf ( n397879 , n397878 );
nand ( n50453 , n50280 , n397879 );
buf ( n397881 , n50453 );
not ( n50455 , n397881 );
or ( n50456 , n50182 , n50455 );
buf ( n397884 , n397607 );
not ( n50458 , n397884 );
buf ( n397886 , n397600 );
nand ( n50460 , n50458 , n397886 );
buf ( n397888 , n50460 );
nand ( n50462 , n50456 , n397888 );
buf ( n397890 , n50462 );
not ( n50464 , n397890 );
buf ( n397892 , n396474 );
buf ( n397893 , n396334 );
xor ( n50467 , n397892 , n397893 );
buf ( n397895 , n396682 );
xnor ( n50469 , n50467 , n397895 );
buf ( n397897 , n50469 );
buf ( n397898 , n397897 );
not ( n50472 , n397898 );
and ( n50473 , n49761 , n397316 );
not ( n50474 , n49761 );
and ( n50475 , n50474 , n397313 );
nor ( n50476 , n50473 , n50475 );
xor ( n50477 , n396923 , n50476 );
buf ( n397905 , n50477 );
not ( n50479 , n397905 );
or ( n50480 , n50472 , n50479 );
buf ( n397908 , n395362 );
not ( n50482 , n397908 );
buf ( n397910 , n396941 );
not ( n50484 , n397910 );
or ( n50485 , n50482 , n50484 );
buf ( n397913 , n47863 );
buf ( n397914 , n35519 );
and ( n50488 , n397913 , n397914 );
not ( n50489 , n397913 );
buf ( n397917 , n392144 );
and ( n50491 , n50489 , n397917 );
nor ( n50492 , n50488 , n50491 );
buf ( n397920 , n50492 );
buf ( n397921 , n397920 );
buf ( n397922 , n395349 );
nand ( n50496 , n397921 , n397922 );
buf ( n397924 , n50496 );
buf ( n397925 , n397924 );
nand ( n50499 , n50485 , n397925 );
buf ( n397927 , n50499 );
not ( n50501 , n397927 );
buf ( n397929 , n396964 );
buf ( n397930 , n388809 );
and ( n50504 , n397929 , n397930 );
buf ( n397932 , n388760 );
not ( n50506 , n397932 );
buf ( n397934 , n45893 );
not ( n50508 , n397934 );
or ( n50509 , n50506 , n50508 );
buf ( n397937 , n36216 );
buf ( n397938 , n388757 );
nand ( n50512 , n397937 , n397938 );
buf ( n397940 , n50512 );
buf ( n397941 , n397940 );
nand ( n50515 , n50509 , n397941 );
buf ( n397943 , n50515 );
buf ( n397944 , n397943 );
not ( n50518 , n397944 );
buf ( n397946 , n388743 );
nor ( n50520 , n50518 , n397946 );
buf ( n397948 , n50520 );
buf ( n397949 , n397948 );
nor ( n50523 , n50504 , n397949 );
buf ( n397951 , n50523 );
nand ( n50525 , n50501 , n397951 );
not ( n50526 , n50525 );
buf ( n397954 , n370059 );
nand ( n50530 , C1 , n397954 );
buf ( n397956 , n50530 );
not ( n50532 , n397956 );
not ( n50533 , n22497 );
and ( n50547 , n50533 , C1 );
or ( n50553 , n50547 , C0 );
and ( n50554 , n50532 , n50553 );
not ( n50555 , n50532 );
and ( n50557 , n22497 , C1 );
or ( n50561 , n50557 , C0 );
and ( n50562 , n50555 , n50561 );
or ( n50563 , n50554 , n50562 );
not ( n50564 , n50563 );
buf ( n397968 , n50564 );
not ( n50566 , n397968 );
not ( n50567 , n50564 );
not ( n50568 , n22497 );
not ( n50569 , n50532 );
or ( n50570 , n50568 , n50569 );
nand ( n50571 , n397956 , n50533 );
nand ( n50572 , n50570 , n50571 );
not ( n50573 , n50572 );
and ( n50574 , n23551 , n50573 );
not ( n50575 , n23551 );
and ( n50576 , n50575 , n50572 );
or ( n50577 , n50574 , n50576 );
nor ( n50578 , n50567 , n50577 );
buf ( n50579 , n50578 );
not ( n50580 , n50579 );
buf ( n397984 , n50580 );
not ( n50582 , n397984 );
or ( n50583 , n50566 , n50582 );
not ( n50584 , n47891 );
buf ( n397988 , n50584 );
not ( n50586 , n397988 );
buf ( n397990 , n50586 );
buf ( n397991 , n397990 );
not ( n50589 , n397991 );
buf ( n397993 , n388113 );
not ( n50591 , n397993 );
or ( n50592 , n50589 , n50591 );
buf ( n397996 , n385499 );
buf ( n397997 , n50584 );
nand ( n50595 , n397996 , n397997 );
buf ( n397999 , n50595 );
buf ( n398000 , n397999 );
nand ( n50598 , n50592 , n398000 );
buf ( n398002 , n50598 );
buf ( n398003 , n398002 );
nand ( n50601 , n50583 , n398003 );
buf ( n398005 , n50601 );
not ( n50603 , n398005 );
or ( n50604 , n50526 , n50603 );
buf ( n398008 , n397951 );
not ( n50606 , n398008 );
buf ( n398010 , n397927 );
nand ( n50608 , n50606 , n398010 );
buf ( n398012 , n50608 );
nand ( n50610 , n50604 , n398012 );
buf ( n398014 , n50610 );
not ( n50612 , n398014 );
buf ( n398016 , n396676 );
buf ( n398017 , n49050 );
xor ( n50615 , n398016 , n398017 );
buf ( n398019 , n396514 );
xnor ( n50617 , n50615 , n398019 );
buf ( n398021 , n50617 );
buf ( n398022 , n398021 );
not ( n50620 , n398022 );
buf ( n398024 , n50620 );
buf ( n398025 , n398024 );
not ( n50623 , n398025 );
or ( n50624 , n50612 , n50623 );
buf ( n398028 , n50610 );
not ( n50626 , n398028 );
buf ( n398030 , n50626 );
buf ( n398031 , n398030 );
not ( n50629 , n398031 );
buf ( n398033 , n398021 );
not ( n50631 , n398033 );
or ( n50632 , n50629 , n50631 );
xor ( n50633 , n397302 , n397305 );
xor ( n50634 , n50633 , n397309 );
buf ( n398038 , n50634 );
buf ( n398039 , n398038 );
nand ( n50637 , n50632 , n398039 );
buf ( n398041 , n50637 );
buf ( n398042 , n398041 );
nand ( n50640 , n50624 , n398042 );
buf ( n398044 , n50640 );
buf ( n398045 , n398044 );
nand ( n50643 , n50480 , n398045 );
buf ( n398047 , n50643 );
not ( n50645 , n397897 );
buf ( n398049 , n50477 );
not ( n50647 , n398049 );
buf ( n398051 , n50647 );
nand ( n50649 , n50645 , n398051 );
nand ( n50650 , n398047 , n50649 );
buf ( n398054 , n50650 );
not ( n50652 , n398054 );
buf ( n398056 , n50652 );
buf ( n398057 , n398056 );
nand ( n50655 , n50464 , n398057 );
buf ( n398059 , n50655 );
buf ( n398060 , n398059 );
xor ( n50658 , n396825 , n397323 );
xor ( n50659 , n50658 , n397333 );
buf ( n398063 , n50659 );
buf ( n398064 , n398063 );
and ( n50662 , n398060 , n398064 );
buf ( n398066 , n50462 );
buf ( n398067 , n50650 );
and ( n50665 , n398066 , n398067 );
buf ( n398069 , n50665 );
buf ( n398070 , n398069 );
nor ( n50668 , n50662 , n398070 );
buf ( n398072 , n50668 );
buf ( n398073 , n398072 );
and ( n50671 , n50170 , n398073 );
and ( n50672 , n397352 , n397596 );
or ( n50673 , n50671 , n50672 );
buf ( n398077 , n50673 );
xor ( n50675 , n49913 , n398077 );
buf ( n398079 , n49367 );
buf ( n398080 , n397337 );
xor ( n50678 , n398079 , n398080 );
buf ( n398082 , n49380 );
xor ( n50680 , n50678 , n398082 );
buf ( n398084 , n50680 );
not ( n50682 , n398084 );
xor ( n50683 , n397352 , n397596 );
xor ( n50684 , n50683 , n398073 );
buf ( n398088 , n50684 );
not ( n50686 , n398088 );
not ( n50687 , n50686 );
or ( n50688 , n50682 , n50687 );
not ( n50689 , n398084 );
not ( n50690 , n50689 );
not ( n50691 , n398088 );
or ( n50692 , n50690 , n50691 );
buf ( n398096 , n397567 );
buf ( n398097 , n50160 );
xor ( n50695 , n398096 , n398097 );
buf ( n398099 , n397574 );
xnor ( n50697 , n50695 , n398099 );
buf ( n398101 , n50697 );
not ( n50699 , n398101 );
xor ( n50700 , n396948 , n396977 );
xnor ( n50701 , n50700 , n397186 );
buf ( n398105 , n50701 );
buf ( n398106 , n396839 );
not ( n50704 , n398106 );
buf ( n398108 , n50704 );
buf ( n398109 , n398108 );
not ( n50707 , n398109 );
buf ( n398111 , n393409 );
not ( n50709 , n398111 );
and ( n50710 , n50707 , n50709 );
buf ( n398114 , n393384 );
not ( n50712 , n398114 );
buf ( n398116 , n50712 );
buf ( n398117 , n398116 );
not ( n50715 , n398117 );
buf ( n398119 , n386561 );
not ( n50717 , n398119 );
or ( n50718 , n50715 , n50717 );
buf ( n398122 , n382921 );
buf ( n398123 , n393381 );
nand ( n50721 , n398122 , n398123 );
buf ( n398125 , n50721 );
buf ( n398126 , n398125 );
nand ( n50724 , n50718 , n398126 );
buf ( n398128 , n50724 );
buf ( n398129 , n398128 );
buf ( n398130 , n393825 );
and ( n50728 , n398129 , n398130 );
nor ( n50729 , n50710 , n50728 );
buf ( n398133 , n50729 );
buf ( n398134 , n398133 );
not ( n50732 , n398134 );
buf ( n398136 , n391027 );
not ( n50734 , n398136 );
buf ( n398138 , n385774 );
not ( n50736 , n398138 );
or ( n50737 , n50734 , n50736 );
buf ( n398141 , n389423 );
buf ( n398142 , n391024 );
nand ( n50740 , n398141 , n398142 );
buf ( n398144 , n50740 );
buf ( n398145 , n398144 );
nand ( n50743 , n50737 , n398145 );
buf ( n398147 , n50743 );
buf ( n398148 , n398147 );
not ( n50746 , n398148 );
buf ( n398150 , n50746 );
not ( n50748 , n398150 );
not ( n50749 , n43537 );
and ( n50750 , n50748 , n50749 );
and ( n50751 , n49942 , n43515 );
nor ( n50752 , n50750 , n50751 );
buf ( n398156 , n50752 );
not ( n50754 , n398156 );
or ( n50755 , n50732 , n50754 );
buf ( n398159 , n392740 );
not ( n50757 , n398159 );
buf ( n398161 , n49963 );
not ( n50759 , n398161 );
or ( n50760 , n50757 , n50759 );
buf ( n398164 , n392247 );
not ( n50762 , n398164 );
buf ( n398166 , n37027 );
not ( n50764 , n398166 );
or ( n50765 , n50762 , n50764 );
buf ( n398169 , n385834 );
buf ( n398170 , n392244 );
nand ( n50768 , n398169 , n398170 );
buf ( n398172 , n50768 );
buf ( n398173 , n398172 );
nand ( n50771 , n50765 , n398173 );
buf ( n398175 , n50771 );
buf ( n398176 , n398175 );
buf ( n398177 , n45260 );
nand ( n50775 , n398176 , n398177 );
buf ( n398179 , n50775 );
buf ( n398180 , n398179 );
nand ( n50778 , n50760 , n398180 );
buf ( n398182 , n50778 );
buf ( n398183 , n398182 );
nand ( n50781 , n50755 , n398183 );
buf ( n398185 , n50781 );
buf ( n398186 , n398185 );
not ( n50784 , n50752 );
buf ( n398188 , n398133 );
not ( n50786 , n398188 );
buf ( n398190 , n50786 );
nand ( n50788 , n50784 , n398190 );
buf ( n398192 , n50788 );
nand ( n50790 , n398186 , n398192 );
buf ( n398194 , n50790 );
buf ( n398195 , n398194 );
or ( n50793 , n398105 , n398195 );
buf ( n398197 , n50793 );
buf ( n398198 , n398197 );
xor ( n50796 , n396855 , n396879 );
xor ( n50797 , n50796 , n396905 );
buf ( n398201 , n50797 );
buf ( n398202 , n398201 );
xor ( n50800 , n397244 , n397266 );
xor ( n50801 , n50800 , n397295 );
buf ( n398205 , n50801 );
buf ( n398206 , n398205 );
buf ( n398207 , n392788 );
not ( n50805 , n398207 );
buf ( n398209 , n397284 );
not ( n50807 , n398209 );
or ( n50808 , n50805 , n50807 );
buf ( n398212 , n47412 );
not ( n50810 , n398212 );
buf ( n398214 , n27612 );
not ( n50812 , n398214 );
or ( n50813 , n50810 , n50812 );
buf ( n398217 , n40758 );
buf ( n398218 , n49102 );
nand ( n50816 , n398217 , n398218 );
buf ( n398220 , n50816 );
buf ( n398221 , n398220 );
nand ( n50819 , n50813 , n398221 );
buf ( n398223 , n50819 );
buf ( n398224 , n398223 );
buf ( n398225 , n390432 );
nand ( n50823 , n398224 , n398225 );
buf ( n398227 , n50823 );
buf ( n398228 , n398227 );
nand ( n50826 , n50808 , n398228 );
buf ( n398230 , n50826 );
buf ( n398231 , n398230 );
buf ( n50829 , n36792 );
buf ( n398233 , n50829 );
buf ( n398234 , n42073 );
not ( n50832 , n398234 );
buf ( n398236 , n36809 );
not ( n50834 , n398236 );
or ( n50835 , n50832 , n50834 );
buf ( n398239 , n40885 );
buf ( n398240 , n42074 );
nand ( n50838 , n398239 , n398240 );
buf ( n398242 , n50838 );
buf ( n398243 , n398242 );
nand ( n50841 , n50835 , n398243 );
buf ( n398245 , n50841 );
buf ( n398246 , n398245 );
nand ( n50844 , n398233 , n398246 );
buf ( n398248 , n50844 );
or ( n50846 , n398248 , n40901 );
nand ( n50847 , n397050 , n40901 );
nand ( n50848 , n50846 , n50847 );
buf ( n398252 , n50848 );
xor ( n50850 , n398231 , n398252 );
buf ( n398254 , n49672 );
not ( n50852 , n398254 );
buf ( n398256 , n50852 );
buf ( n398257 , n398256 );
buf ( n398258 , n394666 );
not ( n50856 , n398258 );
buf ( n398260 , n393525 );
not ( n50858 , n398260 );
or ( n50859 , n50856 , n50858 );
buf ( n398263 , n385473 );
buf ( n398264 , n388566 );
nand ( n50862 , n398263 , n398264 );
buf ( n398266 , n50862 );
buf ( n398267 , n398266 );
nand ( n50865 , n50859 , n398267 );
buf ( n398269 , n50865 );
buf ( n398270 , n398269 );
not ( n50868 , n398270 );
buf ( n398272 , n46056 );
not ( n50870 , n398272 );
or ( n50871 , n50868 , n50870 );
buf ( n398275 , n397130 );
buf ( n398276 , n49166 );
nand ( n50874 , n398275 , n398276 );
buf ( n398278 , n50874 );
buf ( n398279 , n398278 );
nand ( n50877 , n50871 , n398279 );
buf ( n398281 , n50877 );
buf ( n398282 , n398281 );
xor ( n50880 , n398257 , n398282 );
buf ( n398284 , n397754 );
not ( n50882 , n398284 );
buf ( n398286 , n46921 );
not ( n50884 , n398286 );
or ( n50885 , n50882 , n50884 );
not ( n50886 , n24049 );
buf ( n398290 , n28248 );
not ( n50888 , n398290 );
buf ( n398292 , n50888 );
not ( n50890 , n398292 );
or ( n50891 , n50886 , n50890 );
buf ( n398295 , n28250 );
buf ( n398296 , n24049 );
not ( n50894 , n398296 );
buf ( n398298 , n50894 );
buf ( n398299 , n398298 );
nand ( n50897 , n398295 , n398299 );
buf ( n398301 , n50897 );
nand ( n50899 , n50891 , n398301 );
buf ( n398303 , n50899 );
buf ( n398304 , n389125 );
nand ( n50902 , n398303 , n398304 );
buf ( n398306 , n50902 );
buf ( n398307 , n398306 );
nand ( n50905 , n50885 , n398307 );
buf ( n398309 , n50905 );
buf ( n398310 , n398309 );
and ( n50908 , n50880 , n398310 );
and ( n50909 , n398257 , n398282 );
or ( n50910 , n50908 , n50909 );
buf ( n398314 , n50910 );
buf ( n398315 , n398314 );
and ( n50913 , n50850 , n398315 );
and ( n50914 , n398231 , n398252 );
or ( n50915 , n50913 , n50914 );
buf ( n398319 , n50915 );
buf ( n398320 , n398319 );
xor ( n50918 , n398206 , n398320 );
buf ( n398322 , n41711 );
not ( n50920 , n398322 );
buf ( n398324 , n41671 );
buf ( n398325 , n389467 );
not ( n50923 , n398325 );
buf ( n398327 , n50923 );
buf ( n398328 , n398327 );
and ( n50926 , n398324 , n398328 );
not ( n50927 , n398324 );
buf ( n398331 , n389289 );
and ( n50929 , n50927 , n398331 );
nor ( n50930 , n50926 , n50929 );
buf ( n398334 , n50930 );
buf ( n398335 , n398334 );
not ( n50933 , n398335 );
or ( n50934 , n50920 , n50933 );
buf ( n398338 , n397429 );
buf ( n398339 , n389162 );
nand ( n50937 , n398338 , n398339 );
buf ( n398341 , n50937 );
buf ( n398342 , n398341 );
nand ( n50940 , n50934 , n398342 );
buf ( n398344 , n50940 );
buf ( n398345 , n398344 );
and ( n50943 , n50918 , n398345 );
and ( n50944 , n398206 , n398320 );
or ( n50945 , n50943 , n50944 );
buf ( n398349 , n50945 );
buf ( n398350 , n398349 );
or ( n50948 , n398202 , n398350 );
not ( n50949 , n397148 );
xor ( n50950 , n397175 , n50949 );
not ( n50951 , n397063 );
xor ( n50952 , n50950 , n50951 );
buf ( n398356 , n50952 );
not ( n50954 , n398356 );
not ( n50955 , n388746 );
buf ( n398359 , n388760 );
not ( n50957 , n398359 );
buf ( n398361 , n385734 );
not ( n50959 , n398361 );
or ( n50960 , n50957 , n50959 );
buf ( n398364 , n384180 );
buf ( n50962 , n398364 );
buf ( n398366 , n50962 );
buf ( n398367 , n398366 );
buf ( n398368 , n388757 );
nand ( n50966 , n398367 , n398368 );
buf ( n398370 , n50966 );
buf ( n398371 , n398370 );
nand ( n50969 , n50960 , n398371 );
buf ( n398373 , n50969 );
not ( n50971 , n398373 );
or ( n50972 , n50955 , n50971 );
buf ( n398376 , n397943 );
buf ( n398377 , n388809 );
nand ( n50975 , n398376 , n398377 );
buf ( n398379 , n50975 );
nand ( n50977 , n50972 , n398379 );
buf ( n398381 , n50977 );
not ( n50979 , n398381 );
or ( n50980 , n50954 , n50979 );
buf ( n398384 , n50977 );
buf ( n398385 , n50952 );
or ( n50983 , n398384 , n398385 );
xor ( n50984 , n397105 , n397115 );
xor ( n50985 , n50984 , n397144 );
buf ( n398389 , n50985 );
buf ( n398390 , n388502 );
not ( n50988 , n398390 );
buf ( n398392 , n36395 );
not ( n50990 , n398392 );
or ( n50991 , n50988 , n50990 );
not ( n50992 , n36395 );
buf ( n398396 , n50992 );
buf ( n398397 , n388511 );
nand ( n50995 , n398396 , n398397 );
buf ( n398399 , n50995 );
buf ( n398400 , n398399 );
nand ( n398401 , n50991 , n398400 );
buf ( n398402 , n398401 );
not ( n51000 , n398402 );
buf ( n398404 , n384008 );
not ( n51002 , n398404 );
buf ( n398406 , n51002 );
not ( n51004 , n398406 );
or ( n51005 , n51000 , n51004 );
buf ( n398409 , n397160 );
buf ( n398410 , n383940 );
nand ( n51008 , n398409 , n398410 );
buf ( n398412 , n51008 );
nand ( n51010 , n51005 , n398412 );
xor ( n51011 , n398389 , n51010 );
buf ( n398415 , n394210 );
not ( n51013 , n398415 );
buf ( n398417 , n385987 );
not ( n51015 , n398417 );
or ( n51016 , n51013 , n51015 );
buf ( n398420 , n389997 );
buf ( n398421 , n394219 );
nand ( n51019 , n398420 , n398421 );
buf ( n398423 , n51019 );
buf ( n398424 , n398423 );
nand ( n51022 , n51016 , n398424 );
buf ( n398426 , n51022 );
buf ( n398427 , n398426 );
not ( n51025 , n398427 );
buf ( n398429 , n382592 );
not ( n51027 , n398429 );
buf ( n398431 , n51027 );
buf ( n398432 , n398431 );
not ( n51030 , n398432 );
or ( n51031 , n51025 , n51030 );
buf ( n398435 , n379463 );
buf ( n398436 , n50099 );
nand ( n51034 , n398435 , n398436 );
buf ( n398438 , n51034 );
buf ( n398439 , n398438 );
nand ( n51037 , n51031 , n398439 );
buf ( n398441 , n51037 );
and ( n51039 , n51011 , n398441 );
and ( n51040 , n398389 , n51010 );
or ( n51041 , n51039 , n51040 );
buf ( n398445 , n51041 );
nand ( n51043 , n50983 , n398445 );
buf ( n398447 , n51043 );
buf ( n398448 , n398447 );
nand ( n51046 , n50980 , n398448 );
buf ( n398450 , n51046 );
buf ( n398451 , n398450 );
nand ( n51049 , n50948 , n398451 );
buf ( n398453 , n51049 );
buf ( n398454 , n398453 );
buf ( n398455 , n398201 );
buf ( n398456 , n398349 );
nand ( n51054 , n398455 , n398456 );
buf ( n398458 , n51054 );
buf ( n398459 , n398458 );
nand ( n51057 , n398454 , n398459 );
buf ( n398461 , n51057 );
buf ( n398462 , n398461 );
and ( n51060 , n398198 , n398462 );
buf ( n398464 , n398194 );
buf ( n398465 , n50701 );
and ( n51063 , n398464 , n398465 );
buf ( n398467 , n51063 );
buf ( n398468 , n398467 );
nor ( n51066 , n51060 , n398468 );
buf ( n398470 , n51066 );
buf ( n398471 , n398470 );
buf ( n398472 , n397551 );
buf ( n398473 , n397556 );
nand ( n51071 , n398472 , n398473 );
buf ( n398475 , n51071 );
and ( n51073 , n50136 , n49926 );
not ( n51074 , n50136 );
and ( n51075 , n51074 , n397357 );
nor ( n51076 , n51073 , n51075 );
xor ( n51077 , n398475 , n51076 );
buf ( n398481 , n51077 );
xor ( n51079 , n398471 , n398481 );
xor ( n51080 , n396849 , n396909 );
buf ( n398484 , n51080 );
buf ( n398485 , n49485 );
not ( n51083 , n398485 );
buf ( n398487 , n51083 );
buf ( n398488 , n398487 );
and ( n51086 , n398484 , n398488 );
not ( n51087 , n398484 );
buf ( n398491 , n49485 );
and ( n51089 , n51087 , n398491 );
nor ( n51090 , n51086 , n51089 );
buf ( n398494 , n51090 );
buf ( n398495 , n397384 );
not ( n51093 , n398495 );
buf ( n398497 , n50118 );
not ( n51095 , n398497 );
buf ( n398499 , n51095 );
buf ( n398500 , n398499 );
not ( n51098 , n398500 );
or ( n51099 , n51093 , n51098 );
buf ( n398503 , n397387 );
buf ( n398504 , n50118 );
nand ( n51102 , n398503 , n398504 );
buf ( n398506 , n51102 );
buf ( n398507 , n398506 );
nand ( n51105 , n51099 , n398507 );
buf ( n398509 , n51105 );
buf ( n398510 , n398509 );
buf ( n398511 , n49974 );
and ( n51109 , n398510 , n398511 );
not ( n51110 , n398510 );
buf ( n398514 , n397405 );
and ( n51112 , n51110 , n398514 );
nor ( n51113 , n51109 , n51112 );
buf ( n398517 , n51113 );
xor ( n51115 , n398494 , n398517 );
xor ( n51116 , n397710 , n397704 );
xnor ( n51117 , n51116 , n50445 );
and ( n51118 , n51115 , n51117 );
and ( n51119 , n398494 , n398517 );
or ( n51120 , n51118 , n51119 );
buf ( n398524 , n51120 );
and ( n51122 , n51079 , n398524 );
and ( n51123 , n398471 , n398481 );
or ( n51124 , n51122 , n51123 );
buf ( n398528 , n51124 );
not ( n51126 , n398528 );
and ( n51127 , n50699 , n51126 );
buf ( n398531 , n397443 );
buf ( n51129 , n398531 );
buf ( n398533 , n51129 );
buf ( n398534 , n398533 );
buf ( n398535 , n397543 );
not ( n51133 , n398535 );
buf ( n398537 , n397451 );
not ( n51135 , n398537 );
or ( n51136 , n51133 , n51135 );
buf ( n398540 , n397543 );
not ( n51138 , n398540 );
buf ( n398542 , n51138 );
buf ( n398543 , n398542 );
buf ( n398544 , n397436 );
nand ( n51142 , n398543 , n398544 );
buf ( n398546 , n51142 );
buf ( n398547 , n398546 );
nand ( n51145 , n51136 , n398547 );
buf ( n398549 , n51145 );
buf ( n398550 , n398549 );
xor ( n51148 , n398534 , n398550 );
buf ( n398552 , n51148 );
buf ( n398553 , n398552 );
not ( n51151 , n398553 );
buf ( n398555 , n51151 );
buf ( n398556 , n398555 );
not ( n51154 , n398556 );
xor ( n51155 , n397483 , n397518 );
xor ( n51156 , n51155 , n397539 );
buf ( n398560 , n51156 );
not ( n51158 , n43727 );
not ( n51159 , n391027 );
not ( n51160 , n38357 );
or ( n51161 , n51159 , n51160 );
not ( n51162 , n391027 );
not ( n51163 , n37147 );
nand ( n51164 , n51162 , n51163 );
nand ( n51165 , n51161 , n51164 );
not ( n51166 , n51165 );
or ( n51167 , n51158 , n51166 );
buf ( n398571 , n398147 );
buf ( n398572 , n43515 );
nand ( n51170 , n398571 , n398572 );
buf ( n398574 , n51170 );
nand ( n51172 , n51167 , n398574 );
or ( n51173 , n398560 , n51172 );
not ( n51174 , n11366 );
nand ( n51175 , n51174 , n359022 );
not ( n51176 , n359036 );
nor ( n51177 , n51176 , n359039 );
nand ( n51178 , n51177 , n11347 );
nand ( n51179 , n359022 , n11364 );
not ( n51180 , n359039 );
nor ( n51181 , n51180 , n359036 );
nand ( n51182 , n11347 , n51181 );
nand ( n51183 , n51175 , n51178 , n51179 , n51182 );
not ( n51184 , n51183 );
buf ( n51185 , n51184 );
buf ( n398589 , n51185 );
buf ( n398590 , n385328 );
and ( n51188 , n398589 , n398590 );
not ( n51189 , n398589 );
buf ( n398593 , n384143 );
and ( n51191 , n51189 , n398593 );
nor ( n51192 , n51188 , n51191 );
buf ( n398596 , n51192 );
buf ( n398597 , n382938 );
buf ( n398598 , n397510 );
nand ( n51202 , n398597 , n398598 );
buf ( n398600 , n51202 );
buf ( n398601 , n398600 );
nand ( n51205 , C1 , n398601 );
buf ( n398603 , n51205 );
buf ( n398604 , n398603 );
buf ( n398605 , n388141 );
not ( n51209 , n398605 );
buf ( n398607 , n397471 );
not ( n51211 , n398607 );
or ( n51212 , n51209 , n51211 );
not ( n51213 , n388154 );
not ( n51214 , n389940 );
or ( n51215 , n51213 , n51214 );
nand ( n51216 , n396534 , n394884 );
nand ( n51217 , n51215 , n51216 );
buf ( n398615 , n51217 );
buf ( n398616 , n397476 );
nand ( n51220 , n398615 , n398616 );
buf ( n398618 , n51220 );
buf ( n398619 , n398618 );
nand ( n51223 , n51212 , n398619 );
buf ( n398621 , n51223 );
buf ( n398622 , n398621 );
xor ( n51226 , n398604 , n398622 );
buf ( n398624 , n390432 );
not ( n51228 , n398624 );
buf ( n398626 , n49102 );
buf ( n398627 , n41118 );
and ( n51231 , n398626 , n398627 );
not ( n51232 , n398626 );
buf ( n398630 , n27195 );
and ( n51234 , n51232 , n398630 );
nor ( n51235 , n51231 , n51234 );
buf ( n398633 , n51235 );
buf ( n398634 , n398633 );
not ( n51238 , n398634 );
or ( n51239 , n51228 , n51238 );
buf ( n398637 , n398223 );
buf ( n398638 , n392788 );
nand ( n51242 , n398637 , n398638 );
buf ( n398640 , n51242 );
buf ( n398641 , n398640 );
nand ( n51245 , n51239 , n398641 );
buf ( n398643 , n51245 );
buf ( n398644 , n398643 );
buf ( n398645 , n37338 );
not ( n51249 , n398645 );
buf ( n398647 , n389602 );
not ( n51251 , n398647 );
buf ( n398649 , n37345 );
not ( n51253 , n398649 );
or ( n51254 , n51251 , n51253 );
buf ( n398652 , n393562 );
buf ( n398653 , n389593 );
nand ( n51257 , n398652 , n398653 );
buf ( n398655 , n51257 );
buf ( n398656 , n398655 );
nand ( n51260 , n51254 , n398656 );
buf ( n398658 , n51260 );
buf ( n398659 , n398658 );
not ( n51263 , n398659 );
or ( n51264 , n51249 , n51263 );
buf ( n398662 , n397774 );
buf ( n398663 , n393100 );
not ( n51267 , n398663 );
buf ( n398665 , n51267 );
buf ( n398666 , n398665 );
not ( n51270 , n398666 );
buf ( n398668 , n51270 );
buf ( n398669 , n398668 );
nand ( n51273 , n398662 , n398669 );
buf ( n398671 , n51273 );
buf ( n398672 , n398671 );
nand ( n51276 , n51264 , n398672 );
buf ( n398674 , n51276 );
buf ( n398675 , n398674 );
xor ( n51279 , n398644 , n398675 );
buf ( n398677 , n397476 );
not ( n51281 , n398677 );
buf ( n398679 , n394884 );
not ( n51283 , n398679 );
buf ( n398681 , n393135 );
not ( n51285 , n398681 );
or ( n51286 , n51283 , n51285 );
buf ( n398684 , n388892 );
buf ( n398685 , n388154 );
nand ( n51289 , n398684 , n398685 );
buf ( n398687 , n51289 );
buf ( n398688 , n398687 );
nand ( n51292 , n51286 , n398688 );
buf ( n398690 , n51292 );
buf ( n398691 , n398690 );
not ( n51295 , n398691 );
or ( n51296 , n51281 , n51295 );
nand ( n51297 , n51217 , n47726 );
buf ( n398695 , n51297 );
nand ( n51299 , n51296 , n398695 );
buf ( n398697 , n51299 );
buf ( n398698 , n398697 );
and ( n51302 , n51279 , n398698 );
and ( n51303 , n398644 , n398675 );
or ( n51304 , n51302 , n51303 );
buf ( n398702 , n51304 );
buf ( n398703 , n398702 );
and ( n51307 , n51226 , n398703 );
and ( n51308 , n398604 , n398622 );
or ( n51309 , n51307 , n51308 );
buf ( n398707 , n51309 );
nand ( n51311 , n51173 , n398707 );
buf ( n398709 , n51311 );
nand ( n51313 , n51172 , n398560 );
buf ( n398711 , n51313 );
nand ( n51315 , n398709 , n398711 );
buf ( n398713 , n51315 );
buf ( n398714 , n398713 );
not ( n51318 , n398714 );
or ( n51319 , n51154 , n51318 );
buf ( n398717 , n398555 );
buf ( n398718 , n398713 );
or ( n51322 , n398717 , n398718 );
not ( n51323 , n388102 );
buf ( n398721 , n49525 );
not ( n51325 , n398721 );
buf ( n398723 , n51325 );
not ( n51327 , n398723 );
or ( n51328 , n51323 , n51327 );
buf ( n398726 , n49525 );
buf ( n398727 , n388105 );
nand ( n51331 , n398726 , n398727 );
buf ( n398729 , n51331 );
nand ( n51333 , n51328 , n398729 );
and ( n51334 , n51333 , n43286 );
and ( n51335 , n50202 , n390362 );
nor ( n51336 , n51334 , n51335 );
not ( n51337 , n51336 );
not ( n51338 , n51337 );
buf ( n398736 , n49117 );
not ( n51340 , n398736 );
buf ( n398738 , n35435 );
not ( n51342 , n398738 );
buf ( n398740 , n51342 );
buf ( n398741 , n398740 );
not ( n51345 , n398741 );
or ( n51346 , n51340 , n51345 );
nand ( n51347 , n49124 , n40711 );
buf ( n398745 , n51347 );
nand ( n51349 , n51346 , n398745 );
buf ( n398747 , n51349 );
buf ( n398748 , n398747 );
not ( n51352 , n398748 );
buf ( n398750 , n396868 );
not ( n51354 , n398750 );
or ( n51355 , n51352 , n51354 );
buf ( n398753 , n383137 );
buf ( n398754 , n397839 );
nand ( n51358 , n398753 , n398754 );
buf ( n398756 , n51358 );
buf ( n398757 , n398756 );
nand ( n51361 , n51355 , n398757 );
buf ( n398759 , n51361 );
buf ( n398760 , n398759 );
or ( n51364 , n50248 , n391176 );
buf ( n398762 , n392611 );
buf ( n398763 , n388576 );
and ( n51367 , n398762 , n398763 );
not ( n51368 , n398762 );
buf ( n398766 , n388556 );
and ( n51370 , n51368 , n398766 );
nor ( n51371 , n51367 , n51370 );
buf ( n398769 , n51371 );
or ( n51373 , n398769 , n391164 );
nand ( n51374 , n51364 , n51373 );
buf ( n398772 , n51374 );
or ( n51376 , n398760 , n398772 );
buf ( n398774 , n51376 );
buf ( n398775 , n398774 );
and ( n51379 , n388263 , n388215 );
not ( n51380 , n388263 );
and ( n51381 , n51380 , n388998 );
or ( n51382 , n51379 , n51381 );
not ( n51383 , n51382 );
not ( n51384 , n383891 );
or ( n51385 , n51383 , n51384 );
buf ( n398783 , n388626 );
not ( n51387 , n398783 );
buf ( n398785 , n397797 );
nand ( n51389 , n51387 , n398785 );
buf ( n398787 , n51389 );
nand ( n51391 , n51385 , n398787 );
buf ( n398789 , n51391 );
not ( n51393 , n398789 );
buf ( n398791 , n40839 );
buf ( n398792 , n390460 );
nand ( n51396 , n398791 , n398792 );
buf ( n398794 , n51396 );
nand ( n51398 , n40990 , n36395 );
nand ( n51399 , n398794 , n51398 );
not ( n51400 , n51399 );
not ( n51401 , n397165 );
or ( n51402 , n51400 , n51401 );
nand ( n51403 , n36363 , n398402 );
nand ( n51404 , n51402 , n51403 );
buf ( n398802 , n51404 );
not ( n51406 , n398802 );
or ( n51407 , n51393 , n51406 );
buf ( n398805 , n51391 );
not ( n51409 , n398805 );
buf ( n398807 , n51409 );
buf ( n398808 , n398807 );
not ( n51412 , n398808 );
buf ( n398810 , n51404 );
not ( n51414 , n398810 );
buf ( n398812 , n51414 );
buf ( n398813 , n398812 );
not ( n51417 , n398813 );
or ( n51418 , n51412 , n51417 );
not ( n51419 , n40858 );
buf ( n398817 , n51419 );
not ( n51421 , n398817 );
buf ( n398819 , n389356 );
buf ( n398820 , n40943 );
and ( n51424 , n398819 , n398820 );
not ( n51425 , n398819 );
buf ( n398823 , n40890 );
and ( n51427 , n51425 , n398823 );
nor ( n51428 , n51424 , n51427 );
buf ( n398826 , n51428 );
buf ( n398827 , n398826 );
not ( n51431 , n398827 );
and ( n51432 , n51421 , n51431 );
buf ( n398830 , n398245 );
not ( n51434 , n398830 );
buf ( n398832 , n36845 );
nor ( n51436 , n51434 , n398832 );
buf ( n398834 , n51436 );
buf ( n398835 , n398834 );
nor ( n51439 , n51432 , n398835 );
buf ( n398837 , n51439 );
not ( n51441 , n398837 );
buf ( n398839 , n51441 );
nand ( n51443 , n51418 , n398839 );
buf ( n398841 , n51443 );
buf ( n398842 , n398841 );
nand ( n51446 , n51407 , n398842 );
buf ( n398844 , n51446 );
buf ( n398845 , n398844 );
and ( n51449 , n398775 , n398845 );
buf ( n398847 , n398759 );
buf ( n398848 , n51374 );
and ( n51452 , n398847 , n398848 );
buf ( n398850 , n51452 );
buf ( n398851 , n398850 );
nor ( n51455 , n51449 , n398851 );
buf ( n398853 , n51455 );
buf ( n398854 , n398853 );
not ( n51458 , n398854 );
buf ( n398856 , n51458 );
not ( n51460 , n398856 );
or ( n51461 , n51338 , n51460 );
buf ( n398859 , n51336 );
not ( n51463 , n398859 );
buf ( n398861 , n398853 );
not ( n51465 , n398861 );
or ( n51466 , n51463 , n51465 );
xor ( n51467 , n397662 , n397669 );
xor ( n51468 , n51467 , n397686 );
buf ( n398866 , n51468 );
buf ( n398867 , n398866 );
nand ( n51471 , n51466 , n398867 );
buf ( n398869 , n51471 );
nand ( n51473 , n51461 , n398869 );
buf ( n398871 , n51473 );
nand ( n51475 , n51322 , n398871 );
buf ( n398873 , n51475 );
buf ( n398874 , n398873 );
nand ( n51478 , n51319 , n398874 );
buf ( n398876 , n51478 );
buf ( n398877 , n389341 );
not ( n51481 , n398877 );
buf ( n398879 , n42390 );
not ( n51483 , n398879 );
or ( n51484 , n51481 , n51483 );
buf ( n398882 , n390498 );
buf ( n398883 , n393185 );
nand ( n51487 , n398882 , n398883 );
buf ( n398885 , n51487 );
buf ( n398886 , n398885 );
nand ( n51490 , n51484 , n398886 );
buf ( n398888 , n51490 );
buf ( n398889 , n398888 );
not ( n51493 , n398889 );
buf ( n398891 , n392659 );
not ( n51495 , n398891 );
or ( n51496 , n51493 , n51495 );
not ( n51497 , n397648 );
nand ( n51498 , n51497 , n384554 );
buf ( n398896 , n51498 );
nand ( n51500 , n51496 , n398896 );
buf ( n398898 , n51500 );
not ( n51502 , n388833 );
not ( n51503 , n50394 );
or ( n51504 , n51502 , n51503 );
buf ( n398902 , n388872 );
not ( n51506 , n41349 );
not ( n51507 , n37763 );
or ( n51508 , n51506 , n51507 );
nand ( n51509 , n41342 , n394426 );
nand ( n51510 , n51508 , n51509 );
buf ( n398908 , n51510 );
nand ( n51512 , n398902 , n398908 );
buf ( n398910 , n51512 );
nand ( n51514 , n51504 , n398910 );
or ( n51515 , n398898 , n51514 );
and ( n51516 , n50332 , n397781 );
not ( n51517 , n50332 );
and ( n51518 , n51517 , n50351 );
or ( n51519 , n51516 , n51518 );
and ( n51520 , n51519 , n50377 );
not ( n51521 , n51519 );
not ( n51522 , n50377 );
and ( n51523 , n51521 , n51522 );
nor ( n51524 , n51520 , n51523 );
and ( n51525 , n51515 , n51524 );
buf ( n398923 , n51514 );
buf ( n398924 , n398898 );
and ( n51528 , n398923 , n398924 );
buf ( n398926 , n51528 );
nor ( n51530 , n51525 , n398926 );
buf ( n398928 , n51530 );
buf ( n398929 , n50579 );
not ( n51533 , n398929 );
buf ( n398931 , n47891 );
not ( n51535 , n398931 );
buf ( n398933 , n382529 );
not ( n51537 , n398933 );
or ( n51538 , n51535 , n51537 );
buf ( n398936 , n390351 );
not ( n51540 , n398936 );
buf ( n398938 , n51540 );
buf ( n398939 , n398938 );
buf ( n398940 , n50584 );
nand ( n51544 , n398939 , n398940 );
buf ( n398942 , n51544 );
buf ( n398943 , n398942 );
nand ( n51547 , n51538 , n398943 );
buf ( n398945 , n51547 );
buf ( n398946 , n398945 );
not ( n51550 , n398946 );
or ( n51551 , n51533 , n51550 );
buf ( n398949 , n398002 );
not ( n51553 , n50564 );
buf ( n398951 , n51553 );
nand ( n51555 , n398949 , n398951 );
buf ( n398953 , n51555 );
buf ( n398954 , n398953 );
nand ( n398955 , n51551 , n398954 );
buf ( n398956 , n398955 );
buf ( n398957 , n398956 );
not ( n51561 , n398957 );
buf ( n398959 , n51561 );
buf ( n398960 , n398959 );
xor ( n51564 , n398928 , n398960 );
xor ( n51565 , n50383 , n397826 );
xor ( n51566 , n51565 , n397852 );
buf ( n398964 , n51566 );
and ( n51568 , n51564 , n398964 );
and ( n51569 , n398928 , n398960 );
or ( n51570 , n51568 , n51569 );
buf ( n398968 , n51570 );
buf ( n398969 , n398968 );
not ( n51573 , n398969 );
buf ( n398971 , n51573 );
buf ( n398972 , n398971 );
not ( n51576 , n398972 );
buf ( n398974 , n397617 );
buf ( n398975 , n397697 );
xor ( n51579 , n398974 , n398975 );
buf ( n398977 , n397690 );
xor ( n51581 , n51579 , n398977 );
buf ( n398979 , n51581 );
buf ( n398980 , n398979 );
not ( n51584 , n398980 );
or ( n51585 , n51576 , n51584 );
buf ( n398983 , n398968 );
not ( n51587 , n398983 );
buf ( n398985 , n398979 );
not ( n51589 , n398985 );
buf ( n398987 , n51589 );
buf ( n398988 , n398987 );
not ( n51592 , n398988 );
or ( n51593 , n51587 , n51592 );
xor ( n51594 , n398206 , n398320 );
xor ( n51595 , n51594 , n398345 );
buf ( n398993 , n51595 );
not ( n51597 , n392740 );
not ( n51598 , n398175 );
or ( n51599 , n51597 , n51598 );
buf ( n398997 , n392247 );
not ( n51601 , n398997 );
buf ( n398999 , n49933 );
not ( n51603 , n398999 );
or ( n51604 , n51601 , n51603 );
buf ( n399002 , n49938 );
buf ( n399003 , n392244 );
nand ( n51607 , n399002 , n399003 );
buf ( n399005 , n51607 );
buf ( n399006 , n399005 );
nand ( n51610 , n51604 , n399006 );
buf ( n399008 , n51610 );
buf ( n399009 , n399008 );
buf ( n399010 , n45260 );
nand ( n51614 , n399009 , n399010 );
buf ( n399012 , n51614 );
nand ( n51616 , n51599 , n399012 );
xor ( n51617 , n398993 , n51616 );
buf ( n399015 , n49686 );
not ( n51619 , n399015 );
buf ( n399017 , n49661 );
not ( n51621 , n399017 );
or ( n51622 , n51619 , n51621 );
buf ( n399020 , n49653 );
buf ( n399021 , n46478 );
nand ( n51625 , n399020 , n399021 );
buf ( n399023 , n51625 );
buf ( n399024 , n399023 );
nand ( n51628 , n51622 , n399024 );
buf ( n399026 , n51628 );
buf ( n399027 , n399026 );
not ( n51631 , n399027 );
buf ( n399029 , n38960 );
not ( n51633 , n399029 );
buf ( n399031 , n51633 );
buf ( n399032 , n399031 );
not ( n51636 , n399032 );
or ( n51637 , n51631 , n51636 );
buf ( n399035 , n397099 );
buf ( n399036 , n395199 );
nand ( n51640 , n399035 , n399036 );
buf ( n399038 , n51640 );
buf ( n399039 , n399038 );
nand ( n51643 , n51637 , n399039 );
buf ( n399041 , n51643 );
not ( n51645 , n399041 );
buf ( n399043 , n394666 );
not ( n51647 , n399043 );
not ( n51648 , n22982 );
buf ( n399046 , n51648 );
not ( n51650 , n399046 );
or ( n51651 , n51647 , n51650 );
nand ( n51652 , n49660 , n388566 );
buf ( n399050 , n51652 );
nand ( n51654 , n51651 , n399050 );
buf ( n399052 , n51654 );
buf ( n399053 , n399052 );
not ( n51657 , n399053 );
buf ( n399055 , n399031 );
not ( n51659 , n399055 );
or ( n51660 , n51657 , n51659 );
buf ( n399058 , n399026 );
buf ( n399059 , n395199 );
nand ( n51663 , n399058 , n399059 );
buf ( n399061 , n51663 );
buf ( n399062 , n399061 );
nand ( n51666 , n51660 , n399062 );
buf ( n399064 , n51666 );
buf ( n399065 , n399064 );
not ( n51669 , n399065 );
buf ( n399067 , n51669 );
nand ( n51671 , n51645 , n399067 );
not ( n51672 , n51671 );
buf ( n399070 , n388543 );
not ( n51674 , n399070 );
buf ( n399072 , n393525 );
not ( n51676 , n399072 );
or ( n51677 , n51674 , n51676 );
buf ( n399075 , n388962 );
buf ( n399076 , n388546 );
nand ( n51680 , n399075 , n399076 );
buf ( n399078 , n51680 );
buf ( n399079 , n399078 );
nand ( n51683 , n51677 , n399079 );
buf ( n399081 , n51683 );
buf ( n399082 , n399081 );
not ( n51686 , n399082 );
buf ( n399084 , n393544 );
not ( n51688 , n399084 );
or ( n51689 , n51686 , n51688 );
buf ( n399087 , n398269 );
not ( n51691 , n46060 );
not ( n51692 , n51691 );
buf ( n399090 , n51692 );
nand ( n51694 , n399087 , n399090 );
buf ( n399092 , n51694 );
buf ( n399093 , n399092 );
nand ( n51697 , n51689 , n399093 );
buf ( n399095 , n51697 );
not ( n51699 , n399095 );
or ( n51700 , n51672 , n51699 );
buf ( n399098 , n399041 );
buf ( n399099 , n399064 );
nand ( n51703 , n399098 , n399099 );
buf ( n399101 , n51703 );
nand ( n51705 , n51700 , n399101 );
buf ( n399103 , n388872 );
not ( n51707 , n399103 );
buf ( n399105 , n41342 );
buf ( n399106 , n29077 );
and ( n51710 , n399105 , n399106 );
not ( n51711 , n399105 );
buf ( n399109 , n389802 );
and ( n51713 , n51711 , n399109 );
nor ( n51714 , n51710 , n51713 );
buf ( n399112 , n51714 );
buf ( n399113 , n399112 );
not ( n51717 , n399113 );
or ( n51718 , n51707 , n51717 );
buf ( n399116 , n51510 );
buf ( n399117 , n388833 );
nand ( n51721 , n399116 , n399117 );
buf ( n399119 , n51721 );
buf ( n399120 , n399119 );
nand ( n51724 , n51718 , n399120 );
buf ( n399122 , n51724 );
xor ( n51726 , n51705 , n399122 );
xor ( n51727 , n398257 , n398282 );
xor ( n51728 , n51727 , n398310 );
buf ( n399126 , n51728 );
and ( n51730 , n51726 , n399126 );
and ( n51731 , n51705 , n399122 );
or ( n51732 , n51730 , n51731 );
buf ( n399130 , n51732 );
buf ( n399131 , n388809 );
not ( n51735 , n399131 );
buf ( n399133 , n398373 );
not ( n51737 , n399133 );
or ( n51738 , n51735 , n51737 );
buf ( n399136 , n388760 );
not ( n51740 , n399136 );
buf ( n399138 , n386012 );
not ( n51742 , n399138 );
or ( n51743 , n51740 , n51742 );
buf ( n399141 , n38472 );
buf ( n399142 , n388757 );
nand ( n51746 , n399141 , n399142 );
buf ( n399144 , n51746 );
buf ( n399145 , n399144 );
nand ( n51749 , n51743 , n399145 );
buf ( n399147 , n51749 );
buf ( n399148 , n399147 );
buf ( n399149 , n388746 );
nand ( n51753 , n399148 , n399149 );
buf ( n399151 , n51753 );
buf ( n399152 , n399151 );
nand ( n51756 , n51738 , n399152 );
buf ( n399154 , n51756 );
buf ( n399155 , n399154 );
xor ( n51759 , n399130 , n399155 );
buf ( n399157 , n46921 );
not ( n51761 , n399157 );
buf ( n399159 , n50899 );
not ( n51763 , n399159 );
or ( n51764 , n51761 , n51763 );
buf ( n399162 , n38935 );
not ( n51766 , n399162 );
buf ( n399164 , n51766 );
buf ( n399165 , n399164 );
not ( n51769 , n399165 );
buf ( n399167 , n51769 );
not ( n51771 , n399167 );
not ( n51772 , n46114 );
or ( n51773 , n51771 , n51772 );
nand ( n51774 , n397069 , n398298 );
nand ( n51775 , n51773 , n51774 );
buf ( n399173 , n51775 );
buf ( n399174 , n396622 );
nand ( n51778 , n399173 , n399174 );
buf ( n399176 , n51778 );
buf ( n399177 , n399176 );
nand ( n51781 , n51764 , n399177 );
buf ( n399179 , n51781 );
buf ( n399180 , n399179 );
buf ( n399181 , n388230 );
not ( n51785 , n399181 );
buf ( n399183 , n391563 );
not ( n51787 , n399183 );
or ( n51788 , n51785 , n51787 );
buf ( n399186 , n393562 );
buf ( n399187 , n388242 );
nand ( n51791 , n399186 , n399187 );
buf ( n399189 , n51791 );
buf ( n399190 , n399189 );
nand ( n51794 , n51788 , n399190 );
buf ( n399192 , n51794 );
buf ( n399193 , n399192 );
not ( n51797 , n399193 );
buf ( n399195 , n37338 );
not ( n51799 , n399195 );
or ( n51800 , n51797 , n51799 );
buf ( n399198 , n398658 );
buf ( n399199 , n393100 );
nand ( n51803 , n399198 , n399199 );
buf ( n399201 , n51803 );
buf ( n399202 , n399201 );
nand ( n51806 , n51800 , n399202 );
buf ( n399204 , n51806 );
buf ( n399205 , n399204 );
or ( n51809 , n399180 , n399205 );
buf ( n399207 , n392788 );
not ( n51811 , n399207 );
buf ( n399209 , n398633 );
not ( n51813 , n399209 );
or ( n51814 , n51811 , n51813 );
buf ( n399212 , n47412 );
not ( n51816 , n399212 );
buf ( n399214 , n28215 );
not ( n51818 , n399214 );
or ( n51819 , n51816 , n51818 );
buf ( n399217 , n375822 );
not ( n51821 , n41558 );
not ( n51822 , n51821 );
buf ( n399220 , n51822 );
nand ( n51824 , n399217 , n399220 );
buf ( n399222 , n51824 );
buf ( n399223 , n399222 );
nand ( n51827 , n51819 , n399223 );
buf ( n399225 , n51827 );
buf ( n399226 , n399225 );
buf ( n399227 , n390432 );
nand ( n51831 , n399226 , n399227 );
buf ( n399229 , n51831 );
buf ( n399230 , n399229 );
nand ( n51834 , n51814 , n399230 );
buf ( n399232 , n51834 );
buf ( n399233 , n399232 );
nand ( n51837 , n51809 , n399233 );
buf ( n399235 , n51837 );
buf ( n399236 , n399235 );
buf ( n399237 , n399204 );
buf ( n399238 , n399179 );
nand ( n51842 , n399237 , n399238 );
buf ( n399240 , n51842 );
buf ( n399241 , n399240 );
nand ( n51845 , n399236 , n399241 );
buf ( n399243 , n51845 );
buf ( n399244 , n394817 );
not ( n51848 , n399244 );
buf ( n399246 , n385987 );
not ( n51850 , n399246 );
or ( n51851 , n51848 , n51850 );
buf ( n399249 , n389759 );
buf ( n399250 , n394814 );
nand ( n51854 , n399249 , n399250 );
buf ( n399252 , n51854 );
buf ( n399253 , n399252 );
nand ( n51857 , n51851 , n399253 );
buf ( n399255 , n51857 );
buf ( n399256 , n399255 );
not ( n51860 , n399256 );
buf ( n399258 , n382595 );
not ( n51862 , n399258 );
or ( n51863 , n51860 , n51862 );
buf ( n399261 , n389024 );
buf ( n399262 , n398426 );
nand ( n51866 , n399261 , n399262 );
buf ( n399264 , n51866 );
buf ( n399265 , n399264 );
nand ( n51869 , n51863 , n399265 );
buf ( n399267 , n51869 );
xor ( n51871 , n399243 , n399267 );
xor ( n51872 , n358933 , n359000 );
xor ( n51873 , n51872 , n359018 );
buf ( n399271 , n51873 );
buf ( n399272 , n399271 );
buf ( n51876 , n399272 );
buf ( n399274 , n51876 );
buf ( n399275 , n399274 );
not ( n51879 , n399275 );
buf ( n399277 , n385331 );
not ( n51881 , n399277 );
or ( n51882 , n51879 , n51881 );
buf ( n399280 , n385292 );
buf ( n399281 , n399274 );
not ( n51885 , n399281 );
buf ( n399283 , n51885 );
buf ( n399284 , n399283 );
nand ( n51888 , n399280 , n399284 );
buf ( n399286 , n51888 );
buf ( n399287 , n399286 );
nand ( n51891 , n51882 , n399287 );
buf ( n399289 , n51891 );
buf ( n399290 , n388498 );
buf ( n399291 , n398596 );
or ( n51900 , n399290 , n399291 );
nand ( n51901 , C1 , n51900 );
buf ( n399294 , n51901 );
and ( n51903 , n51871 , n399294 );
and ( n51904 , n399243 , n399267 );
or ( n51905 , n51903 , n51904 );
buf ( n399298 , n51905 );
and ( n51907 , n51759 , n399298 );
and ( n51908 , n399130 , n399155 );
or ( n51909 , n51907 , n51908 );
buf ( n399302 , n51909 );
and ( n51911 , n51617 , n399302 );
and ( n51912 , n398993 , n51616 );
or ( n51913 , n51911 , n51912 );
buf ( n399306 , n51913 );
nand ( n51915 , n51593 , n399306 );
buf ( n399308 , n51915 );
buf ( n399309 , n399308 );
nand ( n51918 , n51585 , n399309 );
buf ( n399311 , n51918 );
xor ( n51920 , n398876 , n399311 );
buf ( n399313 , n50610 );
buf ( n399314 , n398038 );
xor ( n51923 , n399313 , n399314 );
buf ( n399316 , n398024 );
xor ( n51925 , n51923 , n399316 );
buf ( n399318 , n51925 );
and ( n51927 , n51920 , n399318 );
and ( n51928 , n398876 , n399311 );
or ( n51929 , n51927 , n51928 );
not ( n51930 , n51929 );
xor ( n51931 , n398044 , n397897 );
xor ( n51932 , n51931 , n398051 );
buf ( n399325 , n397600 );
buf ( n399326 , n397607 );
xor ( n51935 , n399325 , n399326 );
buf ( n399328 , n397881 );
xor ( n51937 , n51935 , n399328 );
buf ( n399330 , n51937 );
nand ( n51939 , n51932 , n399330 );
not ( n51940 , n51939 );
or ( n51941 , n51930 , n51940 );
buf ( n399334 , n399330 );
not ( n51943 , n399334 );
not ( n51944 , n51932 );
buf ( n399337 , n51944 );
nand ( n51946 , n51943 , n399337 );
buf ( n399339 , n51946 );
nand ( n51948 , n51941 , n399339 );
buf ( n399341 , n398101 );
buf ( n399342 , n398528 );
nand ( n51951 , n399341 , n399342 );
buf ( n399344 , n51951 );
and ( n51953 , n51948 , n399344 );
nor ( n51954 , n51127 , n51953 );
buf ( n399347 , n51954 );
not ( n51956 , n399347 );
buf ( n399349 , n51956 );
nand ( n51958 , n50692 , n399349 );
nand ( n51959 , n50688 , n51958 );
not ( n51960 , n51959 );
nand ( n51961 , n50675 , n51960 );
xor ( n51962 , n398066 , n398067 );
buf ( n399355 , n51962 );
buf ( n399356 , n399355 );
buf ( n399357 , n398063 );
xor ( n51966 , n399356 , n399357 );
buf ( n399359 , n51966 );
buf ( n399360 , n399359 );
xor ( n51969 , n398471 , n398481 );
xor ( n51970 , n51969 , n398524 );
buf ( n399363 , n51970 );
not ( n51972 , n399363 );
xor ( n51973 , n398464 , n398465 );
buf ( n399366 , n51973 );
xnor ( n51975 , n399366 , n398461 );
buf ( n399368 , n51975 );
not ( n51977 , n399368 );
buf ( n399370 , n51977 );
buf ( n399371 , n399370 );
not ( n51980 , n399371 );
xor ( n51981 , n398494 , n398517 );
xor ( n51982 , n51981 , n51117 );
not ( n51983 , n51982 );
buf ( n399376 , n51983 );
not ( n51985 , n399376 );
or ( n51986 , n51980 , n51985 );
buf ( n399379 , n51975 );
not ( n51988 , n399379 );
buf ( n399381 , n51982 );
not ( n51990 , n399381 );
or ( n51991 , n51988 , n51990 );
xor ( n51992 , n397927 , n398005 );
not ( n51993 , n397951 );
xor ( n51994 , n51992 , n51993 );
buf ( n399387 , n51994 );
xor ( n51996 , n50443 , n397737 );
xor ( n51997 , n51996 , n50428 );
buf ( n399390 , n51997 );
xor ( n51999 , n399387 , n399390 );
xor ( n52000 , n398231 , n398252 );
xor ( n52001 , n52000 , n398315 );
buf ( n399394 , n52001 );
buf ( n399395 , n399394 );
buf ( n399396 , n389162 );
not ( n52005 , n399396 );
buf ( n399398 , n398334 );
not ( n52007 , n399398 );
or ( n52008 , n52005 , n52007 );
buf ( n399401 , n41671 );
not ( n52010 , n399401 );
buf ( n399403 , n384089 );
not ( n52012 , n399403 );
or ( n52013 , n52010 , n52012 );
buf ( n399406 , n36509 );
buf ( n399407 , n41678 );
nand ( n52016 , n399406 , n399407 );
buf ( n399409 , n52016 );
buf ( n399410 , n399409 );
nand ( n52019 , n52013 , n399410 );
buf ( n399412 , n52019 );
buf ( n399413 , n399412 );
buf ( n399414 , n41711 );
nand ( n52023 , n399413 , n399414 );
buf ( n399416 , n52023 );
buf ( n399417 , n399416 );
nand ( n52026 , n52008 , n399417 );
buf ( n399419 , n52026 );
buf ( n399420 , n399419 );
xor ( n52029 , n399395 , n399420 );
xor ( n52030 , n398604 , n398622 );
xor ( n52031 , n52030 , n398703 );
buf ( n399424 , n52031 );
buf ( n399425 , n399424 );
and ( n52034 , n52029 , n399425 );
and ( n52035 , n399395 , n399420 );
or ( n52036 , n52034 , n52035 );
buf ( n399429 , n52036 );
buf ( n399430 , n399429 );
buf ( n399431 , n395349 );
not ( n52040 , n399431 );
buf ( n399433 , n47863 );
not ( n52042 , n399433 );
buf ( n399435 , n386424 );
not ( n52044 , n399435 );
or ( n52045 , n52042 , n52044 );
buf ( n399438 , n386418 );
buf ( n399439 , n395312 );
nand ( n52048 , n399438 , n399439 );
buf ( n399441 , n52048 );
buf ( n399442 , n399441 );
nand ( n52051 , n52045 , n399442 );
buf ( n399444 , n52051 );
buf ( n399445 , n399444 );
not ( n52054 , n399445 );
or ( n52055 , n52040 , n52054 );
buf ( n399448 , n397920 );
buf ( n399449 , n395362 );
nand ( n52058 , n399448 , n399449 );
buf ( n399451 , n52058 );
buf ( n399452 , n399451 );
nand ( n52061 , n52055 , n399452 );
buf ( n399454 , n52061 );
buf ( n399455 , n399454 );
xor ( n52064 , n399430 , n399455 );
buf ( n399457 , n391446 );
buf ( n399458 , n42390 );
and ( n52067 , n399457 , n399458 );
not ( n52068 , n399457 );
buf ( n399461 , n391870 );
and ( n52070 , n52068 , n399461 );
nor ( n52071 , n52067 , n52070 );
buf ( n399464 , n52071 );
buf ( n399465 , n399464 );
not ( n52074 , n399465 );
buf ( n399467 , n52074 );
buf ( n399468 , n399467 );
not ( n52077 , n399468 );
buf ( n399470 , n389880 );
not ( n52079 , n399470 );
or ( n52080 , n52077 , n52079 );
buf ( n399473 , n398888 );
buf ( n399474 , n391638 );
nand ( n52083 , n399473 , n399474 );
buf ( n399476 , n52083 );
buf ( n399477 , n399476 );
nand ( n52086 , n52080 , n399477 );
buf ( n399479 , n52086 );
buf ( n399480 , n399479 );
not ( n52089 , n399480 );
buf ( n399482 , n52089 );
buf ( n399483 , n399482 );
not ( n52092 , n399483 );
not ( n52093 , n41711 );
buf ( n399486 , n41671 );
not ( n52095 , n399486 );
buf ( n399488 , n38660 );
not ( n52097 , n399488 );
or ( n52098 , n52095 , n52097 );
buf ( n399491 , n36564 );
buf ( n399492 , n41678 );
nand ( n52101 , n399491 , n399492 );
buf ( n399494 , n52101 );
buf ( n399495 , n399494 );
nand ( n52104 , n52098 , n399495 );
buf ( n399497 , n52104 );
not ( n52106 , n399497 );
or ( n52107 , n52093 , n52106 );
buf ( n399500 , n399412 );
buf ( n399501 , n389162 );
nand ( n52110 , n399500 , n399501 );
buf ( n399503 , n52110 );
nand ( n399504 , n52107 , n399503 );
not ( n52113 , n399504 );
buf ( n399506 , n52113 );
not ( n52115 , n399506 );
or ( n52116 , n52092 , n52115 );
xor ( n52117 , n398644 , n398675 );
xor ( n52118 , n52117 , n398698 );
buf ( n399511 , n52118 );
buf ( n399512 , n399511 );
nand ( n52121 , n52116 , n399512 );
buf ( n399514 , n52121 );
buf ( n399515 , n399514 );
buf ( n399516 , n399504 );
buf ( n399517 , n399479 );
nand ( n52126 , n399516 , n399517 );
buf ( n399519 , n52126 );
buf ( n399520 , n399519 );
nand ( n52129 , n399515 , n399520 );
buf ( n399522 , n52129 );
buf ( n399523 , n399522 );
xor ( n52132 , n398389 , n51010 );
xor ( n52133 , n52132 , n398441 );
buf ( n399526 , n52133 );
xor ( n52135 , n399523 , n399526 );
not ( n52136 , n43515 );
not ( n52137 , n51165 );
or ( n52138 , n52136 , n52137 );
not ( n52139 , n43537 );
buf ( n399532 , n391027 );
buf ( n399533 , n384741 );
and ( n52142 , n399532 , n399533 );
not ( n52143 , n399532 );
buf ( n399536 , n384741 );
not ( n52145 , n399536 );
buf ( n399538 , n52145 );
buf ( n399539 , n399538 );
and ( n52148 , n52143 , n399539 );
nor ( n52149 , n52142 , n52148 );
buf ( n399542 , n52149 );
nand ( n52151 , n52139 , n399542 );
nand ( n52152 , n52138 , n52151 );
buf ( n399545 , n52152 );
and ( n52154 , n52135 , n399545 );
and ( n52155 , n399523 , n399526 );
or ( n52156 , n52154 , n52155 );
buf ( n399549 , n52156 );
buf ( n399550 , n399549 );
and ( n52159 , n52064 , n399550 );
and ( n52160 , n399430 , n399455 );
or ( n52161 , n52159 , n52160 );
buf ( n399554 , n52161 );
buf ( n399555 , n399554 );
and ( n52164 , n51999 , n399555 );
and ( n52165 , n399387 , n399390 );
or ( n52166 , n52164 , n52165 );
buf ( n399559 , n52166 );
buf ( n399560 , n399559 );
nand ( n52169 , n51991 , n399560 );
buf ( n399562 , n52169 );
buf ( n399563 , n399562 );
nand ( n52172 , n51986 , n399563 );
buf ( n399565 , n52172 );
buf ( n399566 , n399565 );
not ( n52175 , n399566 );
buf ( n399568 , n52175 );
not ( n52177 , n399568 );
or ( n52178 , n51972 , n52177 );
buf ( n399571 , n398349 );
buf ( n399572 , n398201 );
xor ( n52181 , n399571 , n399572 );
buf ( n399574 , n398450 );
xnor ( n52183 , n52181 , n399574 );
buf ( n399576 , n52183 );
buf ( n399577 , n399576 );
xor ( n52186 , n398707 , n398560 );
xnor ( n52187 , n52186 , n51172 );
not ( n52188 , n52187 );
not ( n52189 , n393825 );
buf ( n399582 , n35301 );
buf ( n399583 , n393384 );
nand ( n52192 , n399582 , n399583 );
buf ( n399585 , n52192 );
nand ( n52194 , n398116 , n386385 );
nand ( n52195 , n399585 , n52194 );
not ( n52196 , n52195 );
or ( n52197 , n52189 , n52196 );
buf ( n399590 , n398128 );
buf ( n399591 , n45954 );
nand ( n52200 , n399590 , n399591 );
buf ( n399593 , n52200 );
nand ( n52202 , n52197 , n399593 );
not ( n52203 , n52202 );
not ( n52204 , n52203 );
and ( n52205 , n52188 , n52204 );
buf ( n399598 , n52187 );
buf ( n399599 , n52203 );
nand ( n52208 , n399598 , n399599 );
buf ( n399601 , n52208 );
and ( n52210 , n50977 , n50952 );
not ( n52211 , n50977 );
not ( n52212 , n50952 );
and ( n52213 , n52211 , n52212 );
nor ( n52214 , n52210 , n52213 );
and ( n52215 , n52214 , n51041 );
not ( n52216 , n52214 );
not ( n52217 , n51041 );
and ( n52218 , n52216 , n52217 );
nor ( n52219 , n52215 , n52218 );
not ( n52220 , n52219 );
not ( n52221 , n52220 );
and ( n52222 , n399601 , n52221 );
nor ( n52223 , n52205 , n52222 );
buf ( n399616 , n52223 );
xor ( n52225 , n399577 , n399616 );
xor ( n52226 , n398713 , n398552 );
xor ( n52227 , n52226 , n51473 );
buf ( n399620 , n52227 );
and ( n52229 , n52225 , n399620 );
and ( n52230 , n399577 , n399616 );
or ( n52231 , n52229 , n52230 );
buf ( n399624 , n52231 );
not ( n52233 , n399624 );
xor ( n52234 , n50752 , n398190 );
xor ( n52235 , n52234 , n398182 );
buf ( n399628 , n52235 );
xor ( n52237 , n398928 , n398960 );
xor ( n52238 , n52237 , n398964 );
buf ( n399631 , n52238 );
not ( n52240 , n399631 );
buf ( n399633 , n51553 );
not ( n52242 , n399633 );
buf ( n399635 , n398945 );
not ( n52244 , n399635 );
or ( n52245 , n52242 , n52244 );
not ( n52246 , n397990 );
not ( n52247 , n38532 );
or ( n52248 , n52246 , n52247 );
buf ( n399641 , n35519 );
buf ( n399642 , n50584 );
nand ( n52251 , n399641 , n399642 );
buf ( n399644 , n52251 );
nand ( n52253 , n52248 , n399644 );
nand ( n52254 , n52253 , n50579 );
buf ( n399647 , n52254 );
nand ( n52256 , n52245 , n399647 );
buf ( n399649 , n52256 );
not ( n52258 , n399649 );
buf ( n399651 , n391032 );
not ( n52274 , n399651 );
buf ( n399653 , n52274 );
buf ( n399654 , C1 );
or ( n52339 , n52258 , C0 );
xor ( n52343 , n398847 , n398848 );
buf ( n399657 , n52343 );
xor ( n52345 , n398844 , n399657 );
nand ( n52346 , C1 , n52345 );
nand ( n52347 , n52339 , n52346 );
not ( n52348 , n52347 );
not ( n52349 , n52348 );
or ( n52350 , n52240 , n52349 );
nor ( n52351 , n52348 , n399631 );
not ( n52352 , n390362 );
not ( n52353 , n51333 );
or ( n52354 , n52352 , n52353 );
buf ( n399668 , n388102 );
not ( n52356 , n399668 );
buf ( n399670 , n37215 );
not ( n52358 , n399670 );
or ( n52359 , n52356 , n52358 );
buf ( n399673 , n36216 );
buf ( n399674 , n388105 );
nand ( n52362 , n399673 , n399674 );
buf ( n399676 , n52362 );
buf ( n399677 , n399676 );
nand ( n52365 , n52359 , n399677 );
buf ( n399679 , n52365 );
buf ( n399680 , n399679 );
buf ( n399681 , n43286 );
nand ( n52369 , n399680 , n399681 );
buf ( n399683 , n52369 );
nand ( n52371 , n52354 , n399683 );
buf ( n399685 , n52371 );
xor ( n52373 , n398923 , n398924 );
buf ( n399687 , n52373 );
and ( n52375 , n399687 , n51524 );
not ( n52376 , n399687 );
not ( n52377 , n51524 );
and ( n52378 , n52376 , n52377 );
nor ( n52379 , n52375 , n52378 );
buf ( n399693 , n52379 );
xor ( n52381 , n399685 , n399693 );
not ( n52382 , n390635 );
not ( n52383 , n398747 );
or ( n52384 , n52382 , n52383 );
and ( n52385 , n397498 , n390453 );
not ( n52386 , n397498 );
and ( n52387 , n52386 , n35435 );
or ( n52388 , n52385 , n52387 );
nand ( n52389 , n38765 , n52388 );
nand ( n52390 , n52384 , n52389 );
buf ( n399704 , n52390 );
buf ( n399705 , n392884 );
buf ( n399706 , n388556 );
not ( n52394 , n399706 );
xor ( n52395 , n399705 , n52394 );
buf ( n399709 , n52395 );
buf ( n399710 , n399709 );
not ( n52398 , n399710 );
buf ( n399712 , n52398 );
buf ( n399713 , n399712 );
not ( n52401 , n399713 );
buf ( n399715 , n391652 );
not ( n52403 , n399715 );
or ( n52404 , n52401 , n52403 );
buf ( n399718 , n398769 );
not ( n52406 , n399718 );
buf ( n399720 , n391173 );
nand ( n52408 , n52406 , n399720 );
buf ( n399722 , n52408 );
buf ( n399723 , n399722 );
nand ( n52411 , n52404 , n399723 );
buf ( n399725 , n52411 );
buf ( n399726 , n399725 );
xor ( n52414 , n399704 , n399726 );
buf ( n399728 , n388502 );
not ( n52416 , n399728 );
buf ( n399730 , n389936 );
not ( n52418 , n399730 );
or ( n52419 , n52416 , n52418 );
buf ( n399733 , n40775 );
buf ( n399734 , n388511 );
nand ( n52422 , n399733 , n399734 );
buf ( n399736 , n52422 );
buf ( n399737 , n399736 );
nand ( n52425 , n52419 , n399737 );
buf ( n399739 , n52425 );
buf ( n399740 , n399739 );
not ( n52428 , n399740 );
buf ( n399742 , n383891 );
not ( n52430 , n399742 );
or ( n52431 , n52428 , n52430 );
nand ( n52432 , n391602 , n51382 );
buf ( n399746 , n52432 );
nand ( n52434 , n52431 , n399746 );
buf ( n399748 , n52434 );
buf ( n399749 , n399748 );
buf ( n399750 , n47726 );
not ( n52438 , n399750 );
buf ( n399752 , n398690 );
not ( n52440 , n399752 );
or ( n52441 , n52438 , n52440 );
buf ( n399755 , n40758 );
not ( n52443 , n399755 );
buf ( n399757 , n388154 );
not ( n52445 , n399757 );
and ( n52446 , n52443 , n52445 );
buf ( n399760 , n40778 );
buf ( n399761 , n388154 );
and ( n52449 , n399760 , n399761 );
nor ( n52450 , n52446 , n52449 );
buf ( n399764 , n52450 );
buf ( n399765 , n399764 );
not ( n52453 , n399765 );
buf ( n399767 , n397476 );
nand ( n52455 , n52453 , n399767 );
buf ( n399769 , n52455 );
buf ( n399770 , n399769 );
nand ( n52458 , n52441 , n399770 );
buf ( n399772 , n52458 );
buf ( n399773 , n399772 );
xor ( n52461 , n399749 , n399773 );
buf ( n399775 , n42073 );
not ( n52463 , n399775 );
buf ( n399777 , n47256 );
not ( n52465 , n399777 );
or ( n52466 , n52463 , n52465 );
buf ( n399780 , n36396 );
buf ( n399781 , n42074 );
nand ( n52469 , n399780 , n399781 );
buf ( n399783 , n52469 );
buf ( n399784 , n399783 );
nand ( n52472 , n52466 , n399784 );
buf ( n399786 , n52472 );
buf ( n399787 , n399786 );
not ( n52475 , n399787 );
buf ( n399789 , n390832 );
not ( n52477 , n399789 );
or ( n52478 , n52475 , n52477 );
nand ( n52479 , n51399 , n388346 );
buf ( n399793 , n52479 );
nand ( n52481 , n52478 , n399793 );
buf ( n399795 , n52481 );
buf ( n399796 , n399795 );
and ( n52484 , n52461 , n399796 );
and ( n52485 , n399749 , n399773 );
or ( n52486 , n52484 , n52485 );
buf ( n399800 , n52486 );
buf ( n399801 , n399800 );
and ( n52489 , n52414 , n399801 );
and ( n52490 , n399704 , n399726 );
or ( n52491 , n52489 , n52490 );
buf ( n399805 , n52491 );
buf ( n399806 , n399805 );
and ( n52494 , n52381 , n399806 );
and ( n52495 , n399685 , n399693 );
or ( n52496 , n52494 , n52495 );
buf ( n399810 , n52496 );
or ( n52498 , n52351 , n399810 );
nand ( n52499 , n52350 , n52498 );
buf ( n399813 , n52499 );
xor ( n52501 , n399628 , n399813 );
buf ( n399815 , n398979 );
buf ( n399816 , n398971 );
and ( n52504 , n399815 , n399816 );
not ( n52505 , n399815 );
buf ( n399819 , n398968 );
and ( n52507 , n52505 , n399819 );
nor ( n52508 , n52504 , n52507 );
buf ( n399822 , n52508 );
xnor ( n52510 , n399822 , n51913 );
buf ( n399824 , n52510 );
and ( n52512 , n52501 , n399824 );
and ( n52513 , n399628 , n399813 );
or ( n52514 , n52512 , n52513 );
buf ( n399828 , n52514 );
not ( n52516 , n399828 );
or ( n52517 , n52233 , n52516 );
xor ( n52518 , n398876 , n399311 );
xor ( n52519 , n52518 , n399318 );
nand ( n52520 , n52517 , n52519 );
not ( n52521 , n399624 );
buf ( n399835 , n399828 );
not ( n52523 , n399835 );
buf ( n399837 , n52523 );
nand ( n52525 , n52521 , n399837 );
nand ( n52526 , n52520 , n52525 );
nand ( n52527 , n52178 , n52526 );
buf ( n399841 , n52527 );
buf ( n399842 , n399363 );
not ( n52530 , n399842 );
buf ( n399844 , n399565 );
nand ( n52532 , n52530 , n399844 );
buf ( n399846 , n52532 );
buf ( n399847 , n399846 );
nand ( n52535 , n399841 , n399847 );
buf ( n399849 , n52535 );
buf ( n399850 , n399849 );
xor ( n52538 , n399360 , n399850 );
buf ( n399852 , n51948 );
not ( n52540 , n399852 );
xnor ( n52541 , n398101 , n398528 );
buf ( n399855 , n52541 );
not ( n52543 , n399855 );
or ( n52544 , n52540 , n52543 );
buf ( n399858 , n51948 );
buf ( n399859 , n52541 );
or ( n52547 , n399858 , n399859 );
nand ( n52548 , n52544 , n52547 );
buf ( n399862 , n52548 );
buf ( n399863 , n399862 );
and ( n52551 , n52538 , n399863 );
and ( n52552 , n399360 , n399850 );
or ( n52553 , n52551 , n52552 );
buf ( n399867 , n52553 );
buf ( n399868 , n399867 );
not ( n52556 , n399868 );
buf ( n399870 , n52556 );
not ( n52558 , n398084 );
not ( n52559 , n51954 );
not ( n52560 , n52559 );
or ( n52561 , n52558 , n52560 );
nand ( n52562 , n50689 , n51954 );
nand ( n52563 , n52561 , n52562 );
not ( n52564 , n398088 );
and ( n52565 , n52563 , n52564 );
not ( n52566 , n52563 );
not ( n52567 , n50686 );
and ( n52568 , n52566 , n52567 );
nor ( n52569 , n52565 , n52568 );
nand ( n52570 , n399870 , n52569 );
nand ( n52571 , n51961 , n52570 );
not ( n52572 , n52571 );
buf ( n399886 , n52572 );
buf ( n399887 , n393732 );
buf ( n399888 , n393864 );
xor ( n52576 , n399887 , n399888 );
buf ( n399890 , n393737 );
xnor ( n52578 , n52576 , n399890 );
buf ( n399892 , n52578 );
buf ( n399893 , n399892 );
buf ( n399894 , n49281 );
not ( n52582 , n399894 );
buf ( n399896 , n48772 );
not ( n52584 , n399896 );
or ( n52585 , n52582 , n52584 );
buf ( n399899 , n49907 );
buf ( n399900 , n48772 );
not ( n52588 , n399900 );
buf ( n399902 , n396718 );
nand ( n52590 , n52588 , n399902 );
buf ( n399904 , n52590 );
buf ( n399905 , n399904 );
nand ( n52593 , n399899 , n399905 );
buf ( n399907 , n52593 );
buf ( n399908 , n399907 );
nand ( n52596 , n52585 , n399908 );
buf ( n399910 , n52596 );
buf ( n399911 , n399910 );
not ( n52599 , n399911 );
buf ( n399913 , n52599 );
buf ( n399914 , n399913 );
xor ( n52602 , n399893 , n399914 );
xor ( n52603 , n394637 , n395060 );
xor ( n52604 , n52603 , n395613 );
buf ( n399918 , n52604 );
buf ( n399919 , n399918 );
xor ( n52607 , n52602 , n399919 );
buf ( n399921 , n52607 );
xor ( n52609 , n48753 , n49912 );
and ( n52610 , n52609 , n398077 );
and ( n52611 , n48753 , n49912 );
or ( n52612 , n52610 , n52611 );
nand ( n52613 , n399921 , n52612 );
xor ( n52614 , n394619 , n394629 );
xor ( n52615 , n52614 , n395618 );
buf ( n399929 , n52615 );
xor ( n52617 , n399893 , n399914 );
and ( n52618 , n52617 , n399919 );
and ( n52619 , n399893 , n399914 );
or ( n52620 , n52618 , n52619 );
buf ( n399934 , n52620 );
nand ( n52622 , n399929 , n399934 );
and ( n52623 , n52613 , n52622 );
buf ( n399937 , n52623 );
and ( n52625 , n399886 , n399937 );
buf ( n399939 , n52625 );
nand ( n52627 , n396187 , n399939 );
not ( n52628 , n52627 );
not ( n52629 , n399330 );
and ( n52630 , n51929 , n52629 );
not ( n52631 , n51929 );
and ( n52632 , n52631 , n399330 );
nor ( n52633 , n52630 , n52632 );
buf ( n399947 , n52633 );
not ( n52635 , n51944 );
buf ( n399949 , n52635 );
and ( n52637 , n399947 , n399949 );
not ( n52638 , n399947 );
buf ( n399952 , n51944 );
and ( n52640 , n52638 , n399952 );
nor ( n52641 , n52637 , n52640 );
buf ( n399955 , n52641 );
not ( n52643 , n399363 );
not ( n52644 , n52643 );
not ( n52645 , n399568 );
or ( n52646 , n52644 , n52645 );
nand ( n52647 , n399363 , n399565 );
nand ( n52648 , n52646 , n52647 );
not ( n52649 , n52526 );
and ( n52650 , n52648 , n52649 );
not ( n52651 , n52648 );
and ( n52652 , n52651 , n52526 );
nor ( n52653 , n52650 , n52652 );
xor ( n52654 , n399955 , n52653 );
xor ( n52655 , n399387 , n399390 );
xor ( n52656 , n52655 , n399555 );
buf ( n399970 , n52656 );
buf ( n399971 , n399970 );
xor ( n52659 , n51336 , n398866 );
xnor ( n399973 , n52659 , n398856 );
buf ( n399974 , n399973 );
xor ( n52662 , n398993 , n51616 );
xor ( n52663 , n52662 , n399302 );
buf ( n399977 , n52663 );
xor ( n52665 , n399974 , n399977 );
buf ( n399979 , n392740 );
not ( n52667 , n399979 );
buf ( n399981 , n399008 );
not ( n52669 , n399981 );
or ( n52670 , n52667 , n52669 );
buf ( n399984 , n44776 );
not ( n52672 , n399984 );
buf ( n399986 , n52672 );
buf ( n399987 , n399986 );
not ( n52675 , n399987 );
buf ( n399989 , n389420 );
not ( n52677 , n399989 );
or ( n52678 , n52675 , n52677 );
buf ( n399992 , n396298 );
buf ( n399993 , n44776 );
nand ( n52681 , n399992 , n399993 );
buf ( n399995 , n52681 );
buf ( n399996 , n399995 );
nand ( n52684 , n52678 , n399996 );
buf ( n399998 , n52684 );
buf ( n399999 , n399998 );
buf ( n400000 , n45260 );
nand ( n52688 , n399999 , n400000 );
buf ( n400002 , n52688 );
buf ( n400003 , n400002 );
nand ( n52691 , n52670 , n400003 );
buf ( n400005 , n52691 );
buf ( n400006 , n400005 );
not ( n52694 , n388833 );
not ( n52695 , n399112 );
or ( n52696 , n52694 , n52695 );
buf ( n400010 , n41342 );
not ( n52698 , n400010 );
buf ( n400012 , n388931 );
not ( n52700 , n400012 );
or ( n52701 , n52698 , n52700 );
buf ( n400015 , n389940 );
buf ( n400016 , n45897 );
nand ( n52704 , n400015 , n400016 );
buf ( n400018 , n52704 );
buf ( n400019 , n400018 );
nand ( n52707 , n52701 , n400019 );
buf ( n400021 , n52707 );
buf ( n400022 , n400021 );
buf ( n400023 , n388872 );
nand ( n52711 , n400022 , n400023 );
buf ( n400025 , n52711 );
nand ( n52713 , n52696 , n400025 );
not ( n52714 , n52713 );
xor ( n52715 , n358941 , n358983 );
xor ( n52716 , n52715 , n358996 );
buf ( n400030 , n52716 );
buf ( n400031 , n400030 );
buf ( n52719 , n400031 );
buf ( n400033 , n52719 );
buf ( n400034 , n400033 );
not ( n52722 , n400034 );
buf ( n400036 , n385331 );
not ( n52724 , n400036 );
or ( n52725 , n52722 , n52724 );
buf ( n400039 , n382854 );
buf ( n400040 , n400033 );
not ( n52728 , n400040 );
buf ( n400042 , n52728 );
buf ( n400043 , n400042 );
nand ( n52731 , n400039 , n400043 );
buf ( n400045 , n52731 );
buf ( n400046 , n400045 );
nand ( n52734 , n52725 , n400046 );
buf ( n400048 , n52734 );
buf ( n400049 , n382938 );
buf ( n400050 , n399289 );
nand ( n52741 , n400049 , n400050 );
buf ( n400052 , n52741 );
nand ( n52743 , C1 , n400052 );
not ( n52744 , n52743 );
or ( n52745 , n52714 , n52744 );
or ( n52746 , n52713 , n52743 );
and ( n52747 , n399041 , n399064 );
not ( n52748 , n399041 );
and ( n52749 , n52748 , n399067 );
or ( n52750 , n52747 , n52749 );
not ( n52751 , n399095 );
and ( n52752 , n52750 , n52751 );
not ( n52753 , n52750 );
and ( n52754 , n52753 , n399095 );
nor ( n52755 , n52752 , n52754 );
nand ( n52756 , n52746 , n52755 );
nand ( n52757 , n52745 , n52756 );
buf ( n400068 , n52757 );
buf ( n400069 , n396622 );
not ( n52760 , n400069 );
buf ( n400071 , n24049 );
not ( n52762 , n400071 );
not ( n52763 , n41145 );
buf ( n400074 , n52763 );
not ( n52765 , n400074 );
or ( n52766 , n52762 , n52765 );
buf ( n400077 , n41145 );
buf ( n400078 , n399164 );
nand ( n52769 , n400077 , n400078 );
buf ( n400080 , n52769 );
buf ( n400081 , n400080 );
nand ( n52772 , n52766 , n400081 );
buf ( n400083 , n52772 );
buf ( n400084 , n400083 );
not ( n52775 , n400084 );
or ( n52776 , n52760 , n52775 );
buf ( n400087 , n51775 );
buf ( n400088 , n41563 );
nand ( n52779 , n400087 , n400088 );
buf ( n400090 , n52779 );
buf ( n400091 , n400090 );
nand ( n52782 , n52776 , n400091 );
buf ( n400093 , n52782 );
buf ( n400094 , n400093 );
buf ( n400095 , n12471 );
not ( n52786 , n400095 );
buf ( n400097 , n393525 );
not ( n52788 , n400097 );
or ( n52789 , n52786 , n52788 );
buf ( n400100 , n388962 );
buf ( n400101 , n389593 );
nand ( n52792 , n400100 , n400101 );
buf ( n400103 , n52792 );
buf ( n400104 , n400103 );
nand ( n52795 , n52789 , n400104 );
buf ( n400106 , n52795 );
buf ( n400107 , n400106 );
not ( n52798 , n400107 );
buf ( n400109 , n46056 );
not ( n52800 , n400109 );
or ( n52801 , n52798 , n52800 );
buf ( n400112 , n46061 );
not ( n52803 , n400112 );
buf ( n400114 , n399081 );
nand ( n52805 , n52803 , n400114 );
buf ( n400116 , n52805 );
buf ( n400117 , n400116 );
nand ( n52808 , n52801 , n400117 );
buf ( n400119 , n52808 );
buf ( n400120 , n400119 );
or ( n52811 , n400094 , n400120 );
not ( n52812 , n42950 );
buf ( n400123 , n52812 );
not ( n52814 , n400123 );
buf ( n400125 , n51821 );
not ( n52816 , n400125 );
buf ( n400127 , n46043 );
not ( n52818 , n400127 );
or ( n52819 , n52816 , n52818 );
buf ( n400130 , n28248 );
buf ( n400131 , n51822 );
nand ( n52822 , n400130 , n400131 );
buf ( n400133 , n52822 );
buf ( n400134 , n400133 );
nand ( n52825 , n52819 , n400134 );
buf ( n400136 , n52825 );
buf ( n400137 , n400136 );
not ( n52828 , n400137 );
or ( n52829 , n52814 , n52828 );
buf ( n400140 , n399225 );
buf ( n400141 , n42923 );
not ( n52832 , n400141 );
buf ( n400143 , n52832 );
buf ( n400144 , n400143 );
nand ( n52835 , n400140 , n400144 );
buf ( n400146 , n52835 );
buf ( n400147 , n400146 );
nand ( n52838 , n52829 , n400147 );
buf ( n400149 , n52838 );
buf ( n400150 , n400149 );
nand ( n52841 , n52811 , n400150 );
buf ( n400152 , n52841 );
buf ( n400153 , n400152 );
buf ( n400154 , n400119 );
buf ( n400155 , n400093 );
nand ( n52846 , n400154 , n400155 );
buf ( n400157 , n52846 );
buf ( n400158 , n400157 );
nand ( n52849 , n400153 , n400158 );
buf ( n400160 , n52849 );
buf ( n400161 , n400160 );
buf ( n400162 , n389341 );
not ( n52853 , n400162 );
buf ( n400164 , n388419 );
not ( n52855 , n400164 );
or ( n52856 , n52853 , n52855 );
nand ( n52857 , n40891 , n393185 );
buf ( n400168 , n52857 );
nand ( n52859 , n52856 , n400168 );
buf ( n400170 , n52859 );
buf ( n400171 , n400170 );
not ( n52862 , n400171 );
buf ( n400173 , n36801 );
not ( n52864 , n400173 );
or ( n52865 , n52862 , n52864 );
buf ( n400176 , n398826 );
not ( n52867 , n400176 );
buf ( n400178 , n392111 );
nand ( n52869 , n52867 , n400178 );
buf ( n400180 , n52869 );
buf ( n400181 , n400180 );
nand ( n52872 , n52865 , n400181 );
buf ( n400183 , n52872 );
buf ( n400184 , n400183 );
xor ( n52875 , n400161 , n400184 );
buf ( n400186 , n49117 );
not ( n52877 , n400186 );
buf ( n400188 , n385972 );
not ( n52879 , n400188 );
or ( n52880 , n52877 , n52879 );
buf ( n400191 , n31963 );
buf ( n400192 , n49124 );
nand ( n52883 , n400191 , n400192 );
buf ( n400194 , n52883 );
buf ( n400195 , n400194 );
nand ( n52886 , n52880 , n400195 );
buf ( n400197 , n52886 );
buf ( n400198 , n400197 );
not ( n52889 , n400198 );
buf ( n400200 , n389015 );
not ( n52891 , n400200 );
or ( n52892 , n52889 , n52891 );
buf ( n400203 , n399255 );
buf ( n400204 , n389024 );
nand ( n52895 , n400203 , n400204 );
buf ( n400206 , n52895 );
buf ( n400207 , n400206 );
nand ( n52898 , n52892 , n400207 );
buf ( n400209 , n52898 );
buf ( n400210 , n400209 );
and ( n52901 , n52875 , n400210 );
and ( n52902 , n400161 , n400184 );
or ( n52903 , n52901 , n52902 );
buf ( n400214 , n52903 );
buf ( n400215 , n400214 );
xor ( n52906 , n400068 , n400215 );
buf ( n400217 , n388746 );
not ( n52908 , n400217 );
buf ( n400219 , n388760 );
not ( n52910 , n400219 );
buf ( n400221 , n394120 );
not ( n52912 , n400221 );
or ( n52913 , n52910 , n52912 );
buf ( n400224 , n36709 );
buf ( n400225 , n388757 );
nand ( n52916 , n400224 , n400225 );
buf ( n400227 , n52916 );
buf ( n400228 , n400227 );
nand ( n52919 , n52913 , n400228 );
buf ( n400230 , n52919 );
buf ( n400231 , n400230 );
not ( n52922 , n400231 );
or ( n52923 , n52908 , n52922 );
buf ( n400234 , n399147 );
buf ( n400235 , n388809 );
nand ( n52926 , n400234 , n400235 );
buf ( n400237 , n52926 );
buf ( n400238 , n400237 );
nand ( n52929 , n52923 , n400238 );
buf ( n400240 , n52929 );
buf ( n400241 , n400240 );
and ( n52932 , n52906 , n400241 );
and ( n52933 , n400068 , n400215 );
or ( n52934 , n52932 , n52933 );
buf ( n400245 , n52934 );
buf ( n400246 , n400245 );
xor ( n52937 , n400006 , n400246 );
buf ( n400248 , n45954 );
not ( n52939 , n400248 );
buf ( n400250 , n52195 );
not ( n52941 , n400250 );
or ( n52942 , n52939 , n52941 );
buf ( n400253 , n398116 );
not ( n52944 , n400253 );
buf ( n400255 , n37027 );
not ( n52946 , n400255 );
or ( n52947 , n52944 , n52946 );
buf ( n400258 , n37027 );
not ( n52949 , n400258 );
buf ( n400260 , n393384 );
nand ( n52951 , n52949 , n400260 );
buf ( n400262 , n52951 );
buf ( n400263 , n400262 );
nand ( n52954 , n52947 , n400263 );
buf ( n400265 , n52954 );
buf ( n400266 , n400265 );
buf ( n400267 , n393825 );
nand ( n52958 , n400266 , n400267 );
buf ( n400269 , n52958 );
buf ( n400270 , n400269 );
nand ( n52961 , n52942 , n400270 );
buf ( n400272 , n52961 );
buf ( n400273 , n400272 );
and ( n52964 , n52937 , n400273 );
and ( n52965 , n400006 , n400246 );
or ( n52966 , n52964 , n52965 );
buf ( n400277 , n52966 );
buf ( n400278 , n400277 );
and ( n52969 , n52665 , n400278 );
and ( n52970 , n399974 , n399977 );
or ( n52971 , n52969 , n52970 );
buf ( n400282 , n52971 );
buf ( n400283 , n400282 );
xor ( n52974 , n399971 , n400283 );
xor ( n52975 , n399395 , n399420 );
xor ( n52976 , n52975 , n399425 );
buf ( n400287 , n52976 );
buf ( n400288 , n400287 );
xor ( n52979 , n51705 , n399122 );
xor ( n52980 , n52979 , n399126 );
not ( n52981 , n399464 );
not ( n52982 , n384551 );
and ( n52983 , n52981 , n52982 );
buf ( n400294 , n392611 );
not ( n52985 , n400294 );
buf ( n400296 , n384562 );
not ( n52987 , n400296 );
or ( n52988 , n52985 , n52987 );
buf ( n400299 , n389894 );
buf ( n400300 , n392620 );
nand ( n52991 , n400299 , n400300 );
buf ( n400302 , n52991 );
buf ( n400303 , n400302 );
nand ( n52994 , n52988 , n400303 );
buf ( n400305 , n52994 );
not ( n52996 , n400305 );
buf ( n400307 , n37050 );
buf ( n400308 , n384609 );
buf ( n400309 , n384545 );
nand ( n53000 , n400307 , n400308 , n400309 );
buf ( n400311 , n53000 );
nor ( n53002 , n52996 , n400311 );
nor ( n53003 , n52983 , n53002 );
buf ( n400314 , n53003 );
not ( n53005 , n400314 );
buf ( n400316 , n53005 );
not ( n53007 , n400316 );
buf ( n400318 , n399179 );
buf ( n400319 , n399232 );
xor ( n53010 , n400318 , n400319 );
buf ( n400321 , n399204 );
xnor ( n53012 , n53010 , n400321 );
buf ( n400323 , n53012 );
buf ( n400324 , n400323 );
not ( n53015 , n400324 );
buf ( n400326 , n53015 );
not ( n53017 , n400326 );
or ( n53018 , n53007 , n53017 );
buf ( n400329 , n400323 );
not ( n53020 , n400329 );
buf ( n400331 , n53003 );
not ( n53022 , n400331 );
or ( n53023 , n53020 , n53022 );
not ( n53024 , n399764 );
not ( n53025 , n40640 );
and ( n53026 , n53024 , n53025 );
buf ( n400337 , n394884 );
not ( n53028 , n400337 );
buf ( n400339 , n43044 );
not ( n53030 , n400339 );
or ( n53031 , n53028 , n53030 );
buf ( n400342 , n27196 );
buf ( n400343 , n388154 );
nand ( n53034 , n400342 , n400343 );
buf ( n400345 , n53034 );
buf ( n400346 , n400345 );
nand ( n53037 , n53031 , n400346 );
buf ( n400348 , n53037 );
and ( n53039 , n400348 , n397476 );
nor ( n53040 , n53026 , n53039 );
not ( n53041 , n53040 );
not ( n53042 , n53041 );
buf ( n400353 , n36250 );
buf ( n53044 , n400353 );
buf ( n400355 , n53044 );
and ( n53046 , n400355 , n390460 );
not ( n53047 , n400355 );
and ( n53048 , n53047 , n40990 );
or ( n53049 , n53046 , n53048 );
not ( n53050 , n53049 );
not ( n53051 , n383891 );
or ( n53052 , n53050 , n53051 );
buf ( n400363 , n388626 );
not ( n53054 , n400363 );
buf ( n400365 , n399739 );
nand ( n53056 , n53054 , n400365 );
buf ( n400367 , n53056 );
nand ( n53058 , n53052 , n400367 );
not ( n53059 , n53058 );
or ( n53060 , n53042 , n53059 );
buf ( n400371 , n53040 );
not ( n53062 , n400371 );
buf ( n400373 , n53058 );
not ( n53064 , n400373 );
buf ( n400375 , n53064 );
buf ( n400376 , n400375 );
not ( n53067 , n400376 );
or ( n53068 , n53062 , n53067 );
not ( n53069 , n388872 );
buf ( n400380 , n41342 );
not ( n53071 , n400380 );
buf ( n400382 , n386150 );
not ( n53073 , n400382 );
or ( n53074 , n53071 , n53073 );
buf ( n400385 , n386147 );
buf ( n400386 , n45897 );
nand ( n53077 , n400385 , n400386 );
buf ( n400388 , n53077 );
buf ( n400389 , n400388 );
nand ( n53080 , n53074 , n400389 );
buf ( n400391 , n53080 );
not ( n53082 , n400391 );
or ( n53083 , n53069 , n53082 );
buf ( n400394 , n400021 );
buf ( n400395 , n388833 );
nand ( n53086 , n400394 , n400395 );
buf ( n400397 , n53086 );
nand ( n53088 , n53083 , n400397 );
buf ( n400399 , n53088 );
nand ( n53090 , n53068 , n400399 );
buf ( n400401 , n53090 );
nand ( n53092 , n53060 , n400401 );
buf ( n400403 , n53092 );
nand ( n53094 , n53023 , n400403 );
buf ( n400405 , n53094 );
nand ( n53096 , n53018 , n400405 );
xor ( n53097 , n52980 , n53096 );
not ( n53098 , n45260 );
buf ( n400409 , n399986 );
not ( n53100 , n400409 );
buf ( n400411 , n38356 );
not ( n53102 , n400411 );
or ( n53103 , n53100 , n53102 );
not ( n53104 , n37147 );
not ( n53105 , n392247 );
nand ( n53106 , n53104 , n53105 );
buf ( n400417 , n53106 );
nand ( n53108 , n53103 , n400417 );
buf ( n400419 , n53108 );
not ( n53110 , n400419 );
or ( n53111 , n53098 , n53110 );
buf ( n400422 , n399998 );
buf ( n400423 , n392740 );
nand ( n53114 , n400422 , n400423 );
buf ( n400425 , n53114 );
nand ( n53116 , n53111 , n400425 );
and ( n53117 , n53097 , n53116 );
and ( n53118 , n52980 , n53096 );
or ( n53119 , n53117 , n53118 );
buf ( n400430 , n53119 );
xor ( n53121 , n400288 , n400430 );
xor ( n53122 , n399749 , n399773 );
xor ( n53123 , n53122 , n399796 );
buf ( n400434 , n53123 );
buf ( n400435 , n400434 );
buf ( n400436 , n38765 );
not ( n53127 , n400436 );
buf ( n400438 , n51185 );
not ( n53129 , n400438 );
buf ( n400440 , n53129 );
not ( n53131 , n400440 );
xor ( n53132 , n38685 , n53131 );
buf ( n400443 , n53132 );
not ( n53134 , n400443 );
or ( n53135 , n53127 , n53134 );
nand ( n53136 , n52388 , n390476 );
buf ( n400447 , n53136 );
nand ( n53138 , n53135 , n400447 );
buf ( n400449 , n53138 );
buf ( n400450 , n400449 );
or ( n53141 , n400435 , n400450 );
buf ( n400452 , n53141 );
buf ( n400453 , n389359 );
not ( n53144 , n400453 );
buf ( n400455 , n40973 );
not ( n53146 , n400455 );
or ( n53147 , n53144 , n53146 );
buf ( n400458 , n50992 );
buf ( n400459 , n389356 );
nand ( n53150 , n400458 , n400459 );
buf ( n400461 , n53150 );
buf ( n400462 , n400461 );
nand ( n53153 , n53147 , n400462 );
buf ( n400464 , n53153 );
buf ( n400465 , n400464 );
not ( n53156 , n400465 );
buf ( n400467 , n388460 );
not ( n53158 , n400467 );
or ( n53159 , n53156 , n53158 );
buf ( n400470 , n399786 );
buf ( n400471 , n383940 );
nand ( n53162 , n400470 , n400471 );
buf ( n400473 , n53162 );
buf ( n400474 , n400473 );
nand ( n53165 , n53159 , n400474 );
buf ( n400476 , n53165 );
buf ( n400477 , n400476 );
not ( n53168 , n400477 );
and ( n53169 , n391443 , n40943 );
not ( n53170 , n391443 );
and ( n53171 , n53170 , n390875 );
or ( n53172 , n53169 , n53171 );
not ( n53173 , n53172 );
not ( n53174 , n36801 );
or ( n53175 , n53173 , n53174 );
buf ( n400486 , n392111 );
buf ( n400487 , n400170 );
nand ( n53178 , n400486 , n400487 );
buf ( n400489 , n53178 );
nand ( n53180 , n53175 , n400489 );
buf ( n400491 , n53180 );
not ( n53182 , n400491 );
or ( n53183 , n53168 , n53182 );
buf ( n400494 , n400476 );
buf ( n400495 , n53180 );
or ( n53186 , n400494 , n400495 );
buf ( n400497 , n388543 );
not ( n53188 , n400497 );
buf ( n400499 , n49661 );
not ( n53190 , n400499 );
or ( n53191 , n53188 , n53190 );
buf ( n400502 , n49653 );
buf ( n400503 , n388546 );
nand ( n53194 , n400502 , n400503 );
buf ( n400505 , n53194 );
buf ( n400506 , n400505 );
nand ( n53197 , n53191 , n400506 );
buf ( n400508 , n53197 );
buf ( n400509 , n400508 );
not ( n53200 , n400509 );
buf ( n400511 , n397102 );
not ( n400512 , n400511 );
or ( n53203 , n53200 , n400512 );
buf ( n400514 , n399052 );
buf ( n400515 , n393127 );
nand ( n53206 , n400514 , n400515 );
buf ( n400517 , n53206 );
buf ( n400518 , n400517 );
nand ( n53209 , n53203 , n400518 );
buf ( n400520 , n53209 );
buf ( n400521 , n400520 );
not ( n53212 , n400521 );
buf ( n400523 , n388230 );
not ( n53214 , n400523 );
buf ( n400525 , n388965 );
not ( n53216 , n400525 );
or ( n53217 , n53214 , n53216 );
buf ( n400528 , n388962 );
buf ( n400529 , n388227 );
nand ( n53220 , n400528 , n400529 );
buf ( n400531 , n53220 );
buf ( n400532 , n400531 );
nand ( n53223 , n53217 , n400532 );
buf ( n400534 , n53223 );
buf ( n400535 , n400534 );
not ( n53226 , n400535 );
buf ( n400537 , n393544 );
not ( n53228 , n400537 );
or ( n53229 , n53226 , n53228 );
buf ( n400540 , n400106 );
buf ( n400541 , n49166 );
nand ( n53232 , n400540 , n400541 );
buf ( n400543 , n53232 );
buf ( n400544 , n400543 );
nand ( n53235 , n53229 , n400544 );
buf ( n400546 , n53235 );
buf ( n400547 , n400546 );
not ( n53238 , n400547 );
or ( n53239 , n53212 , n53238 );
buf ( n400550 , n400546 );
buf ( n400551 , n400520 );
or ( n53242 , n400550 , n400551 );
buf ( n400553 , n400143 );
not ( n53244 , n400553 );
buf ( n400555 , n400136 );
not ( n53246 , n400555 );
or ( n53247 , n53244 , n53246 );
not ( n53248 , n51822 );
not ( n53249 , n393557 );
or ( n53250 , n53248 , n53249 );
buf ( n53251 , n41558 );
not ( n53252 , n53251 );
nand ( n53253 , n53252 , n46114 );
nand ( n53254 , n53250 , n53253 );
nand ( n53255 , n53254 , n390432 );
buf ( n400566 , n53255 );
nand ( n53257 , n53247 , n400566 );
buf ( n400568 , n53257 );
buf ( n400569 , n400568 );
nand ( n53260 , n53242 , n400569 );
buf ( n400571 , n53260 );
buf ( n400572 , n400571 );
nand ( n53263 , n53239 , n400572 );
buf ( n400574 , n53263 );
buf ( n400575 , n400574 );
nand ( n53266 , n53186 , n400575 );
buf ( n400577 , n53266 );
buf ( n400578 , n400577 );
nand ( n53269 , n53183 , n400578 );
buf ( n400580 , n53269 );
and ( n53271 , n400452 , n400580 );
buf ( n400582 , n400449 );
buf ( n400583 , n400434 );
and ( n53274 , n400582 , n400583 );
buf ( n400585 , n53274 );
nor ( n53276 , n53271 , n400585 );
buf ( n400587 , n53276 );
not ( n53278 , n400587 );
not ( n53279 , n399479 );
not ( n53280 , n52113 );
or ( n53281 , n53279 , n53280 );
buf ( n400592 , n399482 );
buf ( n400593 , n399504 );
nand ( n53284 , n400592 , n400593 );
buf ( n400595 , n53284 );
nand ( n53286 , n53281 , n400595 );
buf ( n400597 , n399511 );
not ( n53288 , n400597 );
buf ( n400599 , n53288 );
and ( n53290 , n53286 , n400599 );
not ( n53291 , n53286 );
and ( n53292 , n53291 , n399511 );
nor ( n53293 , n53290 , n53292 );
buf ( n400604 , n53293 );
not ( n53295 , n400604 );
buf ( n400606 , n53295 );
buf ( n400607 , n400606 );
nand ( n53298 , n53278 , n400607 );
buf ( n400609 , n53298 );
not ( n53300 , n53293 );
not ( n53301 , n53276 );
or ( n53302 , n53300 , n53301 );
buf ( n400613 , n399067 );
buf ( n400614 , n400083 );
not ( n53305 , n400614 );
buf ( n400616 , n41562 );
nor ( n53307 , n53305 , n400616 );
buf ( n400618 , n53307 );
not ( n53309 , n400618 );
buf ( n400620 , n24049 );
buf ( n400621 , n389856 );
and ( n53312 , n400620 , n400621 );
not ( n53313 , n400620 );
buf ( n400624 , n49686 );
and ( n53315 , n53313 , n400624 );
nor ( n53316 , n53312 , n53315 );
buf ( n400627 , n53316 );
nor ( n53318 , n389119 , n400627 );
nand ( n53319 , n611 , n613 );
nand ( n53320 , n610 , n614 );
and ( n53321 , n53319 , n53320 );
not ( n53322 , n53319 );
not ( n53323 , n53320 );
and ( n53324 , n53322 , n53323 );
nor ( n53325 , n53321 , n53324 );
nand ( n53326 , n608 , n616 );
and ( n53327 , n53325 , n53326 );
nor ( n53328 , n53325 , n53326 );
nor ( n53329 , n53327 , n53328 );
nand ( n53330 , n609 , n615 );
nand ( n53331 , n610 , n615 );
not ( n53332 , n53331 );
nand ( n53333 , n612 , n53332 );
nand ( n53334 , n612 , n613 );
and ( n53335 , n53333 , n53334 );
xor ( n53336 , n53330 , n53335 );
nand ( n53337 , n611 , n614 );
nand ( n53338 , n609 , n616 );
xor ( n53339 , n53337 , n53338 );
nand ( n53340 , n608 , n617 );
and ( n53341 , n53339 , n53340 );
and ( n53342 , n53337 , n53338 );
or ( n53343 , n53341 , n53342 );
xor ( n53344 , n53336 , n53343 );
xor ( n53345 , n53329 , n53344 );
nand ( n53346 , n612 , n614 );
nand ( n53347 , n611 , n615 );
xor ( n53348 , n53346 , n53347 );
nand ( n53349 , n609 , n617 );
and ( n53350 , n53348 , n53349 );
and ( n53351 , n53346 , n53347 );
or ( n53352 , n53350 , n53351 );
and ( n53353 , n53334 , n612 );
nor ( n53354 , C0 , n53353 );
and ( n53355 , n53354 , n53332 );
not ( n53356 , n53354 );
and ( n53357 , n53356 , n53331 );
nor ( n53358 , n53355 , n53357 );
xor ( n53359 , n53352 , n53358 );
xor ( n53360 , n53337 , n53338 );
xor ( n53361 , n53360 , n53340 );
and ( n53362 , n53359 , n53361 );
and ( n53363 , n53352 , n53358 );
or ( n53364 , n53362 , n53363 );
and ( n53365 , n53345 , n53364 );
and ( n53366 , n53329 , n53344 );
or ( n53367 , n53365 , n53366 );
nand ( n53368 , n610 , n613 );
nand ( n53369 , n608 , n615 );
xor ( n53370 , n53368 , n53369 );
not ( n53371 , n53323 );
not ( n53372 , n53319 );
not ( n53373 , n53372 );
or ( n53374 , n53371 , n53373 );
not ( n53375 , n53320 );
not ( n53376 , n53319 );
or ( n53377 , n53375 , n53376 );
not ( n53378 , n53326 );
nand ( n53379 , n53377 , n53378 );
nand ( n53380 , n53374 , n53379 );
not ( n53381 , n53380 );
xor ( n53382 , n53370 , n53381 );
nand ( n53383 , n609 , n614 );
nand ( n53384 , n611 , n612 );
xor ( n53385 , n53383 , n53384 );
not ( n53386 , n611 );
xor ( n53387 , n53385 , n53386 );
xor ( n53388 , n53330 , n53335 );
and ( n53389 , n53388 , n53343 );
and ( n53390 , n53330 , n53335 );
or ( n53391 , n53389 , n53390 );
xor ( n53392 , n53387 , n53391 );
xor ( n53393 , n53382 , n53392 );
nand ( n53394 , n53367 , n53393 );
xor ( n53395 , n53368 , n53369 );
xor ( n53396 , n53395 , n53381 );
and ( n53397 , n53387 , n53396 );
xor ( n53398 , n53368 , n53369 );
xor ( n53399 , n53398 , n53381 );
and ( n53400 , n53391 , n53399 );
and ( n53401 , n53387 , n53391 );
or ( n53402 , n53397 , n53400 , n53401 );
nand ( n53403 , n609 , n613 );
nand ( n53404 , n610 , n612 );
xor ( n53405 , n53403 , n53404 );
nand ( n53406 , n608 , n614 );
xor ( n53407 , n53405 , n53406 );
xor ( n53408 , n53383 , n53384 );
and ( n53409 , n53408 , n53386 );
and ( n53410 , n53383 , n53384 );
or ( n53411 , n53409 , n53410 );
xor ( n53412 , n53368 , n53369 );
and ( n53413 , n53412 , n53381 );
and ( n53414 , n53368 , n53369 );
or ( n53415 , n53413 , n53414 );
xor ( n53416 , n53411 , n53415 );
xor ( n53417 , n53407 , n53416 );
nand ( n53418 , n53402 , n53417 );
and ( n53419 , n53394 , n53418 );
xor ( n53420 , n53403 , n53404 );
and ( n53421 , n53420 , n53406 );
and ( n53422 , n53403 , n53404 );
or ( n53423 , n53421 , n53422 );
nand ( n53424 , n609 , n612 );
xor ( n53425 , n53423 , n53424 );
nand ( n53426 , n608 , n613 );
nand ( n53427 , n610 , n611 );
xor ( n53428 , n53426 , n53427 );
not ( n53429 , n610 );
xor ( n53430 , n53428 , n53429 );
and ( n53431 , n53425 , n53430 );
and ( n53432 , n53423 , n53424 );
or ( n53433 , n53431 , n53432 );
nand ( n53434 , n609 , n611 );
nand ( n53435 , n608 , n612 );
xor ( n53436 , n53434 , n53435 );
xor ( n53437 , n53426 , n53427 );
and ( n53438 , n53437 , n53429 );
and ( n53439 , n53426 , n53427 );
or ( n53440 , n53438 , n53439 );
xor ( n53441 , n53436 , n53440 );
nand ( n53442 , n53433 , n53441 );
not ( n53443 , n53442 );
xor ( n53444 , n53434 , n53435 );
and ( n53445 , n53444 , n53440 );
and ( n53446 , n53434 , n53435 );
or ( n53447 , n53445 , n53446 );
nand ( n53448 , n608 , n611 );
nand ( n53449 , n609 , n610 );
xor ( n53450 , n53448 , n53449 );
not ( n53451 , n609 );
xor ( n53452 , n53450 , n53451 );
nand ( n53453 , n53447 , n53452 );
xor ( n53454 , n53448 , n53449 );
and ( n53455 , n53454 , n53451 );
and ( n53456 , n53448 , n53449 );
or ( n53457 , n53455 , n53456 );
nand ( n53458 , n608 , n610 );
nand ( n53459 , n53457 , n53458 );
nand ( n53460 , n53453 , n53459 );
nor ( n53461 , n53443 , n53460 );
xor ( n53462 , n53403 , n53404 );
xor ( n53463 , n53462 , n53406 );
and ( n53464 , n53411 , n53463 );
xor ( n53465 , n53403 , n53404 );
xor ( n53466 , n53465 , n53406 );
and ( n53467 , n53415 , n53466 );
and ( n53468 , n53411 , n53415 );
or ( n53469 , n53464 , n53467 , n53468 );
xor ( n53470 , n53423 , n53424 );
xor ( n53471 , n53470 , n53430 );
nand ( n53472 , n53469 , n53471 );
and ( n53473 , n53419 , n53461 , n53472 );
not ( n53474 , n53473 );
nand ( n53475 , n610 , n616 );
nand ( n53476 , n608 , n618 );
xor ( n53477 , n53475 , n53476 );
nand ( n53478 , n612 , n615 );
nand ( n53479 , n610 , n617 );
xor ( n53480 , n53478 , n53479 );
nand ( n53481 , n609 , n618 );
and ( n53482 , n53480 , n53481 );
and ( n53483 , n53478 , n53479 );
or ( n53484 , n53482 , n53483 );
xor ( n53485 , n53477 , n53484 );
and ( n53486 , n608 , n619 );
not ( n53487 , n53486 );
nand ( n53488 , n609 , n619 );
not ( n53489 , n53488 );
nand ( n53490 , n611 , n617 );
not ( n53491 , n53490 );
or ( n53492 , n53489 , n53491 );
nand ( n53493 , n608 , n620 );
not ( n53494 , n53493 );
nand ( n53495 , n53492 , n53494 );
not ( n53496 , n53488 );
not ( n53497 , n53490 );
nand ( n53498 , n53496 , n53497 );
nand ( n53499 , n53495 , n53498 );
not ( n53500 , n53499 );
or ( n53501 , n53487 , n53500 );
or ( n53502 , n53499 , n53486 );
nand ( n53503 , n612 , n616 );
nand ( n53504 , n613 , n615 );
xor ( n53505 , n53503 , n53504 );
nand ( n53506 , n610 , n618 );
and ( n53507 , n53505 , n53506 );
and ( n53508 , n53503 , n53504 );
nor ( n53509 , n53507 , n53508 );
nand ( n53510 , n53502 , n53509 );
nand ( n53511 , n53501 , n53510 );
nand ( n53512 , n613 , n614 );
and ( n53513 , n611 , n616 );
nand ( n53514 , n613 , n53513 );
nand ( n53515 , n53512 , n53514 );
not ( n53516 , n53515 );
xor ( n53517 , n53346 , n53347 );
xor ( n53518 , n53517 , n53349 );
not ( n53519 , n53518 );
or ( n53520 , n53516 , n53519 );
or ( n53521 , n53518 , n53515 );
nand ( n53522 , n53520 , n53521 );
xnor ( n53523 , n53511 , n53522 );
and ( n53524 , n53512 , n613 );
nor ( n53525 , C0 , n53524 );
xor ( n53526 , n53525 , n53513 );
xor ( n53527 , n53478 , n53479 );
xor ( n53528 , n53527 , n53481 );
xor ( n53529 , n53526 , n53528 );
xor ( n53530 , n53486 , n53509 );
xnor ( n53531 , n53530 , n53499 );
and ( n53532 , n53529 , n53531 );
and ( n53533 , n53526 , n53528 );
or ( n53534 , n53532 , n53533 );
xor ( n53535 , n53523 , n53534 );
xor ( n53536 , n53485 , n53535 );
nand ( n53537 , n611 , n618 );
nand ( n53538 , n608 , n621 );
xor ( n53539 , n53537 , n53538 );
nand ( n53540 , n613 , n616 );
and ( n53541 , n53539 , n53540 );
and ( n53542 , n53537 , n53538 );
or ( n53543 , n53541 , n53542 );
nand ( n53544 , n614 , n615 );
nand ( n53545 , n612 , n617 );
xor ( n53546 , n53544 , n53545 );
not ( n53547 , n614 );
and ( n53548 , n53546 , n53547 );
and ( n53549 , n53544 , n53545 );
or ( n53550 , n53548 , n53549 );
xor ( n53551 , n53543 , n53550 );
xor ( n53552 , n53503 , n53504 );
xor ( n53553 , n53552 , n53506 );
and ( n53554 , n53551 , n53553 );
and ( n53555 , n53543 , n53550 );
or ( n53556 , n53554 , n53555 );
xor ( n53557 , n53526 , n53528 );
xor ( n53558 , n53557 , n53531 );
xor ( n53559 , n53556 , n53558 );
xor ( n53560 , n53544 , n53545 );
xor ( n53561 , n53560 , n53547 );
not ( n53562 , n53561 );
nand ( n53563 , n612 , n618 );
nand ( n53564 , n610 , n620 );
xor ( n53565 , n53563 , n53564 );
nand ( n53566 , n609 , n621 );
and ( n53567 , n53565 , n53566 );
and ( n53568 , n53563 , n53564 );
or ( n53569 , n53567 , n53568 );
not ( n53570 , n53569 );
or ( n53571 , n53562 , n53570 );
not ( n53572 , n53569 );
not ( n53573 , n53572 );
not ( n53574 , n53561 );
not ( n53575 , n53574 );
or ( n53576 , n53573 , n53575 );
xor ( n53577 , n53537 , n53538 );
xor ( n53578 , n53577 , n53540 );
nand ( n53579 , n53576 , n53578 );
nand ( n53580 , n53571 , n53579 );
not ( n53581 , n53580 );
nand ( n53582 , n610 , n619 );
nand ( n53583 , n609 , n620 );
xor ( n53584 , n53582 , n53583 );
nand ( n53585 , n614 , n616 );
nand ( n53586 , n611 , n619 );
xor ( n53587 , n53585 , n53586 );
nand ( n53588 , n613 , n617 );
and ( n53589 , n53587 , n53588 );
and ( n53590 , n53585 , n53586 );
or ( n53591 , n53589 , n53590 );
and ( n53592 , n53584 , n53591 );
and ( n53593 , n53582 , n53583 );
or ( n53594 , n53592 , n53593 );
not ( n53595 , n53594 );
not ( n53596 , n53488 );
not ( n53597 , n53497 );
or ( n53598 , n53596 , n53597 );
or ( n53599 , n53488 , n53497 );
nand ( n53600 , n53598 , n53599 );
not ( n53601 , n53600 );
not ( n53602 , n53493 );
and ( n53603 , n53601 , n53602 );
and ( n53604 , n53600 , n53493 );
nor ( n53605 , n53603 , n53604 );
not ( n53606 , n53605 );
nand ( n53607 , n53595 , n53606 );
not ( n53608 , n53607 );
or ( n53609 , n53581 , n53608 );
nand ( n53610 , n53594 , n53605 );
nand ( n53611 , n53609 , n53610 );
and ( n53612 , n53559 , n53611 );
and ( n53613 , n53556 , n53558 );
or ( n53614 , n53612 , n53613 );
nand ( n53615 , n53536 , n53614 );
xor ( n53616 , n53475 , n53476 );
xor ( n53617 , n53616 , n53484 );
and ( n53618 , n53523 , n53617 );
xor ( n53619 , n53475 , n53476 );
xor ( n53620 , n53619 , n53484 );
and ( n53621 , n53534 , n53620 );
and ( n53622 , n53523 , n53534 );
or ( n53623 , n53618 , n53621 , n53622 );
xor ( n53624 , n53352 , n53358 );
xor ( n53625 , n53624 , n53361 );
xor ( n53626 , n53475 , n53476 );
and ( n53627 , n53626 , n53484 );
and ( n53628 , n53475 , n53476 );
or ( n53629 , n53627 , n53628 );
not ( n53630 , n53515 );
nand ( n53631 , n53630 , n53518 );
not ( n53632 , n53631 );
not ( n53633 , n53511 );
or ( n53634 , n53632 , n53633 );
not ( n53635 , n53518 );
nand ( n53636 , n53635 , n53515 );
nand ( n53637 , n53634 , n53636 );
not ( n53638 , n53637 );
xor ( n53639 , n53629 , n53638 );
xor ( n53640 , n53625 , n53639 );
nand ( n53641 , n53623 , n53640 );
and ( n53642 , n53615 , n53641 );
xor ( n53643 , n53352 , n53358 );
xor ( n53644 , n53643 , n53361 );
and ( n53645 , n53629 , n53644 );
xor ( n53646 , n53352 , n53358 );
xor ( n53647 , n53646 , n53361 );
and ( n53648 , n53638 , n53647 );
and ( n53649 , n53629 , n53638 );
or ( n53650 , n53645 , n53648 , n53649 );
xor ( n53651 , n53329 , n53344 );
xor ( n53652 , n53651 , n53364 );
nand ( n53653 , n53650 , n53652 );
and ( n53654 , n53642 , n53653 );
not ( n53655 , n53654 );
not ( n53656 , n53580 );
not ( n53657 , n53594 );
not ( n53658 , n53606 );
or ( n53659 , n53657 , n53658 );
nand ( n53660 , n53595 , n53605 );
nand ( n53661 , n53659 , n53660 );
nand ( n53662 , n53656 , n53661 );
nand ( n53663 , n53594 , n53580 , n53605 );
nand ( n53664 , n53595 , n53580 , n53606 );
nand ( n53665 , n53662 , n53663 , n53664 );
xor ( n53666 , n53543 , n53550 );
xor ( n53667 , n53666 , n53553 );
and ( n53668 , n53665 , n53667 );
xor ( n53669 , n53582 , n53583 );
xor ( n53670 , n53669 , n53591 );
nand ( n53671 , n608 , n622 );
nand ( n53672 , n615 , n616 );
xor ( n53673 , n53671 , n53672 );
nand ( n53674 , n609 , n622 );
nand ( n53675 , n608 , n623 );
xor ( n53676 , n53674 , n53675 );
nand ( n53677 , n613 , n618 );
and ( n53678 , n53676 , n53677 );
and ( n53679 , n53674 , n53675 );
or ( n53680 , n53678 , n53679 );
and ( n53681 , n53673 , n53680 );
and ( n53682 , n53671 , n53672 );
or ( n53683 , n53681 , n53682 );
xor ( n53684 , n53670 , n53683 );
nand ( n53685 , n614 , n617 );
nand ( n53686 , n611 , n620 );
xor ( n53687 , n53685 , n53686 );
nand ( n53688 , n612 , n619 );
and ( n53689 , n53687 , n53688 );
and ( n53690 , n53685 , n53686 );
or ( n53691 , n53689 , n53690 );
xor ( n53692 , n53563 , n53564 );
xor ( n53693 , n53692 , n53566 );
xor ( n53694 , n53691 , n53693 );
xor ( n53695 , n53585 , n53586 );
xor ( n53696 , n53695 , n53588 );
and ( n53697 , n53694 , n53696 );
and ( n53698 , n53691 , n53693 );
or ( n53699 , n53697 , n53698 );
and ( n53700 , n53684 , n53699 );
and ( n53701 , n53670 , n53683 );
or ( n53702 , n53700 , n53701 );
xor ( n53703 , n53543 , n53550 );
xor ( n53704 , n53703 , n53553 );
and ( n53705 , n53702 , n53704 );
and ( n53706 , n53665 , n53702 );
or ( n53707 , n53668 , n53705 , n53706 );
xor ( n53708 , n53556 , n53558 );
xor ( n53709 , n53708 , n53611 );
nand ( n53710 , n53707 , n53709 );
xor ( n53711 , n53543 , n53550 );
xor ( n53712 , n53711 , n53553 );
xor ( n53713 , n53665 , n53702 );
xor ( n53714 , n53712 , n53713 );
and ( n53715 , n53574 , n53578 , n53572 );
and ( n53716 , n53561 , n53569 , n53578 );
nor ( n53717 , n53715 , n53716 );
nor ( n53718 , n53578 , n53569 );
and ( n53719 , n53718 , n53561 );
nor ( n53720 , n53561 , n53572 , n53578 );
nor ( n53721 , n53719 , n53720 );
nand ( n53722 , n53717 , n53721 );
nand ( n53723 , n610 , n621 );
nand ( n53724 , n615 , n617 , n614 , n618 );
xor ( n53725 , n53723 , n53724 );
not ( n53726 , n616 );
nand ( n53727 , n53726 , n615 );
and ( n53728 , n53725 , n53727 );
and ( n53729 , n53723 , n53724 );
or ( n53730 , n53728 , n53729 );
xor ( n53731 , n53671 , n53672 );
xor ( n53732 , n53731 , n53680 );
xor ( n53733 , n53730 , n53732 );
nand ( n53734 , n613 , n619 );
nand ( n53735 , n611 , n621 );
xor ( n53736 , n53734 , n53735 );
nand ( n53737 , n612 , n620 );
and ( n401048 , n53736 , n53737 );
and ( n53739 , n53734 , n53735 );
or ( n53740 , n401048 , n53739 );
xor ( n53741 , n53685 , n53686 );
xor ( n53742 , n53741 , n53688 );
xor ( n53743 , n53740 , n53742 );
xor ( n53744 , n53674 , n53675 );
xor ( n53745 , n53744 , n53677 );
and ( n53746 , n53743 , n53745 );
and ( n53747 , n53740 , n53742 );
or ( n53748 , n53746 , n53747 );
and ( n53749 , n53733 , n53748 );
and ( n53750 , n53730 , n53732 );
or ( n53751 , n53749 , n53750 );
xor ( n53752 , n53722 , n53751 );
xor ( n53753 , n53670 , n53683 );
xor ( n53754 , n53753 , n53699 );
and ( n53755 , n53752 , n53754 );
and ( n53756 , n53722 , n53751 );
or ( n53757 , n53755 , n53756 );
nand ( n53758 , n53714 , n53757 );
and ( n53759 , n53710 , n53758 );
not ( n53760 , n53759 );
nand ( n53761 , n610 , n622 );
nand ( n53762 , n609 , n623 );
xor ( n53763 , n53761 , n53762 );
and ( n53764 , n614 , n618 );
not ( n53765 , n53764 );
nand ( n53766 , n615 , n617 );
not ( n53767 , n53766 );
and ( n53768 , n53765 , n53767 );
and ( n53769 , n53766 , n53764 );
nor ( n53770 , n53768 , n53769 );
xor ( n53771 , n53763 , n53770 );
xor ( n53772 , n53734 , n53735 );
xor ( n53773 , n53772 , n53737 );
and ( n53774 , n53771 , n53773 );
nand ( n53775 , n615 , n619 );
not ( n53776 , n53775 );
and ( n53777 , n616 , n618 );
nand ( n53778 , n53776 , n53777 );
nand ( n53779 , n616 , n617 );
and ( n53780 , n53779 , n616 );
nor ( n53781 , C0 , n53780 );
xor ( n53782 , n53778 , n53781 );
nand ( n53783 , n612 , n622 );
not ( n53784 , n53783 );
nand ( n53785 , n614 , n620 );
not ( n53786 , n53785 );
or ( n53787 , n53784 , n53786 );
and ( n53788 , n613 , n621 );
nand ( n53789 , n53787 , n53788 );
not ( n53790 , n53783 );
not ( n53791 , n53785 );
nand ( n53792 , n53790 , n53791 );
and ( n53793 , n53789 , n53792 );
and ( n53794 , n53782 , n53793 );
and ( n53795 , n53778 , n53781 );
or ( n53796 , n53794 , n53795 );
xor ( n53797 , n53734 , n53735 );
xor ( n53798 , n53797 , n53737 );
and ( n53799 , n53796 , n53798 );
and ( n53800 , n53771 , n53796 );
or ( n53801 , n53774 , n53799 , n53800 );
xor ( n53802 , n53740 , n53742 );
xor ( n53803 , n53802 , n53745 );
xor ( n53804 , n53801 , n53803 );
xor ( n53805 , n53761 , n53762 );
and ( n53806 , n53805 , n53770 );
and ( n53807 , n53761 , n53762 );
or ( n53808 , n53806 , n53807 );
xor ( n53809 , n53723 , n53724 );
xor ( n53810 , n53809 , n53727 );
xor ( n53811 , n53808 , n53810 );
nand ( n53812 , n611 , n622 );
not ( n53813 , n53812 );
not ( n53814 , n53813 );
nand ( n53815 , n612 , n621 );
not ( n53816 , n53815 );
not ( n53817 , n53816 );
or ( n53818 , n53814 , n53817 );
not ( n53819 , n53812 );
not ( n53820 , n53815 );
or ( n53821 , n53819 , n53820 );
and ( n53822 , n615 , n618 );
nand ( n53823 , n53821 , n53822 );
nand ( n53824 , n53818 , n53823 );
not ( n53825 , n53824 );
xor ( n53826 , n53779 , n53825 );
nand ( n53827 , n610 , n623 );
not ( n53828 , n53827 );
not ( n53829 , n53828 );
nand ( n53830 , n613 , n620 );
not ( n53831 , n53830 );
not ( n53832 , n53831 );
or ( n53833 , n53829 , n53832 );
not ( n53834 , n53827 );
not ( n53835 , n53830 );
or ( n53836 , n53834 , n53835 );
and ( n53837 , n614 , n619 );
nand ( n53838 , n53836 , n53837 );
nand ( n53839 , n53833 , n53838 );
not ( n53840 , n53839 );
and ( n53841 , n53826 , n53840 );
and ( n53842 , n53779 , n53825 );
or ( n53843 , n53841 , n53842 );
xor ( n53844 , n53811 , n53843 );
xor ( n53845 , n53804 , n53844 );
xor ( n53846 , n53779 , n53825 );
xor ( n53847 , n53846 , n53840 );
not ( n53848 , n53827 );
not ( n53849 , n53837 );
or ( n53850 , n53848 , n53849 );
or ( n53851 , n53827 , n53837 );
nand ( n53852 , n53850 , n53851 );
and ( n53853 , n53852 , n53831 );
not ( n53854 , n53852 );
and ( n53855 , n53854 , n53830 );
nor ( n53856 , n53853 , n53855 );
not ( n53857 , n53856 );
not ( n53858 , n53857 );
not ( n53859 , n53815 );
not ( n53860 , n53822 );
or ( n53861 , n53859 , n53860 );
or ( n53862 , n53815 , n53822 );
nand ( n53863 , n53861 , n53862 );
and ( n53864 , n53863 , n53812 );
not ( n53865 , n53863 );
and ( n53866 , n53865 , n53813 );
nor ( n53867 , n53864 , n53866 );
not ( n53868 , n53867 );
or ( n53869 , n53858 , n53868 );
nand ( n53870 , n611 , n623 );
nand ( n53871 , n617 , n618 );
xor ( n53872 , n53870 , n53871 );
not ( n53873 , n53775 );
not ( n53874 , n53777 );
or ( n53875 , n53873 , n53874 );
or ( n53876 , n53775 , n53777 );
nand ( n53877 , n53875 , n53876 );
not ( n53878 , n53877 );
and ( n53879 , n53872 , n53878 );
and ( n53880 , n53870 , n53871 );
or ( n53881 , n53879 , n53880 );
not ( n53882 , n53881 );
nand ( n53883 , n53869 , n53882 );
not ( n53884 , n53867 );
nand ( n53885 , n53884 , n53856 );
and ( n53886 , n53883 , n53885 );
xor ( n53887 , n53847 , n53886 );
xor ( n53888 , n53734 , n53735 );
xor ( n53889 , n53888 , n53737 );
xor ( n53890 , n53771 , n53796 );
xor ( n53891 , n53889 , n53890 );
and ( n53892 , n53887 , n53891 );
and ( n53893 , n53847 , n53886 );
or ( n53894 , n53892 , n53893 );
nand ( n53895 , n53845 , n53894 );
xor ( n53896 , n53801 , n53803 );
and ( n53897 , n53896 , n53844 );
and ( n53898 , n53801 , n53803 );
or ( n53899 , n53897 , n53898 );
xor ( n53900 , n53691 , n53693 );
xor ( n53901 , n53900 , n53696 );
xor ( n53902 , n53730 , n53732 );
xor ( n53903 , n53902 , n53748 );
xor ( n53904 , n53901 , n53903 );
xor ( n53905 , n53808 , n53810 );
and ( n53906 , n53905 , n53843 );
and ( n53907 , n53808 , n53810 );
or ( n53908 , n53906 , n53907 );
xor ( n53909 , n53904 , n53908 );
nand ( n53910 , n53899 , n53909 );
xor ( n53911 , n53722 , n53751 );
xor ( n53912 , n53911 , n53754 );
xor ( n53913 , n53901 , n53903 );
and ( n53914 , n53913 , n53908 );
and ( n53915 , n53901 , n53903 );
or ( n53916 , n53914 , n53915 );
nand ( n53917 , n53912 , n53916 );
and ( n53918 , n53895 , n53910 , n53917 );
not ( n53919 , n53918 );
xor ( n53920 , n53847 , n53886 );
xor ( n53921 , n53920 , n53891 );
xor ( n53922 , n53778 , n53781 );
xor ( n53923 , n53922 , n53793 );
nand ( n53924 , n616 , n619 );
nand ( n53925 , n614 , n621 );
xor ( n53926 , n53924 , n53925 );
nand ( n53927 , n615 , n620 );
and ( n53928 , n53926 , n53927 );
and ( n53929 , n53924 , n53925 );
or ( n53930 , n53928 , n53929 );
not ( n53931 , n53783 );
not ( n53932 , n53788 );
or ( n53933 , n53931 , n53932 );
or ( n53934 , n53783 , n53788 );
nand ( n53935 , n53933 , n53934 );
and ( n53936 , n53935 , n53785 );
not ( n53937 , n53935 );
and ( n53938 , n53937 , n53791 );
nor ( n53939 , n53936 , n53938 );
xor ( n53940 , n53930 , n53939 );
nand ( n53941 , n613 , n622 );
nand ( n53942 , n612 , n623 );
nand ( n53943 , n53941 , n53942 );
not ( n53944 , n53943 );
nand ( n53945 , n616 , n620 );
nand ( n53946 , n617 , n619 );
nor ( n53947 , n53945 , n53946 );
not ( n53948 , n53947 );
or ( n53949 , n53944 , n53948 );
not ( n53950 , n53942 );
not ( n53951 , n53941 );
nand ( n53952 , n53950 , n53951 );
nand ( n53953 , n53949 , n53952 );
not ( n53954 , n53953 );
and ( n53955 , n53940 , n53954 );
and ( n53956 , n53930 , n53939 );
or ( n53957 , n53955 , n53956 );
xor ( n53958 , n53923 , n53957 );
not ( n53959 , n53867 );
not ( n53960 , n53856 );
or ( n53961 , n53959 , n53960 );
or ( n53962 , n53867 , n53856 );
nand ( n53963 , n53961 , n53962 );
xnor ( n53964 , n53963 , n53882 );
and ( n53965 , n53958 , n53964 );
and ( n53966 , n53923 , n53957 );
or ( n53967 , n53965 , n53966 );
nand ( n53968 , n53921 , n53967 );
not ( n53969 , n53968 );
xor ( n53970 , n53923 , n53957 );
xor ( n53971 , n53970 , n53964 );
xor ( n53972 , n53870 , n53871 );
not ( n53973 , n53877 );
xor ( n53974 , n53972 , n53973 );
and ( n53975 , n53871 , n617 );
nor ( n53976 , C0 , n53975 );
nand ( n53977 , n613 , n623 );
not ( n53978 , n53977 );
nand ( n53979 , n615 , n621 );
not ( n53980 , n53979 );
or ( n53981 , n53978 , n53980 );
and ( n53982 , n614 , n622 );
nand ( n53983 , n53981 , n53982 );
not ( n53984 , n53977 );
not ( n53985 , n53979 );
nand ( n53986 , n53984 , n53985 );
and ( n53987 , n53983 , n53986 );
xor ( n53988 , n53976 , n53987 );
xor ( n53989 , n53924 , n53925 );
xor ( n53990 , n53989 , n53927 );
and ( n53991 , n53988 , n53990 );
and ( n53992 , n53976 , n53987 );
or ( n53993 , n53991 , n53992 );
xor ( n53994 , n53974 , n53993 );
xor ( n53995 , n53930 , n53939 );
xor ( n53996 , n53995 , n53954 );
and ( n53997 , n53994 , n53996 );
and ( n53998 , n53974 , n53993 );
or ( n53999 , n53997 , n53998 );
and ( n54000 , n53971 , n53999 );
nor ( n54001 , n53969 , n54000 );
not ( n54002 , n54001 );
xor ( n54003 , n53974 , n53993 );
xor ( n54004 , n54003 , n53996 );
not ( n54005 , n53951 );
not ( n54006 , n53942 );
and ( n54007 , n54005 , n54006 );
and ( n54008 , n53942 , n53951 );
nor ( n54009 , n54007 , n54008 );
not ( n54010 , n54009 );
not ( n54011 , n53947 );
and ( n54012 , n54010 , n54011 );
and ( n54013 , n53947 , n54009 );
nor ( n54014 , n54012 , n54013 );
nand ( n54015 , n618 , n619 );
xnor ( n54016 , n53946 , n53945 );
xor ( n54017 , n54015 , n54016 );
nand ( n54018 , n616 , n621 );
nand ( n54019 , n615 , n622 );
xor ( n54020 , n54018 , n54019 );
nand ( n54021 , n617 , n620 );
and ( n54022 , n54020 , n54021 );
and ( n54023 , n54018 , n54019 );
or ( n54024 , n54022 , n54023 );
and ( n54025 , n54017 , n54024 );
and ( n54026 , n54015 , n54016 );
or ( n54027 , n54025 , n54026 );
xor ( n54028 , n54014 , n54027 );
xor ( n54029 , n53976 , n53987 );
xor ( n54030 , n54029 , n53990 );
and ( n54031 , n54028 , n54030 );
and ( n54032 , n54014 , n54027 );
or ( n54033 , n54031 , n54032 );
nand ( n54034 , n54004 , n54033 );
not ( n54035 , n54034 );
xor ( n54036 , n54014 , n54027 );
xor ( n54037 , n54036 , n54030 );
not ( n54038 , n53977 );
not ( n54039 , n53982 );
or ( n54040 , n54038 , n54039 );
or ( n54041 , n53977 , n53982 );
nand ( n54042 , n54040 , n54041 );
and ( n54043 , n54042 , n53979 );
not ( n54044 , n54042 );
and ( n54045 , n54044 , n53985 );
nor ( n54046 , n54043 , n54045 );
nand ( n54047 , n614 , n623 );
not ( n54048 , n54047 );
nand ( n54049 , n618 , n620 );
nand ( n54050 , n617 , n621 );
nor ( n54051 , n54049 , n54050 );
not ( n54052 , n54051 );
not ( n54053 , n54052 );
or ( n54054 , n54048 , n54053 );
and ( n54055 , n54015 , n618 );
nor ( n54056 , C0 , n54055 );
not ( n54057 , n54056 );
nand ( n54058 , n54054 , n54057 );
not ( n54059 , n54047 );
nand ( n54060 , n54059 , n54051 );
and ( n54061 , n54058 , n54060 );
xor ( n54062 , n54046 , n54061 );
xor ( n54063 , n54015 , n54016 );
xor ( n54064 , n54063 , n54024 );
and ( n54065 , n54062 , n54064 );
and ( n54066 , n54046 , n54061 );
or ( n54067 , n54065 , n54066 );
and ( n54068 , n54037 , n54067 );
nor ( n54069 , n54035 , n54068 );
not ( n54070 , n54069 );
xor ( n54071 , n54046 , n54061 );
xor ( n54072 , n54071 , n54064 );
nand ( n54073 , n616 , n622 );
nand ( n54074 , n615 , n623 );
xor ( n54075 , n54073 , n54074 );
nand ( n54076 , n619 , n620 );
and ( n54077 , n54075 , n54076 );
and ( n54078 , n54073 , n54074 );
or ( n54079 , n54077 , n54078 );
xor ( n54080 , n54018 , n54019 );
xor ( n54081 , n54080 , n54021 );
xor ( n54082 , n54079 , n54081 );
xor ( n54083 , n54047 , n54051 );
xnor ( n54084 , n54083 , n54056 );
and ( n54085 , n54082 , n54084 );
and ( n54086 , n54079 , n54081 );
or ( n54087 , n54085 , n54086 );
nand ( n54088 , n54072 , n54087 );
xor ( n54089 , n54079 , n54081 );
xor ( n54090 , n54089 , n54084 );
xnor ( n54091 , n54049 , n54050 );
nand ( n54092 , n616 , n623 );
not ( n54093 , n54092 );
nand ( n54094 , n617 , n622 );
not ( n54095 , n54094 );
or ( n54096 , n54093 , n54095 );
nand ( n54097 , n618 , n621 );
not ( n54098 , n54097 );
nand ( n54099 , n54096 , n54098 );
not ( n54100 , n54092 );
not ( n54101 , n54094 );
nand ( n54102 , n54100 , n54101 );
and ( n54103 , n54099 , n54102 );
xor ( n54104 , n54091 , n54103 );
xor ( n54105 , n54073 , n54074 );
xor ( n54106 , n54105 , n54076 );
and ( n54107 , n54104 , n54106 );
and ( n54108 , n54091 , n54103 );
or ( n54109 , n54107 , n54108 );
nand ( n54110 , n54090 , n54109 );
and ( n54111 , n54088 , n54110 );
not ( n54112 , n54111 );
and ( n54113 , n618 , n622 );
and ( n54114 , n619 , n621 );
and ( n54115 , n54113 , n54114 );
not ( n54116 , n619 );
not ( n54117 , n54076 );
or ( n54118 , n54116 , n54117 );
nand ( n54119 , n54118 , C1 );
xor ( n54120 , n54115 , n54119 );
not ( n54121 , n54092 );
not ( n54122 , n54101 );
or ( n54123 , n54121 , n54122 );
or ( n54124 , n54092 , n54101 );
nand ( n54125 , n54123 , n54124 );
and ( n54126 , n54125 , n54098 );
not ( n54127 , n54125 );
and ( n54128 , n54127 , n54097 );
nor ( n54129 , n54126 , n54128 );
and ( n54130 , n54120 , n54129 );
and ( n54131 , n54115 , n54119 );
or ( n54132 , n54130 , n54131 );
not ( n54133 , n54132 );
xor ( n54134 , n54091 , n54103 );
xor ( n54135 , n54134 , n54106 );
nand ( n54136 , n54133 , n54135 );
not ( n54137 , n54136 );
nand ( n54138 , n617 , n623 );
not ( n54139 , n54138 );
not ( n54140 , n54139 );
nand ( n54141 , n620 , n621 );
not ( n54142 , n54141 );
not ( n54143 , n54142 );
or ( n54144 , n54140 , n54143 );
not ( n54145 , n54138 );
not ( n54146 , n54141 );
or ( n54147 , n54145 , n54146 );
xor ( n54148 , n54113 , n54114 );
nand ( n54149 , n54147 , n54148 );
nand ( n54150 , n54144 , n54149 );
xor ( n54151 , n54115 , n54119 );
xor ( n54152 , n54151 , n54129 );
xor ( n54153 , n54150 , n54152 );
and ( n54154 , n54148 , n54138 );
not ( n54155 , n54148 );
and ( n54156 , n54155 , n54139 );
or ( n54157 , n54154 , n54156 );
xnor ( n54158 , n54142 , n54157 );
and ( n54159 , n619 , n622 );
and ( n54160 , n618 , n623 );
xor ( n54161 , n54159 , n54160 );
not ( n54162 , n620 );
not ( n54163 , n54141 );
or ( n54164 , n54162 , n54163 );
nand ( n54165 , n54164 , C1 );
and ( n54166 , n54161 , n54165 );
and ( n54167 , n54159 , n54160 );
or ( n54168 , n54166 , n54167 );
not ( n54169 , n54168 );
nand ( n54170 , n54158 , n54169 );
not ( n54171 , n54170 );
nand ( n54172 , n621 , n623 );
nand ( n54173 , n622 , n623 );
nor ( n54174 , n54172 , n54173 );
not ( n54175 , n54174 );
not ( n54176 , n54175 );
not ( n54177 , n54141 );
nand ( n54178 , n54177 , n623 );
not ( n54179 , n54178 );
and ( n54180 , n620 , n622 );
not ( n54181 , n54180 );
nand ( n54182 , n619 , n623 );
not ( n54183 , n54182 );
and ( n54184 , n54181 , n54183 );
and ( n54185 , n54180 , n54182 );
nor ( n54186 , n54184 , n54185 );
not ( n54187 , n54186 );
nor ( n54188 , n54179 , n54187 );
not ( n54189 , n54188 );
and ( n54190 , n54176 , n54189 );
not ( n54191 , n54186 );
nand ( n54192 , n620 , n623 );
nand ( n54193 , n54192 , n621 );
nand ( n54194 , n621 , n622 );
nor ( n54195 , n54193 , n54194 );
nand ( n54196 , n54191 , n54195 );
nand ( n54197 , n54187 , n54179 );
nand ( n54198 , n54196 , n54197 );
nor ( n54199 , n54190 , n54198 );
xor ( n54200 , n54159 , n54160 );
xor ( n54201 , n54200 , n54165 );
nor ( n54202 , n54076 , n54173 );
nor ( n54203 , n54201 , n54202 );
or ( n54204 , n54199 , n54203 );
nand ( n54205 , n54201 , n54202 );
nand ( n54206 , n54204 , n54205 );
not ( n54207 , n54206 );
or ( n54208 , n54171 , n54207 );
nor ( n54209 , n54158 , n54169 );
not ( n54210 , n54209 );
nand ( n54211 , n54208 , n54210 );
and ( n54212 , n54153 , n54211 );
and ( n54213 , n54150 , n54152 );
or ( n54214 , n54212 , n54213 );
not ( n54215 , n54214 );
or ( n54216 , n54137 , n54215 );
not ( n54217 , n54135 );
nand ( n54218 , n54217 , n54132 );
nand ( n54219 , n54216 , n54218 );
not ( n54220 , n54219 );
or ( n54221 , n54112 , n54220 );
nor ( n54222 , n54090 , n54109 );
nand ( n54223 , n54088 , n54222 );
or ( n54224 , n54072 , n54087 );
and ( n54225 , n54223 , n54224 );
nand ( n54226 , n54221 , n54225 );
not ( n54227 , n54226 );
or ( n54228 , n54070 , n54227 );
nor ( n54229 , n54067 , n54037 );
nand ( n54230 , n54034 , n54229 );
or ( n54231 , n54004 , n54033 );
and ( n54232 , n54230 , n54231 );
nand ( n54233 , n54228 , n54232 );
not ( n54234 , n54233 );
or ( n54235 , n54002 , n54234 );
nor ( n54236 , n53971 , n53999 );
nand ( n54237 , n54236 , n53968 );
or ( n54238 , n53967 , n53921 );
and ( n54239 , n54237 , n54238 );
nand ( n54240 , n54235 , n54239 );
not ( n54241 , n54240 );
or ( n54242 , n53919 , n54241 );
not ( n54243 , n53910 );
nor ( n54244 , n53845 , n53894 );
not ( n54245 , n54244 );
or ( n54246 , n54243 , n54245 );
or ( n54247 , n53899 , n53909 );
nand ( n54248 , n54246 , n54247 );
and ( n54249 , n53917 , n54248 );
nor ( n54250 , n53912 , n53916 );
nor ( n54251 , n54249 , n54250 );
nand ( n54252 , n54242 , n54251 );
not ( n54253 , n54252 );
or ( n54254 , n53760 , n54253 );
nor ( n54255 , n53714 , n53757 );
and ( n54256 , n53710 , n54255 );
nor ( n54257 , n53707 , n53709 );
nor ( n54258 , n54256 , n54257 );
nand ( n54259 , n54254 , n54258 );
not ( n54260 , n54259 );
or ( n54261 , n53655 , n54260 );
nor ( n54262 , n53536 , n53614 );
and ( n54263 , n54262 , n53641 );
nor ( n54264 , n53623 , n53640 );
nor ( n54265 , n54263 , n54264 );
not ( n54266 , n54265 );
and ( n54267 , n54266 , n53653 );
nor ( n401578 , n53650 , n53652 );
nor ( n54269 , n54267 , n401578 );
nand ( n54270 , n54261 , n54269 );
not ( n54271 , n54270 );
or ( n54272 , n53474 , n54271 );
nor ( n54273 , n53367 , n53393 );
and ( n54274 , n54273 , n53418 );
nor ( n54275 , n53402 , n53417 );
nor ( n54276 , n54274 , n54275 );
not ( n54277 , n53472 );
or ( n54278 , n54276 , n54277 );
nor ( n54279 , n53469 , n53471 );
not ( n54280 , n54279 );
nand ( n54281 , n54278 , n54280 );
and ( n54282 , n54281 , n53461 );
nor ( n54283 , n53433 , n53441 );
and ( n54284 , n54283 , n53453 );
nor ( n54285 , n53447 , n53452 );
nor ( n54286 , n54284 , n54285 );
not ( n54287 , n53459 );
or ( n54288 , n54286 , n54287 );
or ( n54289 , n53457 , n53458 );
nand ( n54290 , n54288 , n54289 );
nor ( n54291 , n54282 , n54290 );
nand ( n54292 , n54272 , n54291 );
nand ( n54293 , n53451 , n608 );
nor ( n54294 , n54292 , n54293 );
not ( n54295 , n54294 );
nand ( n54296 , n54292 , n54293 );
nand ( n54297 , n54295 , n54296 );
buf ( n401608 , n54297 );
buf ( n401609 , n14549 );
buf ( n401610 , n14087 );
not ( n54301 , n401610 );
buf ( n401612 , n54301 );
buf ( n401613 , n401612 );
and ( n54304 , n401609 , n401613 );
not ( n54305 , n401609 );
buf ( n401616 , n14087 );
and ( n54307 , n54305 , n401616 );
nor ( n54308 , n54304 , n54307 );
buf ( n401619 , n54308 );
buf ( n401620 , n401619 );
buf ( n401621 , n14549 );
nand ( n54312 , n401620 , n401621 );
buf ( n401623 , n54312 );
buf ( n401624 , n401623 );
not ( n54315 , n401624 );
buf ( n401626 , n54315 );
buf ( n401627 , n401626 );
and ( n54318 , n401608 , n401627 );
not ( n54319 , n608 );
nor ( n54320 , n54319 , n53460 );
not ( n54321 , n54320 );
and ( n54322 , n53419 , n53472 , n53442 );
not ( n54323 , n54322 );
not ( n54324 , n54270 );
or ( n54325 , n54323 , n54324 );
and ( n54326 , n54281 , n53442 );
nor ( n54327 , n54326 , n54283 );
nand ( n54328 , n54325 , n54327 );
not ( n54329 , n54328 );
or ( n54330 , n54321 , n54329 );
and ( n54331 , n54285 , n53459 );
not ( n54332 , n54289 );
nor ( n54333 , n54331 , n54332 , n609 );
not ( n54334 , n54333 );
nand ( n54335 , n54334 , n608 );
nand ( n54336 , n54330 , n54335 );
buf ( n401647 , n54336 );
buf ( n401648 , n401619 );
not ( n54339 , n401648 );
buf ( n401650 , n54339 );
buf ( n401651 , n401650 );
and ( n54342 , n401647 , n401651 );
nor ( n54343 , n54318 , n54342 );
buf ( n401654 , n54343 );
buf ( n401655 , n401654 );
buf ( n54346 , n6088 );
buf ( n401657 , n54346 );
buf ( n401658 , n15290 );
xnor ( n54349 , n401657 , n401658 );
buf ( n401660 , n54349 );
buf ( n401661 , n401660 );
buf ( n401662 , n401612 );
nor ( n54353 , n401661 , n401662 );
buf ( n401664 , n54353 );
buf ( n401665 , n401664 );
not ( n54356 , n401665 );
buf ( n401667 , n401660 );
buf ( n401668 , n54346 );
buf ( n401669 , n14087 );
xor ( n54360 , n401668 , n401669 );
buf ( n401671 , n54360 );
buf ( n401672 , n401671 );
and ( n54363 , n401667 , n401672 );
buf ( n401674 , n54363 );
buf ( n401675 , n401674 );
buf ( n401676 , n14087 );
buf ( n54367 , n401676 );
buf ( n401678 , n54367 );
buf ( n401679 , n401678 );
nand ( n54370 , n401675 , n401679 );
buf ( n401681 , n54370 );
buf ( n401682 , n401681 );
nand ( n54373 , n54356 , n401682 );
buf ( n401684 , n54373 );
buf ( n401685 , n401684 );
xor ( n54376 , n401655 , n401685 );
buf ( n401687 , n401612 );
buf ( n54378 , n401687 );
buf ( n401689 , n54378 );
buf ( n401690 , n401689 );
not ( n54381 , n401690 );
buf ( n401692 , n54381 );
buf ( n401693 , n401692 );
buf ( n54384 , n401693 );
buf ( n401695 , n54384 );
buf ( n401696 , n401695 );
buf ( n401697 , n54336 );
not ( n54388 , n401697 );
buf ( n401699 , n54388 );
buf ( n401700 , n401699 );
and ( n54391 , n401696 , n401700 );
not ( n54392 , n401696 );
buf ( n401703 , n54336 );
and ( n54394 , n54392 , n401703 );
nor ( n54395 , n54391 , n54394 );
buf ( n401706 , n54395 );
buf ( n401707 , n401706 );
not ( n54398 , n401707 );
buf ( n401709 , n54398 );
buf ( n401710 , n401709 );
buf ( n401711 , n401674 );
and ( n54402 , n401710 , n401711 );
buf ( n401713 , n401664 );
nor ( n54404 , n54402 , n401713 );
buf ( n401715 , n54404 );
buf ( n401716 , n401715 );
not ( n54407 , n53453 );
nor ( n54408 , n53443 , n54277 , n54407 );
and ( n54409 , n53653 , n53419 , n54408 );
not ( n54410 , n54409 );
not ( n54411 , n53642 );
not ( n54412 , n54259 );
or ( n54413 , n54411 , n54412 );
nand ( n54414 , n54413 , n54265 );
not ( n54415 , n54414 );
or ( n54416 , n54410 , n54415 );
not ( n54417 , n53419 );
not ( n54418 , n401578 );
or ( n54419 , n54417 , n54418 );
nand ( n54420 , n54419 , n54276 );
and ( n54421 , n54420 , n54408 );
and ( n54422 , n54279 , n53442 );
nor ( n54423 , n54422 , n54283 );
or ( n54424 , n54423 , n54407 );
not ( n54425 , n54285 );
nand ( n54426 , n54424 , n54425 );
nor ( n54427 , n54421 , n54426 );
nand ( n54428 , n54416 , n54427 );
nand ( n54429 , n53459 , n54289 );
nor ( n54430 , n54428 , n54429 );
not ( n54431 , n54430 );
nand ( n54432 , n54428 , n54429 );
nand ( n54433 , n54431 , n54432 );
buf ( n401744 , n54433 );
buf ( n401745 , n401626 );
and ( n54436 , n401744 , n401745 );
buf ( n401747 , n54297 );
buf ( n401748 , n401650 );
and ( n54439 , n401747 , n401748 );
nor ( n54440 , n54436 , n54439 );
buf ( n401751 , n54440 );
buf ( n401752 , n401751 );
nand ( n54443 , n401716 , n401752 );
buf ( n401754 , n54443 );
buf ( n401755 , n401754 );
not ( n54446 , n401755 );
buf ( n401757 , n54446 );
buf ( n401758 , n401757 );
and ( n54449 , n54376 , n401758 );
and ( n54450 , n401655 , n401685 );
or ( n54451 , n54449 , n54450 );
buf ( n401762 , n54451 );
buf ( n401763 , n401762 );
buf ( n401764 , n54336 );
buf ( n401765 , n401626 );
nand ( n54456 , n401764 , n401765 );
buf ( n401767 , n54456 );
buf ( n401768 , n401767 );
nand ( n54459 , n401763 , n401768 );
buf ( n401770 , n54459 );
nor ( n54461 , n53318 , n401770 );
nand ( n54462 , n53309 , n54461 );
buf ( n401773 , n54462 );
xor ( n54464 , n400613 , n401773 );
buf ( n401775 , n43058 );
buf ( n401776 , n388998 );
buf ( n401777 , n37346 );
and ( n54468 , n401776 , n401777 );
not ( n54469 , n401776 );
buf ( n401780 , n393117 );
and ( n54471 , n54469 , n401780 );
nor ( n54472 , n54468 , n54471 );
buf ( n401783 , n54472 );
buf ( n401784 , n401783 );
or ( n54475 , n401775 , n401784 );
buf ( n401786 , n399192 );
not ( n54477 , n401786 );
buf ( n401788 , n54477 );
buf ( n401789 , n401788 );
buf ( n401790 , n398665 );
or ( n54481 , n401789 , n401790 );
nand ( n54482 , n54475 , n54481 );
buf ( n401793 , n54482 );
buf ( n401794 , n401793 );
and ( n54485 , n54464 , n401794 );
and ( n54486 , n400613 , n401773 );
or ( n54487 , n54485 , n54486 );
buf ( n401798 , n54487 );
buf ( n401799 , n401798 );
buf ( n401800 , n389162 );
not ( n54491 , n401800 );
buf ( n401802 , n399497 );
not ( n54493 , n401802 );
or ( n54494 , n54491 , n54493 );
buf ( n401805 , n41671 );
not ( n54496 , n401805 );
buf ( n401807 , n394426 );
not ( n54498 , n401807 );
or ( n54499 , n54496 , n54498 );
buf ( n401810 , n37763 );
buf ( n401811 , n41670 );
nand ( n54502 , n401810 , n401811 );
buf ( n401813 , n54502 );
buf ( n401814 , n401813 );
nand ( n54505 , n54499 , n401814 );
buf ( n401816 , n54505 );
buf ( n401817 , n401816 );
buf ( n401818 , n41711 );
nand ( n54509 , n401817 , n401818 );
buf ( n401820 , n54509 );
buf ( n401821 , n401820 );
nand ( n54512 , n54494 , n401821 );
buf ( n401823 , n54512 );
buf ( n401824 , n401823 );
xor ( n54515 , n401799 , n401824 );
buf ( n401826 , n394210 );
buf ( n401827 , n388556 );
and ( n54518 , n401826 , n401827 );
not ( n54519 , n401826 );
buf ( n401830 , n395919 );
and ( n54521 , n54519 , n401830 );
nor ( n54522 , n54518 , n54521 );
buf ( n401833 , n54522 );
buf ( n401834 , n401833 );
not ( n54525 , n401834 );
buf ( n401836 , n391270 );
not ( n54527 , n401836 );
or ( n54528 , n54525 , n54527 );
buf ( n401839 , n399709 );
not ( n54530 , n401839 );
buf ( n401841 , n383406 );
nand ( n54532 , n54530 , n401841 );
buf ( n401843 , n54532 );
buf ( n401844 , n401843 );
nand ( n54535 , n54528 , n401844 );
buf ( n401846 , n54535 );
buf ( n401847 , n401846 );
and ( n54538 , n54515 , n401847 );
and ( n54539 , n401799 , n401824 );
or ( n54540 , n54538 , n54539 );
buf ( n401851 , n54540 );
nand ( n54542 , n53302 , n401851 );
nand ( n54543 , n400609 , n54542 );
buf ( n401854 , n54543 );
and ( n54545 , n53121 , n401854 );
and ( n54546 , n400288 , n400430 );
or ( n54547 , n54545 , n54546 );
buf ( n401858 , n54547 );
buf ( n401859 , n401858 );
buf ( n401860 , n395349 );
not ( n54551 , n401860 );
buf ( n401862 , n47863 );
not ( n54553 , n401862 );
buf ( n401864 , n382924 );
not ( n54555 , n401864 );
or ( n54556 , n54553 , n54555 );
buf ( n401867 , n386561 );
not ( n54558 , n401867 );
buf ( n401869 , n395312 );
nand ( n54560 , n54558 , n401869 );
buf ( n401871 , n54560 );
buf ( n401872 , n401871 );
nand ( n54563 , n54556 , n401872 );
buf ( n401874 , n54563 );
buf ( n401875 , n401874 );
not ( n54566 , n401875 );
or ( n54567 , n54551 , n54566 );
buf ( n401878 , n399444 );
buf ( n401879 , n395362 );
nand ( n54570 , n401878 , n401879 );
buf ( n401881 , n54570 );
buf ( n401882 , n401881 );
nand ( n54573 , n54567 , n401882 );
buf ( n401884 , n54573 );
buf ( n401885 , n401884 );
xor ( n54576 , n399130 , n399155 );
xor ( n54577 , n54576 , n399298 );
buf ( n401888 , n54577 );
buf ( n401889 , n401888 );
xor ( n54580 , n401885 , n401889 );
not ( n54581 , n398837 );
buf ( n401892 , n51391 );
buf ( n401893 , n51404 );
and ( n54584 , n401892 , n401893 );
not ( n54585 , n401892 );
buf ( n401896 , n398812 );
and ( n54587 , n54585 , n401896 );
nor ( n54588 , n54584 , n54587 );
buf ( n401899 , n54588 );
not ( n54590 , n401899 );
not ( n54591 , n54590 );
or ( n54592 , n54581 , n54591 );
nand ( n54593 , n401899 , n51441 );
nand ( n54594 , n54592 , n54593 );
buf ( n401905 , n54594 );
not ( n54596 , n401905 );
buf ( n401907 , n54596 );
buf ( n401908 , n401907 );
not ( n54599 , n401908 );
not ( n54600 , n43286 );
not ( n54601 , n384180 );
not ( n54602 , n388105 );
or ( n54603 , n54601 , n54602 );
nand ( n54604 , n388102 , n384202 );
nand ( n54605 , n54603 , n54604 );
not ( n54606 , n54605 );
or ( n54607 , n54600 , n54606 );
buf ( n401918 , n399679 );
buf ( n401919 , n390362 );
nand ( n54610 , n401918 , n401919 );
buf ( n401921 , n54610 );
nand ( n54612 , n54607 , n401921 );
buf ( n401923 , n54612 );
not ( n54614 , n401923 );
or ( n54615 , n54599 , n54614 );
xor ( n54616 , n399243 , n399267 );
xor ( n54617 , n54616 , n399294 );
buf ( n401928 , n54617 );
buf ( n401929 , n54612 );
not ( n54620 , n401929 );
buf ( n401931 , n54594 );
nand ( n54622 , n54620 , n401931 );
buf ( n401933 , n54622 );
buf ( n401934 , n401933 );
nand ( n54625 , n401928 , n401934 );
buf ( n401936 , n54625 );
buf ( n401937 , n401936 );
nand ( n54628 , n54615 , n401937 );
buf ( n401939 , n54628 );
buf ( n401940 , n401939 );
and ( n54631 , n54580 , n401940 );
and ( n54632 , n401885 , n401889 );
or ( n54633 , n54631 , n54632 );
buf ( n401944 , n54633 );
buf ( n401945 , n401944 );
xor ( n54636 , n401859 , n401945 );
not ( n54637 , n52220 );
not ( n54638 , n52202 );
and ( n54639 , n54637 , n54638 );
and ( n54640 , n52220 , n52202 );
nor ( n54641 , n54639 , n54640 );
and ( n54642 , n54641 , n52187 );
not ( n54643 , n54641 );
not ( n54644 , n52187 );
and ( n54645 , n54643 , n54644 );
nor ( n54646 , n54642 , n54645 );
buf ( n401957 , n54646 );
and ( n54648 , n54636 , n401957 );
and ( n54649 , n401859 , n401945 );
or ( n54650 , n54648 , n54649 );
buf ( n401961 , n54650 );
buf ( n401962 , n401961 );
and ( n54653 , n52974 , n401962 );
and ( n54654 , n399971 , n400283 );
or ( n54655 , n54653 , n54654 );
buf ( n401966 , n54655 );
buf ( n401967 , n401966 );
not ( n54658 , n401967 );
buf ( n401969 , n54658 );
buf ( n401970 , n401969 );
buf ( n401971 , n399559 );
buf ( n401972 , n51975 );
and ( n54663 , n401971 , n401972 );
not ( n54664 , n401971 );
buf ( n401975 , n399370 );
and ( n54666 , n54664 , n401975 );
nor ( n54667 , n54663 , n54666 );
buf ( n401978 , n54667 );
buf ( n54669 , n51983 );
and ( n54670 , n401978 , n54669 );
not ( n54671 , n401978 );
not ( n54672 , n54669 );
and ( n54673 , n54671 , n54672 );
nor ( n54674 , n54670 , n54673 );
buf ( n401985 , n54674 );
xor ( n54676 , n401970 , n401985 );
xor ( n54677 , n399624 , n52519 );
xor ( n54678 , n54677 , n399837 );
buf ( n401989 , n54678 );
and ( n54680 , n54676 , n401989 );
and ( n54681 , n401970 , n401985 );
or ( n54682 , n54680 , n54681 );
buf ( n401993 , n54682 );
xor ( n54684 , n52654 , n401993 );
xor ( n54685 , n399577 , n399616 );
xor ( n54686 , n54685 , n399620 );
buf ( n401997 , n54686 );
buf ( n401998 , n401997 );
xor ( n54689 , n399628 , n399813 );
xor ( n54690 , n54689 , n399824 );
buf ( n402001 , n54690 );
buf ( n402002 , n402001 );
xor ( n54693 , n401998 , n402002 );
buf ( n402004 , n52347 );
buf ( n402005 , n399810 );
xor ( n54696 , n402004 , n402005 );
buf ( n402007 , n399631 );
xnor ( n54698 , n54696 , n402007 );
buf ( n402009 , n54698 );
xor ( n54700 , n399430 , n399455 );
xor ( n54701 , n54700 , n399550 );
buf ( n402012 , n54701 );
or ( n54703 , n402009 , n402012 );
xor ( n54704 , n399523 , n399526 );
xor ( n54705 , n54704 , n399545 );
buf ( n402016 , n54705 );
buf ( n402017 , n402016 );
buf ( n402018 , n43727 );
not ( n54709 , n402018 );
buf ( n402020 , n391027 );
not ( n54711 , n402020 );
buf ( n402022 , n383762 );
not ( n54713 , n402022 );
or ( n54714 , n54711 , n54713 );
buf ( n402025 , n49525 );
buf ( n402026 , n391024 );
nand ( n54717 , n402025 , n402026 );
buf ( n402028 , n54717 );
buf ( n402029 , n402028 );
nand ( n54720 , n54714 , n402029 );
buf ( n402031 , n54720 );
buf ( n402032 , n402031 );
not ( n54723 , n402032 );
or ( n54724 , n54709 , n54723 );
buf ( n402035 , n399542 );
buf ( n402036 , n43515 );
nand ( n54727 , n402035 , n402036 );
buf ( n402038 , n54727 );
buf ( n402039 , n402038 );
nand ( n54730 , n54724 , n402039 );
buf ( n402041 , n54730 );
buf ( n402042 , n402041 );
buf ( n402043 , C0 );
buf ( n402044 , n402043 );
xor ( n54764 , n402042 , n402044 );
buf ( n402046 , n45954 );
not ( n54766 , n402046 );
buf ( n402048 , n400265 );
not ( n54768 , n402048 );
or ( n54769 , n54766 , n54768 );
buf ( n402051 , n398116 );
not ( n54771 , n402051 );
buf ( n402053 , n49933 );
not ( n54773 , n402053 );
or ( n54774 , n54771 , n54773 );
buf ( n402056 , n49938 );
buf ( n402057 , n393384 );
nand ( n54777 , n402056 , n402057 );
buf ( n402059 , n54777 );
buf ( n402060 , n402059 );
nand ( n54780 , n54774 , n402060 );
buf ( n402062 , n54780 );
buf ( n402063 , n402062 );
buf ( n402064 , n393825 );
nand ( n54784 , n402063 , n402064 );
buf ( n402066 , n54784 );
buf ( n402067 , n402066 );
nand ( n54787 , n54769 , n402067 );
buf ( n402069 , n54787 );
buf ( n402070 , n402069 );
and ( n54790 , n54764 , n402070 );
or ( n402072 , n54790 , C0 );
buf ( n402073 , n402072 );
buf ( n402074 , n402073 );
xor ( n54795 , n402017 , n402074 );
xor ( n54796 , n399654 , n52258 );
xnor ( n54797 , n54796 , n52345 );
buf ( n402078 , n54797 );
and ( n54799 , n54795 , n402078 );
and ( n54800 , n402017 , n402074 );
or ( n54801 , n54799 , n54800 );
buf ( n402082 , n54801 );
nand ( n54803 , n54703 , n402082 );
buf ( n402084 , n402009 );
buf ( n402085 , n402012 );
nand ( n54806 , n402084 , n402085 );
buf ( n402087 , n54806 );
and ( n54808 , n54803 , n402087 );
buf ( n402089 , n54808 );
and ( n54810 , n54693 , n402089 );
and ( n54811 , n401998 , n402002 );
or ( n54812 , n54810 , n54811 );
buf ( n402093 , n54812 );
buf ( n402094 , n402093 );
xor ( n54815 , n399971 , n400283 );
xor ( n54816 , n54815 , n401962 );
buf ( n402097 , n54816 );
buf ( n402098 , n402097 );
not ( n54819 , n402098 );
xor ( n54820 , n399685 , n399693 );
xor ( n54821 , n54820 , n399806 );
buf ( n402102 , n54821 );
buf ( n402103 , n402102 );
not ( n54824 , n52253 );
not ( n54825 , n54824 );
not ( n54826 , n50564 );
and ( n54827 , n54825 , n54826 );
and ( n54828 , n50584 , n388774 );
not ( n54829 , n50584 );
and ( n54830 , n54829 , n386421 );
or ( n54831 , n54828 , n54830 );
and ( n54832 , n54831 , n50579 );
nor ( n54833 , n54827 , n54832 );
not ( n54834 , n54833 );
not ( n54835 , n54834 );
xor ( n54836 , n399704 , n399726 );
xor ( n54837 , n54836 , n399801 );
buf ( n402118 , n54837 );
not ( n54839 , n402118 );
or ( n54840 , n54835 , n54839 );
not ( n54841 , n402118 );
buf ( n402122 , n54841 );
not ( n54843 , n402122 );
buf ( n402124 , n54833 );
not ( n54845 , n402124 );
or ( n54846 , n54843 , n54845 );
not ( n54847 , n390362 );
not ( n54848 , n54605 );
or ( n54849 , n54847 , n54848 );
buf ( n402130 , n388102 );
not ( n54851 , n402130 );
buf ( n402132 , n384239 );
not ( n54853 , n402132 );
or ( n54854 , n54851 , n54853 );
buf ( n402135 , n41595 );
buf ( n402136 , n388105 );
nand ( n54857 , n402135 , n402136 );
buf ( n402138 , n54857 );
buf ( n402139 , n402138 );
nand ( n54860 , n54854 , n402139 );
buf ( n402141 , n54860 );
buf ( n402142 , n402141 );
buf ( n402143 , n43286 );
nand ( n54864 , n402142 , n402143 );
buf ( n402145 , n54864 );
nand ( n54866 , n54849 , n402145 );
buf ( n402147 , n54866 );
buf ( n402148 , n388809 );
not ( n54869 , n402148 );
buf ( n402150 , n400230 );
not ( n54871 , n402150 );
or ( n54872 , n54869 , n54871 );
xor ( n54873 , n36509 , n388757 );
buf ( n402154 , n54873 );
not ( n54875 , n402154 );
buf ( n402156 , n388746 );
nand ( n54877 , n54875 , n402156 );
buf ( n402158 , n54877 );
buf ( n402159 , n402158 );
nand ( n54880 , n54872 , n402159 );
buf ( n402161 , n54880 );
buf ( n402162 , n402161 );
xor ( n54883 , n402147 , n402162 );
buf ( n402164 , n400093 );
buf ( n402165 , n400149 );
xor ( n54886 , n402164 , n402165 );
buf ( n402167 , n400119 );
xnor ( n54888 , n54886 , n402167 );
buf ( n402169 , n54888 );
not ( n54890 , n402169 );
not ( n54891 , n54890 );
not ( n54892 , n389162 );
not ( n54893 , n401816 );
or ( n54894 , n54892 , n54893 );
buf ( n402175 , n41671 );
not ( n54896 , n402175 );
buf ( n402177 , n388979 );
not ( n54898 , n402177 );
or ( n54899 , n54896 , n54898 );
buf ( n402180 , n29077 );
buf ( n402181 , n41670 );
nand ( n54902 , n402180 , n402181 );
buf ( n402183 , n54902 );
buf ( n402184 , n402183 );
nand ( n54905 , n54899 , n402184 );
buf ( n402186 , n54905 );
buf ( n402187 , n402186 );
buf ( n402188 , n41711 );
nand ( n54909 , n402187 , n402188 );
buf ( n402190 , n54909 );
nand ( n54911 , n54894 , n402190 );
not ( n54912 , n54911 );
or ( n54913 , n54891 , n54912 );
not ( n54914 , n402169 );
not ( n54915 , n54911 );
not ( n54916 , n54915 );
or ( n54917 , n54914 , n54916 );
or ( n54918 , n53318 , n400618 );
nand ( n54919 , n54918 , n401770 );
nand ( n54920 , n54919 , n54462 );
buf ( n402201 , n54920 );
not ( n54922 , n388502 );
and ( n54923 , n54922 , n393562 );
not ( n54924 , n54922 );
and ( n54925 , n54924 , n388897 );
or ( n54926 , n54923 , n54925 );
not ( n54927 , n54926 );
not ( n54928 , n45662 );
or ( n54929 , n54927 , n54928 );
not ( n54930 , n401783 );
nand ( n54931 , n54930 , n398668 );
nand ( n54932 , n54929 , n54931 );
buf ( n402213 , n54932 );
xor ( n54934 , n402201 , n402213 );
buf ( n402215 , n401762 );
buf ( n402216 , n401767 );
or ( n54937 , n402215 , n402216 );
buf ( n402218 , n401770 );
nand ( n54939 , n54937 , n402218 );
buf ( n402220 , n54939 );
not ( n54941 , n400143 );
not ( n54942 , n53254 );
or ( n54943 , n54941 , n54942 );
not ( n54944 , n47412 );
not ( n54945 , n52763 );
or ( n54946 , n54944 , n54945 );
buf ( n402227 , n388643 );
buf ( n402228 , n53251 );
nand ( n54949 , n402227 , n402228 );
buf ( n402230 , n54949 );
nand ( n54951 , n54946 , n402230 );
nand ( n54952 , n54951 , n52812 );
nand ( n54953 , n54943 , n54952 );
xor ( n54954 , n402220 , n54953 );
buf ( n402235 , n12471 );
not ( n54956 , n402235 );
not ( n54957 , n49653 );
buf ( n402238 , n54957 );
not ( n54959 , n402238 );
or ( n54960 , n54956 , n54959 );
buf ( n402241 , n49653 );
buf ( n402242 , n389593 );
nand ( n54963 , n402241 , n402242 );
buf ( n402244 , n54963 );
buf ( n402245 , n402244 );
nand ( n54966 , n54960 , n402245 );
buf ( n402247 , n54966 );
buf ( n402248 , n402247 );
not ( n54969 , n402248 );
buf ( n402250 , n38961 );
not ( n54971 , n402250 );
or ( n54972 , n54969 , n54971 );
buf ( n402253 , n400508 );
buf ( n402254 , n395199 );
nand ( n54975 , n402253 , n402254 );
buf ( n402256 , n54975 );
buf ( n402257 , n402256 );
nand ( n54978 , n54972 , n402257 );
buf ( n402259 , n54978 );
and ( n54980 , n54954 , n402259 );
and ( n54981 , n402220 , n54953 );
or ( n54982 , n54980 , n54981 );
buf ( n402263 , n54982 );
and ( n54984 , n54934 , n402263 );
and ( n54985 , n402201 , n402213 );
or ( n54986 , n54984 , n54985 );
buf ( n402267 , n54986 );
nand ( n54988 , n54917 , n402267 );
nand ( n54989 , n54913 , n54988 );
buf ( n402270 , n54989 );
and ( n54991 , n54883 , n402270 );
and ( n54992 , n402147 , n402162 );
or ( n54993 , n54991 , n54992 );
buf ( n402274 , n54993 );
buf ( n402275 , n402274 );
nand ( n54996 , n54846 , n402275 );
buf ( n402277 , n54996 );
nand ( n54998 , n54840 , n402277 );
buf ( n402279 , n54998 );
xor ( n55000 , n402103 , n402279 );
xor ( n55001 , n400006 , n400246 );
xor ( n55002 , n55001 , n400273 );
buf ( n402283 , n55002 );
buf ( n402284 , n402283 );
and ( n55005 , n55000 , n402284 );
and ( n55006 , n402103 , n402279 );
or ( n55007 , n55005 , n55006 );
buf ( n402288 , n55007 );
buf ( n402289 , n402288 );
xor ( n55010 , n400068 , n400215 );
xor ( n55011 , n55010 , n400241 );
buf ( n402292 , n55011 );
buf ( n402293 , n402292 );
not ( n55014 , n402293 );
buf ( n402295 , n395362 );
not ( n55016 , n402295 );
buf ( n402297 , n401874 );
not ( n55018 , n402297 );
or ( n55019 , n55016 , n55018 );
buf ( n402300 , n47863 );
not ( n55021 , n402300 );
buf ( n402302 , n386385 );
not ( n55023 , n402302 );
or ( n55024 , n55021 , n55023 );
buf ( n402305 , n386385 );
not ( n55026 , n402305 );
buf ( n402307 , n55026 );
buf ( n402308 , n402307 );
buf ( n402309 , n395312 );
nand ( n55030 , n402308 , n402309 );
buf ( n402311 , n55030 );
buf ( n402312 , n402311 );
nand ( n55033 , n55024 , n402312 );
buf ( n402314 , n55033 );
buf ( n402315 , n402314 );
buf ( n402316 , n395349 );
nand ( n55037 , n402315 , n402316 );
buf ( n402318 , n55037 );
buf ( n402319 , n402318 );
nand ( n55040 , n55019 , n402319 );
buf ( n402321 , n55040 );
buf ( n402322 , n402321 );
not ( n55043 , n402322 );
or ( n55044 , n55014 , n55043 );
buf ( n402325 , n402292 );
buf ( n402326 , n402321 );
or ( n55047 , n402325 , n402326 );
not ( n55048 , n358982 );
buf ( n402329 , n358979 );
buf ( n402330 , n358964 );
nand ( n55051 , n402329 , n402330 );
buf ( n402332 , n55051 );
nand ( n55053 , n55048 , n402332 );
buf ( n55054 , n55053 );
not ( n55055 , n55054 );
buf ( n402336 , n55055 );
not ( n55057 , n402336 );
buf ( n402338 , n384096 );
not ( n55059 , n402338 );
or ( n55060 , n55057 , n55059 );
buf ( n402341 , n382854 );
buf ( n402342 , n55054 );
nand ( n55063 , n402341 , n402342 );
buf ( n402344 , n55063 );
buf ( n402345 , n402344 );
nand ( n55066 , n55060 , n402345 );
buf ( n402347 , n55066 );
buf ( n402348 , n389547 );
buf ( n402349 , n400048 );
nand ( n55075 , n402348 , n402349 );
buf ( n402351 , n55075 );
buf ( n402352 , n402351 );
nand ( n55078 , C1 , n402352 );
buf ( n402354 , n55078 );
buf ( n402355 , n402354 );
not ( n55081 , n402355 );
buf ( n402357 , n55081 );
not ( n55083 , n402357 );
buf ( n402359 , n392884 );
not ( n55085 , n402359 );
buf ( n402361 , n384562 );
not ( n55087 , n402361 );
or ( n55088 , n55085 , n55087 );
buf ( n402364 , n389894 );
buf ( n402365 , n392887 );
nand ( n55091 , n402364 , n402365 );
buf ( n402367 , n55091 );
buf ( n402368 , n402367 );
nand ( n55094 , n55088 , n402368 );
buf ( n402370 , n55094 );
buf ( n402371 , n402370 );
not ( n55097 , n402371 );
buf ( n402373 , n400311 );
not ( n55099 , n402373 );
buf ( n402375 , n55099 );
buf ( n402376 , n402375 );
not ( n55102 , n402376 );
or ( n55103 , n55097 , n55102 );
buf ( n402379 , n400305 );
buf ( n402380 , n384548 );
nand ( n55106 , n402379 , n402380 );
buf ( n402382 , n55106 );
buf ( n402383 , n402382 );
nand ( n55109 , n55103 , n402383 );
buf ( n402385 , n55109 );
buf ( n402386 , n402385 );
not ( n55112 , n402386 );
buf ( n402388 , n55112 );
not ( n55114 , n402388 );
and ( n55115 , n55083 , n55114 );
buf ( n402391 , n402357 );
buf ( n402392 , n402388 );
nand ( n55118 , n402391 , n402392 );
buf ( n402394 , n55118 );
buf ( n402395 , n397498 );
not ( n55121 , n402395 );
buf ( n402397 , n382994 );
not ( n55123 , n402397 );
or ( n55124 , n55121 , n55123 );
buf ( n402400 , n31963 );
buf ( n402401 , n397495 );
nand ( n55127 , n402400 , n402401 );
buf ( n402403 , n55127 );
buf ( n402404 , n402403 );
nand ( n55130 , n55124 , n402404 );
buf ( n402406 , n55130 );
not ( n55132 , n402406 );
not ( n55133 , n389744 );
or ( n55134 , n55132 , n55133 );
buf ( n402410 , n400197 );
buf ( n402411 , n389021 );
nand ( n55137 , n402410 , n402411 );
buf ( n402413 , n55137 );
nand ( n55139 , n55134 , n402413 );
buf ( n55140 , n55139 );
and ( n55141 , n402394 , n55140 );
nor ( n55142 , n55115 , n55141 );
buf ( n402418 , n55142 );
not ( n55144 , n402418 );
xor ( n55145 , n400161 , n400184 );
xor ( n55146 , n55145 , n400210 );
buf ( n402422 , n55146 );
buf ( n402423 , n402422 );
not ( n55149 , n402423 );
buf ( n402425 , n55149 );
buf ( n402426 , n402425 );
not ( n55152 , n402426 );
or ( n55153 , n55144 , n55152 );
not ( n55154 , n52713 );
not ( n55155 , n52755 );
and ( n55156 , n55154 , n55155 );
and ( n55157 , n52713 , n52755 );
nor ( n55158 , n55156 , n55157 );
not ( n55159 , n52743 );
and ( n55160 , n55158 , n55159 );
not ( n55161 , n55158 );
and ( n55162 , n55161 , n52743 );
nor ( n55163 , n55160 , n55162 );
buf ( n402439 , n55163 );
not ( n55165 , n402439 );
buf ( n402441 , n55165 );
buf ( n402442 , n402441 );
nand ( n55168 , n55153 , n402442 );
buf ( n402444 , n55168 );
buf ( n402445 , n402444 );
buf ( n402446 , n55142 );
not ( n55172 , n402446 );
buf ( n402448 , n402422 );
nand ( n55174 , n55172 , n402448 );
buf ( n402450 , n55174 );
buf ( n402451 , n402450 );
nand ( n55177 , n402445 , n402451 );
buf ( n402453 , n55177 );
buf ( n402454 , n402453 );
nand ( n55180 , n55047 , n402454 );
buf ( n402456 , n55180 );
buf ( n402457 , n402456 );
nand ( n55183 , n55044 , n402457 );
buf ( n402459 , n55183 );
buf ( n402460 , n402459 );
not ( n55186 , n402460 );
xor ( n55187 , n400288 , n400430 );
xor ( n55188 , n55187 , n401854 );
buf ( n402464 , n55188 );
buf ( n402465 , n402464 );
not ( n55191 , n402465 );
or ( n55192 , n55186 , n55191 );
buf ( n402468 , n402464 );
buf ( n402469 , n402459 );
or ( n55195 , n402468 , n402469 );
not ( n55196 , n54612 );
not ( n55197 , n54594 );
or ( n55198 , n55196 , n55197 );
or ( n55199 , n54612 , n54594 );
nand ( n55200 , n55198 , n55199 );
not ( n55201 , n54617 );
and ( n55202 , n55200 , n55201 );
not ( n55203 , n55200 );
and ( n55204 , n55203 , n54617 );
nor ( n55205 , n55202 , n55204 );
buf ( n402481 , n55205 );
not ( n55207 , n402481 );
buf ( n402483 , n55207 );
buf ( n402484 , n402483 );
not ( n55210 , n402484 );
xor ( n55211 , n52980 , n53096 );
xor ( n55212 , n55211 , n53116 );
not ( n55213 , n55212 );
not ( n55214 , n55213 );
buf ( n402490 , n55214 );
not ( n55216 , n402490 );
or ( n55217 , n55210 , n55216 );
buf ( n402493 , n55205 );
not ( n55219 , n402493 );
buf ( n402495 , n55213 );
not ( n55221 , n402495 );
or ( n55222 , n55219 , n55221 );
buf ( n402498 , C1 );
not ( n55259 , n53003 );
not ( n55260 , n400326 );
or ( n55261 , n55259 , n55260 );
buf ( n402502 , n400323 );
buf ( n402503 , n400316 );
nand ( n55264 , n402502 , n402503 );
buf ( n402505 , n55264 );
nand ( n55266 , n55261 , n402505 );
buf ( n402507 , n53092 );
not ( n55268 , n402507 );
buf ( n402509 , n55268 );
not ( n55270 , n402509 );
and ( n55271 , n55266 , n55270 );
not ( n55272 , n55266 );
and ( n55273 , n55272 , n402509 );
nor ( n55274 , n55271 , n55273 );
xor ( n55275 , n402498 , n55274 );
xor ( n55276 , n400613 , n401773 );
xor ( n55277 , n55276 , n401794 );
buf ( n402518 , n55277 );
buf ( n402519 , n399274 );
not ( n55280 , n402519 );
buf ( n402521 , n40714 );
not ( n55282 , n402521 );
or ( n55283 , n55280 , n55282 );
buf ( n402524 , n40711 );
buf ( n402525 , n399283 );
nand ( n55286 , n402524 , n402525 );
buf ( n402527 , n55286 );
buf ( n402528 , n402527 );
nand ( n55289 , n55283 , n402528 );
buf ( n402530 , n55289 );
buf ( n402531 , n402530 );
not ( n55292 , n402531 );
buf ( n402533 , n396868 );
not ( n55294 , n402533 );
or ( n55295 , n55292 , n55294 );
buf ( n402536 , n383137 );
buf ( n402537 , n53132 );
nand ( n55298 , n402536 , n402537 );
buf ( n402539 , n55298 );
buf ( n402540 , n402539 );
nand ( n55301 , n55295 , n402540 );
buf ( n402542 , n55301 );
xor ( n55303 , n402518 , n402542 );
xor ( n55304 , n53040 , n53058 );
xnor ( n55305 , n55304 , n53088 );
and ( n55306 , n55303 , n55305 );
and ( n55307 , n402518 , n402542 );
or ( n55308 , n55306 , n55307 );
and ( n55309 , n55275 , n55308 );
and ( n402550 , n402498 , n55274 );
or ( n55311 , n55309 , n402550 );
buf ( n402552 , n55311 );
nand ( n55313 , n55222 , n402552 );
buf ( n402554 , n55313 );
buf ( n402555 , n402554 );
nand ( n55316 , n55217 , n402555 );
buf ( n402557 , n55316 );
buf ( n402558 , n402557 );
nand ( n55319 , n55195 , n402558 );
buf ( n402560 , n55319 );
buf ( n402561 , n402560 );
nand ( n55322 , n55192 , n402561 );
buf ( n402563 , n55322 );
buf ( n402564 , n402563 );
xor ( n55325 , n402289 , n402564 );
xor ( n55326 , n399974 , n399977 );
xor ( n55327 , n55326 , n400278 );
buf ( n402568 , n55327 );
buf ( n402569 , n402568 );
and ( n55330 , n55325 , n402569 );
and ( n55331 , n402289 , n402564 );
or ( n55332 , n55330 , n55331 );
buf ( n402573 , n55332 );
buf ( n402574 , n402573 );
not ( n55335 , n402574 );
or ( n55336 , n54819 , n55335 );
buf ( n402577 , n402573 );
not ( n55338 , n402577 );
buf ( n402579 , n55338 );
buf ( n402580 , n402579 );
not ( n55341 , n402580 );
buf ( n402582 , n402097 );
not ( n55343 , n402582 );
buf ( n402584 , n55343 );
buf ( n402585 , n402584 );
not ( n55346 , n402585 );
or ( n55347 , n55341 , n55346 );
xor ( n55348 , n401859 , n401945 );
xor ( n55349 , n55348 , n401957 );
buf ( n402590 , n55349 );
xor ( n55351 , n401885 , n401889 );
xor ( n55352 , n55351 , n401940 );
buf ( n402593 , n55352 );
not ( n55354 , n402593 );
buf ( n402595 , n400419 );
buf ( n402596 , n392740 );
and ( n55357 , n402595 , n402596 );
and ( n55358 , n37173 , n44776 );
not ( n55359 , n37173 );
and ( n55360 , n55359 , n392247 );
or ( n55361 , n55358 , n55360 );
buf ( n402602 , n55361 );
buf ( n402603 , n45260 );
and ( n55364 , n402602 , n402603 );
buf ( n402605 , n55364 );
buf ( n402606 , n402605 );
nor ( n55367 , n55357 , n402606 );
buf ( n402608 , n55367 );
buf ( n402609 , n402608 );
buf ( n402610 , n47726 );
not ( n55371 , n402610 );
buf ( n402612 , n400348 );
not ( n55373 , n402612 );
or ( n55374 , n55371 , n55373 );
not ( n55375 , n40817 );
not ( n55376 , n388154 );
or ( n55377 , n55375 , n55376 );
nand ( n55378 , n28215 , n394884 );
nand ( n55379 , n55377 , n55378 );
buf ( n402620 , n55379 );
buf ( n402621 , n397476 );
nand ( n55382 , n402620 , n402621 );
buf ( n402623 , n55382 );
buf ( n402624 , n402623 );
nand ( n55385 , n55374 , n402624 );
buf ( n402626 , n55385 );
buf ( n402627 , n402626 );
not ( n55388 , n35225 );
not ( n55389 , n55388 );
nand ( n55390 , n55389 , n382989 );
buf ( n402631 , n55390 );
buf ( n402632 , n358975 );
and ( n55393 , n402631 , n402632 );
not ( n55394 , n55388 );
not ( n55395 , n35400 );
or ( n55396 , n55394 , n55395 );
nand ( n55397 , n55396 , n385328 );
buf ( n402638 , n55397 );
nor ( n55399 , n55393 , n402638 );
buf ( n402640 , n55399 );
buf ( n402641 , n402640 );
xor ( n55402 , n402627 , n402641 );
buf ( n402643 , n42073 );
not ( n55404 , n402643 );
buf ( n402645 , n388272 );
not ( n55406 , n402645 );
or ( n55407 , n55404 , n55406 );
buf ( n402648 , n388263 );
buf ( n402649 , n42074 );
nand ( n55410 , n402648 , n402649 );
buf ( n402651 , n55410 );
buf ( n402652 , n402651 );
nand ( n55413 , n55407 , n402652 );
buf ( n402654 , n55413 );
buf ( n402655 , n402654 );
not ( n55416 , n402655 );
buf ( n402657 , n383894 );
not ( n55418 , n402657 );
or ( n55419 , n55416 , n55418 );
buf ( n402660 , n53049 );
buf ( n402661 , n383907 );
nand ( n55422 , n402660 , n402661 );
buf ( n402663 , n55422 );
buf ( n402664 , n402663 );
nand ( n55425 , n55419 , n402664 );
buf ( n402666 , n55425 );
buf ( n402667 , n402666 );
and ( n55428 , n55402 , n402667 );
and ( n55429 , n402627 , n402641 );
or ( n55430 , n55428 , n55429 );
buf ( n402671 , n55430 );
not ( n55432 , n402671 );
buf ( n402673 , n54873 );
not ( n55434 , n402673 );
buf ( n402675 , n388806 );
not ( n55436 , n402675 );
and ( n55437 , n55434 , n55436 );
buf ( n402678 , n388757 );
not ( n55439 , n402678 );
buf ( n402680 , n38155 );
not ( n55441 , n402680 );
or ( n55442 , n55439 , n55441 );
buf ( n402683 , n36564 );
buf ( n402684 , n388757 );
or ( n55445 , n402683 , n402684 );
buf ( n402686 , n55445 );
buf ( n402687 , n402686 );
nand ( n55448 , n55442 , n402687 );
buf ( n402689 , n55448 );
buf ( n402690 , n402689 );
buf ( n402691 , n388746 );
and ( n55452 , n402690 , n402691 );
nor ( n55453 , n55437 , n55452 );
buf ( n402694 , n55453 );
buf ( n402695 , n394817 );
not ( n55456 , n402695 );
buf ( n402697 , n395919 );
not ( n55458 , n402697 );
or ( n55459 , n55456 , n55458 );
buf ( n402700 , n385630 );
buf ( n402701 , n394814 );
nand ( n55462 , n402700 , n402701 );
buf ( n402703 , n55462 );
buf ( n402704 , n402703 );
nand ( n55465 , n55459 , n402704 );
buf ( n402706 , n55465 );
buf ( n402707 , n402706 );
not ( n55468 , n402707 );
buf ( n402709 , n383470 );
not ( n55470 , n402709 );
or ( n55471 , n55468 , n55470 );
buf ( n402712 , n391170 );
buf ( n402713 , n401833 );
nand ( n55474 , n402712 , n402713 );
buf ( n402715 , n55474 );
buf ( n402716 , n402715 );
nand ( n55477 , n55471 , n402716 );
buf ( n402718 , n55477 );
not ( n55479 , n402718 );
nand ( n55480 , n402694 , n55479 );
not ( n55481 , n55480 );
or ( n55482 , n55432 , n55481 );
buf ( n402723 , n402718 );
buf ( n402724 , n402694 );
not ( n55485 , n402724 );
buf ( n402726 , n55485 );
buf ( n402727 , n402726 );
nand ( n55488 , n402723 , n402727 );
buf ( n402729 , n55488 );
nand ( n55490 , n55482 , n402729 );
not ( n55491 , n55490 );
buf ( n402732 , n55491 );
and ( n55493 , n402609 , n402732 );
buf ( n402734 , n55493 );
buf ( n402735 , n402734 );
xor ( n55496 , n401799 , n401824 );
xor ( n55497 , n55496 , n401847 );
buf ( n402738 , n55497 );
buf ( n402739 , n402738 );
not ( n55500 , n402739 );
buf ( n402741 , n55500 );
buf ( n402742 , n402741 );
or ( n55503 , n402735 , n402742 );
buf ( n402744 , n55491 );
buf ( n402745 , n402608 );
or ( n55506 , n402744 , n402745 );
buf ( n402747 , n55506 );
buf ( n402748 , n402747 );
nand ( n55509 , n55503 , n402748 );
buf ( n402750 , n55509 );
buf ( n402751 , n402750 );
xor ( n55512 , n402042 , n402044 );
xor ( n55513 , n55512 , n402070 );
buf ( n402754 , n55513 );
buf ( n402755 , n402754 );
xor ( n55516 , n402751 , n402755 );
xor ( n55517 , n400582 , n400583 );
buf ( n402758 , n55517 );
xor ( n55519 , n400580 , n402758 );
buf ( n402760 , n55519 );
buf ( n402761 , n44945 );
not ( n55522 , n402761 );
buf ( n402763 , n388105 );
not ( n55524 , n402763 );
and ( n55525 , n55522 , n55524 );
buf ( n402766 , n44945 );
buf ( n402767 , n388105 );
and ( n55528 , n402766 , n402767 );
nor ( n55529 , n55525 , n55528 );
buf ( n402770 , n55529 );
buf ( n402771 , n402770 );
not ( n55532 , n402771 );
buf ( n402773 , n388093 );
not ( n55534 , n402773 );
and ( n55535 , n55532 , n55534 );
buf ( n402776 , n402141 );
buf ( n402777 , n388068 );
and ( n55538 , n402776 , n402777 );
nor ( n55539 , n55535 , n55538 );
buf ( n402780 , n55539 );
buf ( n402781 , n402780 );
not ( n55542 , n402781 );
not ( n55543 , n51184 );
buf ( n402784 , n55543 );
not ( n55545 , n402784 );
buf ( n402786 , n382994 );
not ( n55547 , n402786 );
or ( n55548 , n55545 , n55547 );
buf ( n402789 , n389759 );
buf ( n402790 , n51185 );
nand ( n55551 , n402789 , n402790 );
buf ( n402792 , n55551 );
buf ( n402793 , n402792 );
nand ( n55554 , n55548 , n402793 );
buf ( n402795 , n55554 );
buf ( n402796 , n402795 );
not ( n55557 , n402796 );
buf ( n402798 , n392834 );
not ( n55559 , n402798 );
or ( n55560 , n55557 , n55559 );
buf ( n402801 , n402406 );
buf ( n402802 , n389021 );
nand ( n55563 , n402801 , n402802 );
buf ( n402804 , n55563 );
buf ( n402805 , n402804 );
nand ( n55566 , n55560 , n402805 );
buf ( n402807 , n55566 );
buf ( n402808 , n402807 );
not ( n55569 , n402808 );
buf ( n402810 , n55569 );
not ( n55571 , n402810 );
not ( n55572 , n389348 );
not ( n55573 , n55572 );
not ( n55574 , n402347 );
not ( n55575 , n55574 );
or ( n55576 , n55573 , n55575 );
buf ( n402817 , n358975 );
not ( n55583 , n402817 );
buf ( n402819 , n55583 );
nand ( n55590 , C1 , n389348 );
nand ( n55591 , n55576 , n55590 );
not ( n55592 , n55591 );
and ( n55593 , n55571 , n55592 );
buf ( n402824 , n402810 );
buf ( n402825 , n55591 );
nand ( n55596 , n402824 , n402825 );
buf ( n402827 , n55596 );
buf ( n402828 , n394666 );
not ( n55599 , n402828 );
buf ( n402830 , n398298 );
not ( n55601 , n402830 );
or ( n55602 , n55599 , n55601 );
buf ( n402833 , n24049 );
buf ( n402834 , n27258 );
not ( n55605 , n402834 );
buf ( n402836 , n55605 );
buf ( n402837 , n402836 );
nand ( n55608 , n402833 , n402837 );
buf ( n402839 , n55608 );
buf ( n402840 , n402839 );
nand ( n55611 , n55602 , n402840 );
buf ( n402842 , n55611 );
buf ( n402843 , n402842 );
not ( n55614 , n402843 );
buf ( n402845 , n396622 );
not ( n55616 , n402845 );
or ( n55617 , n55614 , n55616 );
buf ( n402848 , n400627 );
not ( n55619 , n402848 );
buf ( n402850 , n41563 );
nand ( n55621 , n55619 , n402850 );
buf ( n402852 , n55621 );
buf ( n402853 , n402852 );
nand ( n55624 , n55617 , n402853 );
buf ( n402855 , n55624 );
buf ( n402856 , n402855 );
buf ( n402857 , n388998 );
not ( n55628 , n402857 );
buf ( n402859 , n388965 );
not ( n55630 , n402859 );
or ( n55631 , n55628 , n55630 );
buf ( n402862 , n388962 );
buf ( n402863 , n388215 );
nand ( n55634 , n402862 , n402863 );
buf ( n402865 , n55634 );
buf ( n402866 , n402865 );
nand ( n55637 , n55631 , n402866 );
buf ( n402868 , n55637 );
buf ( n402869 , n402868 );
not ( n55640 , n402869 );
buf ( n402871 , n46056 );
not ( n55642 , n402871 );
or ( n55643 , n55640 , n55642 );
buf ( n402874 , n37923 );
not ( n55645 , n402874 );
buf ( n402876 , n400534 );
nand ( n55647 , n55645 , n402876 );
buf ( n402878 , n55647 );
buf ( n402879 , n402878 );
nand ( n55650 , n55643 , n402879 );
buf ( n402881 , n55650 );
buf ( n402882 , n402881 );
xor ( n55653 , n402856 , n402882 );
buf ( n402884 , n397476 );
not ( n55655 , n402884 );
not ( n55656 , n388406 );
not ( n55657 , n388154 );
or ( n55658 , n55656 , n55657 );
nand ( n55659 , n46043 , n394884 );
nand ( n55660 , n55658 , n55659 );
buf ( n402891 , n55660 );
not ( n55662 , n402891 );
or ( n55663 , n55655 , n55662 );
buf ( n402894 , n55379 );
buf ( n402895 , n47726 );
nand ( n55666 , n402894 , n402895 );
buf ( n402897 , n55666 );
buf ( n402898 , n402897 );
nand ( n55669 , n55663 , n402898 );
buf ( n402900 , n55669 );
buf ( n402901 , n402900 );
and ( n55672 , n55653 , n402901 );
and ( n55673 , n402856 , n402882 );
or ( n55674 , n55672 , n55673 );
buf ( n402905 , n55674 );
and ( n55676 , n402827 , n402905 );
nor ( n55677 , n55593 , n55676 );
buf ( n402908 , n55677 );
not ( n55679 , n402908 );
or ( n55680 , n55542 , n55679 );
buf ( n402911 , n392611 );
not ( n55682 , n402911 );
buf ( n402913 , n390875 );
not ( n55684 , n402913 );
or ( n55685 , n55682 , n55684 );
buf ( n402916 , n40885 );
buf ( n402917 , n392620 );
nand ( n55688 , n402916 , n402917 );
buf ( n402919 , n55688 );
buf ( n402920 , n402919 );
nand ( n55691 , n55685 , n402920 );
buf ( n402922 , n55691 );
buf ( n402923 , n402922 );
not ( n55694 , n402923 );
buf ( n402925 , n40858 );
not ( n55696 , n402925 );
or ( n55697 , n55694 , n55696 );
nand ( n55698 , n392111 , n53172 );
buf ( n402929 , n55698 );
nand ( n55700 , n55697 , n402929 );
buf ( n402931 , n55700 );
not ( n55702 , n402931 );
and ( n55703 , n389341 , n40972 );
not ( n55704 , n389341 );
and ( n55705 , n55704 , n36395 );
nor ( n55706 , n55703 , n55705 );
buf ( n402937 , n55706 );
not ( n55708 , n402937 );
buf ( n402939 , n397165 );
not ( n55710 , n402939 );
or ( n55711 , n55708 , n55710 );
buf ( n402942 , n400464 );
buf ( n402943 , n388346 );
nand ( n55714 , n402942 , n402943 );
buf ( n402945 , n55714 );
buf ( n402946 , n402945 );
nand ( n55717 , n55711 , n402946 );
buf ( n402948 , n55717 );
not ( n55719 , n402948 );
or ( n55720 , n55702 , n55719 );
buf ( n402951 , n402931 );
buf ( n402952 , n402948 );
nor ( n55723 , n402951 , n402952 );
buf ( n402954 , n55723 );
buf ( n402955 , n388833 );
not ( n55726 , n402955 );
buf ( n402957 , n400391 );
not ( n55728 , n402957 );
or ( n55729 , n55726 , n55728 );
buf ( n402960 , n41342 );
not ( n55731 , n402960 );
buf ( n402962 , n40759 );
not ( n55733 , n402962 );
or ( n55734 , n55731 , n55733 );
buf ( n402965 , n40758 );
buf ( n402966 , n45897 );
nand ( n55737 , n402965 , n402966 );
buf ( n402968 , n55737 );
buf ( n402969 , n402968 );
nand ( n55740 , n55734 , n402969 );
buf ( n402971 , n55740 );
buf ( n402972 , n402971 );
buf ( n402973 , n388872 );
nand ( n55744 , n402972 , n402973 );
buf ( n402975 , n55744 );
buf ( n402976 , n402975 );
nand ( n55747 , n55729 , n402976 );
buf ( n402978 , n55747 );
buf ( n402979 , n402978 );
not ( n55750 , n402979 );
buf ( n402981 , n55750 );
or ( n55752 , n402954 , n402981 );
nand ( n55753 , n55720 , n55752 );
buf ( n402984 , n55753 );
nand ( n55755 , n55680 , n402984 );
buf ( n402986 , n55755 );
buf ( n402987 , n402986 );
buf ( n402988 , n402780 );
not ( n55759 , n402988 );
buf ( n402990 , n55677 );
not ( n55761 , n402990 );
buf ( n402992 , n55761 );
buf ( n402993 , n402992 );
nand ( n55764 , n55759 , n402993 );
buf ( n402995 , n55764 );
buf ( n402996 , n402995 );
nand ( n55767 , n402987 , n402996 );
buf ( n402998 , n55767 );
buf ( n402999 , n402998 );
xor ( n55770 , n402760 , n402999 );
buf ( n403001 , n400520 );
buf ( n403002 , n400568 );
xor ( n55773 , n403001 , n403002 );
buf ( n403004 , n400546 );
xnor ( n55775 , n55773 , n403004 );
buf ( n403006 , n55775 );
buf ( n403007 , n403006 );
buf ( n403008 , n389162 );
not ( n55779 , n403008 );
buf ( n403010 , n402186 );
not ( n55781 , n403010 );
or ( n55782 , n55779 , n55781 );
and ( n55783 , n28159 , n24117 );
not ( n55784 , n28159 );
and ( n55785 , n55784 , n24116 );
or ( n55786 , n55783 , n55785 );
buf ( n403017 , n55786 );
buf ( n403018 , n41711 );
nand ( n55789 , n403017 , n403018 );
buf ( n403020 , n55789 );
buf ( n403021 , n403020 );
nand ( n55792 , n55782 , n403021 );
buf ( n403023 , n55792 );
buf ( n403024 , n403023 );
not ( n55795 , n403024 );
buf ( n403026 , n55795 );
buf ( n403027 , n403026 );
nand ( n55798 , n403007 , n403027 );
buf ( n403029 , n55798 );
buf ( n403030 , n403029 );
not ( n55801 , n403030 );
xor ( n55802 , n401655 , n401685 );
xor ( n55803 , n55802 , n401758 );
buf ( n403034 , n55803 );
buf ( n403035 , n403034 );
not ( n55806 , n403035 );
buf ( n403037 , n28644 );
not ( n55808 , n403037 );
buf ( n403039 , n55808 );
buf ( n403040 , n403039 );
not ( n55811 , n403040 );
buf ( n403042 , n55811 );
buf ( n403043 , n403042 );
not ( n55814 , n403043 );
buf ( n403045 , n399164 );
not ( n55816 , n403045 );
or ( n55817 , n55814 , n55816 );
buf ( n403048 , n28644 );
not ( n55819 , n403048 );
buf ( n403050 , n24049 );
nand ( n55821 , n55819 , n403050 );
buf ( n403052 , n55821 );
buf ( n403053 , n403052 );
nand ( n55824 , n55817 , n403053 );
buf ( n403055 , n55824 );
buf ( n403056 , n403055 );
not ( n55827 , n403056 );
buf ( n403058 , n396622 );
not ( n55829 , n403058 );
or ( n55830 , n55827 , n55829 );
not ( n55831 , n41562 );
buf ( n403062 , n55831 );
buf ( n403063 , n402842 );
nand ( n55834 , n403062 , n403063 );
buf ( n403065 , n55834 );
buf ( n403066 , n403065 );
nand ( n55837 , n55830 , n403066 );
buf ( n403068 , n55837 );
buf ( n403069 , n403068 );
not ( n55840 , n403069 );
buf ( n403071 , n55840 );
buf ( n403072 , n403071 );
not ( n55843 , n403072 );
or ( n55844 , n55806 , n55843 );
nand ( n55845 , n53453 , n54425 );
xnor ( n55846 , n55845 , n54328 );
buf ( n403077 , n55846 );
not ( n55848 , n403077 );
buf ( n403079 , n55848 );
buf ( n403080 , n403079 );
buf ( n403081 , n401626 );
not ( n55852 , n403081 );
buf ( n403083 , n55852 );
buf ( n403084 , n403083 );
or ( n55855 , n403080 , n403084 );
buf ( n403086 , n54433 );
not ( n55857 , n403086 );
buf ( n403088 , n55857 );
buf ( n403089 , n403088 );
buf ( n403090 , n401650 );
not ( n55861 , n403090 );
buf ( n403092 , n55861 );
buf ( n403093 , n403092 );
or ( n55864 , n403089 , n403093 );
nand ( n55865 , n55855 , n55864 );
buf ( n403096 , n55865 );
not ( n55867 , n4031 );
not ( n55868 , n351734 );
or ( n55869 , n55867 , n55868 );
nand ( n55870 , n55869 , n351739 );
not ( n55871 , n55870 );
not ( n55872 , n353695 );
or ( n55873 , n55871 , n55872 );
or ( n55874 , n353695 , n55870 );
nand ( n55875 , n55873 , n55874 );
buf ( n403106 , n55875 );
not ( n55877 , n403106 );
buf ( n403108 , n55877 );
buf ( n403109 , n403108 );
buf ( n403110 , n15287 );
buf ( n403111 , n353695 );
and ( n55882 , n403110 , n403111 );
buf ( n403113 , n15290 );
buf ( n403114 , n353618 );
and ( n55885 , n403113 , n403114 );
nor ( n55886 , n55882 , n55885 );
buf ( n403117 , n55886 );
buf ( n403118 , n403117 );
nand ( n55889 , n403109 , n403118 );
buf ( n403120 , n55889 );
buf ( n403121 , n403120 );
not ( n55892 , n403121 );
buf ( n403123 , n55892 );
buf ( n403124 , n403123 );
not ( n55895 , n15287 );
buf ( n403126 , n55895 );
nand ( n55897 , n403124 , n403126 );
buf ( n403128 , n55897 );
buf ( n403129 , n403128 );
not ( n55900 , n403129 );
buf ( n403131 , n55875 );
not ( n55902 , n403131 );
buf ( n403133 , n55902 );
buf ( n403134 , n403133 );
not ( n55905 , n55895 );
buf ( n403136 , n55905 );
nor ( n55907 , n403134 , n403136 );
buf ( n403138 , n55907 );
buf ( n403139 , n403138 );
nor ( n55910 , n55900 , n403139 );
buf ( n403141 , n55910 );
xor ( n55912 , n403096 , n403141 );
buf ( n403143 , n54297 );
buf ( n403144 , n401695 );
not ( n55915 , n403144 );
buf ( n403146 , n55915 );
buf ( n403147 , n403146 );
and ( n55918 , n403143 , n403147 );
not ( n55919 , n54297 );
buf ( n403150 , n55919 );
buf ( n403151 , n401695 );
and ( n55922 , n403150 , n403151 );
nor ( n55923 , n55918 , n55922 );
buf ( n403154 , n55923 );
buf ( n403155 , n403154 );
buf ( n403156 , n401674 );
not ( n55927 , n403156 );
buf ( n403158 , n55927 );
buf ( n403159 , n403158 );
or ( n55930 , n403155 , n403159 );
buf ( n403161 , n401706 );
buf ( n403162 , n401660 );
not ( n55933 , n403162 );
buf ( n403164 , n55933 );
buf ( n403165 , n403164 );
not ( n55936 , n403165 );
buf ( n403167 , n55936 );
buf ( n403168 , n403167 );
or ( n55939 , n403161 , n403168 );
nand ( n55940 , n55930 , n55939 );
buf ( n403171 , n55940 );
and ( n55942 , n55912 , n403171 );
and ( n55943 , n403096 , n403141 );
or ( n55944 , n55942 , n55943 );
buf ( n403175 , n55944 );
buf ( n403176 , n401715 );
buf ( n403177 , n401751 );
or ( n55948 , n403176 , n403177 );
buf ( n403179 , n401754 );
nand ( n55950 , n55948 , n403179 );
buf ( n403181 , n55950 );
buf ( n403182 , n403181 );
xor ( n55953 , n403175 , n403182 );
buf ( n403184 , n55905 );
buf ( n403185 , n54336 );
and ( n55956 , n403184 , n403185 );
not ( n55957 , n403184 );
buf ( n403188 , n401699 );
and ( n55959 , n55957 , n403188 );
nor ( n55960 , n55956 , n55959 );
buf ( n403191 , n55960 );
buf ( n403192 , n403191 );
not ( n55963 , n403192 );
buf ( n403194 , n55963 );
buf ( n403195 , n403194 );
buf ( n403196 , n403123 );
and ( n55967 , n403195 , n403196 );
buf ( n403198 , n403138 );
nor ( n55969 , n55967 , n403198 );
buf ( n403200 , n55969 );
buf ( n403201 , n403200 );
and ( n55972 , n53653 , n53419 , n53472 );
not ( n55973 , n55972 );
not ( n55974 , n54414 );
or ( n55975 , n55973 , n55974 );
and ( n55976 , n54420 , n53472 );
nor ( n55977 , n55976 , n54279 );
nand ( n55978 , n55975 , n55977 );
not ( n55979 , n54283 );
nand ( n55980 , n55979 , n53442 );
nor ( n55981 , n55978 , n55980 );
not ( n55982 , n55981 );
nand ( n55983 , n55978 , n55980 );
nand ( n55984 , n55982 , n55983 );
buf ( n403215 , n55984 );
buf ( n403216 , n401626 );
and ( n55987 , n403215 , n403216 );
buf ( n403218 , n55846 );
buf ( n403219 , n401650 );
and ( n55990 , n403218 , n403219 );
nor ( n55991 , n55987 , n55990 );
buf ( n403222 , n55991 );
buf ( n403223 , n403222 );
nand ( n55994 , n403201 , n403223 );
buf ( n403225 , n55994 );
xor ( n55996 , n403096 , n403141 );
xor ( n55997 , n55996 , n403171 );
and ( n55998 , n403225 , n55997 );
buf ( n403229 , n403200 );
buf ( n403230 , n403222 );
or ( n56001 , n403229 , n403230 );
buf ( n403232 , n403225 );
nand ( n56003 , n56001 , n403232 );
buf ( n403234 , n56003 );
buf ( n403235 , n403234 );
buf ( n403236 , n403146 );
buf ( n403237 , n54433 );
and ( n56008 , n403236 , n403237 );
not ( n56009 , n403236 );
buf ( n403240 , n403088 );
and ( n56011 , n56009 , n403240 );
nor ( n56012 , n56008 , n56011 );
buf ( n403243 , n56012 );
buf ( n403244 , n403243 );
buf ( n403245 , n403158 );
or ( n56016 , n403244 , n403245 );
buf ( n403247 , n403154 );
buf ( n403248 , n403167 );
or ( n56019 , n403247 , n403248 );
nand ( n56020 , n56016 , n56019 );
buf ( n403251 , n56020 );
buf ( n403252 , n403251 );
xor ( n56023 , n403235 , n403252 );
buf ( n403254 , n54297 );
buf ( n403255 , n55905 );
and ( n56026 , n403254 , n403255 );
buf ( n403257 , n55919 );
buf ( n403258 , n55895 );
and ( n56029 , n403257 , n403258 );
nor ( n56030 , n56026 , n56029 );
buf ( n403261 , n56030 );
buf ( n403262 , n403261 );
buf ( n403263 , n403120 );
or ( n56034 , n403262 , n403263 );
buf ( n403265 , n403191 );
buf ( n403266 , n403133 );
or ( n56037 , n403265 , n403266 );
nand ( n56038 , n56034 , n56037 );
buf ( n403269 , n56038 );
buf ( n403270 , n403269 );
not ( n56041 , n55870 );
not ( n56042 , n56041 );
not ( n56043 , n5730 );
or ( n56044 , n56042 , n56043 );
buf ( n56045 , n2071 );
or ( n56046 , n56045 , n56041 );
nand ( n56047 , n56044 , n56046 );
buf ( n403278 , n56047 );
buf ( n403279 , n56045 );
buf ( n56050 , n5720 );
buf ( n403281 , n56050 );
not ( n56052 , n403281 );
buf ( n403283 , n56052 );
buf ( n403284 , n403283 );
and ( n56055 , n403279 , n403284 );
not ( n56056 , n403279 );
buf ( n403287 , n56050 );
and ( n56058 , n56056 , n403287 );
nor ( n56059 , n56055 , n56058 );
buf ( n403290 , n56059 );
buf ( n403291 , n403290 );
nand ( n56062 , n403278 , n403291 );
buf ( n403293 , n56062 );
not ( n56064 , n403293 );
buf ( n403295 , n56064 );
buf ( n403296 , n56041 );
not ( n56067 , n403296 );
buf ( n403298 , n56067 );
buf ( n403299 , n403298 );
nand ( n56070 , n403295 , n403299 );
buf ( n403301 , n56070 );
buf ( n403302 , n403301 );
buf ( n403303 , n403290 );
not ( n56074 , n403303 );
buf ( n403305 , n56074 );
buf ( n403306 , n403305 );
buf ( n403307 , n403298 );
nand ( n56078 , n403306 , n403307 );
buf ( n403309 , n56078 );
buf ( n403310 , n403309 );
and ( n56081 , n403302 , n403310 );
buf ( n403312 , n56081 );
buf ( n403313 , n403312 );
xor ( n56084 , n403270 , n403313 );
buf ( n403315 , n55846 );
buf ( n403316 , n403146 );
and ( n56087 , n403315 , n403316 );
buf ( n403318 , n403079 );
buf ( n403319 , n401695 );
and ( n56090 , n403318 , n403319 );
nor ( n56091 , n56087 , n56090 );
buf ( n403322 , n56091 );
buf ( n403323 , n403322 );
buf ( n403324 , n403158 );
or ( n56095 , n403323 , n403324 );
buf ( n403326 , n403243 );
buf ( n403327 , n403167 );
or ( n56098 , n403326 , n403327 );
nand ( n56099 , n56095 , n56098 );
buf ( n403330 , n56099 );
buf ( n403331 , n403330 );
and ( n56102 , n56084 , n403331 );
and ( n56103 , n403270 , n403313 );
or ( n56104 , n56102 , n56103 );
buf ( n403335 , n56104 );
buf ( n403336 , n403335 );
and ( n56107 , n56023 , n403336 );
and ( n56108 , n403235 , n403252 );
or ( n56109 , n56107 , n56108 );
buf ( n403340 , n56109 );
xor ( n56111 , n403096 , n403141 );
xor ( n56112 , n56111 , n403171 );
and ( n56113 , n403340 , n56112 );
and ( n56114 , n403225 , n403340 );
or ( n56115 , n55998 , n56113 , n56114 );
buf ( n403346 , n56115 );
and ( n56117 , n55953 , n403346 );
and ( n56118 , n403175 , n403182 );
or ( n56119 , n56117 , n56118 );
buf ( n403350 , n56119 );
buf ( n403351 , n403350 );
nand ( n56122 , n55844 , n403351 );
buf ( n403353 , n56122 );
buf ( n403354 , n403353 );
buf ( n403355 , n403034 );
not ( n56126 , n403355 );
buf ( n403357 , n403068 );
nand ( n56128 , n56126 , n403357 );
buf ( n403359 , n56128 );
buf ( n403360 , n403359 );
nand ( n56131 , n403354 , n403360 );
buf ( n403362 , n56131 );
buf ( n403363 , n403362 );
buf ( n403364 , n388872 );
not ( n56135 , n403364 );
buf ( n403366 , n41342 );
not ( n56137 , n403366 );
buf ( n403368 , n40831 );
not ( n56139 , n403368 );
or ( n56140 , n56137 , n56139 );
buf ( n403371 , n27195 );
buf ( n403372 , n45897 );
nand ( n56143 , n403371 , n403372 );
buf ( n403374 , n56143 );
buf ( n403375 , n403374 );
nand ( n56146 , n56140 , n403375 );
buf ( n403377 , n56146 );
buf ( n403378 , n403377 );
not ( n56149 , n403378 );
or ( n56150 , n56135 , n56149 );
buf ( n403381 , n402971 );
buf ( n403382 , n388833 );
nand ( n56153 , n403381 , n403382 );
buf ( n403384 , n56153 );
buf ( n403385 , n403384 );
nand ( n56156 , n56150 , n403385 );
buf ( n403387 , n56156 );
buf ( n403388 , n403387 );
xor ( n56159 , n403363 , n403388 );
buf ( n403390 , n40990 );
not ( n56161 , n403390 );
buf ( n403392 , n390548 );
not ( n56163 , n403392 );
or ( n56164 , n56161 , n56163 );
buf ( n403395 , n388905 );
buf ( n403396 , n390460 );
nand ( n56167 , n403395 , n403396 );
buf ( n403398 , n56167 );
buf ( n403399 , n403398 );
nand ( n56170 , n56164 , n403399 );
buf ( n403401 , n56170 );
buf ( n403402 , n403401 );
not ( n56173 , n403402 );
buf ( n403404 , n56173 );
or ( n56175 , n403404 , n43058 );
nand ( n56176 , n37316 , n54926 );
nand ( n56177 , n56175 , n56176 );
buf ( n403408 , n56177 );
and ( n56179 , n56159 , n403408 );
and ( n56180 , n403363 , n403388 );
or ( n56181 , n56179 , n56180 );
buf ( n403412 , n56181 );
buf ( n403413 , n403412 );
not ( n56184 , n403413 );
or ( n56185 , n55801 , n56184 );
buf ( n403416 , n403006 );
not ( n56187 , n403416 );
buf ( n403418 , n56187 );
buf ( n403419 , n403418 );
buf ( n403420 , n403023 );
nand ( n56191 , n403419 , n403420 );
buf ( n403422 , n56191 );
buf ( n403423 , n403422 );
nand ( n56194 , n56185 , n403423 );
buf ( n403425 , n56194 );
buf ( n403426 , n403425 );
buf ( n403427 , n43727 );
not ( n56198 , n403427 );
buf ( n403429 , n391027 );
not ( n56200 , n403429 );
buf ( n403431 , n384183 );
not ( n56202 , n403431 );
or ( n56203 , n56200 , n56202 );
buf ( n403434 , n390119 );
buf ( n403435 , n391024 );
nand ( n56206 , n403434 , n403435 );
buf ( n403437 , n56206 );
buf ( n403438 , n403437 );
nand ( n56209 , n56203 , n403438 );
buf ( n403440 , n56209 );
buf ( n403441 , n403440 );
not ( n56212 , n403441 );
or ( n56213 , n56198 , n56212 );
buf ( n403444 , n391027 );
not ( n56215 , n403444 );
buf ( n403446 , n42234 );
not ( n56217 , n403446 );
or ( n56218 , n56215 , n56217 );
buf ( n403449 , n36217 );
buf ( n403450 , n391024 );
nand ( n56221 , n403449 , n403450 );
buf ( n403452 , n56221 );
buf ( n403453 , n403452 );
nand ( n56224 , n56218 , n403453 );
buf ( n403455 , n56224 );
buf ( n403456 , n403455 );
buf ( n403457 , n43515 );
nand ( n56228 , n403456 , n403457 );
buf ( n403459 , n56228 );
buf ( n403460 , n403459 );
nand ( n56231 , n56213 , n403460 );
buf ( n403462 , n56231 );
buf ( n403463 , n403462 );
xor ( n56234 , n403426 , n403463 );
buf ( n403465 , n400574 );
buf ( n403466 , n400476 );
xor ( n56237 , n403465 , n403466 );
buf ( n403468 , n53180 );
xor ( n56239 , n56237 , n403468 );
buf ( n403470 , n56239 );
buf ( n403471 , n403470 );
and ( n56242 , n56234 , n403471 );
and ( n56243 , n403426 , n403463 );
or ( n56244 , n56242 , n56243 );
buf ( n403475 , n56244 );
buf ( n403476 , n403475 );
and ( n56247 , n55770 , n403476 );
and ( n56248 , n402760 , n402999 );
or ( n56249 , n56247 , n56248 );
buf ( n403480 , n56249 );
buf ( n403481 , n403480 );
and ( n56252 , n55516 , n403481 );
and ( n56253 , n402751 , n402755 );
or ( n56254 , n56252 , n56253 );
buf ( n403485 , n56254 );
not ( n56256 , n403485 );
or ( n56257 , n55354 , n56256 );
or ( n56258 , n402593 , n403485 );
xor ( n56259 , n402017 , n402074 );
xor ( n56260 , n56259 , n402078 );
buf ( n403491 , n56260 );
nand ( n56262 , n56258 , n403491 );
nand ( n56263 , n56257 , n56262 );
xor ( n56264 , n402590 , n56263 );
buf ( n403495 , n402012 );
buf ( n403496 , n402082 );
xor ( n56267 , n403495 , n403496 );
buf ( n403498 , n402009 );
xor ( n56269 , n56267 , n403498 );
buf ( n403500 , n56269 );
and ( n56271 , n56264 , n403500 );
and ( n56272 , n402590 , n56263 );
or ( n56273 , n56271 , n56272 );
buf ( n403504 , n56273 );
nand ( n56275 , n55347 , n403504 );
buf ( n403506 , n56275 );
buf ( n403507 , n403506 );
nand ( n56278 , n55336 , n403507 );
buf ( n403509 , n56278 );
buf ( n403510 , n403509 );
not ( n56281 , n403510 );
buf ( n403512 , n56281 );
buf ( n403513 , n403512 );
xor ( n56284 , n402094 , n403513 );
xor ( n56285 , n401970 , n401985 );
xor ( n56286 , n56285 , n401989 );
buf ( n403517 , n56286 );
buf ( n403518 , n403517 );
and ( n56289 , n56284 , n403518 );
and ( n56290 , n402094 , n403513 );
or ( n56291 , n56289 , n56290 );
buf ( n403522 , n56291 );
nand ( n56293 , n54684 , n403522 );
buf ( n403524 , n56293 );
xor ( n56295 , n399360 , n399850 );
xor ( n56296 , n56295 , n399863 );
buf ( n403527 , n56296 );
not ( n56298 , n403527 );
xor ( n56299 , n399955 , n52653 );
and ( n56300 , n56299 , n401993 );
and ( n56301 , n399955 , n52653 );
or ( n56302 , n56300 , n56301 );
nand ( n56303 , n56298 , n56302 );
buf ( n403534 , n56303 );
and ( n56305 , n403524 , n403534 );
buf ( n403536 , n56305 );
buf ( n403537 , n403536 );
xor ( n56308 , n401998 , n402002 );
xor ( n56309 , n56308 , n402089 );
buf ( n403540 , n56309 );
buf ( n403541 , n403540 );
buf ( n403542 , C0 );
buf ( n403543 , n403542 );
buf ( n403544 , n43515 );
not ( n56335 , n403544 );
buf ( n403546 , n402031 );
not ( n56337 , n403546 );
or ( n56338 , n56335 , n56337 );
buf ( n403549 , n403455 );
buf ( n403550 , n43727 );
nand ( n56341 , n403549 , n403550 );
buf ( n403552 , n56341 );
buf ( n403553 , n403552 );
nand ( n56344 , n56338 , n403553 );
buf ( n403555 , n56344 );
buf ( n403556 , n403555 );
xor ( n56347 , n403543 , n403556 );
buf ( n403558 , n45954 );
not ( n56349 , n403558 );
buf ( n403560 , n402062 );
not ( n56351 , n403560 );
or ( n56352 , n56349 , n56351 );
buf ( n403563 , n393369 );
not ( n56354 , n403563 );
buf ( n403565 , n396298 );
not ( n56356 , n403565 );
buf ( n403567 , n56356 );
buf ( n403568 , n403567 );
not ( n56359 , n403568 );
or ( n56360 , n56354 , n56359 );
buf ( n403571 , n389423 );
buf ( n403572 , n393381 );
nand ( n56363 , n403571 , n403572 );
buf ( n403574 , n56363 );
buf ( n403575 , n403574 );
nand ( n56366 , n56360 , n403575 );
buf ( n403577 , n56366 );
buf ( n403578 , n403577 );
buf ( n403579 , n393825 );
nand ( n56370 , n403578 , n403579 );
buf ( n403581 , n56370 );
buf ( n403582 , n403581 );
nand ( n56373 , n56352 , n403582 );
buf ( n403584 , n56373 );
buf ( n403585 , n403584 );
and ( n56376 , n56347 , n403585 );
or ( n56378 , n56376 , C0 );
buf ( n403588 , n56378 );
buf ( n403589 , n403588 );
buf ( n56381 , n53276 );
buf ( n403591 , n400606 );
not ( n56383 , n403591 );
buf ( n403593 , n401851 );
not ( n56385 , n403593 );
buf ( n403595 , n56385 );
buf ( n403596 , n403595 );
not ( n56388 , n403596 );
or ( n56389 , n56383 , n56388 );
buf ( n403599 , n401851 );
buf ( n403600 , n53293 );
nand ( n56392 , n403599 , n403600 );
buf ( n403602 , n56392 );
buf ( n403603 , n403602 );
nand ( n56395 , n56389 , n403603 );
buf ( n403605 , n56395 );
xnor ( n56397 , n56381 , n403605 );
buf ( n403607 , n56397 );
xor ( n56399 , n403589 , n403607 );
and ( n56400 , n54841 , n54833 );
not ( n56401 , n54841 );
and ( n56402 , n56401 , n54834 );
nor ( n56403 , n56400 , n56402 );
xor ( n56404 , n56403 , n402274 );
buf ( n403614 , n56404 );
and ( n56406 , n56399 , n403614 );
and ( n56407 , n403589 , n403607 );
or ( n56408 , n56406 , n56407 );
buf ( n403618 , n56408 );
buf ( n403619 , n403618 );
xor ( n56411 , n402103 , n402279 );
xor ( n56412 , n56411 , n402284 );
buf ( n403622 , n56412 );
buf ( n403623 , n403622 );
xor ( n56415 , n403619 , n403623 );
not ( n56416 , n45954 );
not ( n56417 , n403577 );
or ( n56418 , n56416 , n56417 );
buf ( n403628 , n393369 );
not ( n56420 , n403628 );
buf ( n403630 , n37147 );
not ( n56422 , n403630 );
or ( n56423 , n56420 , n56422 );
buf ( n403633 , n394463 );
buf ( n403634 , n393381 );
nand ( n56426 , n403633 , n403634 );
buf ( n403636 , n56426 );
buf ( n403637 , n403636 );
nand ( n56429 , n56423 , n403637 );
buf ( n403639 , n56429 );
nand ( n56431 , n403639 , n393825 );
nand ( n56432 , n56418 , n56431 );
or ( n56449 , C0 , n56432 );
not ( n56450 , n402726 );
not ( n56451 , n55479 );
or ( n56452 , n56450 , n56451 );
nand ( n56453 , n402718 , n402694 );
nand ( n56454 , n56452 , n56453 );
and ( n56455 , n56454 , n402671 );
not ( n56456 , n56454 );
buf ( n403650 , n402671 );
not ( n56458 , n403650 );
buf ( n403652 , n56458 );
and ( n56460 , n56456 , n403652 );
nor ( n56461 , n56455 , n56460 );
nand ( n56462 , n56449 , n56461 );
nand ( n56463 , C1 , n56462 );
not ( n56464 , n56463 );
buf ( n403658 , n50579 );
not ( n56466 , n403658 );
buf ( n403660 , n47891 );
not ( n56468 , n403660 );
buf ( n403662 , n386561 );
not ( n56470 , n403662 );
or ( n56471 , n56468 , n56470 );
buf ( n403665 , n382921 );
buf ( n403666 , n47891 );
not ( n56474 , n403666 );
buf ( n403668 , n56474 );
buf ( n403669 , n403668 );
nand ( n56477 , n403665 , n403669 );
buf ( n403671 , n56477 );
buf ( n403672 , n403671 );
nand ( n56480 , n56471 , n403672 );
buf ( n403674 , n56480 );
buf ( n403675 , n403674 );
not ( n56483 , n403675 );
or ( n56484 , n56466 , n56483 );
buf ( n403678 , n54831 );
buf ( n403679 , n51553 );
nand ( n56487 , n403678 , n403679 );
buf ( n403681 , n56487 );
buf ( n403682 , n403681 );
nand ( n56490 , n56484 , n403682 );
buf ( n403684 , n56490 );
buf ( n403685 , n403684 );
not ( n56493 , n403685 );
buf ( n403687 , n56493 );
nand ( n56495 , n56464 , n403687 );
not ( n56496 , n56495 );
buf ( n403690 , n402441 );
not ( n56498 , n403690 );
buf ( n403692 , n402425 );
not ( n56500 , n403692 );
or ( n56501 , n56498 , n56500 );
buf ( n403695 , n402422 );
buf ( n403696 , n55163 );
nand ( n56504 , n403695 , n403696 );
buf ( n403698 , n56504 );
buf ( n403699 , n403698 );
nand ( n56507 , n56501 , n403699 );
buf ( n403701 , n56507 );
not ( n56509 , n55142 );
and ( n56510 , n403701 , n56509 );
not ( n56511 , n403701 );
not ( n56512 , n56509 );
and ( n56513 , n56511 , n56512 );
nor ( n56514 , n56510 , n56513 );
not ( n56515 , n56514 );
or ( n56516 , n56496 , n56515 );
buf ( n403710 , n403687 );
not ( n56518 , n403710 );
buf ( n403712 , n56463 );
nand ( n56520 , n56518 , n403712 );
buf ( n403714 , n56520 );
nand ( n56522 , n56516 , n403714 );
buf ( n403716 , n56522 );
not ( n56524 , n403716 );
buf ( n403718 , n402453 );
buf ( n403719 , n402292 );
xor ( n56527 , n403718 , n403719 );
buf ( n403721 , n402321 );
xnor ( n56529 , n56527 , n403721 );
buf ( n403723 , n56529 );
not ( n56531 , n403723 );
buf ( n403725 , n56531 );
not ( n56533 , n403725 );
or ( n56534 , n56524 , n56533 );
buf ( n403728 , n403723 );
not ( n56536 , n403728 );
buf ( n403730 , n56522 );
not ( n56538 , n403730 );
buf ( n403732 , n56538 );
buf ( n403733 , n403732 );
not ( n56541 , n403733 );
or ( n56542 , n56536 , n56541 );
xor ( n56543 , n402147 , n402162 );
xor ( n56544 , n56543 , n402270 );
buf ( n403738 , n56544 );
buf ( n403739 , n395362 );
not ( n56547 , n403739 );
buf ( n403741 , n402314 );
not ( n56549 , n403741 );
or ( n56550 , n56547 , n56549 );
xor ( n56551 , n35991 , n47863 );
xnor ( n56552 , n56551 , n35990 );
buf ( n403746 , n56552 );
buf ( n403747 , n395349 );
nand ( n56555 , n403746 , n403747 );
buf ( n403749 , n56555 );
buf ( n403750 , n403749 );
nand ( n56558 , n56550 , n403750 );
buf ( n403752 , n56558 );
or ( n56560 , n403738 , n403752 );
xor ( n56561 , n402169 , n54911 );
xor ( n56562 , n56561 , n402267 );
buf ( n403756 , n56562 );
not ( n56564 , n403756 );
buf ( n403758 , n56564 );
buf ( n403759 , n403758 );
not ( n56567 , n403759 );
and ( n56568 , n55139 , n402385 );
not ( n56569 , n55139 );
and ( n56570 , n56569 , n402388 );
nor ( n56571 , n56568 , n56570 );
buf ( n403765 , n56571 );
buf ( n403766 , n402354 );
and ( n56574 , n403765 , n403766 );
not ( n56575 , n403765 );
buf ( n403769 , n402357 );
and ( n56577 , n56575 , n403769 );
nor ( n56578 , n56574 , n56577 );
buf ( n403772 , n56578 );
buf ( n403773 , n403772 );
not ( n56581 , n403773 );
buf ( n403775 , n56581 );
buf ( n403776 , n403775 );
not ( n56584 , n403776 );
buf ( n403778 , n56584 );
buf ( n403779 , n403778 );
not ( n56587 , n403779 );
or ( n56588 , n56567 , n56587 );
buf ( n403782 , n56562 );
not ( n56590 , n403782 );
buf ( n403784 , n403775 );
not ( n56592 , n403784 );
or ( n56593 , n56590 , n56592 );
not ( n56594 , n402375 );
buf ( n403788 , n394210 );
not ( n56596 , n403788 );
buf ( n403790 , n42390 );
not ( n56598 , n403790 );
or ( n56599 , n56596 , n56598 );
buf ( n403793 , n37037 );
buf ( n403794 , n394219 );
nand ( n56602 , n403793 , n403794 );
buf ( n403796 , n56602 );
buf ( n403797 , n403796 );
nand ( n56605 , n56599 , n403797 );
buf ( n403799 , n56605 );
not ( n56607 , n403799 );
or ( n56608 , n56594 , n56607 );
not ( n56609 , n402370 );
or ( n56610 , n56609 , n384551 );
nand ( n56611 , n56608 , n56610 );
buf ( n403805 , n56611 );
not ( n56613 , n403805 );
buf ( n403807 , n49117 );
not ( n56615 , n403807 );
buf ( n403809 , n388576 );
not ( n56617 , n403809 );
or ( n56618 , n56615 , n56617 );
buf ( n403812 , n385630 );
buf ( n403813 , n49124 );
nand ( n56621 , n403812 , n403813 );
buf ( n403815 , n56621 );
buf ( n403816 , n403815 );
nand ( n56624 , n56618 , n403816 );
buf ( n403818 , n56624 );
buf ( n56626 , n403818 );
not ( n56627 , n56626 );
not ( n56628 , n391270 );
or ( n56629 , n56627 , n56628 );
nand ( n56630 , n383406 , n402706 );
nand ( n56631 , n56629 , n56630 );
buf ( n403825 , n56631 );
not ( n56633 , n403825 );
or ( n56634 , n56613 , n56633 );
or ( n56635 , n56631 , n56611 );
buf ( n403829 , n389359 );
not ( n56637 , n403829 );
buf ( n403831 , n388272 );
not ( n56639 , n403831 );
or ( n56640 , n56637 , n56639 );
buf ( n403834 , n36250 );
buf ( n403835 , n389356 );
nand ( n56643 , n403834 , n403835 );
buf ( n403837 , n56643 );
buf ( n403838 , n403837 );
nand ( n56646 , n56640 , n403838 );
buf ( n403840 , n56646 );
buf ( n403841 , n403840 );
not ( n56649 , n403841 );
buf ( n403843 , n36317 );
not ( n56651 , n403843 );
or ( n56652 , n56649 , n56651 );
buf ( n403846 , n402654 );
buf ( n403847 , n383904 );
nand ( n56655 , n403846 , n403847 );
buf ( n403849 , n56655 );
buf ( n403850 , n403849 );
nand ( n56658 , n56652 , n403850 );
buf ( n403852 , n56658 );
not ( n56660 , n403852 );
not ( n56661 , n389162 );
not ( n56662 , n55786 );
or ( n56663 , n56661 , n56662 );
buf ( n403857 , n375781 );
not ( n56665 , n403857 );
buf ( n403859 , n24117 );
not ( n56667 , n403859 );
and ( n56668 , n56665 , n56667 );
buf ( n403862 , n375781 );
buf ( n403863 , n24117 );
and ( n56671 , n403862 , n403863 );
nor ( n56672 , n56668 , n56671 );
buf ( n403866 , n56672 );
or ( n56674 , n403866 , n41710 );
nand ( n56675 , n56663 , n56674 );
not ( n56676 , n56675 );
or ( n56677 , n56660 , n56676 );
buf ( n403871 , n403852 );
buf ( n403872 , n56675 );
or ( n56680 , n403871 , n403872 );
xor ( n56681 , n402220 , n54953 );
xor ( n56682 , n56681 , n402259 );
buf ( n403876 , n56682 );
nand ( n56684 , n56680 , n403876 );
buf ( n403878 , n56684 );
nand ( n56686 , n56677 , n403878 );
nand ( n56687 , n56635 , n56686 );
buf ( n403881 , n56687 );
nand ( n56689 , n56634 , n403881 );
buf ( n403883 , n56689 );
buf ( n403884 , n403883 );
nand ( n56692 , n56593 , n403884 );
buf ( n403886 , n56692 );
buf ( n403887 , n403886 );
nand ( n56695 , n56588 , n403887 );
buf ( n403889 , n56695 );
and ( n56697 , n56560 , n403889 );
and ( n56698 , n403738 , n403752 );
nor ( n56699 , n56697 , n56698 );
buf ( n403893 , n56699 );
not ( n56701 , n403893 );
buf ( n403895 , n56701 );
buf ( n403896 , n403895 );
nand ( n56704 , n56542 , n403896 );
buf ( n403898 , n56704 );
buf ( n403899 , n403898 );
nand ( n56707 , n56534 , n403899 );
buf ( n403901 , n56707 );
buf ( n403902 , n403901 );
and ( n56710 , n56415 , n403902 );
and ( n56711 , n403619 , n403623 );
or ( n56712 , n56710 , n56711 );
buf ( n403906 , n56712 );
buf ( n403907 , n403906 );
not ( n56715 , n403907 );
buf ( n403909 , n56715 );
buf ( n403910 , n403909 );
not ( n56718 , n403910 );
xor ( n56719 , n402289 , n402564 );
xor ( n56720 , n56719 , n402569 );
buf ( n403914 , n56720 );
not ( n56722 , n403914 );
buf ( n403916 , n56722 );
not ( n56724 , n403916 );
or ( n56725 , n56718 , n56724 );
buf ( n403919 , n402557 );
buf ( n403920 , n402459 );
xor ( n56728 , n403919 , n403920 );
buf ( n403922 , n56728 );
buf ( n56730 , n402464 );
not ( n56731 , n56730 );
and ( n56732 , n403922 , n56731 );
not ( n56733 , n403922 );
and ( n56734 , n56733 , n56730 );
nor ( n56735 , n56732 , n56734 );
not ( n56736 , n56735 );
not ( n56737 , n56736 );
not ( n56738 , n402483 );
not ( n56739 , n55213 );
or ( n56740 , n56738 , n56739 );
nand ( n56741 , n55212 , n55205 );
nand ( n56742 , n56740 , n56741 );
and ( n56743 , n56742 , n55311 );
not ( n56744 , n56742 );
buf ( n403938 , n55311 );
not ( n56746 , n403938 );
buf ( n403940 , n56746 );
and ( n56748 , n56744 , n403940 );
nor ( n56749 , n56743 , n56748 );
buf ( n56750 , n56749 );
not ( n56751 , n56750 );
xor ( n56752 , n402609 , n402732 );
buf ( n403946 , n56752 );
buf ( n403947 , n403946 );
buf ( n403948 , n402741 );
and ( n56756 , n403947 , n403948 );
not ( n56757 , n403947 );
buf ( n403951 , n402738 );
and ( n56759 , n56757 , n403951 );
nor ( n56760 , n56756 , n56759 );
buf ( n403954 , n56760 );
buf ( n403955 , n403954 );
not ( n56763 , n403955 );
buf ( n403957 , n56763 );
not ( n56765 , n403957 );
xor ( n56766 , n402518 , n402542 );
xor ( n56767 , n56766 , n55305 );
not ( n56768 , n56767 );
not ( n56769 , n395349 );
buf ( n403963 , n395315 );
buf ( n403964 , n36067 );
and ( n56772 , n403963 , n403964 );
not ( n56773 , n403963 );
buf ( n403967 , n36066 );
and ( n56775 , n56773 , n403967 );
nor ( n56776 , n56772 , n56775 );
buf ( n403970 , n56776 );
not ( n56778 , n403970 );
or ( n56779 , n56769 , n56778 );
buf ( n403973 , n56552 );
buf ( n403974 , n395362 );
nand ( n56782 , n403973 , n403974 );
buf ( n403976 , n56782 );
nand ( n56784 , n56779 , n403976 );
not ( n56785 , n56784 );
nand ( n56803 , n56785 , C1 );
not ( n56804 , n56803 );
or ( n56805 , n56768 , n56804 );
nand ( n56808 , n56805 , C1 );
not ( n56809 , n56808 );
or ( n56810 , n56765 , n56809 );
buf ( n403985 , n56808 );
not ( n56812 , n403985 );
buf ( n403987 , n56812 );
not ( n56814 , n403987 );
not ( n56815 , n403954 );
or ( n56816 , n56814 , n56815 );
not ( n56817 , n388760 );
not ( n56818 , n41904 );
or ( n56819 , n56817 , n56818 );
buf ( n403994 , n37763 );
buf ( n403995 , n388757 );
nand ( n56822 , n403994 , n403995 );
buf ( n403997 , n56822 );
nand ( n56824 , n56819 , n403997 );
buf ( n403999 , n56824 );
not ( n56826 , n403999 );
buf ( n404001 , n56826 );
buf ( n404002 , n404001 );
not ( n56829 , n404002 );
buf ( n404004 , n388743 );
not ( n56831 , n404004 );
and ( n56832 , n56829 , n56831 );
buf ( n404007 , n402689 );
buf ( n404008 , n388809 );
and ( n56835 , n404007 , n404008 );
nor ( n56836 , n56832 , n56835 );
buf ( n404011 , n56836 );
buf ( n404012 , n382938 );
buf ( n404013 , n358975 );
nand ( n56840 , n404012 , n404013 );
buf ( n404015 , n56840 );
buf ( n56842 , n46531 );
not ( n56843 , n56842 );
buf ( n404018 , n391443 );
buf ( n404019 , n36395 );
and ( n56846 , n404018 , n404019 );
not ( n56847 , n404018 );
buf ( n404022 , n50992 );
and ( n56849 , n56847 , n404022 );
or ( n56850 , n56846 , n56849 );
buf ( n404025 , n56850 );
nor ( n56852 , n56843 , n404025 );
nand ( n56853 , n56852 , n388349 );
not ( n56854 , n383937 );
nand ( n56855 , n56854 , n55706 );
nand ( n56856 , n404015 , n56853 , n56855 );
buf ( n404031 , n388230 );
not ( n56858 , n404031 );
buf ( n404033 , n51648 );
not ( n56860 , n404033 );
or ( n56861 , n56858 , n56860 );
buf ( n404036 , n22982 );
buf ( n404037 , n388227 );
nand ( n56864 , n404036 , n404037 );
buf ( n404039 , n56864 );
buf ( n404040 , n404039 );
nand ( n56867 , n56861 , n404040 );
buf ( n404042 , n56867 );
buf ( n404043 , n404042 );
not ( n56870 , n404043 );
buf ( n404045 , n399031 );
not ( n56872 , n404045 );
or ( n56873 , n56870 , n56872 );
buf ( n404048 , n402247 );
buf ( n404049 , n386477 );
nand ( n56876 , n404048 , n404049 );
buf ( n404051 , n56876 );
buf ( n404052 , n404051 );
nand ( n56879 , n56873 , n404052 );
buf ( n404054 , n56879 );
not ( n56881 , n404054 );
buf ( n404056 , n388502 );
not ( n56883 , n404056 );
buf ( n404058 , n393525 );
not ( n56885 , n404058 );
or ( n56886 , n56883 , n56885 );
buf ( n404061 , n385473 );
buf ( n404062 , n388511 );
nand ( n56889 , n404061 , n404062 );
buf ( n404064 , n56889 );
buf ( n404065 , n404064 );
nand ( n56892 , n56886 , n404065 );
buf ( n404067 , n56892 );
buf ( n404068 , n404067 );
not ( n56895 , n404068 );
buf ( n404070 , n393544 );
not ( n56897 , n404070 );
or ( n56898 , n56895 , n56897 );
buf ( n404073 , n46061 );
not ( n56900 , n404073 );
buf ( n404075 , n402868 );
nand ( n56902 , n56900 , n404075 );
buf ( n404077 , n56902 );
buf ( n404078 , n404077 );
nand ( n56905 , n56898 , n404078 );
buf ( n404080 , n56905 );
not ( n56907 , n404080 );
or ( n56908 , n56881 , n56907 );
or ( n56909 , n404080 , n404054 );
buf ( n404084 , n54951 );
buf ( n404085 , n392788 );
and ( n56912 , n404084 , n404085 );
buf ( n404087 , n53252 );
not ( n56914 , n404087 );
buf ( n404089 , n389856 );
not ( n56916 , n404089 );
or ( n56917 , n56914 , n56916 );
buf ( n404092 , n49686 );
not ( n56919 , n41559 );
buf ( n404094 , n56919 );
nand ( n56921 , n404092 , n404094 );
buf ( n404096 , n56921 );
buf ( n404097 , n404096 );
nand ( n56924 , n56917 , n404097 );
buf ( n404099 , n56924 );
buf ( n404100 , n404099 );
buf ( n404101 , n390432 );
and ( n56928 , n404100 , n404101 );
buf ( n404103 , n56928 );
buf ( n404104 , n404103 );
nor ( n56931 , n56912 , n404104 );
buf ( n404106 , n56931 );
buf ( n404107 , n404106 );
not ( n56934 , n404107 );
buf ( n404109 , n56934 );
nand ( n56936 , n56909 , n404109 );
nand ( n56937 , n56908 , n56936 );
nand ( n56938 , n56856 , n56937 );
not ( n56939 , n388349 );
not ( n56940 , n56852 );
or ( n56941 , n56939 , n56940 );
nand ( n56942 , n56941 , n56855 );
not ( n56943 , n404015 );
nand ( n56944 , n56942 , n56943 );
nand ( n56945 , n404011 , n56938 , n56944 );
not ( n56946 , n56945 );
xor ( n56947 , n402201 , n402213 );
xor ( n56948 , n56947 , n402263 );
buf ( n404123 , n56948 );
not ( n56950 , n404123 );
or ( n56951 , n56946 , n56950 );
not ( n56952 , n404011 );
nand ( n56953 , n56938 , n56944 );
nand ( n56954 , n56952 , n56953 );
nand ( n56955 , n56951 , n56954 );
buf ( n404130 , n56955 );
buf ( n404131 , n45260 );
not ( n56958 , n404131 );
buf ( n404133 , n392247 );
not ( n56960 , n404133 );
buf ( n404135 , n398723 );
not ( n56962 , n404135 );
or ( n56963 , n56960 , n56962 );
buf ( n404138 , n49525 );
buf ( n404139 , n392244 );
nand ( n56966 , n404138 , n404139 );
buf ( n404141 , n56966 );
buf ( n404142 , n404141 );
nand ( n56969 , n56963 , n404142 );
buf ( n404144 , n56969 );
buf ( n404145 , n404144 );
not ( n56972 , n404145 );
or ( n56973 , n56958 , n56972 );
buf ( n404148 , n55361 );
buf ( n404149 , n392740 );
nand ( n56976 , n404148 , n404149 );
buf ( n404151 , n56976 );
buf ( n404152 , n404151 );
nand ( n56979 , n56973 , n404152 );
buf ( n404154 , n56979 );
buf ( n404155 , n404154 );
xor ( n56982 , n404130 , n404155 );
buf ( n404157 , n400033 );
not ( n56984 , n404157 );
buf ( n404159 , n40714 );
not ( n56986 , n404159 );
or ( n56987 , n56984 , n56986 );
buf ( n404162 , n40711 );
buf ( n404163 , n400042 );
nand ( n56990 , n404162 , n404163 );
buf ( n404165 , n56990 );
buf ( n404166 , n404165 );
nand ( n56993 , n56987 , n404166 );
buf ( n404168 , n56993 );
buf ( n404169 , n404168 );
not ( n56996 , n404169 );
buf ( n404171 , n38765 );
not ( n56998 , n404171 );
or ( n56999 , n56996 , n56998 );
buf ( n404174 , n390635 );
buf ( n404175 , n402530 );
nand ( n57002 , n404174 , n404175 );
buf ( n404177 , n57002 );
buf ( n404178 , n404177 );
nand ( n57005 , n56999 , n404178 );
buf ( n404180 , n57005 );
buf ( n404181 , n404180 );
xor ( n57008 , n402627 , n402641 );
xor ( n57009 , n57008 , n402667 );
buf ( n404184 , n57009 );
buf ( n404185 , n404184 );
xor ( n57012 , n404181 , n404185 );
not ( n57013 , n388746 );
buf ( n404188 , n388760 );
not ( n57015 , n404188 );
buf ( n404190 , n388979 );
not ( n57017 , n404190 );
or ( n57018 , n57015 , n57017 );
buf ( n404193 , n385342 );
buf ( n404194 , n388757 );
nand ( n57021 , n404193 , n404194 );
buf ( n404196 , n57021 );
buf ( n404197 , n404196 );
nand ( n57024 , n57018 , n404197 );
buf ( n404199 , n57024 );
not ( n57026 , n404199 );
or ( n57027 , n57013 , n57026 );
nand ( n57028 , n56824 , n388809 );
nand ( n57029 , n57027 , n57028 );
buf ( n404204 , n392884 );
not ( n57031 , n404204 );
buf ( n404206 , n40886 );
not ( n57033 , n404206 );
or ( n57034 , n57031 , n57033 );
buf ( n404209 , n40885 );
buf ( n404210 , n392887 );
nand ( n57037 , n404209 , n404210 );
buf ( n404212 , n57037 );
buf ( n404213 , n404212 );
nand ( n57040 , n57034 , n404213 );
buf ( n404215 , n57040 );
not ( n57042 , n404215 );
not ( n57043 , n36801 );
or ( n57044 , n57042 , n57043 );
buf ( n404219 , n388669 );
buf ( n404220 , n402922 );
nand ( n57047 , n404219 , n404220 );
buf ( n404222 , n57047 );
nand ( n57049 , n57044 , n404222 );
or ( n57050 , n57029 , n57049 );
buf ( n404225 , n399274 );
not ( n57052 , n404225 );
buf ( n404227 , n389753 );
not ( n57054 , n404227 );
or ( n57055 , n57052 , n57054 );
buf ( n404230 , n31964 );
buf ( n404231 , n399283 );
nand ( n57058 , n404230 , n404231 );
buf ( n404233 , n57058 );
buf ( n404234 , n404233 );
nand ( n57061 , n57055 , n404234 );
buf ( n404236 , n57061 );
buf ( n404237 , n404236 );
not ( n57064 , n404237 );
buf ( n404239 , n398431 );
not ( n57066 , n404239 );
or ( n57067 , n57064 , n57066 );
buf ( n404242 , n389024 );
buf ( n404243 , n402795 );
nand ( n57070 , n404242 , n404243 );
buf ( n404245 , n57070 );
buf ( n404246 , n404245 );
nand ( n57073 , n57067 , n404246 );
buf ( n404248 , n57073 );
nand ( n57075 , n57050 , n404248 );
buf ( n404250 , n57075 );
nand ( n57077 , n57029 , n57049 );
buf ( n404252 , n57077 );
nand ( n57079 , n404250 , n404252 );
buf ( n404254 , n57079 );
buf ( n404255 , n404254 );
and ( n57082 , n57012 , n404255 );
and ( n57083 , n404181 , n404185 );
or ( n57084 , n57082 , n57083 );
buf ( n404259 , n57084 );
buf ( n404260 , n404259 );
and ( n57087 , n56982 , n404260 );
and ( n57088 , n404130 , n404155 );
or ( n57089 , n57087 , n57088 );
buf ( n404264 , n57089 );
nand ( n57091 , n56816 , n404264 );
nand ( n57092 , n56810 , n57091 );
not ( n57093 , n57092 );
or ( n57094 , n56751 , n57093 );
buf ( n404269 , n57092 );
not ( n57096 , n404269 );
buf ( n404271 , n57096 );
not ( n57098 , n404271 );
not ( n57099 , n56750 );
not ( n57100 , n57099 );
or ( n57101 , n57098 , n57100 );
xor ( n57102 , n402498 , n55274 );
xor ( n57103 , n57102 , n55308 );
buf ( n404278 , n57103 );
xor ( n57105 , n403543 , n403556 );
xor ( n57106 , n57105 , n403585 );
buf ( n404281 , n57106 );
buf ( n404282 , n404281 );
xor ( n57109 , n404278 , n404282 );
buf ( n404284 , n50579 );
not ( n57111 , n404284 );
buf ( n404286 , n47891 );
not ( n57113 , n404286 );
buf ( n404288 , n386391 );
not ( n57115 , n404288 );
or ( n57116 , n57113 , n57115 );
buf ( n404291 , n35301 );
buf ( n404292 , n50584 );
nand ( n57119 , n404291 , n404292 );
buf ( n404294 , n57119 );
buf ( n404295 , n404294 );
nand ( n57122 , n57116 , n404295 );
buf ( n404297 , n57122 );
buf ( n404298 , n404297 );
not ( n57125 , n404298 );
or ( n57126 , n57111 , n57125 );
buf ( n404301 , n403674 );
buf ( n404302 , n51553 );
nand ( n57129 , n404301 , n404302 );
buf ( n404304 , n57129 );
buf ( n404305 , n404304 );
nand ( n57132 , n57126 , n404305 );
buf ( n404307 , n57132 );
buf ( n404308 , n389692 );
not ( n57135 , n404308 );
buf ( n404310 , n391024 );
not ( n57137 , n404310 );
and ( n57138 , n57135 , n57137 );
buf ( n404313 , n38472 );
buf ( n404314 , n391024 );
and ( n57141 , n404313 , n404314 );
nor ( n57142 , n57138 , n57141 );
buf ( n404317 , n57142 );
not ( n57144 , n404317 );
not ( n57145 , n43537 );
and ( n57146 , n57144 , n57145 );
and ( n57147 , n403440 , n43515 );
nor ( n57148 , n57146 , n57147 );
not ( n57149 , n57148 );
not ( n57150 , n57149 );
buf ( n404325 , n402770 );
not ( n57152 , n404325 );
buf ( n404327 , n57152 );
buf ( n404328 , n404327 );
buf ( n404329 , n390362 );
and ( n57156 , n404328 , n404329 );
buf ( n404331 , n388102 );
not ( n57158 , n404331 );
buf ( n404333 , n384083 );
not ( n57160 , n404333 );
or ( n57161 , n57158 , n57160 );
buf ( n404336 , n390657 );
buf ( n404337 , n388105 );
nand ( n57164 , n404336 , n404337 );
buf ( n404339 , n57164 );
buf ( n404340 , n404339 );
nand ( n57167 , n57161 , n404340 );
buf ( n404342 , n57167 );
buf ( n404343 , n404342 );
not ( n57170 , n404343 );
buf ( n404345 , n388093 );
nor ( n57172 , n57170 , n404345 );
buf ( n404347 , n57172 );
buf ( n404348 , n404347 );
nor ( n57175 , n57156 , n404348 );
buf ( n404350 , n57175 );
buf ( n404351 , n404350 );
not ( n57178 , n404351 );
buf ( n404353 , n57178 );
not ( n57180 , n404353 );
or ( n57181 , n57150 , n57180 );
not ( n57182 , n404350 );
not ( n57183 , n57148 );
or ( n57184 , n57182 , n57183 );
and ( n57185 , n402948 , n402981 );
not ( n57186 , n402948 );
and ( n57187 , n57186 , n402978 );
or ( n57188 , n57185 , n57187 );
buf ( n57189 , n402931 );
and ( n57190 , n57188 , n57189 );
not ( n57191 , n57188 );
not ( n57192 , n57189 );
and ( n57193 , n57191 , n57192 );
nor ( n57194 , n57190 , n57193 );
nand ( n57195 , n57184 , n57194 );
nand ( n57196 , n57181 , n57195 );
or ( n57197 , n404307 , n57196 );
xor ( n57198 , n403426 , n403463 );
xor ( n57199 , n57198 , n403471 );
buf ( n404374 , n57199 );
nand ( n57201 , n57197 , n404374 );
buf ( n404376 , n57201 );
nand ( n57203 , n57196 , n404307 );
buf ( n404378 , n57203 );
nand ( n57205 , n404376 , n404378 );
buf ( n404380 , n57205 );
buf ( n404381 , n404380 );
and ( n57208 , n57109 , n404381 );
and ( n57209 , n404278 , n404282 );
or ( n57210 , n57208 , n57209 );
buf ( n404385 , n57210 );
buf ( n57212 , n404385 );
nand ( n57213 , n57101 , n57212 );
nand ( n57214 , n57094 , n57213 );
not ( n57215 , n57214 );
or ( n57216 , n56737 , n57215 );
or ( n57217 , n57214 , n56736 );
xor ( n57218 , n402593 , n403485 );
xor ( n57219 , n57218 , n403491 );
nand ( n57220 , n57217 , n57219 );
nand ( n57221 , n57216 , n57220 );
buf ( n404396 , n57221 );
nand ( n57223 , n56725 , n404396 );
buf ( n404398 , n57223 );
buf ( n404399 , n404398 );
buf ( n404400 , n403914 );
buf ( n404401 , n403906 );
nand ( n57228 , n404400 , n404401 );
buf ( n404403 , n57228 );
buf ( n404404 , n404403 );
and ( n57231 , n404399 , n404404 );
buf ( n404406 , n57231 );
buf ( n404407 , n404406 );
xor ( n57234 , n403541 , n404407 );
buf ( n404409 , n402573 );
not ( n57236 , n404409 );
buf ( n404411 , n402584 );
not ( n57238 , n404411 );
or ( n57239 , n57236 , n57238 );
buf ( n404414 , n402097 );
buf ( n404415 , n402579 );
nand ( n57242 , n404414 , n404415 );
buf ( n404417 , n57242 );
buf ( n404418 , n404417 );
nand ( n57245 , n57239 , n404418 );
buf ( n404420 , n57245 );
buf ( n404421 , n404420 );
buf ( n404422 , n56273 );
not ( n57249 , n404422 );
buf ( n404424 , n57249 );
buf ( n404425 , n404424 );
and ( n57252 , n404421 , n404425 );
not ( n57253 , n404421 );
buf ( n404428 , n56273 );
and ( n57255 , n57253 , n404428 );
nor ( n57256 , n57252 , n57255 );
buf ( n404431 , n57256 );
buf ( n404432 , n404431 );
and ( n57259 , n57234 , n404432 );
and ( n57260 , n403541 , n404407 );
or ( n57261 , n57259 , n57260 );
buf ( n404436 , n57261 );
not ( n57263 , n404436 );
xor ( n57264 , n402094 , n403513 );
xor ( n57265 , n57264 , n403518 );
buf ( n404440 , n57265 );
not ( n57267 , n404440 );
or ( n57268 , n57263 , n57267 );
xor ( n57269 , n403541 , n404407 );
xor ( n57270 , n57269 , n404432 );
buf ( n404445 , n57270 );
buf ( n404446 , n404445 );
xor ( n57273 , n402751 , n402755 );
xor ( n57274 , n57273 , n403481 );
buf ( n404449 , n57274 );
buf ( n404450 , n404449 );
xor ( n57277 , n403589 , n403607 );
xor ( n57278 , n57277 , n403614 );
buf ( n404453 , n57278 );
buf ( n404454 , n404453 );
xor ( n57281 , n404450 , n404454 );
buf ( n404456 , n403738 );
buf ( n404457 , n403752 );
xor ( n57284 , n404456 , n404457 );
buf ( n404459 , n403889 );
xor ( n57286 , n57284 , n404459 );
buf ( n404461 , n57286 );
not ( n57288 , n404461 );
xor ( n57289 , n402760 , n402999 );
xor ( n57290 , n57289 , n403476 );
buf ( n404465 , n57290 );
not ( n57292 , n404465 );
or ( n57293 , n57288 , n57292 );
or ( n57294 , n404465 , n404461 );
xor ( n57295 , n402905 , n402807 );
xnor ( n57296 , n57295 , n55591 );
buf ( n404471 , n57296 );
not ( n57298 , n404471 );
buf ( n404473 , n403026 );
not ( n57300 , n404473 );
buf ( n404475 , n403418 );
not ( n57302 , n404475 );
or ( n57303 , n57300 , n57302 );
buf ( n404478 , n403006 );
buf ( n404479 , n403023 );
nand ( n57306 , n404478 , n404479 );
buf ( n404481 , n57306 );
buf ( n404482 , n404481 );
nand ( n57309 , n57303 , n404482 );
buf ( n404484 , n57309 );
buf ( n404485 , n404484 );
buf ( n404486 , n403412 );
not ( n57313 , n404486 );
buf ( n404488 , n57313 );
buf ( n404489 , n404488 );
and ( n57316 , n404485 , n404489 );
not ( n57317 , n404485 );
buf ( n404492 , n403412 );
and ( n57319 , n57317 , n404492 );
nor ( n57320 , n57316 , n57319 );
buf ( n404495 , n57320 );
buf ( n404496 , n404495 );
not ( n57323 , n404496 );
buf ( n404498 , n57323 );
buf ( n404499 , n404498 );
not ( n57326 , n404499 );
or ( n57327 , n57298 , n57326 );
not ( n57328 , n57296 );
nand ( n57329 , n57328 , n404495 );
buf ( n404504 , n394817 );
not ( n57331 , n404504 );
buf ( n404506 , n42390 );
not ( n57333 , n404506 );
or ( n57334 , n57331 , n57333 );
buf ( n404509 , n391870 );
buf ( n404510 , n394814 );
nand ( n57337 , n404509 , n404510 );
buf ( n404512 , n57337 );
buf ( n404513 , n404512 );
nand ( n57340 , n57334 , n404513 );
buf ( n404515 , n57340 );
buf ( n404516 , n404515 );
not ( n57343 , n404516 );
buf ( n404518 , n389880 );
not ( n57345 , n404518 );
or ( n57346 , n57343 , n57345 );
buf ( n404521 , n403799 );
buf ( n404522 , n391638 );
nand ( n57349 , n404521 , n404522 );
buf ( n404524 , n57349 );
buf ( n404525 , n404524 );
nand ( n57352 , n57346 , n404525 );
buf ( n404527 , n57352 );
buf ( n404528 , n404527 );
xor ( n57355 , n403363 , n403388 );
xor ( n57356 , n57355 , n403408 );
buf ( n404531 , n57356 );
buf ( n404532 , n404531 );
xor ( n57359 , n404528 , n404532 );
buf ( n404534 , n43286 );
not ( n57361 , n404534 );
buf ( n404536 , n388102 );
not ( n57363 , n404536 );
buf ( n404538 , n41896 );
not ( n57365 , n404538 );
or ( n57366 , n57363 , n57365 );
buf ( n404541 , n36564 );
buf ( n404542 , n388105 );
nand ( n57369 , n404541 , n404542 );
buf ( n404544 , n57369 );
buf ( n404545 , n404544 );
nand ( n57372 , n57366 , n404545 );
buf ( n404547 , n57372 );
buf ( n404548 , n404547 );
not ( n57375 , n404548 );
or ( n57376 , n57361 , n57375 );
buf ( n404551 , n404342 );
buf ( n404552 , n388068 );
nand ( n57379 , n404551 , n404552 );
buf ( n404554 , n57379 );
buf ( n404555 , n404554 );
nand ( n57382 , n57376 , n404555 );
buf ( n404557 , n57382 );
buf ( n404558 , n404557 );
and ( n57385 , n57359 , n404558 );
and ( n57386 , n404528 , n404532 );
or ( n57387 , n57385 , n57386 );
buf ( n404562 , n57387 );
nand ( n57389 , n57329 , n404562 );
buf ( n404564 , n57389 );
nand ( n57391 , n57327 , n404564 );
buf ( n404566 , n57391 );
not ( n57393 , n404566 );
or ( n57394 , n402780 , n55753 );
nand ( n57395 , n55753 , n402780 );
nand ( n57396 , n57394 , n57395 );
buf ( n57397 , n55677 );
and ( n57398 , n57396 , n57397 );
not ( n57399 , n57396 );
and ( n57400 , n57399 , n402992 );
nor ( n57401 , n57398 , n57400 );
buf ( n404576 , n57401 );
not ( n57403 , n404576 );
buf ( n404578 , n57403 );
not ( n57405 , n404578 );
or ( n57406 , n57393 , n57405 );
buf ( n404581 , n404566 );
not ( n57408 , n404581 );
buf ( n404583 , n57408 );
not ( n57410 , n404583 );
not ( n57411 , n57401 );
or ( n57412 , n57410 , n57411 );
xor ( n57413 , n402856 , n402882 );
xor ( n57414 , n57413 , n402901 );
buf ( n404589 , n57414 );
not ( n57416 , n404589 );
buf ( n404591 , n47726 );
not ( n57418 , n404591 );
buf ( n404593 , n55660 );
not ( n57420 , n404593 );
or ( n57421 , n57418 , n57420 );
nand ( n57422 , n394884 , n388367 );
not ( n57423 , n57422 );
buf ( n404598 , n397069 );
buf ( n404599 , n388192 );
not ( n57426 , n404599 );
buf ( n404601 , n57426 );
buf ( n404602 , n404601 );
nand ( n57429 , n404598 , n404602 );
buf ( n404604 , n57429 );
not ( n57431 , n404604 );
or ( n57432 , n57423 , n57431 );
nand ( n57433 , n57432 , n397476 );
buf ( n404608 , n57433 );
nand ( n57435 , n57421 , n404608 );
buf ( n404610 , n57435 );
buf ( n404611 , n404610 );
not ( n57438 , n404611 );
buf ( n404613 , n42073 );
not ( n57440 , n404613 );
buf ( n404615 , n390548 );
not ( n57442 , n404615 );
or ( n57443 , n57440 , n57442 );
buf ( n404618 , n388905 );
buf ( n404619 , n42074 );
nand ( n57446 , n404618 , n404619 );
buf ( n404621 , n57446 );
buf ( n404622 , n404621 );
nand ( n57449 , n57443 , n404622 );
buf ( n404624 , n57449 );
not ( n57451 , n404624 );
not ( n57452 , n45662 );
or ( n57453 , n57451 , n57452 );
buf ( n404628 , n403401 );
buf ( n404629 , n37314 );
nand ( n57456 , n404628 , n404629 );
buf ( n404631 , n57456 );
nand ( n57458 , n57453 , n404631 );
buf ( n404633 , n57458 );
not ( n57460 , n404633 );
or ( n57461 , n57438 , n57460 );
buf ( n404636 , n57458 );
buf ( n404637 , n404610 );
or ( n57464 , n404636 , n404637 );
buf ( n404639 , n388833 );
not ( n57466 , n404639 );
buf ( n404641 , n403377 );
not ( n57468 , n404641 );
or ( n57469 , n57466 , n57468 );
not ( n57470 , n41342 );
not ( n57471 , n50317 );
or ( n57472 , n57470 , n57471 );
buf ( n404647 , n40818 );
buf ( n404648 , n45897 );
nand ( n57475 , n404647 , n404648 );
buf ( n404650 , n57475 );
nand ( n57477 , n57472 , n404650 );
buf ( n404652 , n57477 );
buf ( n404653 , n388872 );
nand ( n57480 , n404652 , n404653 );
buf ( n404655 , n57480 );
buf ( n404656 , n404655 );
nand ( n57483 , n57469 , n404656 );
buf ( n404658 , n57483 );
buf ( n404659 , n404658 );
nand ( n57486 , n57464 , n404659 );
buf ( n404661 , n57486 );
buf ( n404662 , n404661 );
nand ( n57489 , n57461 , n404662 );
buf ( n404664 , n57489 );
not ( n57491 , n404664 );
nand ( n57492 , n57416 , n57491 );
not ( n57493 , n57492 );
xor ( n57494 , n403175 , n403182 );
xor ( n57495 , n57494 , n403346 );
buf ( n404670 , n57495 );
buf ( n404671 , n404670 );
buf ( n404672 , n42924 );
not ( n57499 , n404672 );
buf ( n404674 , n404099 );
not ( n57501 , n404674 );
or ( n57502 , n57499 , n57501 );
and ( n57503 , n27258 , n24071 );
not ( n57504 , n27258 );
buf ( n57505 , n24070 );
and ( n57506 , n57504 , n57505 );
or ( n57507 , n57503 , n57506 );
buf ( n404682 , n57507 );
buf ( n404683 , n390429 );
nand ( n57510 , n404682 , n404683 );
buf ( n404685 , n57510 );
buf ( n404686 , n404685 );
nand ( n57513 , n57502 , n404686 );
buf ( n404688 , n57513 );
buf ( n404689 , n404688 );
xor ( n57516 , n404671 , n404689 );
buf ( n404691 , n388998 );
not ( n57518 , n404691 );
buf ( n404693 , n46906 );
not ( n57520 , n404693 );
or ( n57521 , n57518 , n57520 );
buf ( n404696 , n22982 );
buf ( n404697 , n388215 );
nand ( n57524 , n404696 , n404697 );
buf ( n404699 , n57524 );
buf ( n404700 , n404699 );
nand ( n57527 , n57521 , n404700 );
buf ( n404702 , n57527 );
buf ( n404703 , n404702 );
not ( n57530 , n404703 );
buf ( n404705 , n38961 );
not ( n57532 , n404705 );
or ( n57533 , n57530 , n57532 );
buf ( n404708 , n404042 );
buf ( n404709 , n393127 );
nand ( n57536 , n404708 , n404709 );
buf ( n404711 , n57536 );
buf ( n404712 , n404711 );
nand ( n57539 , n57533 , n404712 );
buf ( n404714 , n57539 );
buf ( n404715 , n404714 );
and ( n57542 , n57516 , n404715 );
and ( n57543 , n404671 , n404689 );
or ( n57544 , n57542 , n57543 );
buf ( n404719 , n57544 );
buf ( n404720 , n404719 );
not ( n57547 , n404720 );
buf ( n404722 , n389162 );
not ( n57549 , n404722 );
buf ( n404724 , n403866 );
not ( n57551 , n404724 );
buf ( n404726 , n57551 );
buf ( n404727 , n404726 );
not ( n57554 , n404727 );
or ( n57555 , n57549 , n57554 );
buf ( n404730 , n24118 );
not ( n57557 , n404730 );
buf ( n404732 , n40777 );
not ( n57559 , n404732 );
or ( n57560 , n57557 , n57559 );
buf ( n404735 , n40758 );
buf ( n404736 , n24117 );
nand ( n57563 , n404735 , n404736 );
buf ( n404738 , n57563 );
buf ( n404739 , n404738 );
nand ( n57566 , n57560 , n404739 );
buf ( n404741 , n57566 );
buf ( n404742 , n404741 );
buf ( n57569 , n45076 );
buf ( n404744 , n57569 );
nand ( n57571 , n404742 , n404744 );
buf ( n404746 , n57571 );
buf ( n404747 , n404746 );
nand ( n57574 , n57555 , n404747 );
buf ( n404749 , n57574 );
buf ( n404750 , n404749 );
not ( n57577 , n404750 );
or ( n57578 , n57547 , n57577 );
buf ( n404753 , n404749 );
buf ( n404754 , n404719 );
or ( n57581 , n404753 , n404754 );
buf ( n404756 , n403055 );
not ( n57583 , n404756 );
buf ( n404758 , n396622 );
not ( n57585 , n404758 );
or ( n57586 , n57583 , n57585 );
buf ( n404761 , n403065 );
nand ( n57588 , n57586 , n404761 );
buf ( n404763 , n57588 );
buf ( n404764 , n404763 );
not ( n57591 , n404764 );
buf ( n404766 , n403350 );
not ( n57593 , n404766 );
buf ( n404768 , n403034 );
not ( n57595 , n404768 );
and ( n57596 , n57593 , n57595 );
buf ( n404771 , n403350 );
buf ( n404772 , n403034 );
and ( n57599 , n404771 , n404772 );
nor ( n57600 , n57596 , n57599 );
buf ( n404775 , n57600 );
buf ( n404776 , n404775 );
not ( n57603 , n404776 );
and ( n57604 , n57591 , n57603 );
buf ( n404779 , n404763 );
buf ( n404780 , n404775 );
and ( n57607 , n404779 , n404780 );
nor ( n57608 , n57604 , n57607 );
buf ( n404783 , n57608 );
buf ( n404784 , n404783 );
not ( n57611 , n404784 );
buf ( n404786 , n57611 );
buf ( n404787 , n404786 );
nand ( n57614 , n57581 , n404787 );
buf ( n404789 , n57614 );
buf ( n404790 , n404789 );
nand ( n57617 , n57578 , n404790 );
buf ( n404792 , n57617 );
not ( n57619 , n404792 );
or ( n57620 , n57493 , n57619 );
nand ( n57621 , n404664 , n404589 );
nand ( n57622 , n57620 , n57621 );
buf ( n404797 , n57622 );
buf ( n404798 , n45954 );
not ( n57625 , n404798 );
buf ( n404800 , n403639 );
not ( n57627 , n404800 );
or ( n57628 , n57625 , n57627 );
and ( n57629 , n393381 , n384741 );
not ( n57630 , n393381 );
and ( n57631 , n57630 , n389525 );
nor ( n57632 , n57629 , n57631 );
buf ( n404807 , n57632 );
not ( n57634 , n404807 );
buf ( n404809 , n393825 );
nand ( n57636 , n57634 , n404809 );
buf ( n404811 , n57636 );
buf ( n404812 , n404811 );
nand ( n57639 , n57628 , n404812 );
buf ( n404814 , n57639 );
buf ( n404815 , n404814 );
xor ( n57642 , n404797 , n404815 );
buf ( n404817 , n397498 );
not ( n57644 , n404817 );
buf ( n404819 , n395919 );
not ( n57646 , n404819 );
or ( n57647 , n57644 , n57646 );
buf ( n404822 , n385630 );
buf ( n404823 , n397495 );
nand ( n57650 , n404822 , n404823 );
buf ( n404825 , n57650 );
buf ( n404826 , n404825 );
nand ( n57653 , n57647 , n404826 );
buf ( n404828 , n57653 );
not ( n57655 , n404828 );
not ( n57656 , n391649 );
or ( n57657 , n57655 , n57656 );
buf ( n404832 , n403818 );
buf ( n404833 , n391170 );
nand ( n57660 , n404832 , n404833 );
buf ( n404835 , n57660 );
nand ( n57662 , n57657 , n404835 );
not ( n57663 , n57662 );
xor ( n57664 , n403852 , n56675 );
xnor ( n57665 , n57664 , n56682 );
not ( n57666 , n57665 );
not ( n57667 , n57666 );
or ( n57668 , n57663 , n57667 );
not ( n57669 , n57662 );
not ( n57670 , n57669 );
not ( n57671 , n57665 );
or ( n57672 , n57670 , n57671 );
buf ( n404847 , n55055 );
not ( n57674 , n404847 );
buf ( n404849 , n40714 );
not ( n57676 , n404849 );
or ( n57677 , n57674 , n57676 );
buf ( n404852 , n35435 );
buf ( n404853 , n55055 );
not ( n57680 , n404853 );
buf ( n404855 , n57680 );
buf ( n404856 , n404855 );
nand ( n57683 , n404852 , n404856 );
buf ( n404858 , n57683 );
buf ( n404859 , n404858 );
nand ( n57686 , n57677 , n404859 );
buf ( n404861 , n57686 );
buf ( n404862 , n404861 );
not ( n57689 , n404862 );
buf ( n404864 , n386300 );
not ( n57691 , n404864 );
or ( n57692 , n57689 , n57691 );
buf ( n404867 , n383137 );
buf ( n404868 , n404168 );
nand ( n57695 , n404867 , n404868 );
buf ( n404870 , n57695 );
buf ( n404871 , n404870 );
nand ( n57698 , n57692 , n404871 );
buf ( n404873 , n57698 );
nand ( n57700 , n57672 , n404873 );
nand ( n57701 , n57668 , n57700 );
buf ( n404876 , n57701 );
and ( n57703 , n57642 , n404876 );
and ( n57704 , n404797 , n404815 );
or ( n57705 , n57703 , n57704 );
buf ( n404880 , n57705 );
nand ( n57707 , n57412 , n404880 );
nand ( n57708 , n57406 , n57707 );
nand ( n57709 , n57294 , n57708 );
nand ( n57710 , n57293 , n57709 );
buf ( n404885 , n57710 );
and ( n57712 , n57281 , n404885 );
and ( n57713 , n404450 , n404454 );
or ( n57714 , n57712 , n57713 );
buf ( n404889 , n57714 );
buf ( n404890 , n404889 );
xor ( n57717 , n403619 , n403623 );
xor ( n57718 , n57717 , n403902 );
buf ( n404893 , n57718 );
buf ( n404894 , n404893 );
xor ( n57721 , n404890 , n404894 );
not ( n57722 , n403895 );
not ( n57723 , n403732 );
or ( n57724 , n57722 , n57723 );
buf ( n404899 , n56522 );
buf ( n404900 , n56699 );
nand ( n57727 , n404899 , n404900 );
buf ( n404902 , n57727 );
nand ( n57729 , n57724 , n404902 );
not ( n57730 , n56531 );
and ( n57731 , n57729 , n57730 );
not ( n57732 , n57729 );
and ( n57733 , n57732 , n56531 );
nor ( n57734 , n57731 , n57733 );
buf ( n404909 , n57734 );
not ( n57736 , n404909 );
xor ( n57737 , n56749 , n404271 );
xor ( n57738 , n57737 , n404385 );
buf ( n404913 , n57738 );
not ( n57740 , n404913 );
or ( n57741 , n57736 , n57740 );
xor ( n57742 , n403684 , n56463 );
xnor ( n57743 , n57742 , n56514 );
buf ( n404918 , n57743 );
not ( n57745 , n404918 );
buf ( n404920 , n57745 );
buf ( n404921 , n404920 );
not ( n57748 , n404921 );
xor ( n57749 , n56562 , n403772 );
xor ( n57750 , n57749 , n403883 );
not ( n57751 , n56611 );
xor ( n57752 , n56686 , n57751 );
buf ( n57753 , n56631 );
xnor ( n57754 , n57752 , n57753 );
not ( n57755 , n57754 );
or ( n57768 , n57755 , C1 );
xor ( n57769 , n57751 , n56686 );
xor ( n57770 , n57769 , n56631 );
not ( n57771 , n57770 );
or ( n57776 , n57771 , C0 );
xor ( n57777 , n404011 , n404123 );
xor ( n57778 , n57777 , n56953 );
buf ( n404937 , n57778 );
not ( n57780 , n404937 );
buf ( n404939 , n57780 );
nand ( n57782 , n57776 , n404939 );
nand ( n57783 , n57768 , n57782 );
buf ( n404942 , n57783 );
not ( n57785 , n404942 );
buf ( n404944 , n57785 );
xor ( n57787 , n57750 , n404944 );
not ( n57788 , n56432 );
not ( n57789 , n57788 );
not ( n57790 , n56461 );
or ( n57791 , n57789 , n57790 );
or ( n57792 , n57788 , n56461 );
nand ( n57793 , n57791 , n57792 );
buf ( n404952 , C1 );
and ( n57797 , n57793 , n404952 );
nor ( n57800 , n57797 , C0 );
and ( n57801 , n57787 , n57800 );
and ( n57802 , n57750 , n404944 );
or ( n57803 , n57801 , n57802 );
buf ( n404958 , n57803 );
not ( n57805 , n404958 );
buf ( n404960 , n57805 );
buf ( n404961 , n404960 );
not ( n57808 , n404961 );
or ( n57809 , n57748 , n57808 );
buf ( n404964 , n57743 );
not ( n57811 , n404964 );
buf ( n404966 , n57803 );
not ( n57813 , n404966 );
or ( n57814 , n57811 , n57813 );
not ( n57816 , n56785 );
or ( n57817 , C0 , n57816 );
nand ( n57820 , n57817 , C1 );
and ( n57821 , n57820 , n56767 );
not ( n57822 , n57820 );
not ( n57823 , n56767 );
and ( n57824 , n57822 , n57823 );
nor ( n57825 , n57821 , n57824 );
buf ( n404977 , n57825 );
not ( n57827 , n404977 );
buf ( n404979 , n57827 );
not ( n57829 , n404979 );
xor ( n57830 , n404130 , n404155 );
xor ( n57831 , n57830 , n404260 );
buf ( n404983 , n57831 );
not ( n57833 , n404983 );
or ( n57834 , n57829 , n57833 );
buf ( n404986 , n404983 );
not ( n57836 , n404986 );
buf ( n404988 , n57836 );
not ( n57838 , n404988 );
not ( n57839 , n57825 );
or ( n57840 , n57838 , n57839 );
buf ( n404992 , n392740 );
not ( n57842 , n404992 );
buf ( n404994 , n404144 );
not ( n57844 , n404994 );
or ( n57845 , n57842 , n57844 );
buf ( n404997 , n399986 );
not ( n57847 , n404997 );
buf ( n404999 , n48233 );
not ( n57849 , n404999 );
or ( n57850 , n57847 , n57849 );
buf ( n405002 , n36217 );
buf ( n405003 , n392244 );
nand ( n57853 , n405002 , n405003 );
buf ( n405005 , n57853 );
buf ( n405006 , n405005 );
nand ( n57856 , n57850 , n405006 );
buf ( n405008 , n57856 );
buf ( n405009 , n405008 );
buf ( n405010 , n45260 );
nand ( n57860 , n405009 , n405010 );
buf ( n405012 , n57860 );
buf ( n405013 , n405012 );
nand ( n57863 , n57845 , n405013 );
buf ( n405015 , n57863 );
buf ( n405016 , n405015 );
and ( n57866 , n56937 , n404015 );
not ( n57867 , n56937 );
and ( n57868 , n57867 , n56943 );
nor ( n57869 , n57866 , n57868 );
nand ( n57870 , n56853 , n56855 );
and ( n57871 , n57869 , n57870 );
not ( n57872 , n57869 );
not ( n57873 , n57870 );
and ( n57874 , n57872 , n57873 );
nor ( n57875 , n57871 , n57874 );
not ( n57876 , n57875 );
not ( n57877 , n57876 );
not ( n57878 , n392111 );
not ( n57879 , n404215 );
or ( n57880 , n57878 , n57879 );
not ( n57881 , n388359 );
not ( n57882 , n36810 );
not ( n57883 , n394219 );
or ( n57884 , n57882 , n57883 );
nand ( n57885 , n396373 , n394210 );
nand ( n57886 , n57884 , n57885 );
nand ( n57887 , n57881 , n57886 );
nand ( n57888 , n57880 , n57887 );
buf ( n57889 , n382984 );
and ( n57890 , n397524 , n57889 );
nor ( n57891 , n57890 , n37402 );
buf ( n405043 , n57891 );
buf ( n405044 , n397524 );
buf ( n405045 , n382984 );
or ( n57895 , n405044 , n405045 );
buf ( n405047 , n358975 );
nand ( n57897 , n57895 , n405047 );
buf ( n405049 , n57897 );
buf ( n405050 , n405049 );
nand ( n57900 , n405043 , n405050 );
buf ( n405052 , n57900 );
not ( n57902 , n405052 );
or ( n57903 , n57888 , n57902 );
buf ( n405055 , n404080 );
not ( n57905 , n405055 );
buf ( n405057 , n57905 );
buf ( n405058 , n405057 );
not ( n57908 , n405058 );
and ( n57909 , n404054 , n404106 );
not ( n57910 , n404054 );
and ( n57911 , n57910 , n404109 );
or ( n57912 , n57909 , n57911 );
buf ( n405064 , n57912 );
not ( n57914 , n405064 );
or ( n57915 , n57908 , n57914 );
buf ( n405067 , n57912 );
buf ( n405068 , n405057 );
or ( n57918 , n405067 , n405068 );
nand ( n57919 , n57915 , n57918 );
buf ( n405071 , n57919 );
nand ( n57921 , n57903 , n405071 );
buf ( n405073 , n57921 );
nand ( n57923 , n57888 , n57902 );
buf ( n405075 , n57923 );
and ( n57925 , n405073 , n405075 );
buf ( n405077 , n57925 );
buf ( n405078 , n405077 );
not ( n57928 , n405078 );
buf ( n405080 , n57928 );
not ( n57930 , n405080 );
or ( n57931 , n57877 , n57930 );
buf ( n405083 , n57875 );
not ( n57933 , n405083 );
buf ( n405085 , n405077 );
not ( n57935 , n405085 );
or ( n57936 , n57933 , n57935 );
and ( n57937 , n392620 , n36396 );
not ( n57938 , n392620 );
and ( n57939 , n57938 , n47256 );
nor ( n57940 , n57937 , n57939 );
or ( n57941 , n388463 , n57940 );
nor ( n57942 , n388349 , n404025 );
not ( n57943 , n57942 );
nand ( n57944 , n57941 , n57943 );
buf ( n405096 , n389341 );
not ( n57946 , n405096 );
buf ( n405098 , n388266 );
not ( n57948 , n405098 );
or ( n57949 , n57946 , n57948 );
buf ( n405101 , n388263 );
buf ( n405102 , n393185 );
nand ( n57952 , n405101 , n405102 );
buf ( n405104 , n57952 );
buf ( n405105 , n405104 );
nand ( n57955 , n57949 , n405105 );
buf ( n405107 , n57955 );
not ( n57957 , n405107 );
not ( n57958 , n383891 );
or ( n57959 , n57957 , n57958 );
buf ( n405111 , n403840 );
buf ( n405112 , n391602 );
nand ( n57962 , n405111 , n405112 );
buf ( n405114 , n57962 );
nand ( n57964 , n57959 , n405114 );
or ( n57965 , n57944 , n57964 );
not ( n57966 , n396622 );
buf ( n405118 , n12471 );
not ( n57968 , n405118 );
buf ( n405120 , n398298 );
not ( n57970 , n405120 );
or ( n57971 , n57968 , n57970 );
buf ( n405123 , n399167 );
buf ( n405124 , n12471 );
not ( n57974 , n405124 );
buf ( n405126 , n57974 );
buf ( n405127 , n405126 );
nand ( n57977 , n405123 , n405127 );
buf ( n405129 , n57977 );
buf ( n405130 , n405129 );
nand ( n57980 , n57971 , n405130 );
buf ( n405132 , n57980 );
not ( n57982 , n405132 );
or ( n57983 , n57966 , n57982 );
buf ( n405135 , n403055 );
buf ( n405136 , n55831 );
nand ( n57986 , n405135 , n405136 );
buf ( n405138 , n57986 );
nand ( n57988 , n57983 , n405138 );
not ( n57989 , n57988 );
not ( n57990 , n397476 );
and ( n57991 , n388643 , n404601 );
not ( n57992 , n388643 );
and ( n57993 , n57992 , n394884 );
or ( n57994 , n57991 , n57993 );
not ( n57995 , n57994 );
or ( n57996 , n57990 , n57995 );
not ( n57997 , n57422 );
not ( n57998 , n404604 );
or ( n57999 , n57997 , n57998 );
nand ( n58000 , n57999 , n47726 );
nand ( n58001 , n57996 , n58000 );
not ( n58002 , n58001 );
or ( n58003 , n57989 , n58002 );
or ( n58004 , n57988 , n58001 );
buf ( n405156 , n42924 );
not ( n58006 , n405156 );
buf ( n405158 , n57507 );
not ( n58008 , n405158 );
or ( n58009 , n58006 , n58008 );
buf ( n405161 , n41559 );
not ( n58011 , n405161 );
buf ( n405163 , n403039 );
not ( n58013 , n405163 );
or ( n58014 , n58011 , n58013 );
buf ( n405166 , n41558 );
buf ( n405167 , n28644 );
nand ( n58017 , n405166 , n405167 );
buf ( n405169 , n58017 );
buf ( n405170 , n405169 );
nand ( n58020 , n58014 , n405170 );
buf ( n405172 , n58020 );
buf ( n405173 , n405172 );
buf ( n405174 , n52812 );
nand ( n58024 , n405173 , n405174 );
buf ( n405176 , n58024 );
buf ( n405177 , n405176 );
nand ( n58027 , n58009 , n405177 );
buf ( n405179 , n58027 );
not ( n58029 , n405179 );
xor ( n58030 , n403096 , n403141 );
xor ( n58031 , n58030 , n403171 );
xor ( n58032 , n403225 , n403340 );
xor ( n58033 , n58031 , n58032 );
not ( n58034 , n58033 );
or ( n58035 , n58029 , n58034 );
nor ( n58036 , n58033 , n405179 );
xor ( n58037 , n403235 , n403252 );
xor ( n58038 , n58037 , n403336 );
buf ( n405190 , n58038 );
buf ( n405191 , n405190 );
not ( n58041 , n54430 );
nand ( n58042 , n58041 , n54432 );
buf ( n405194 , n58042 );
buf ( n405195 , n55905 );
and ( n58045 , n405194 , n405195 );
buf ( n405197 , n403088 );
buf ( n405198 , n55895 );
and ( n58048 , n405197 , n405198 );
nor ( n58049 , n58045 , n58048 );
buf ( n405201 , n58049 );
buf ( n405202 , n405201 );
buf ( n405203 , n403120 );
or ( n58053 , n405202 , n405203 );
buf ( n405205 , n403261 );
buf ( n405206 , n403133 );
or ( n58056 , n405205 , n405206 );
nand ( n58057 , n58053 , n58056 );
buf ( n405209 , n58057 );
buf ( n405210 , n405209 );
buf ( n405211 , n54336 );
buf ( n58061 , n55870 );
buf ( n405213 , n58061 );
not ( n58063 , n405213 );
buf ( n405215 , n58063 );
buf ( n405216 , n405215 );
and ( n58066 , n405211 , n405216 );
buf ( n405218 , n401699 );
buf ( n405219 , n58061 );
and ( n58069 , n405218 , n405219 );
nor ( n58070 , n58066 , n58069 );
buf ( n405222 , n58070 );
buf ( n405223 , n405222 );
buf ( n405224 , n403293 );
or ( n58074 , n405223 , n405224 );
buf ( n405226 , n403309 );
nand ( n58076 , n58074 , n405226 );
buf ( n405228 , n58076 );
buf ( n405229 , n405228 );
nor ( n58079 , n405210 , n405229 );
buf ( n405231 , n58079 );
buf ( n405232 , n405231 );
not ( n58082 , n53419 );
not ( n58083 , n54270 );
or ( n58084 , n58082 , n58083 );
nand ( n58085 , n58084 , n54276 );
nand ( n58086 , n53472 , n54280 );
nor ( n58087 , n58085 , n58086 );
not ( n58088 , n58087 );
nand ( n58089 , n58085 , n58086 );
nand ( n58090 , n58088 , n58089 );
buf ( n405242 , n58090 );
buf ( n405243 , n401626 );
and ( n58093 , n405242 , n405243 );
buf ( n405245 , n55984 );
buf ( n405246 , n401650 );
and ( n58096 , n405245 , n405246 );
nor ( n58097 , n58093 , n58096 );
buf ( n405249 , n58097 );
buf ( n405250 , n405249 );
or ( n58100 , n405232 , n405250 );
buf ( n405252 , n405249 );
not ( n58102 , n405252 );
buf ( n405254 , n405231 );
not ( n58104 , n405254 );
or ( n58105 , n58102 , n58104 );
xor ( n58106 , n403270 , n403313 );
xor ( n58107 , n58106 , n403331 );
buf ( n405259 , n58107 );
buf ( n405260 , n405259 );
nand ( n58110 , n58105 , n405260 );
buf ( n405262 , n58110 );
buf ( n405263 , n405262 );
nand ( n58113 , n58100 , n405263 );
buf ( n405265 , n58113 );
buf ( n405266 , n405265 );
and ( n58116 , n405191 , n405266 );
buf ( n405268 , n405190 );
not ( n58118 , n405268 );
buf ( n405270 , n405265 );
not ( n58120 , n405270 );
and ( n58121 , n58118 , n58120 );
buf ( n405273 , n405259 );
buf ( n405274 , n405231 );
buf ( n405275 , n405249 );
xor ( n58125 , n405274 , n405275 );
buf ( n405277 , n58125 );
buf ( n405278 , n405277 );
xnor ( n58128 , n405273 , n405278 );
buf ( n405280 , n58128 );
buf ( n405281 , n405280 );
not ( n58131 , n405281 );
buf ( n405283 , n55984 );
buf ( n405284 , n403146 );
and ( n58134 , n405283 , n405284 );
not ( n58135 , n55984 );
buf ( n405287 , n58135 );
buf ( n405288 , n401695 );
and ( n58138 , n405287 , n405288 );
nor ( n58139 , n58134 , n58138 );
buf ( n405291 , n58139 );
buf ( n405292 , n405291 );
not ( n58142 , n405292 );
buf ( n405294 , n58142 );
buf ( n405295 , n405294 );
buf ( n405296 , n401674 );
and ( n58146 , n405295 , n405296 );
buf ( n405298 , n403322 );
not ( n58148 , n405298 );
buf ( n405300 , n58148 );
buf ( n405301 , n405300 );
buf ( n405302 , n403164 );
and ( n58152 , n405301 , n405302 );
nor ( n58153 , n58146 , n58152 );
buf ( n405305 , n58153 );
buf ( n405306 , n405305 );
not ( n58156 , n53394 );
not ( n58157 , n54270 );
or ( n58158 , n58156 , n58157 );
not ( n58159 , n54273 );
nand ( n58160 , n58158 , n58159 );
not ( n58161 , n54275 );
nand ( n58162 , n58161 , n53418 );
nor ( n58163 , n58160 , n58162 );
not ( n58164 , n58163 );
nand ( n58165 , n58160 , n58162 );
nand ( n58166 , n58164 , n58165 );
buf ( n405318 , n58166 );
buf ( n405319 , n401626 );
and ( n58169 , n405318 , n405319 );
buf ( n405321 , n58090 );
buf ( n405322 , n401650 );
and ( n58172 , n405321 , n405322 );
nor ( n58173 , n58169 , n58172 );
buf ( n405325 , n58173 );
buf ( n405326 , n405325 );
xor ( n58176 , n405306 , n405326 );
not ( n58177 , n58087 );
nand ( n58178 , n58177 , n58089 );
buf ( n405330 , n58178 );
buf ( n405331 , n403146 );
and ( n58181 , n405330 , n405331 );
buf ( n405333 , n58090 );
not ( n58183 , n405333 );
buf ( n405335 , n58183 );
buf ( n405336 , n405335 );
buf ( n405337 , n401695 );
and ( n58187 , n405336 , n405337 );
nor ( n58188 , n58181 , n58187 );
buf ( n405340 , n58188 );
buf ( n405341 , n405340 );
buf ( n405342 , n403158 );
or ( n58192 , n405341 , n405342 );
buf ( n405344 , n405291 );
buf ( n405345 , n403167 );
or ( n58195 , n405344 , n405345 );
nand ( n58196 , n58192 , n58195 );
buf ( n405348 , n58196 );
buf ( n405349 , n405348 );
nand ( n58199 , n53394 , n58159 );
xnor ( n58200 , n54270 , n58199 );
not ( n58201 , n58200 );
buf ( n405353 , n58201 );
buf ( n405354 , n403083 );
or ( n58204 , n405353 , n405354 );
not ( n58205 , n58166 );
buf ( n405357 , n58205 );
buf ( n405358 , n403092 );
or ( n58208 , n405357 , n405358 );
nand ( n58209 , n58204 , n58208 );
buf ( n405361 , n58209 );
buf ( n405362 , n405361 );
and ( n58212 , n405349 , n405362 );
buf ( n405364 , n405348 );
not ( n58214 , n405364 );
buf ( n405366 , n405361 );
not ( n58216 , n405366 );
and ( n58217 , n58214 , n58216 );
not ( n58218 , n13935 );
buf ( n405370 , n58218 );
buf ( n405371 , n14083 );
and ( n58221 , n405370 , n405371 );
not ( n58222 , n405370 );
not ( n58223 , n14083 );
buf ( n405375 , n58223 );
and ( n58225 , n58222 , n405375 );
nor ( n58226 , n58221 , n58225 );
buf ( n405378 , n58226 );
buf ( n405379 , n405378 );
not ( n58229 , n405379 );
buf ( n405381 , n58229 );
buf ( n405382 , n405381 );
not ( n58232 , n405382 );
buf ( n405384 , n58232 );
buf ( n405385 , n405384 );
buf ( n405386 , n403283 );
not ( n58236 , n405386 );
buf ( n405388 , n58236 );
buf ( n405389 , n405388 );
not ( n58239 , n405389 );
buf ( n405391 , n58239 );
buf ( n405392 , n405391 );
nor ( n58242 , n405385 , n405392 );
buf ( n405394 , n58242 );
buf ( n405395 , n405394 );
not ( n58245 , n405395 );
buf ( n405397 , n56050 );
buf ( n405398 , n58218 );
or ( n58248 , n405397 , n405398 );
buf ( n405400 , n56050 );
buf ( n405401 , n58218 );
nand ( n58251 , n405400 , n405401 );
buf ( n405403 , n58251 );
buf ( n405404 , n405403 );
buf ( n405405 , n405378 );
nand ( n58255 , n58248 , n405404 , n405405 );
buf ( n405407 , n58255 );
buf ( n405408 , n405407 );
not ( n58258 , n405408 );
buf ( n405410 , n58258 );
buf ( n405411 , n405410 );
buf ( n405412 , n405388 );
nand ( n58262 , n405411 , n405412 );
buf ( n405414 , n58262 );
buf ( n405415 , n405414 );
nand ( n58265 , n58245 , n405415 );
buf ( n405417 , n58265 );
buf ( n405418 , n405417 );
nor ( n58268 , n58217 , n405418 );
buf ( n405420 , n58268 );
buf ( n405421 , n405420 );
nor ( n58271 , n58212 , n405421 );
buf ( n405423 , n58271 );
buf ( n405424 , n405423 );
and ( n58274 , n58176 , n405424 );
and ( n58275 , n405306 , n405326 );
or ( n58276 , n58274 , n58275 );
buf ( n405428 , n58276 );
buf ( n405429 , n405428 );
not ( n58279 , n405429 );
and ( n58280 , n58131 , n58279 );
buf ( n405432 , n405280 );
buf ( n405433 , n405428 );
and ( n58283 , n405432 , n405433 );
buf ( n405435 , n405209 );
buf ( n405436 , n405228 );
and ( n58286 , n405435 , n405436 );
buf ( n405438 , n405231 );
nor ( n58288 , n58286 , n405438 );
buf ( n405440 , n58288 );
buf ( n405441 , n405440 );
not ( n58291 , n405441 );
buf ( n405443 , n58291 );
buf ( n405444 , n405443 );
buf ( n405445 , n55846 );
buf ( n405446 , n55905 );
and ( n58296 , n405445 , n405446 );
buf ( n405448 , n403079 );
buf ( n405449 , n55895 );
and ( n58299 , n405448 , n405449 );
nor ( n58300 , n58296 , n58299 );
buf ( n405452 , n58300 );
buf ( n405453 , n405452 );
buf ( n405454 , n403120 );
or ( n58304 , n405453 , n405454 );
buf ( n405456 , n405201 );
buf ( n405457 , n403133 );
or ( n58307 , n405456 , n405457 );
nand ( n58308 , n58304 , n58307 );
buf ( n405460 , n58308 );
buf ( n405461 , n405460 );
buf ( n405462 , n54297 );
buf ( n405463 , n405215 );
and ( n58313 , n405462 , n405463 );
buf ( n405465 , n55919 );
buf ( n405466 , n58061 );
and ( n58316 , n405465 , n405466 );
nor ( n58317 , n58313 , n58316 );
buf ( n405469 , n58317 );
buf ( n405470 , n405469 );
buf ( n405471 , n403293 );
or ( n58321 , n405470 , n405471 );
buf ( n405473 , n405222 );
buf ( n405474 , n403305 );
not ( n58324 , n405474 );
buf ( n405476 , n58324 );
buf ( n405477 , n405476 );
or ( n58327 , n405473 , n405477 );
nand ( n58328 , n58321 , n58327 );
buf ( n405480 , n58328 );
buf ( n405481 , n405480 );
xor ( n58331 , n405461 , n405481 );
buf ( n405483 , n54336 );
buf ( n405484 , n405391 );
and ( n58334 , n405483 , n405484 );
buf ( n405486 , n401699 );
buf ( n405487 , n405388 );
and ( n58337 , n405486 , n405487 );
nor ( n58338 , n58334 , n58337 );
buf ( n405490 , n58338 );
buf ( n405491 , n405490 );
not ( n58341 , n405491 );
buf ( n405493 , n58341 );
buf ( n405494 , n405493 );
buf ( n405495 , n405410 );
and ( n58345 , n405494 , n405495 );
buf ( n405497 , n405394 );
nor ( n58347 , n58345 , n405497 );
buf ( n405499 , n58347 );
buf ( n405500 , n405499 );
not ( n58350 , n401578 );
nand ( n58351 , n58350 , n53653 );
xnor ( n58352 , n54414 , n58351 );
buf ( n405504 , n58352 );
buf ( n405505 , n401626 );
and ( n58355 , n405504 , n405505 );
buf ( n405507 , n58200 );
buf ( n405508 , n401650 );
and ( n58358 , n405507 , n405508 );
nor ( n58359 , n58355 , n58358 );
buf ( n405511 , n58359 );
buf ( n405512 , n405511 );
nand ( n58362 , n405500 , n405512 );
buf ( n405514 , n58362 );
buf ( n405515 , n405514 );
and ( n58365 , n58331 , n405515 );
and ( n58366 , n405461 , n405481 );
or ( n58367 , n58365 , n58366 );
buf ( n405519 , n58367 );
buf ( n405520 , n405519 );
and ( n58370 , n405444 , n405520 );
buf ( n405522 , n405443 );
not ( n58372 , n405522 );
buf ( n405524 , n405519 );
not ( n58374 , n405524 );
and ( n58375 , n58372 , n58374 );
xor ( n58376 , n405306 , n405326 );
xor ( n58377 , n58376 , n405424 );
buf ( n405529 , n58377 );
buf ( n405530 , n405529 );
nor ( n58380 , n58375 , n405530 );
buf ( n405532 , n58380 );
buf ( n405533 , n405532 );
nor ( n58383 , n58370 , n405533 );
buf ( n405535 , n58383 );
buf ( n405536 , n405535 );
nor ( n58386 , n58283 , n405536 );
buf ( n405538 , n58386 );
buf ( n405539 , n405538 );
nor ( n58389 , n58280 , n405539 );
buf ( n405541 , n58389 );
buf ( n405542 , n405541 );
nor ( n58392 , n58121 , n405542 );
buf ( n405544 , n58392 );
buf ( n405545 , n405544 );
nor ( n58395 , n58116 , n405545 );
buf ( n405547 , n58395 );
or ( n58397 , n58036 , n405547 );
nand ( n58398 , n58035 , n58397 );
nand ( n58399 , n58004 , n58398 );
nand ( n58400 , n58003 , n58399 );
nand ( n58401 , n57965 , n58400 );
nand ( n58402 , n57944 , n57964 );
nand ( n58403 , n58401 , n58402 );
buf ( n405555 , n58403 );
nand ( n58405 , n57936 , n405555 );
buf ( n405557 , n58405 );
nand ( n58407 , n57931 , n405557 );
buf ( n405559 , n58407 );
xor ( n58409 , n405016 , n405559 );
xor ( n58410 , n404181 , n404185 );
xor ( n58411 , n58410 , n404255 );
buf ( n405563 , n58411 );
buf ( n405564 , n405563 );
and ( n58414 , n58409 , n405564 );
and ( n58415 , n405016 , n405559 );
or ( n58416 , n58414 , n58415 );
buf ( n405568 , n58416 );
nand ( n58418 , n57840 , n405568 );
nand ( n58419 , n57834 , n58418 );
buf ( n405571 , n58419 );
nand ( n58421 , n57814 , n405571 );
buf ( n405573 , n58421 );
buf ( n405574 , n405573 );
nand ( n58424 , n57809 , n405574 );
buf ( n405576 , n58424 );
buf ( n405577 , n405576 );
nand ( n58427 , n57741 , n405577 );
buf ( n405579 , n58427 );
buf ( n405580 , n405579 );
buf ( n405581 , n57734 );
not ( n58431 , n405581 );
buf ( n405583 , n57738 );
not ( n58433 , n405583 );
buf ( n405585 , n58433 );
buf ( n405586 , n405585 );
nand ( n58436 , n58431 , n405586 );
buf ( n405588 , n58436 );
buf ( n405589 , n405588 );
nand ( n58439 , n405580 , n405589 );
buf ( n405591 , n58439 );
buf ( n405592 , n405591 );
and ( n58442 , n57721 , n405592 );
and ( n58443 , n404890 , n404894 );
or ( n58444 , n58442 , n58443 );
buf ( n405596 , n58444 );
buf ( n405597 , n405596 );
buf ( n58447 , n405597 );
buf ( n405599 , n58447 );
xor ( n58449 , n402590 , n56263 );
xor ( n58450 , n58449 , n403500 );
not ( n58451 , n58450 );
and ( n58452 , n403909 , n403914 );
not ( n58453 , n403909 );
and ( n58454 , n58453 , n56722 );
nor ( n58455 , n58452 , n58454 );
and ( n58456 , n58455 , n57221 );
not ( n58457 , n58455 );
not ( n58458 , n57221 );
and ( n58459 , n58457 , n58458 );
nor ( n58460 , n58456 , n58459 );
nand ( n58461 , n58451 , n58460 );
and ( n58462 , n405599 , n58461 );
not ( n58463 , n58450 );
nor ( n58464 , n58463 , n58460 );
nor ( n58465 , n58462 , n58464 );
buf ( n405617 , n58465 );
nand ( n58467 , n404446 , n405617 );
buf ( n405619 , n58467 );
nand ( n58469 , n57268 , n405619 );
not ( n58470 , n58469 );
buf ( n405622 , n58470 );
nand ( n58472 , n403537 , n405622 );
buf ( n405624 , n58472 );
buf ( n405625 , n405624 );
not ( n58475 , n405625 );
buf ( n405627 , n58475 );
not ( n58477 , n405576 );
not ( n58478 , n58477 );
not ( n58479 , n57734 );
not ( n58480 , n58479 );
or ( n58481 , n58478 , n58480 );
nand ( n58482 , n57734 , n405576 );
nand ( n58483 , n58481 , n58482 );
and ( n58484 , n58483 , n405585 );
not ( n58485 , n58483 );
buf ( n405637 , n405585 );
not ( n58487 , n405637 );
buf ( n405639 , n58487 );
and ( n58489 , n58485 , n405639 );
nor ( n58490 , n58484 , n58489 );
buf ( n405642 , n58419 );
buf ( n405643 , n404920 );
and ( n58493 , n405642 , n405643 );
not ( n58494 , n405642 );
buf ( n405646 , n57743 );
and ( n58496 , n58494 , n405646 );
nor ( n58497 , n58493 , n58496 );
buf ( n405649 , n58497 );
xnor ( n58499 , n57803 , n405649 );
buf ( n405651 , n58499 );
buf ( n405652 , n56808 );
buf ( n405653 , n403957 );
and ( n58503 , n405652 , n405653 );
not ( n58504 , n405652 );
buf ( n405656 , n403954 );
and ( n58506 , n58504 , n405656 );
nor ( n58507 , n58503 , n58506 );
buf ( n405659 , n58507 );
xor ( n58509 , n404264 , n405659 );
buf ( n405661 , n58509 );
xor ( n58511 , n404278 , n404282 );
xor ( n58512 , n58511 , n404381 );
buf ( n405664 , n58512 );
buf ( n405665 , n405664 );
xor ( n58515 , n405661 , n405665 );
buf ( n405667 , n395362 );
not ( n58517 , n405667 );
buf ( n405669 , n403970 );
not ( n58519 , n405669 );
or ( n58520 , n58517 , n58519 );
buf ( n405672 , n47863 );
not ( n58522 , n405672 );
buf ( n405674 , n385774 );
not ( n58524 , n405674 );
or ( n58525 , n58522 , n58524 );
buf ( n405677 , n389423 );
buf ( n405678 , n395315 );
nand ( n58528 , n405677 , n405678 );
buf ( n405680 , n58528 );
buf ( n405681 , n405680 );
nand ( n58531 , n58525 , n405681 );
buf ( n405683 , n58531 );
buf ( n405684 , n405683 );
buf ( n405685 , n395349 );
nand ( n58535 , n405684 , n405685 );
buf ( n405687 , n58535 );
buf ( n405688 , n405687 );
nand ( n58538 , n58520 , n405688 );
buf ( n405690 , n58538 );
not ( n58540 , n405690 );
not ( n58541 , n43727 );
not ( n58542 , n391027 );
not ( n58543 , n394120 );
or ( n58544 , n58542 , n58543 );
not ( n58545 , n36708 );
buf ( n58546 , n58545 );
buf ( n405698 , n58546 );
buf ( n405699 , n391024 );
nand ( n58549 , n405698 , n405699 );
buf ( n405701 , n58549 );
nand ( n58551 , n58544 , n405701 );
not ( n58552 , n58551 );
or ( n58553 , n58541 , n58552 );
not ( n58554 , n404317 );
nand ( n58555 , n58554 , n43515 );
nand ( n58556 , n58553 , n58555 );
not ( n58557 , n58556 );
not ( n58558 , n45260 );
not ( n58559 , n398366 );
not ( n58560 , n392244 );
or ( n58561 , n58559 , n58560 );
buf ( n405713 , n390119 );
not ( n58563 , n405713 );
buf ( n405715 , n58563 );
nand ( n58565 , n405715 , n399986 );
nand ( n58566 , n58561 , n58565 );
not ( n58567 , n58566 );
or ( n58568 , n58558 , n58567 );
nand ( n58569 , n405008 , n392740 );
nand ( n58570 , n58568 , n58569 );
not ( n58571 , n58570 );
or ( n58572 , n58557 , n58571 );
not ( n58573 , n58556 );
buf ( n405725 , n58573 );
not ( n58575 , n405725 );
not ( n58576 , n58570 );
buf ( n405728 , n58576 );
not ( n58578 , n405728 );
or ( n58579 , n58575 , n58578 );
not ( n58580 , n388809 );
not ( n58581 , n404199 );
or ( n58582 , n58580 , n58581 );
buf ( n405734 , n388754 );
not ( n58584 , n405734 );
buf ( n405736 , n58584 );
buf ( n405737 , n405736 );
not ( n58587 , n405737 );
buf ( n405739 , n388919 );
not ( n58589 , n405739 );
or ( n58590 , n58587 , n58589 );
buf ( n405742 , n389940 );
buf ( n405743 , n388757 );
nand ( n58593 , n405742 , n405743 );
buf ( n405745 , n58593 );
buf ( n405746 , n405745 );
nand ( n58596 , n58590 , n405746 );
buf ( n405748 , n58596 );
buf ( n405749 , n405748 );
buf ( n405750 , n388746 );
nand ( n58600 , n405749 , n405750 );
buf ( n405752 , n58600 );
nand ( n58602 , n58582 , n405752 );
not ( n58603 , n40990 );
not ( n58604 , n388965 );
or ( n58605 , n58603 , n58604 );
buf ( n405757 , n385473 );
buf ( n405758 , n390460 );
nand ( n58608 , n405757 , n405758 );
buf ( n405760 , n58608 );
nand ( n58610 , n58605 , n405760 );
buf ( n405762 , n58610 );
not ( n58612 , n405762 );
buf ( n405764 , n393544 );
not ( n58614 , n405764 );
or ( n58615 , n58612 , n58614 );
buf ( n405767 , n404067 );
buf ( n405768 , n51692 );
nand ( n58618 , n405767 , n405768 );
buf ( n405770 , n58618 );
buf ( n405771 , n405770 );
nand ( n58621 , n58615 , n405771 );
buf ( n405773 , n58621 );
not ( n58623 , n405773 );
not ( n58624 , n388833 );
not ( n58625 , n57477 );
or ( n58626 , n58624 , n58625 );
buf ( n405778 , n41342 );
not ( n58628 , n405778 );
buf ( n405780 , n388409 );
not ( n58630 , n405780 );
or ( n58631 , n58628 , n58630 );
buf ( n405783 , n46043 );
not ( n58633 , n405783 );
buf ( n405785 , n58633 );
buf ( n405786 , n405785 );
buf ( n405787 , n45897 );
nand ( n58637 , n405786 , n405787 );
buf ( n405789 , n58637 );
buf ( n405790 , n405789 );
nand ( n58640 , n58631 , n405790 );
buf ( n405792 , n58640 );
buf ( n405793 , n405792 );
buf ( n405794 , n388872 );
nand ( n58644 , n405793 , n405794 );
buf ( n405796 , n58644 );
nand ( n58646 , n58626 , n405796 );
not ( n58647 , n58646 );
or ( n58648 , n58623 , n58647 );
or ( n58649 , n405773 , n58646 );
xor ( n58650 , n404671 , n404689 );
xor ( n58651 , n58650 , n404715 );
buf ( n405803 , n58651 );
nand ( n58653 , n58649 , n405803 );
nand ( n58654 , n58648 , n58653 );
xor ( n58655 , n58602 , n58654 );
buf ( n405807 , n404741 );
buf ( n405808 , n389162 );
nand ( n58658 , n405807 , n405808 );
buf ( n405810 , n58658 );
buf ( n405811 , n24118 );
not ( n58661 , n405811 );
buf ( n405813 , n41118 );
not ( n58663 , n405813 );
or ( n58664 , n58661 , n58663 );
buf ( n405816 , n27195 );
buf ( n405817 , n24117 );
nand ( n58667 , n405816 , n405817 );
buf ( n405819 , n58667 );
buf ( n405820 , n405819 );
nand ( n58670 , n58664 , n405820 );
buf ( n405822 , n58670 );
nand ( n58672 , n405822 , n41711 );
nand ( n58673 , n405810 , n58672 );
not ( n58674 , n58673 );
not ( n58675 , n58674 );
not ( n58676 , n37338 );
and ( n58677 , n389359 , n393562 );
not ( n58678 , n389359 );
and ( n58679 , n58678 , n388908 );
nor ( n58680 , n58677 , n58679 );
not ( n58681 , n58680 );
or ( n58682 , n58676 , n58681 );
nand ( n58683 , n404624 , n37314 );
nand ( n58684 , n58682 , n58683 );
not ( n58685 , n58684 );
not ( n58686 , n58685 );
or ( n58687 , n58675 , n58686 );
buf ( n405839 , n388230 );
not ( n58689 , n405839 );
buf ( n405841 , n398298 );
not ( n58691 , n405841 );
or ( n58692 , n58689 , n58691 );
buf ( n405844 , n24049 );
buf ( n405845 , n388227 );
nand ( n58695 , n405844 , n405845 );
buf ( n405847 , n58695 );
buf ( n405848 , n405847 );
nand ( n58698 , n58692 , n405848 );
buf ( n405850 , n58698 );
buf ( n405851 , n405850 );
not ( n58701 , n405851 );
buf ( n405853 , n396622 );
not ( n58703 , n405853 );
or ( n58704 , n58701 , n58703 );
buf ( n405856 , n405132 );
buf ( n405857 , n41563 );
nand ( n58707 , n405856 , n405857 );
buf ( n405859 , n58707 );
buf ( n405860 , n405859 );
nand ( n58710 , n58704 , n405860 );
buf ( n405862 , n58710 );
buf ( n405863 , n405862 );
buf ( n405864 , n388502 );
not ( n58714 , n405864 );
buf ( n405866 , n46906 );
not ( n58716 , n405866 );
or ( n58717 , n58714 , n58716 );
buf ( n405869 , n22982 );
buf ( n405870 , n388511 );
nand ( n58720 , n405869 , n405870 );
buf ( n405872 , n58720 );
buf ( n405873 , n405872 );
nand ( n58723 , n58717 , n405873 );
buf ( n405875 , n58723 );
buf ( n405876 , n405875 );
not ( n58726 , n405876 );
buf ( n405878 , n397102 );
not ( n58728 , n405878 );
or ( n58729 , n58726 , n58728 );
buf ( n405881 , n404702 );
buf ( n405882 , n386477 );
nand ( n58732 , n405881 , n405882 );
buf ( n405884 , n58732 );
buf ( n405885 , n405884 );
nand ( n58735 , n58729 , n405885 );
buf ( n405887 , n58735 );
buf ( n405888 , n405887 );
xor ( n58738 , n405863 , n405888 );
buf ( n405890 , n47726 );
not ( n58740 , n405890 );
buf ( n405892 , n57994 );
not ( n58742 , n405892 );
or ( n58743 , n58740 , n58742 );
buf ( n405895 , n404601 );
not ( n58745 , n405895 );
buf ( n405897 , n58745 );
buf ( n405898 , n405897 );
not ( n58748 , n405898 );
buf ( n405900 , n389856 );
not ( n58750 , n405900 );
or ( n58751 , n58748 , n58750 );
buf ( n405903 , n49686 );
buf ( n405904 , n388154 );
nand ( n58754 , n405903 , n405904 );
buf ( n405906 , n58754 );
buf ( n405907 , n405906 );
nand ( n58757 , n58751 , n405907 );
buf ( n405909 , n58757 );
buf ( n405910 , n405909 );
buf ( n405911 , n397476 );
nand ( n58761 , n405910 , n405911 );
buf ( n405913 , n58761 );
buf ( n405914 , n405913 );
nand ( n58764 , n58743 , n405914 );
buf ( n405916 , n58764 );
buf ( n405917 , n405916 );
and ( n58767 , n58738 , n405917 );
and ( n405919 , n405863 , n405888 );
or ( n58769 , n58767 , n405919 );
buf ( n405921 , n58769 );
nand ( n58771 , n58687 , n405921 );
not ( n58772 , n58672 );
not ( n58773 , n405810 );
or ( n58774 , n58772 , n58773 );
nand ( n58775 , n58774 , n58684 );
nand ( n58776 , n58771 , n58775 );
and ( n58777 , n58655 , n58776 );
and ( n58778 , n58602 , n58654 );
or ( n58779 , n58777 , n58778 );
buf ( n405931 , n58779 );
nand ( n58781 , n58579 , n405931 );
buf ( n405933 , n58781 );
nand ( n58783 , n58572 , n405933 );
not ( n58784 , n58783 );
or ( n58785 , n58540 , n58784 );
or ( n58786 , n58783 , n405690 );
and ( n58787 , n404589 , n57491 );
not ( n58788 , n404589 );
and ( n58789 , n58788 , n404664 );
nor ( n58790 , n58787 , n58789 );
xor ( n58791 , n58790 , n404792 );
not ( n58792 , n58791 );
buf ( n405944 , n58792 );
not ( n58794 , n405944 );
xor ( n58795 , n57029 , n57049 );
xor ( n58796 , n58795 , n404248 );
buf ( n405948 , n58796 );
not ( n58798 , n405948 );
or ( n58799 , n58794 , n58798 );
buf ( n405951 , n58792 );
buf ( n405952 , n58796 );
or ( n58802 , n405951 , n405952 );
buf ( n405954 , n404783 );
buf ( n405955 , n404749 );
xor ( n58805 , n405954 , n405955 );
buf ( n405957 , n404719 );
xor ( n58807 , n58805 , n405957 );
buf ( n405959 , n58807 );
buf ( n405960 , n405959 );
not ( n58810 , n405960 );
buf ( n405962 , n58810 );
not ( n58812 , n405962 );
not ( n58813 , n402375 );
buf ( n405965 , n49117 );
not ( n58815 , n405965 );
buf ( n405967 , n42390 );
not ( n58817 , n405967 );
or ( n58818 , n58815 , n58817 );
buf ( n405970 , n389897 );
buf ( n405971 , n49124 );
nand ( n58821 , n405970 , n405971 );
buf ( n405973 , n58821 );
buf ( n405974 , n405973 );
nand ( n58824 , n58818 , n405974 );
buf ( n405976 , n58824 );
not ( n58826 , n405976 );
or ( n58827 , n58813 , n58826 );
buf ( n405979 , n404515 );
buf ( n405980 , n392666 );
nand ( n58830 , n405979 , n405980 );
buf ( n405982 , n58830 );
nand ( n58832 , n58827 , n405982 );
not ( n58833 , n58832 );
or ( n58834 , n58812 , n58833 );
not ( n58835 , n405959 );
not ( n58836 , n58832 );
not ( n58837 , n58836 );
or ( n58838 , n58835 , n58837 );
buf ( n405990 , n405748 );
buf ( n405991 , n388809 );
nand ( n58841 , n405990 , n405991 );
buf ( n405993 , n58841 );
buf ( n405994 , n405736 );
not ( n58844 , n405994 );
buf ( n405996 , n388293 );
not ( n58846 , n405996 );
or ( n58847 , n58844 , n58846 );
buf ( n405999 , n388892 );
buf ( n406000 , n388757 );
nand ( n58850 , n405999 , n406000 );
buf ( n406002 , n58850 );
buf ( n406003 , n406002 );
nand ( n58853 , n58847 , n406003 );
buf ( n406005 , n58853 );
nand ( n58855 , n406005 , n388746 );
nand ( n58856 , n405993 , n58855 );
buf ( n406008 , n391446 );
not ( n58858 , n406008 );
buf ( n406010 , n388299 );
not ( n58860 , n406010 );
or ( n58861 , n58858 , n58860 );
buf ( n406013 , n388263 );
buf ( n406014 , n391455 );
nand ( n58864 , n406013 , n406014 );
buf ( n406016 , n58864 );
buf ( n406017 , n406016 );
nand ( n58867 , n58861 , n406017 );
buf ( n406019 , n58867 );
not ( n58869 , n406019 );
not ( n58870 , n383891 );
or ( n58871 , n58869 , n58870 );
buf ( n406023 , n405107 );
buf ( n406024 , n388629 );
nand ( n58874 , n406023 , n406024 );
buf ( n406026 , n58874 );
nand ( n58876 , n58871 , n406026 );
nor ( n58877 , n58856 , n58876 );
buf ( n406029 , n57988 );
buf ( n406030 , n58001 );
xor ( n58880 , n406029 , n406030 );
buf ( n406032 , n58398 );
xnor ( n58882 , n58880 , n406032 );
buf ( n406034 , n58882 );
or ( n58884 , n58877 , n406034 );
not ( n58885 , n58855 );
not ( n58886 , n405993 );
or ( n58887 , n58885 , n58886 );
nand ( n58888 , n58887 , n58876 );
nand ( n58889 , n58884 , n58888 );
nand ( n58890 , n58838 , n58889 );
nand ( n58891 , n58834 , n58890 );
buf ( n406043 , n58891 );
nand ( n58893 , n58802 , n406043 );
buf ( n406045 , n58893 );
buf ( n406046 , n406045 );
nand ( n58896 , n58799 , n406046 );
buf ( n406048 , n58896 );
nand ( n58898 , n58786 , n406048 );
nand ( n58899 , n58785 , n58898 );
buf ( n406051 , n58899 );
buf ( n406052 , C0 );
buf ( n406053 , n406052 );
buf ( n406054 , n51553 );
not ( n58927 , n406054 );
buf ( n406056 , n404297 );
not ( n58929 , n406056 );
or ( n58930 , n58927 , n58929 );
buf ( n406059 , n47891 );
not ( n58932 , n406059 );
buf ( n406061 , n394307 );
not ( n58934 , n406061 );
or ( n58935 , n58932 , n58934 );
buf ( n406064 , n392333 );
not ( n58937 , n406064 );
buf ( n406066 , n403668 );
nand ( n58939 , n58937 , n406066 );
buf ( n406068 , n58939 );
buf ( n406069 , n406068 );
nand ( n58942 , n58935 , n406069 );
buf ( n406071 , n58942 );
buf ( n406072 , n406071 );
buf ( n406073 , n50579 );
nand ( n58946 , n406072 , n406073 );
buf ( n406075 , n58946 );
buf ( n406076 , n406075 );
nand ( n58949 , n58930 , n406076 );
buf ( n406078 , n58949 );
buf ( n406079 , n406078 );
xor ( n58952 , n406053 , n406079 );
not ( n58953 , n57194 );
not ( n58954 , n58953 );
not ( n58955 , n404353 );
or ( n58956 , n58954 , n58955 );
nand ( n58957 , n57194 , n404350 );
nand ( n58958 , n58956 , n58957 );
buf ( n406087 , n58958 );
buf ( n406088 , n57148 );
buf ( n58961 , n406088 );
buf ( n406090 , n58961 );
buf ( n406091 , n406090 );
not ( n58964 , n406091 );
buf ( n406093 , n58964 );
buf ( n406094 , n406093 );
and ( n58967 , n406087 , n406094 );
not ( n58968 , n406087 );
buf ( n406097 , n406090 );
and ( n58970 , n58968 , n406097 );
nor ( n58971 , n58967 , n58970 );
buf ( n406100 , n58971 );
buf ( n406101 , n406100 );
and ( n58974 , n58952 , n406101 );
or ( n58976 , n58974 , C0 );
buf ( n406104 , n58976 );
buf ( n406105 , n406104 );
xor ( n58979 , n406051 , n406105 );
xor ( n58980 , n57401 , n404566 );
xnor ( n58981 , n58980 , n404880 );
buf ( n406109 , n58981 );
and ( n58983 , n58979 , n406109 );
and ( n58984 , n406051 , n406105 );
or ( n58985 , n58983 , n58984 );
buf ( n406113 , n58985 );
buf ( n406114 , n406113 );
xor ( n58988 , n58515 , n406114 );
buf ( n406116 , n58988 );
buf ( n406117 , n406116 );
xor ( n58991 , n405651 , n406117 );
xor ( n58992 , n406051 , n406105 );
xor ( n58993 , n58992 , n406109 );
buf ( n406121 , n58993 );
buf ( n406122 , n406121 );
xor ( n58996 , n57196 , n404374 );
xnor ( n58997 , n58996 , n404307 );
buf ( n406125 , n388068 );
not ( n58999 , n406125 );
buf ( n406127 , n404547 );
not ( n59001 , n406127 );
or ( n59002 , n58999 , n59001 );
buf ( n406130 , n388105 );
buf ( n406131 , n388952 );
and ( n59005 , n406130 , n406131 );
not ( n59006 , n406130 );
buf ( n406134 , n388949 );
and ( n59008 , n59006 , n406134 );
nor ( n59009 , n59005 , n59008 );
buf ( n406137 , n59009 );
buf ( n406138 , n406137 );
not ( n59012 , n406138 );
buf ( n406140 , n43286 );
nand ( n59014 , n59012 , n406140 );
buf ( n406142 , n59014 );
buf ( n406143 , n406142 );
nand ( n59017 , n59002 , n406143 );
buf ( n406145 , n59017 );
not ( n59019 , n406145 );
buf ( n406147 , n400033 );
not ( n59021 , n406147 );
buf ( n406149 , n385987 );
not ( n59023 , n406149 );
or ( n59024 , n59021 , n59023 );
buf ( n406152 , n31964 );
buf ( n406153 , n400042 );
nand ( n59027 , n406152 , n406153 );
buf ( n406155 , n59027 );
buf ( n406156 , n406155 );
nand ( n59030 , n59024 , n406156 );
buf ( n406158 , n59030 );
buf ( n406159 , n406158 );
not ( n59033 , n406159 );
buf ( n406161 , n389015 );
not ( n59035 , n406161 );
or ( n59036 , n59033 , n59035 );
buf ( n406164 , n389024 );
buf ( n406165 , n404236 );
nand ( n59039 , n406164 , n406165 );
buf ( n406167 , n59039 );
buf ( n406168 , n406167 );
nand ( n59042 , n59036 , n406168 );
buf ( n406170 , n59042 );
not ( n59044 , n406170 );
or ( n59045 , n59019 , n59044 );
buf ( n406173 , n406145 );
buf ( n406174 , n406170 );
nor ( n59048 , n406173 , n406174 );
buf ( n406176 , n59048 );
buf ( n406177 , n404610 );
buf ( n406178 , n57458 );
xor ( n59052 , n406177 , n406178 );
buf ( n406180 , n404658 );
xnor ( n59054 , n59052 , n406180 );
buf ( n406182 , n59054 );
or ( n59056 , n406176 , n406182 );
nand ( n59057 , n59045 , n59056 );
buf ( n406185 , n59057 );
buf ( n406186 , n395349 );
not ( n59060 , n406186 );
buf ( n406188 , n47863 );
not ( n59062 , n406188 );
buf ( n406190 , n38357 );
not ( n59064 , n406190 );
or ( n59065 , n59062 , n59064 );
buf ( n406193 , n391721 );
buf ( n406194 , n395312 );
nand ( n59068 , n406193 , n406194 );
buf ( n406196 , n59068 );
buf ( n406197 , n406196 );
nand ( n59071 , n59065 , n406197 );
buf ( n406199 , n59071 );
buf ( n406200 , n406199 );
not ( n59074 , n406200 );
or ( n59075 , n59060 , n59074 );
buf ( n406203 , n405683 );
buf ( n406204 , n395362 );
nand ( n59078 , n406203 , n406204 );
buf ( n406206 , n59078 );
buf ( n406207 , n406206 );
nand ( n59081 , n59075 , n406207 );
buf ( n406209 , n59081 );
buf ( n406210 , n406209 );
xor ( n59084 , n406185 , n406210 );
xor ( n59085 , n404528 , n404532 );
xor ( n59086 , n59085 , n404558 );
buf ( n406214 , n59086 );
buf ( n406215 , n406214 );
and ( n59089 , n59084 , n406215 );
and ( n59090 , n406185 , n406210 );
or ( n59091 , n59089 , n59090 );
buf ( n406219 , n59091 );
not ( n59093 , n406219 );
buf ( n406221 , n57296 );
buf ( n406222 , n404498 );
xor ( n59096 , n406221 , n406222 );
buf ( n406224 , n404562 );
xnor ( n59098 , n59096 , n406224 );
buf ( n406226 , n59098 );
nand ( n59100 , n59093 , n406226 );
not ( n59101 , n59100 );
xor ( n59102 , n404797 , n404815 );
xor ( n59103 , n59102 , n404876 );
buf ( n406231 , n59103 );
not ( n59105 , n406231 );
or ( n59106 , n59101 , n59105 );
buf ( n406234 , n406226 );
not ( n59108 , n406234 );
buf ( n406236 , n59108 );
nand ( n59110 , n406236 , n406219 );
nand ( n59111 , n59106 , n59110 );
and ( n59112 , n58997 , n59111 );
not ( n59113 , n58997 );
not ( n59114 , n59111 );
and ( n59115 , n59113 , n59114 );
nor ( n59116 , n59112 , n59115 );
xor ( n59117 , n57750 , n404944 );
xor ( n59118 , n59117 , n57800 );
and ( n59119 , n59116 , n59118 );
not ( n59120 , n59116 );
not ( n59121 , n59118 );
and ( n59122 , n59120 , n59121 );
nor ( n59123 , n59119 , n59122 );
buf ( n406251 , n59123 );
or ( n59125 , n406122 , n406251 );
xor ( n59126 , n406053 , n406079 );
xor ( n59127 , n59126 , n406101 );
buf ( n406255 , n59127 );
not ( n59129 , n58403 );
and ( n59130 , n59129 , n57875 );
not ( n59131 , n59129 );
and ( n59132 , n59131 , n57876 );
nor ( n59133 , n59130 , n59132 );
buf ( n406261 , n59133 );
buf ( n406262 , n405080 );
and ( n59136 , n406261 , n406262 );
not ( n59137 , n406261 );
buf ( n406265 , n405077 );
and ( n59139 , n59137 , n406265 );
nor ( n59140 , n59136 , n59139 );
buf ( n406268 , n59140 );
buf ( n406269 , n406268 );
not ( n59143 , n406269 );
buf ( n406271 , n59143 );
buf ( n406272 , n406271 );
not ( n59146 , n406272 );
not ( n59147 , n58779 );
not ( n59148 , n58573 );
not ( n59149 , n58570 );
or ( n59150 , n59148 , n59149 );
or ( n59151 , n58570 , n58573 );
nand ( n59152 , n59150 , n59151 );
not ( n59153 , n59152 );
or ( n59154 , n59147 , n59153 );
or ( n59155 , n59152 , n58779 );
nand ( n59156 , n59154 , n59155 );
buf ( n406284 , n59156 );
not ( n59158 , n406284 );
or ( n59159 , n59146 , n59158 );
buf ( n406287 , n45954 );
not ( n59161 , n406287 );
buf ( n406289 , n393369 );
not ( n59163 , n406289 );
buf ( n406291 , n390373 );
not ( n59165 , n406291 );
or ( n59166 , n59163 , n59165 );
buf ( n406294 , n36187 );
buf ( n406295 , n393381 );
nand ( n59169 , n406294 , n406295 );
buf ( n406297 , n59169 );
buf ( n406298 , n406297 );
nand ( n59172 , n59166 , n406298 );
buf ( n406300 , n59172 );
buf ( n406301 , n406300 );
not ( n59175 , n406301 );
or ( n59176 , n59161 , n59175 );
buf ( n406304 , n393369 );
not ( n59178 , n406304 );
buf ( n406306 , n42234 );
not ( n59180 , n406306 );
or ( n59181 , n59178 , n59180 );
buf ( n406309 , n42234 );
buf ( n406310 , n393369 );
or ( n59184 , n406309 , n406310 );
buf ( n406312 , n59184 );
buf ( n406313 , n406312 );
nand ( n59187 , n59181 , n406313 );
buf ( n406315 , n59187 );
buf ( n406316 , n406315 );
buf ( n406317 , n393825 );
nand ( n59191 , n406316 , n406317 );
buf ( n406319 , n59191 );
buf ( n406320 , n406319 );
nand ( n59194 , n59176 , n406320 );
buf ( n406322 , n59194 );
not ( n59196 , n405962 );
not ( n59197 , n58836 );
or ( n59198 , n59196 , n59197 );
buf ( n406326 , n405959 );
buf ( n406327 , n58832 );
nand ( n59201 , n406326 , n406327 );
buf ( n406329 , n59201 );
nand ( n59203 , n59198 , n406329 );
xor ( n59204 , n59203 , n58889 );
xor ( n59205 , n406322 , n59204 );
not ( n59206 , n34975 );
buf ( n406334 , n59206 );
not ( n59208 , n406334 );
buf ( n406336 , n383414 );
not ( n59210 , n406336 );
or ( n59211 , n59208 , n59210 );
buf ( n406339 , n38425 );
nand ( n59213 , n59211 , n406339 );
buf ( n406341 , n59213 );
buf ( n406342 , n406341 );
not ( n59216 , n406342 );
buf ( n406344 , n34975 );
not ( n59218 , n406344 );
buf ( n406346 , n383417 );
not ( n59220 , n406346 );
or ( n59221 , n59218 , n59220 );
buf ( n406349 , n358975 );
nand ( n59223 , n59221 , n406349 );
buf ( n406351 , n59223 );
buf ( n406352 , n406351 );
nand ( n59226 , n59216 , n406352 );
buf ( n406354 , n59226 );
not ( n59228 , n406354 );
xor ( n59229 , n405863 , n405888 );
xor ( n59230 , n59229 , n405917 );
buf ( n406358 , n59230 );
buf ( n406359 , n406358 );
not ( n59233 , n406359 );
buf ( n406361 , n59233 );
not ( n59235 , n406361 );
or ( n59236 , n59228 , n59235 );
buf ( n406364 , n405190 );
buf ( n406365 , n405265 );
xor ( n59239 , n406364 , n406365 );
buf ( n406367 , n59239 );
buf ( n406368 , n406367 );
not ( n59242 , n406368 );
buf ( n406370 , n405541 );
not ( n59244 , n406370 );
or ( n59245 , n59242 , n59244 );
buf ( n406373 , n405541 );
buf ( n406374 , n406367 );
or ( n59248 , n406373 , n406374 );
nand ( n59249 , n59245 , n59248 );
buf ( n406377 , n59249 );
buf ( n406378 , n406377 );
buf ( n406379 , n12471 );
not ( n59253 , n406379 );
buf ( n406381 , n53251 );
not ( n59255 , n406381 );
or ( n59256 , n59253 , n59255 );
buf ( n406384 , n405126 );
buf ( n406385 , n57505 );
nand ( n59259 , n406384 , n406385 );
buf ( n406387 , n59259 );
buf ( n406388 , n406387 );
nand ( n59262 , n59256 , n406388 );
buf ( n406390 , n59262 );
buf ( n406391 , n406390 );
not ( n59265 , n406391 );
buf ( n406393 , n390429 );
not ( n59267 , n406393 );
or ( n59268 , n59265 , n59267 );
buf ( n406396 , n405172 );
buf ( n406397 , n400143 );
nand ( n59271 , n406396 , n406397 );
buf ( n406399 , n59271 );
buf ( n406400 , n406399 );
nand ( n59274 , n59268 , n406400 );
buf ( n406402 , n59274 );
buf ( n406403 , n406402 );
xor ( n59277 , n406378 , n406403 );
buf ( n406405 , n47726 );
not ( n59279 , n406405 );
buf ( n406407 , n405909 );
not ( n59281 , n406407 );
or ( n59282 , n59279 , n59281 );
not ( n59283 , n388566 );
not ( n59284 , n405897 );
or ( n59285 , n59283 , n59284 );
buf ( n406413 , n402836 );
not ( n59287 , n406413 );
buf ( n406415 , n388154 );
nand ( n59289 , n59287 , n406415 );
buf ( n406417 , n59289 );
nand ( n59291 , n59285 , n406417 );
buf ( n406419 , n59291 );
buf ( n406420 , n50041 );
not ( n59294 , n406420 );
buf ( n406422 , n59294 );
buf ( n406423 , n406422 );
nand ( n59297 , n406419 , n406423 );
buf ( n406425 , n59297 );
buf ( n406426 , n406425 );
nand ( n59300 , n59282 , n406426 );
buf ( n406428 , n59300 );
buf ( n406429 , n406428 );
xor ( n59303 , n59277 , n406429 );
buf ( n406431 , n59303 );
not ( n59305 , n406431 );
buf ( n406433 , n405535 );
not ( n59307 , n406433 );
buf ( n406435 , n405280 );
buf ( n406436 , n405428 );
xor ( n59310 , n406435 , n406436 );
buf ( n406438 , n59310 );
buf ( n406439 , n406438 );
not ( n59313 , n406439 );
or ( n59314 , n59307 , n59313 );
buf ( n406442 , n406438 );
buf ( n406443 , n405535 );
or ( n59317 , n406442 , n406443 );
nand ( n59318 , n59314 , n59317 );
buf ( n406446 , n59318 );
buf ( n406447 , n406446 );
buf ( n406448 , n405529 );
not ( n59322 , n406448 );
buf ( n406450 , n405519 );
buf ( n406451 , n405443 );
and ( n59325 , n406450 , n406451 );
not ( n59326 , n406450 );
buf ( n406454 , n405440 );
and ( n59328 , n59326 , n406454 );
nor ( n59329 , n59325 , n59328 );
buf ( n406457 , n59329 );
buf ( n406458 , n406457 );
not ( n59332 , n406458 );
or ( n59333 , n59322 , n59332 );
buf ( n406461 , n406457 );
buf ( n406462 , n405529 );
or ( n59336 , n406461 , n406462 );
nand ( n59337 , n59333 , n59336 );
buf ( n406465 , n59337 );
buf ( n406466 , n406465 );
buf ( n406467 , n55984 );
buf ( n406468 , n55905 );
and ( n59342 , n406467 , n406468 );
buf ( n406470 , n58135 );
buf ( n406471 , n55895 );
and ( n59345 , n406470 , n406471 );
nor ( n59346 , n59342 , n59345 );
buf ( n406474 , n59346 );
buf ( n406475 , n406474 );
buf ( n406476 , n403120 );
or ( n59350 , n406475 , n406476 );
buf ( n406478 , n405452 );
buf ( n406479 , n403133 );
or ( n59353 , n406478 , n406479 );
nand ( n59354 , n59350 , n59353 );
buf ( n406482 , n59354 );
buf ( n406483 , n406482 );
buf ( n406484 , n58042 );
buf ( n406485 , n405215 );
and ( n59359 , n406484 , n406485 );
buf ( n406487 , n403088 );
buf ( n406488 , n58061 );
and ( n59362 , n406487 , n406488 );
nor ( n59363 , n59359 , n59362 );
buf ( n406491 , n59363 );
buf ( n406492 , n406491 );
buf ( n406493 , n403293 );
or ( n59367 , n406492 , n406493 );
buf ( n406495 , n405469 );
buf ( n406496 , n405476 );
or ( n59370 , n406495 , n406496 );
nand ( n59371 , n59367 , n59370 );
buf ( n406499 , n59371 );
buf ( n406500 , n406499 );
xor ( n59374 , n406483 , n406500 );
buf ( n406502 , n58166 );
buf ( n406503 , n403146 );
and ( n59377 , n406502 , n406503 );
buf ( n406505 , n58205 );
buf ( n406506 , n401695 );
and ( n59380 , n406505 , n406506 );
nor ( n59381 , n59377 , n59380 );
buf ( n406509 , n59381 );
buf ( n406510 , n406509 );
buf ( n406511 , n403158 );
or ( n59385 , n406510 , n406511 );
buf ( n406513 , n405340 );
buf ( n406514 , n403167 );
or ( n59388 , n406513 , n406514 );
nand ( n59389 , n59385 , n59388 );
buf ( n406517 , n59389 );
buf ( n406518 , n406517 );
and ( n59392 , n59374 , n406518 );
and ( n59393 , n406483 , n406500 );
or ( n59394 , n59392 , n59393 );
buf ( n406522 , n59394 );
buf ( n406523 , n405348 );
not ( n59397 , n406523 );
buf ( n406525 , n405361 );
not ( n59399 , n406525 );
buf ( n406527 , n405417 );
not ( n59401 , n406527 );
and ( n59402 , n59399 , n59401 );
buf ( n406530 , n405361 );
buf ( n406531 , n405417 );
and ( n59405 , n406530 , n406531 );
nor ( n59406 , n59402 , n59405 );
buf ( n406534 , n59406 );
buf ( n406535 , n406534 );
not ( n59409 , n406535 );
or ( n59410 , n59397 , n59409 );
buf ( n406538 , n406534 );
buf ( n406539 , n405348 );
or ( n59413 , n406538 , n406539 );
nand ( n59414 , n59410 , n59413 );
buf ( n406542 , n59414 );
xor ( n59416 , n406522 , n406542 );
xor ( n59417 , n405461 , n405481 );
xor ( n59418 , n59417 , n405515 );
buf ( n406546 , n59418 );
and ( n59420 , n59416 , n406546 );
and ( n59421 , n406522 , n406542 );
or ( n59422 , n59420 , n59421 );
buf ( n406550 , n59422 );
xor ( n59424 , n406466 , n406550 );
not ( n59425 , n53615 );
not ( n59426 , n54259 );
or ( n59427 , n59425 , n59426 );
not ( n59428 , n54262 );
nand ( n59429 , n59427 , n59428 );
not ( n59430 , n54264 );
nand ( n59431 , n59430 , n53641 );
nor ( n59432 , n59429 , n59431 );
not ( n59433 , n59432 );
nand ( n59434 , n59429 , n59431 );
nand ( n59435 , n59433 , n59434 );
buf ( n406563 , n59435 );
not ( n59437 , n406563 );
buf ( n406565 , n59437 );
buf ( n406566 , n406565 );
buf ( n406567 , n403083 );
or ( n59441 , n406566 , n406567 );
buf ( n406569 , n58352 );
not ( n59443 , n406569 );
buf ( n406571 , n59443 );
buf ( n406572 , n406571 );
buf ( n406573 , n403092 );
or ( n59447 , n406572 , n406573 );
nand ( n59448 , n59441 , n59447 );
buf ( n406576 , n59448 );
buf ( n406577 , n14083 );
buf ( n59451 , n997 );
buf ( n406579 , n59451 );
not ( n59453 , n406579 );
buf ( n406581 , n59453 );
buf ( n406582 , n406581 );
and ( n59456 , n406577 , n406582 );
not ( n59457 , n14083 );
buf ( n406585 , n59457 );
buf ( n406586 , n59451 );
and ( n59460 , n406585 , n406586 );
nor ( n59461 , n59456 , n59460 );
buf ( n406589 , n59461 );
not ( n59463 , n13091 );
and ( n59464 , n59463 , n406581 );
not ( n59465 , n59463 );
and ( n59466 , n59465 , n59451 );
or ( n59467 , n59464 , n59466 );
and ( n59468 , n406589 , n59467 );
nand ( n59469 , n59468 , n58223 );
buf ( n406597 , n59469 );
not ( n59471 , n59467 );
buf ( n406599 , n59471 );
buf ( n406600 , n58223 );
nand ( n59474 , n406599 , n406600 );
buf ( n406602 , n59474 );
buf ( n406603 , n406602 );
and ( n59477 , n406597 , n406603 );
buf ( n406605 , n59477 );
xor ( n59479 , n406576 , n406605 );
buf ( n406607 , n55846 );
buf ( n406608 , n405215 );
and ( n59482 , n406607 , n406608 );
buf ( n406610 , n403079 );
buf ( n406611 , n58061 );
and ( n59485 , n406610 , n406611 );
nor ( n59486 , n59482 , n59485 );
buf ( n406614 , n59486 );
buf ( n406615 , n406614 );
buf ( n406616 , n403293 );
or ( n59490 , n406615 , n406616 );
buf ( n406618 , n406491 );
buf ( n406619 , n405476 );
or ( n59493 , n406618 , n406619 );
nand ( n59494 , n59490 , n59493 );
buf ( n406622 , n59494 );
and ( n59496 , n59479 , n406622 );
and ( n59497 , n406576 , n406605 );
or ( n59498 , n59496 , n59497 );
buf ( n406626 , n59498 );
buf ( n406627 , n405499 );
buf ( n406628 , n405511 );
or ( n59502 , n406627 , n406628 );
buf ( n406630 , n405514 );
nand ( n59504 , n59502 , n406630 );
buf ( n406632 , n59504 );
buf ( n406633 , n406632 );
xor ( n59507 , n406626 , n406633 );
buf ( n406635 , n58178 );
buf ( n406636 , n55905 );
and ( n59510 , n406635 , n406636 );
buf ( n406638 , n405335 );
buf ( n406639 , n55895 );
and ( n59513 , n406638 , n406639 );
nor ( n59514 , n59510 , n59513 );
buf ( n406642 , n59514 );
buf ( n406643 , n406642 );
buf ( n406644 , n403120 );
or ( n59518 , n406643 , n406644 );
buf ( n406646 , n406474 );
buf ( n406647 , n403133 );
or ( n59521 , n406646 , n406647 );
nand ( n59522 , n59518 , n59521 );
buf ( n406650 , n59522 );
buf ( n406651 , n406650 );
buf ( n406652 , n54297 );
buf ( n406653 , n405391 );
and ( n59527 , n406652 , n406653 );
buf ( n406655 , n55919 );
buf ( n406656 , n405388 );
and ( n59530 , n406655 , n406656 );
nor ( n59531 , n59527 , n59530 );
buf ( n406659 , n59531 );
buf ( n406660 , n406659 );
buf ( n406661 , n405407 );
or ( n59535 , n406660 , n406661 );
buf ( n406663 , n405490 );
buf ( n406664 , n405384 );
or ( n59538 , n406663 , n406664 );
nand ( n59539 , n59535 , n59538 );
buf ( n406667 , n59539 );
buf ( n406668 , n406667 );
xor ( n59542 , n406651 , n406668 );
buf ( n406670 , n58200 );
buf ( n406671 , n403146 );
and ( n59545 , n406670 , n406671 );
buf ( n406673 , n58201 );
buf ( n406674 , n401695 );
and ( n59548 , n406673 , n406674 );
nor ( n59549 , n59545 , n59548 );
buf ( n406677 , n59549 );
buf ( n406678 , n406677 );
buf ( n406679 , n403158 );
or ( n59553 , n406678 , n406679 );
buf ( n406681 , n406509 );
buf ( n406682 , n403167 );
or ( n59556 , n406681 , n406682 );
nand ( n59557 , n59553 , n59556 );
buf ( n406685 , n59557 );
buf ( n406686 , n406685 );
and ( n59560 , n59542 , n406686 );
and ( n59561 , n406651 , n406668 );
or ( n59562 , n59560 , n59561 );
buf ( n406690 , n59562 );
buf ( n406691 , n406690 );
and ( n59565 , n59507 , n406691 );
and ( n59566 , n406626 , n406633 );
or ( n59567 , n59565 , n59566 );
buf ( n406695 , n59567 );
xor ( n59569 , n406522 , n406542 );
xor ( n59570 , n59569 , n406546 );
and ( n59571 , n406695 , n59570 );
buf ( n406699 , n58352 );
buf ( n406700 , n403146 );
and ( n59574 , n406699 , n406700 );
buf ( n406702 , n406571 );
buf ( n406703 , n401695 );
and ( n59577 , n406702 , n406703 );
nor ( n59578 , n59574 , n59577 );
buf ( n406706 , n59578 );
buf ( n406707 , n406706 );
not ( n59581 , n406707 );
buf ( n406709 , n59581 );
buf ( n406710 , n406709 );
buf ( n406711 , n401674 );
and ( n59585 , n406710 , n406711 );
buf ( n406713 , n406677 );
not ( n59587 , n406713 );
buf ( n406715 , n59587 );
buf ( n406716 , n406715 );
buf ( n406717 , n403164 );
and ( n59591 , n406716 , n406717 );
nor ( n59592 , n59585 , n59591 );
buf ( n406720 , n59592 );
buf ( n406721 , n406720 );
nand ( n59595 , n59428 , n53615 );
xnor ( n59596 , n59595 , n54259 );
buf ( n406724 , n59596 );
buf ( n406725 , n401626 );
and ( n59599 , n406724 , n406725 );
buf ( n406727 , n59435 );
buf ( n406728 , n401650 );
and ( n59602 , n406727 , n406728 );
nor ( n59603 , n59599 , n59602 );
buf ( n406731 , n59603 );
buf ( n406732 , n406731 );
nand ( n59606 , n406721 , n406732 );
buf ( n406734 , n59606 );
xor ( n59608 , n406576 , n406605 );
xor ( n59609 , n59608 , n406622 );
and ( n59610 , n406734 , n59609 );
buf ( n406738 , n58042 );
buf ( n406739 , n405391 );
and ( n59613 , n406738 , n406739 );
buf ( n406741 , n403088 );
buf ( n406742 , n405388 );
and ( n59616 , n406741 , n406742 );
nor ( n59617 , n59613 , n59616 );
buf ( n406745 , n59617 );
buf ( n406746 , n406745 );
buf ( n406747 , n405407 );
or ( n59621 , n406746 , n406747 );
buf ( n406749 , n406659 );
buf ( n406750 , n405384 );
or ( n59624 , n406749 , n406750 );
nand ( n59625 , n59621 , n59624 );
buf ( n406753 , n59625 );
buf ( n406754 , n54336 );
not ( n59628 , n59457 );
buf ( n406756 , n59628 );
and ( n59630 , n406754 , n406756 );
buf ( n406758 , n401699 );
buf ( n406759 , n59457 );
and ( n59633 , n406758 , n406759 );
nor ( n59634 , n59630 , n59633 );
buf ( n406762 , n59634 );
buf ( n406763 , n406762 );
not ( n59637 , n59468 );
buf ( n406765 , n59637 );
or ( n59639 , n406763 , n406765 );
buf ( n406767 , n406602 );
nand ( n59641 , n59639 , n406767 );
buf ( n406769 , n59641 );
xor ( n59643 , n406753 , n406769 );
buf ( n406771 , n55984 );
buf ( n406772 , n405215 );
and ( n59646 , n406771 , n406772 );
buf ( n406774 , n58135 );
buf ( n406775 , n58061 );
and ( n59649 , n406774 , n406775 );
nor ( n59650 , n59646 , n59649 );
buf ( n406778 , n59650 );
buf ( n406779 , n406778 );
buf ( n406780 , n403293 );
or ( n59654 , n406779 , n406780 );
buf ( n406782 , n406614 );
buf ( n406783 , n405476 );
or ( n59657 , n406782 , n406783 );
nand ( n59658 , n59654 , n59657 );
buf ( n406786 , n59658 );
and ( n59660 , n59643 , n406786 );
and ( n59661 , n406753 , n406769 );
or ( n59662 , n59660 , n59661 );
xor ( n59663 , n406576 , n406605 );
xor ( n59664 , n59663 , n406622 );
and ( n59665 , n59662 , n59664 );
and ( n59666 , n406734 , n59662 );
or ( n59667 , n59610 , n59665 , n59666 );
xor ( n59668 , n406483 , n406500 );
xor ( n59669 , n59668 , n406518 );
buf ( n406797 , n59669 );
xor ( n59671 , n59667 , n406797 );
xor ( n59672 , n406626 , n406633 );
xor ( n59673 , n59672 , n406691 );
buf ( n406801 , n59673 );
and ( n59675 , n59671 , n406801 );
and ( n59676 , n59667 , n406797 );
or ( n59677 , n59675 , n59676 );
xor ( n59678 , n406522 , n406542 );
xor ( n59679 , n59678 , n406546 );
and ( n59680 , n59677 , n59679 );
and ( n59681 , n406695 , n59677 );
or ( n59682 , n59571 , n59680 , n59681 );
buf ( n406810 , n59682 );
and ( n59684 , n59424 , n406810 );
and ( n59685 , n406466 , n406550 );
or ( n59686 , n59684 , n59685 );
buf ( n406814 , n59686 );
buf ( n406815 , n406814 );
xor ( n59689 , n406447 , n406815 );
buf ( n406817 , n24070 );
not ( n59691 , n406817 );
buf ( n406819 , n27234 );
buf ( n59693 , n406819 );
buf ( n406821 , n59693 );
buf ( n406822 , n406821 );
not ( n59696 , n406822 );
buf ( n406824 , n59696 );
buf ( n406825 , n406824 );
not ( n59699 , n406825 );
and ( n59700 , n59691 , n59699 );
buf ( n406828 , n53252 );
buf ( n406829 , n388227 );
and ( n59703 , n406828 , n406829 );
nor ( n59704 , n59700 , n59703 );
buf ( n406832 , n59704 );
not ( n59706 , n406832 );
buf ( n406834 , n59706 );
not ( n59708 , n406834 );
buf ( n406836 , n390429 );
not ( n59710 , n406836 );
or ( n59711 , n59708 , n59710 );
buf ( n406839 , n406390 );
buf ( n406840 , n42924 );
nand ( n59714 , n406839 , n406840 );
buf ( n406842 , n59714 );
buf ( n406843 , n406842 );
nand ( n59717 , n59711 , n406843 );
buf ( n406845 , n59717 );
buf ( n406846 , n406845 );
and ( n59720 , n59689 , n406846 );
and ( n59721 , n406447 , n406815 );
or ( n59722 , n59720 , n59721 );
buf ( n406850 , n59722 );
not ( n59724 , n406850 );
nand ( n59725 , n59305 , n59724 );
not ( n59726 , n59725 );
buf ( n406854 , n41711 );
not ( n59728 , n406854 );
buf ( n406856 , n24116 );
not ( n59730 , n406856 );
buf ( n406858 , n41194 );
not ( n59732 , n406858 );
or ( n59733 , n59730 , n59732 );
buf ( n406861 , n28250 );
buf ( n406862 , n24117 );
nand ( n59736 , n406861 , n406862 );
buf ( n406864 , n59736 );
buf ( n406865 , n406864 );
nand ( n59739 , n59733 , n406865 );
buf ( n406867 , n59739 );
buf ( n406868 , n406867 );
not ( n59742 , n406868 );
or ( n59743 , n59728 , n59742 );
buf ( n406871 , n24118 );
not ( n59745 , n406871 );
buf ( n406873 , n50317 );
not ( n59747 , n406873 );
or ( n59748 , n59745 , n59747 );
buf ( n406876 , n40818 );
buf ( n406877 , n24117 );
nand ( n59751 , n406876 , n406877 );
buf ( n406879 , n59751 );
buf ( n406880 , n406879 );
nand ( n59754 , n59748 , n406880 );
buf ( n406882 , n59754 );
buf ( n406883 , n406882 );
buf ( n406884 , n389162 );
nand ( n59758 , n406883 , n406884 );
buf ( n406886 , n59758 );
buf ( n406887 , n406886 );
nand ( n59761 , n59743 , n406887 );
buf ( n406889 , n59761 );
not ( n59763 , n406889 );
or ( n59764 , n59726 , n59763 );
nand ( n59765 , n406431 , n406850 );
nand ( n59766 , n59764 , n59765 );
nand ( n59767 , n59236 , n59766 );
buf ( n406895 , n59767 );
buf ( n406896 , n406354 );
not ( n59770 , n406896 );
buf ( n406898 , n406358 );
nand ( n59772 , n59770 , n406898 );
buf ( n406900 , n59772 );
buf ( n406901 , n406900 );
nand ( n59775 , n406895 , n406901 );
buf ( n406903 , n59775 );
buf ( n406904 , n406903 );
xor ( n59778 , n58876 , n406034 );
xnor ( n59779 , n59778 , n58856 );
buf ( n406907 , n59779 );
xor ( n59781 , n406904 , n406907 );
buf ( n406909 , n391164 );
and ( n59783 , n399274 , n395919 );
not ( n59784 , n399274 );
and ( n59785 , n59784 , n389589 );
or ( n59786 , n59783 , n59785 );
buf ( n406914 , n59786 );
not ( n59788 , n406914 );
buf ( n406916 , n59788 );
buf ( n406917 , n406916 );
or ( n59791 , n406909 , n406917 );
buf ( n406919 , n383403 );
buf ( n406920 , n400440 );
buf ( n406921 , n391183 );
and ( n59795 , n406920 , n406921 );
not ( n59796 , n406920 );
buf ( n406924 , n383423 );
and ( n59798 , n59796 , n406924 );
nor ( n59799 , n59795 , n59798 );
buf ( n406927 , n59799 );
buf ( n406928 , n406927 );
or ( n59802 , n406919 , n406928 );
nand ( n59803 , n59791 , n59802 );
buf ( n406931 , n59803 );
buf ( n406932 , n406931 );
and ( n59806 , n59781 , n406932 );
and ( n59807 , n406904 , n406907 );
or ( n59808 , n59806 , n59807 );
buf ( n406936 , n59808 );
and ( n59810 , n59205 , n406936 );
and ( n59811 , n406322 , n59204 );
or ( n59812 , n59810 , n59811 );
buf ( n406940 , n59812 );
nand ( n59814 , n59159 , n406940 );
buf ( n406942 , n59814 );
buf ( n406943 , n406942 );
buf ( n406944 , n59156 );
not ( n59818 , n406944 );
buf ( n406946 , n59818 );
buf ( n406947 , n406946 );
buf ( n406948 , n406268 );
nand ( n59822 , n406947 , n406948 );
buf ( n406950 , n59822 );
buf ( n406951 , n406950 );
nand ( n59825 , n406943 , n406951 );
buf ( n406953 , n59825 );
xor ( n59827 , n406255 , n406953 );
buf ( n406955 , n406219 );
buf ( n406956 , n406231 );
xor ( n59830 , n406955 , n406956 );
buf ( n406958 , n406236 );
xor ( n59832 , n59830 , n406958 );
buf ( n406960 , n59832 );
and ( n59834 , n59827 , n406960 );
and ( n59835 , n406255 , n406953 );
or ( n59836 , n59834 , n59835 );
buf ( n406964 , n59836 );
nand ( n59838 , n59125 , n406964 );
buf ( n406966 , n59838 );
buf ( n406967 , n406966 );
buf ( n406968 , n59123 );
buf ( n406969 , n406121 );
nand ( n59843 , n406968 , n406969 );
buf ( n406971 , n59843 );
buf ( n406972 , n406971 );
nand ( n59846 , n406967 , n406972 );
buf ( n406974 , n59846 );
buf ( n406975 , n406974 );
and ( n59849 , n58991 , n406975 );
and ( n59850 , n405651 , n406117 );
or ( n59851 , n59849 , n59850 );
buf ( n406979 , n59851 );
xor ( n59853 , n58490 , n406979 );
xor ( n59854 , n405661 , n405665 );
and ( n59855 , n59854 , n406114 );
and ( n59856 , n405661 , n405665 );
or ( n59857 , n59855 , n59856 );
buf ( n406985 , n59857 );
xor ( n59859 , n404450 , n404454 );
xor ( n59860 , n59859 , n404885 );
buf ( n406988 , n59860 );
xor ( n59862 , n406985 , n406988 );
not ( n59863 , n59118 );
not ( n59864 , n58997 );
and ( n59865 , n59863 , n59864 );
nand ( n59866 , n58997 , n59118 );
buf ( n59867 , n59111 );
and ( n59868 , n59866 , n59867 );
nor ( n59869 , n59865 , n59868 );
not ( n59870 , n59869 );
not ( n59871 , n59870 );
and ( n59872 , n404465 , n57708 );
not ( n59873 , n404465 );
not ( n59874 , n57708 );
and ( n59875 , n59873 , n59874 );
nor ( n59876 , n59872 , n59875 );
xnor ( n59877 , n59876 , n404461 );
not ( n59878 , n59877 );
not ( n59879 , n59878 );
or ( n59880 , n59871 , n59879 );
not ( n59881 , n59877 );
not ( n59882 , n59869 );
or ( n59883 , n59881 , n59882 );
not ( n59885 , n404939 );
or ( n59886 , C0 , n59885 );
buf ( n407013 , C1 );
nand ( n59891 , n59886 , n407013 );
not ( n59892 , n57754 );
and ( n59893 , n59891 , n59892 );
not ( n59894 , n59891 );
not ( n59895 , n57770 );
and ( n59896 , n59894 , n59895 );
nor ( n59897 , n59893 , n59896 );
not ( n59898 , n59897 );
not ( n59899 , n59898 );
buf ( n407023 , n403668 );
not ( n59901 , n407023 );
buf ( n407025 , n49938 );
not ( n59903 , n407025 );
or ( n59904 , n59901 , n59903 );
buf ( n407028 , n41359 );
buf ( n407029 , n397990 );
nand ( n59907 , n407028 , n407029 );
buf ( n407031 , n59907 );
buf ( n407032 , n407031 );
nand ( n59910 , n59904 , n407032 );
buf ( n407034 , n59910 );
buf ( n407035 , n407034 );
buf ( n407036 , n50579 );
and ( n59914 , n407035 , n407036 );
buf ( n407038 , n406071 );
buf ( n59916 , n51553 );
buf ( n407040 , n59916 );
and ( n59918 , n407038 , n407040 );
nor ( n59919 , n59914 , n59918 );
buf ( n407043 , n59919 );
buf ( n407044 , n407043 );
not ( n59922 , n407044 );
or ( n59945 , n59922 , C0 );
buf ( n407047 , n58551 );
buf ( n407048 , n43515 );
and ( n59948 , n407047 , n407048 );
buf ( n407050 , n391027 );
not ( n59950 , n407050 );
buf ( n407052 , n390651 );
not ( n59952 , n407052 );
or ( n59953 , n59950 , n59952 );
buf ( n407055 , n385983 );
buf ( n407056 , n391024 );
nand ( n59956 , n407055 , n407056 );
buf ( n407058 , n59956 );
buf ( n407059 , n407058 );
nand ( n59959 , n59953 , n407059 );
buf ( n407061 , n59959 );
buf ( n407062 , n407061 );
not ( n59962 , n407062 );
buf ( n407064 , n43537 );
nor ( n59964 , n59962 , n407064 );
buf ( n407066 , n59964 );
buf ( n407067 , n407066 );
nor ( n59967 , n59948 , n407067 );
buf ( n407069 , n59967 );
not ( n59969 , n407069 );
buf ( n407071 , n383014 );
not ( n59971 , n407071 );
buf ( n407073 , n402819 );
buf ( n407074 , n35435 );
and ( n59974 , n407073 , n407074 );
not ( n59975 , n407073 );
buf ( n59976 , n37402 );
buf ( n407078 , n59976 );
and ( n59978 , n59975 , n407078 );
nor ( n59979 , n59974 , n59978 );
buf ( n407081 , n59979 );
buf ( n407082 , n407081 );
not ( n59982 , n407082 );
and ( n59983 , n59971 , n59982 );
buf ( n407085 , n404861 );
not ( n59985 , n407085 );
buf ( n407087 , n386307 );
nor ( n59987 , n59985 , n407087 );
buf ( n407089 , n59987 );
buf ( n407090 , n407089 );
nor ( n59990 , n59983 , n407090 );
buf ( n407092 , n59990 );
not ( n59992 , n407092 );
or ( n59993 , n59969 , n59992 );
xor ( n59994 , n405052 , n405071 );
xnor ( n59995 , n59994 , n57888 );
nand ( n59996 , n59993 , n59995 );
buf ( n407098 , n59996 );
buf ( n407099 , n407069 );
not ( n59999 , n407099 );
buf ( n407101 , n407092 );
not ( n60001 , n407101 );
buf ( n407103 , n60001 );
buf ( n407104 , n407103 );
nand ( n60004 , n59999 , n407104 );
buf ( n407106 , n60004 );
buf ( n407107 , n407106 );
nand ( n60007 , n407098 , n407107 );
buf ( n407109 , n60007 );
buf ( n407110 , n407109 );
nand ( n60010 , n59945 , n407110 );
buf ( n407112 , n60010 );
buf ( n407113 , n407112 );
buf ( n407114 , n407043 );
not ( n60015 , n407114 );
buf ( n407116 , n60015 );
buf ( n407117 , C1 );
buf ( n407118 , n407117 );
nand ( n60021 , n407113 , n407118 );
buf ( n407120 , n60021 );
not ( n60023 , n407120 );
or ( n60024 , n59899 , n60023 );
buf ( n407123 , n57632 );
not ( n60026 , n407123 );
buf ( n407125 , n393409 );
not ( n60028 , n407125 );
and ( n60029 , n60026 , n60028 );
buf ( n407128 , n406300 );
buf ( n407129 , n393825 );
and ( n60032 , n407128 , n407129 );
nor ( n60033 , n60029 , n60032 );
buf ( n407132 , n60033 );
buf ( n60035 , n407132 );
buf ( n407134 , n60035 );
not ( n60037 , n407134 );
and ( n60038 , n57662 , n57665 );
not ( n60039 , n57662 );
and ( n60040 , n60039 , n57666 );
nor ( n60041 , n60038 , n60040 );
and ( n60042 , n60041 , n404873 );
not ( n60043 , n60041 );
buf ( n407142 , n404873 );
not ( n60045 , n407142 );
buf ( n407144 , n60045 );
and ( n60047 , n60043 , n407144 );
nor ( n60048 , n60042 , n60047 );
buf ( n407147 , n60048 );
not ( n60050 , n407147 );
or ( n60051 , n60037 , n60050 );
buf ( n407150 , n383476 );
buf ( n407151 , n406927 );
or ( n60054 , n407150 , n407151 );
buf ( n407153 , n404828 );
not ( n60056 , n407153 );
buf ( n407155 , n60056 );
buf ( n407156 , n407155 );
buf ( n407157 , n383403 );
or ( n60060 , n407156 , n407157 );
nand ( n60061 , n60054 , n60060 );
buf ( n407160 , n60061 );
buf ( n407161 , n407160 );
not ( n60064 , n407161 );
xor ( n60065 , n57964 , n58400 );
not ( n60066 , n60065 );
not ( n60067 , n60066 );
not ( n60068 , n57944 );
or ( n60069 , n60067 , n60068 );
not ( n60070 , n57944 );
nand ( n60071 , n60070 , n60065 );
nand ( n60072 , n60069 , n60071 );
buf ( n407171 , n60072 );
not ( n60074 , n407171 );
or ( n60075 , n60064 , n60074 );
or ( n60076 , n407160 , n60072 );
buf ( n407175 , n405547 );
not ( n60078 , n407175 );
buf ( n407177 , n58033 );
not ( n60080 , n407177 );
and ( n60081 , n60078 , n60080 );
buf ( n407180 , n405547 );
buf ( n407181 , n58033 );
and ( n60084 , n407180 , n407181 );
nor ( n60085 , n60081 , n60084 );
buf ( n407184 , n60085 );
buf ( n407185 , n407184 );
not ( n60088 , n407185 );
buf ( n407187 , n405179 );
not ( n60090 , n407187 );
or ( n60091 , n60088 , n60090 );
buf ( n407190 , n405179 );
buf ( n407191 , n407184 );
or ( n60094 , n407190 , n407191 );
nand ( n60095 , n60091 , n60094 );
buf ( n407194 , n60095 );
buf ( n407195 , n407194 );
not ( n60098 , n46056 );
buf ( n407197 , n42073 );
not ( n60100 , n407197 );
buf ( n407199 , n388965 );
not ( n60102 , n407199 );
or ( n60103 , n60100 , n60102 );
buf ( n407202 , n388962 );
buf ( n407203 , n42074 );
nand ( n60106 , n407202 , n407203 );
buf ( n407205 , n60106 );
buf ( n407206 , n407205 );
nand ( n60109 , n60103 , n407206 );
buf ( n407208 , n60109 );
not ( n60111 , n407208 );
or ( n60112 , n60098 , n60111 );
nand ( n60113 , n51692 , n58610 );
nand ( n60114 , n60112 , n60113 );
buf ( n407213 , n60114 );
xor ( n60116 , n407195 , n407213 );
not ( n60117 , n388830 );
not ( n60118 , n405792 );
or ( n60119 , n60117 , n60118 );
not ( n60120 , n41342 );
not ( n60121 , n388373 );
or ( n60122 , n60120 , n60121 );
nand ( n60123 , n388370 , n45897 );
nand ( n60124 , n60122 , n60123 );
nand ( n60125 , n60124 , n388872 );
nand ( n60126 , n60119 , n60125 );
buf ( n407225 , n60126 );
and ( n60128 , n60116 , n407225 );
and ( n60129 , n407195 , n407213 );
or ( n60130 , n60128 , n60129 );
buf ( n407229 , n60130 );
buf ( n407230 , n407229 );
buf ( n407231 , n57940 );
buf ( n407232 , n383937 );
or ( n60135 , n407231 , n407232 );
buf ( n407234 , n392884 );
buf ( n407235 , n50992 );
and ( n60138 , n407234 , n407235 );
not ( n60139 , n407234 );
buf ( n407238 , n36395 );
and ( n60141 , n60139 , n407238 );
nor ( n60142 , n60138 , n60141 );
buf ( n407241 , n60142 );
nand ( n60144 , n407241 , n383937 , n56842 );
buf ( n407243 , n60144 );
nand ( n60146 , n60135 , n407243 );
buf ( n407245 , n60146 );
buf ( n407246 , n407245 );
xor ( n60149 , n407230 , n407246 );
buf ( n407248 , n394817 );
not ( n60151 , n407248 );
buf ( n407250 , n36809 );
not ( n60153 , n407250 );
or ( n60154 , n60151 , n60153 );
nand ( n60155 , n36810 , n394814 );
buf ( n407254 , n60155 );
nand ( n60157 , n60154 , n407254 );
buf ( n407256 , n60157 );
buf ( n407257 , n407256 );
not ( n407258 , n407257 );
buf ( n407259 , n40858 );
not ( n60162 , n407259 );
or ( n60163 , n407258 , n60162 );
buf ( n407262 , n40901 );
buf ( n407263 , n57886 );
nand ( n60166 , n407262 , n407263 );
buf ( n407265 , n60166 );
buf ( n407266 , n407265 );
nand ( n60169 , n60163 , n407266 );
buf ( n407268 , n60169 );
buf ( n407269 , n407268 );
and ( n60172 , n60149 , n407269 );
and ( n60173 , n407230 , n407246 );
or ( n60174 , n60172 , n60173 );
buf ( n407273 , n60174 );
nand ( n60176 , n60076 , n407273 );
buf ( n407275 , n60176 );
nand ( n60178 , n60075 , n407275 );
buf ( n407277 , n60178 );
buf ( n407278 , n407277 );
nand ( n60181 , n60051 , n407278 );
buf ( n407280 , n60181 );
not ( n60183 , n407280 );
not ( n60184 , n60048 );
buf ( n407283 , n60184 );
not ( n60186 , n407132 );
buf ( n407285 , n60186 );
nand ( n60188 , n407283 , n407285 );
buf ( n407287 , n60188 );
not ( n60190 , n407287 );
or ( n60191 , n60183 , n60190 );
not ( n60192 , n407120 );
nand ( n60193 , n60192 , n59897 );
nand ( n60194 , n60191 , n60193 );
nand ( n60195 , n60024 , n60194 );
buf ( n407294 , n404988 );
not ( n60197 , n407294 );
buf ( n407296 , n404979 );
not ( n60199 , n407296 );
or ( n60200 , n60197 , n60199 );
buf ( n407299 , n57825 );
buf ( n407300 , n404983 );
nand ( n60203 , n407299 , n407300 );
buf ( n407302 , n60203 );
buf ( n407303 , n407302 );
nand ( n60206 , n60200 , n407303 );
buf ( n407305 , n60206 );
buf ( n407306 , n407305 );
buf ( n407307 , n405568 );
and ( n60210 , n407306 , n407307 );
not ( n60211 , n407306 );
buf ( n407310 , n405568 );
not ( n60213 , n407310 );
buf ( n407312 , n60213 );
buf ( n407313 , n407312 );
and ( n60216 , n60211 , n407313 );
nor ( n60217 , n60210 , n60216 );
buf ( n407316 , n60217 );
xor ( n60219 , n60195 , n407316 );
xor ( n60220 , n405690 , n406048 );
xnor ( n60221 , n60220 , n58783 );
buf ( n407320 , n60221 );
not ( n60223 , n407320 );
buf ( n407322 , n60223 );
not ( n60225 , n407322 );
xor ( n60226 , n405016 , n405559 );
xor ( n60227 , n60226 , n405564 );
buf ( n407326 , n60227 );
not ( n60229 , n407326 );
or ( n60230 , n60225 , n60229 );
buf ( n407329 , n407326 );
not ( n60232 , n407329 );
buf ( n407331 , n60232 );
not ( n60234 , n407331 );
not ( n60235 , n60221 );
or ( n60236 , n60234 , n60235 );
buf ( n407335 , C1 );
buf ( n407336 , n395362 );
not ( n60258 , n407336 );
buf ( n407338 , n406199 );
not ( n60260 , n407338 );
or ( n60261 , n60258 , n60260 );
buf ( n407341 , n395349 );
and ( n60263 , n47863 , n389525 );
not ( n60264 , n47863 );
and ( n60265 , n60264 , n37173 );
or ( n60266 , n60263 , n60265 );
buf ( n407346 , n60266 );
nand ( n60268 , n407341 , n407346 );
buf ( n407348 , n60268 );
buf ( n407349 , n407348 );
nand ( n60271 , n60261 , n407349 );
buf ( n407351 , n60271 );
buf ( n407352 , n407351 );
xor ( n60274 , n58602 , n58654 );
xor ( n60275 , n60274 , n58776 );
buf ( n407355 , n60275 );
xor ( n60277 , n407352 , n407355 );
xor ( n60278 , n405773 , n58646 );
xor ( n60279 , n60278 , n405803 );
buf ( n407359 , n60279 );
buf ( n407360 , n389744 );
not ( n60282 , n407360 );
buf ( n407362 , n55055 );
not ( n60284 , n407362 );
buf ( n407364 , n382994 );
not ( n60286 , n407364 );
or ( n60287 , n60284 , n60286 );
buf ( n407367 , n389997 );
buf ( n407368 , n55054 );
nand ( n60290 , n407367 , n407368 );
buf ( n407370 , n60290 );
buf ( n407371 , n407370 );
nand ( n60293 , n60287 , n407371 );
buf ( n407373 , n60293 );
buf ( n407374 , n407373 );
not ( n60296 , n407374 );
or ( n60297 , n60282 , n60296 );
buf ( n407377 , n379463 );
buf ( n407378 , n406158 );
nand ( n60300 , n407377 , n407378 );
buf ( n407380 , n60300 );
buf ( n407381 , n407380 );
nand ( n60303 , n60297 , n407381 );
buf ( n407383 , n60303 );
buf ( n407384 , n407383 );
xor ( n60306 , n407359 , n407384 );
nand ( n60307 , n58673 , n58684 , n405921 );
not ( n60308 , n405921 );
nand ( n60309 , n58684 , n58674 , n60308 );
nand ( n60310 , n58685 , n58674 , n405921 );
nand ( n60311 , n58685 , n58673 , n60308 );
nand ( n60312 , n60307 , n60309 , n60310 , n60311 );
buf ( n407392 , n60312 );
and ( n60314 , n60306 , n407392 );
and ( n60315 , n407359 , n407384 );
or ( n60316 , n60314 , n60315 );
buf ( n407396 , n60316 );
buf ( n407397 , n407396 );
and ( n60319 , n60277 , n407397 );
and ( n60320 , n407352 , n407355 );
or ( n60321 , n60319 , n60320 );
buf ( n407401 , n60321 );
buf ( n407402 , n407401 );
not ( n60324 , n407402 );
buf ( n407404 , n60324 );
not ( n60326 , n407404 );
or ( n60327 , C0 , n60326 );
buf ( n407407 , n406137 );
not ( n60329 , n407407 );
buf ( n407409 , n388071 );
not ( n60331 , n407409 );
and ( n60332 , n60329 , n60331 );
buf ( n407412 , n388102 );
not ( n60334 , n407412 );
buf ( n407414 , n389805 );
not ( n60336 , n407414 );
or ( n60337 , n60334 , n60336 );
buf ( n407417 , n391486 );
buf ( n407418 , n388105 );
nand ( n60340 , n407417 , n407418 );
buf ( n407420 , n60340 );
buf ( n407421 , n407420 );
nand ( n60343 , n60337 , n407421 );
buf ( n407423 , n60343 );
buf ( n407424 , n407423 );
buf ( n407425 , n43286 );
and ( n60347 , n407424 , n407425 );
nor ( n60348 , n60332 , n60347 );
buf ( n407428 , n60348 );
nand ( n60350 , n390635 , n358975 );
or ( n60351 , n407428 , n60350 );
buf ( n407431 , n60350 );
not ( n60353 , n407431 );
buf ( n407433 , n407428 );
not ( n60355 , n407433 );
or ( n60356 , n60353 , n60355 );
xor ( n60357 , n406378 , n406403 );
and ( n60358 , n60357 , n406429 );
and ( n60359 , n406378 , n406403 );
or ( n60360 , n60358 , n60359 );
buf ( n407440 , n60360 );
buf ( n407441 , n407440 );
buf ( n407442 , n40990 );
not ( n60364 , n407442 );
buf ( n407444 , n51648 );
not ( n60366 , n407444 );
or ( n60367 , n60364 , n60366 );
buf ( n407447 , n22982 );
buf ( n407448 , n390460 );
nand ( n60370 , n407447 , n407448 );
buf ( n407450 , n60370 );
buf ( n407451 , n407450 );
nand ( n60373 , n60367 , n407451 );
buf ( n407453 , n60373 );
buf ( n407454 , n407453 );
not ( n60376 , n407454 );
buf ( n407456 , n397102 );
not ( n60378 , n407456 );
or ( n60379 , n60376 , n60378 );
buf ( n407459 , n405875 );
buf ( n407460 , n393127 );
nand ( n60382 , n407459 , n407460 );
buf ( n407462 , n60382 );
buf ( n407463 , n407462 );
nand ( n60385 , n60379 , n407463 );
buf ( n407465 , n60385 );
not ( n60387 , n407465 );
not ( n60388 , n396622 );
buf ( n407468 , n388998 );
not ( n60390 , n407468 );
buf ( n407470 , n398298 );
not ( n60392 , n407470 );
or ( n60393 , n60390 , n60392 );
buf ( n407473 , n24049 );
buf ( n407474 , n388215 );
nand ( n60396 , n407473 , n407474 );
buf ( n407476 , n60396 );
buf ( n407477 , n407476 );
nand ( n60399 , n60393 , n407477 );
buf ( n407479 , n60399 );
not ( n60401 , n407479 );
or ( n60402 , n60388 , n60401 );
nand ( n60403 , n55831 , n405850 );
nand ( n60404 , n60402 , n60403 );
not ( n60405 , n60404 );
nand ( n60406 , n60387 , n60405 );
not ( n60407 , n60406 );
not ( n60408 , n388872 );
buf ( n407488 , n41342 );
not ( n60410 , n407488 );
buf ( n407490 , n394330 );
not ( n60412 , n407490 );
or ( n60413 , n60410 , n60412 );
buf ( n407493 , n388643 );
buf ( n407494 , n45897 );
nand ( n60416 , n407493 , n407494 );
buf ( n407496 , n60416 );
buf ( n407497 , n407496 );
nand ( n60419 , n60413 , n407497 );
buf ( n407499 , n60419 );
not ( n60421 , n407499 );
or ( n60422 , n60408 , n60421 );
buf ( n407502 , n60124 );
buf ( n407503 , n388830 );
nand ( n60425 , n407502 , n407503 );
buf ( n407505 , n60425 );
nand ( n60427 , n60422 , n407505 );
not ( n60428 , n60427 );
or ( n60429 , n60407 , n60428 );
nand ( n60430 , n60404 , n407465 );
nand ( n60431 , n60429 , n60430 );
buf ( n407511 , n60431 );
xor ( n60433 , n407441 , n407511 );
and ( n60434 , n389341 , n390548 );
not ( n60435 , n389341 );
and ( n60436 , n60435 , n393562 );
or ( n60437 , n60434 , n60436 );
not ( n60438 , n60437 );
not ( n60439 , n390536 );
or ( n60440 , n60438 , n60439 );
not ( n60441 , n37313 );
nand ( n60442 , n60441 , n58680 );
nand ( n60443 , n60440 , n60442 );
buf ( n407523 , n60443 );
and ( n60445 , n60433 , n407523 );
and ( n60446 , n407441 , n407511 );
or ( n60447 , n60445 , n60446 );
buf ( n407527 , n60447 );
buf ( n407528 , n407527 );
nand ( n60450 , n60356 , n407528 );
buf ( n407530 , n60450 );
nand ( n60452 , n60351 , n407530 );
buf ( n407532 , n60452 );
buf ( n407533 , n392740 );
not ( n60455 , n407533 );
buf ( n407535 , n58566 );
not ( n60457 , n407535 );
or ( n60458 , n60455 , n60457 );
buf ( n407538 , n392247 );
not ( n60460 , n407538 );
buf ( n407540 , n390810 );
not ( n60462 , n407540 );
or ( n60463 , n60460 , n60462 );
buf ( n407543 , n38472 );
buf ( n407544 , n392244 );
nand ( n60466 , n407543 , n407544 );
buf ( n407546 , n60466 );
buf ( n407547 , n407546 );
nand ( n60469 , n60463 , n407547 );
buf ( n407549 , n60469 );
buf ( n407550 , n407549 );
buf ( n407551 , n45260 );
nand ( n60473 , n407550 , n407551 );
buf ( n407553 , n60473 );
buf ( n407554 , n407553 );
nand ( n60476 , n60458 , n407554 );
buf ( n407556 , n60476 );
buf ( n407557 , n407556 );
xor ( n60479 , n407532 , n407557 );
and ( n60480 , n397498 , n391129 );
not ( n60481 , n397498 );
and ( n60482 , n60481 , n395885 );
or ( n60483 , n60480 , n60482 );
buf ( n407563 , n60483 );
not ( n60485 , n407563 );
buf ( n407565 , n393595 );
not ( n60487 , n407565 );
or ( n60488 , n60485 , n60487 );
buf ( n407568 , n405976 );
buf ( n407569 , n393602 );
nand ( n60491 , n407568 , n407569 );
buf ( n407571 , n60491 );
buf ( n407572 , n407571 );
nand ( n60494 , n60488 , n407572 );
buf ( n407574 , n60494 );
buf ( n407575 , n407574 );
not ( n60497 , n407575 );
buf ( n407577 , n43727 );
not ( n60499 , n407577 );
not ( n60500 , n391027 );
not ( n60501 , n44423 );
or ( n60502 , n60500 , n60501 );
not ( n60503 , n41896 );
nand ( n60504 , n60503 , n391024 );
nand ( n60505 , n60502 , n60504 );
buf ( n407585 , n60505 );
not ( n60507 , n407585 );
or ( n60508 , n60499 , n60507 );
buf ( n407588 , n407061 );
buf ( n407589 , n43515 );
nand ( n60511 , n407588 , n407589 );
buf ( n407591 , n60511 );
buf ( n407592 , n407591 );
nand ( n60514 , n60508 , n407592 );
buf ( n407594 , n60514 );
buf ( n407595 , n407594 );
not ( n60517 , n407595 );
or ( n60518 , n60497 , n60517 );
buf ( n407598 , n407574 );
not ( n60520 , n407598 );
buf ( n407600 , n60520 );
buf ( n407601 , n407600 );
not ( n60523 , n407601 );
buf ( n407603 , n407594 );
not ( n60525 , n407603 );
buf ( n407605 , n60525 );
buf ( n407606 , n407605 );
not ( n60528 , n407606 );
or ( n60529 , n60523 , n60528 );
buf ( n407609 , n389162 );
not ( n60531 , n407609 );
buf ( n407611 , n405822 );
not ( n60533 , n407611 );
or ( n60534 , n60531 , n60533 );
buf ( n407614 , n406882 );
buf ( n407615 , n57569 );
nand ( n60537 , n407614 , n407615 );
buf ( n407617 , n60537 );
buf ( n407618 , n407617 );
nand ( n60540 , n60534 , n407618 );
buf ( n407620 , n60540 );
buf ( n407621 , n392611 );
not ( n60543 , n407621 );
buf ( n407623 , n388299 );
not ( n60545 , n407623 );
or ( n60546 , n60543 , n60545 );
buf ( n407626 , n388263 );
buf ( n407627 , n392620 );
nand ( n60549 , n407626 , n407627 );
buf ( n407629 , n60549 );
buf ( n407630 , n407629 );
nand ( n60552 , n60546 , n407630 );
buf ( n407632 , n60552 );
buf ( n407633 , n407632 );
not ( n60555 , n407633 );
buf ( n407635 , n383891 );
not ( n60557 , n407635 );
or ( n60558 , n60555 , n60557 );
buf ( n407638 , n406019 );
buf ( n407639 , n388629 );
nand ( n60561 , n407638 , n407639 );
buf ( n407641 , n60561 );
buf ( n407642 , n407641 );
nand ( n60564 , n60558 , n407642 );
buf ( n407644 , n60564 );
or ( n60566 , n407620 , n407644 );
buf ( n407646 , n388809 );
not ( n60568 , n407646 );
buf ( n407648 , n406005 );
not ( n60570 , n407648 );
or ( n60571 , n60568 , n60570 );
buf ( n407651 , n405736 );
not ( n60573 , n407651 );
buf ( n407653 , n40759 );
not ( n60575 , n407653 );
or ( n60576 , n60573 , n60575 );
buf ( n407656 , n40758 );
buf ( n407657 , n388757 );
nand ( n60579 , n407656 , n407657 );
buf ( n407659 , n60579 );
buf ( n407660 , n407659 );
nand ( n60582 , n60576 , n407660 );
buf ( n407662 , n60582 );
buf ( n407663 , n407662 );
buf ( n407664 , n388746 );
nand ( n60586 , n407663 , n407664 );
buf ( n407666 , n60586 );
buf ( n407667 , n407666 );
nand ( n60589 , n60571 , n407667 );
buf ( n407669 , n60589 );
nand ( n60591 , n60566 , n407669 );
buf ( n407671 , n60591 );
buf ( n407672 , n407644 );
buf ( n407673 , n407620 );
nand ( n60595 , n407672 , n407673 );
buf ( n407675 , n60595 );
buf ( n407676 , n407675 );
nand ( n60598 , n407671 , n407676 );
buf ( n407678 , n60598 );
buf ( n407679 , n407678 );
nand ( n60601 , n60529 , n407679 );
buf ( n407681 , n60601 );
buf ( n407682 , n407681 );
nand ( n60604 , n60518 , n407682 );
buf ( n407684 , n60604 );
buf ( n407685 , n407684 );
and ( n60607 , n60479 , n407685 );
and ( n60608 , n407532 , n407557 );
or ( n60609 , n60607 , n60608 );
buf ( n407689 , n60609 );
buf ( n60611 , n407689 );
nand ( n407691 , n60327 , n60611 );
buf ( n407692 , C1 );
nand ( n60617 , n407691 , n407692 );
nand ( n60618 , n60236 , n60617 );
nand ( n60619 , n60230 , n60618 );
and ( n60620 , n60219 , n60619 );
and ( n60621 , n60195 , n407316 );
or ( n60622 , n60620 , n60621 );
nand ( n60623 , n59883 , n60622 );
nand ( n60624 , n59880 , n60623 );
xor ( n60625 , n59862 , n60624 );
xor ( n60626 , n59853 , n60625 );
not ( n60627 , n60626 );
not ( n60628 , n59870 );
not ( n60629 , n59878 );
and ( n60630 , n60628 , n60629 );
and ( n60631 , n59870 , n59878 );
nor ( n60632 , n60630 , n60631 );
buf ( n407709 , n60622 );
not ( n60634 , n407709 );
buf ( n407711 , n60634 );
not ( n60636 , n407711 );
and ( n60637 , n60632 , n60636 );
not ( n60638 , n60632 );
and ( n60639 , n60638 , n407711 );
nor ( n60640 , n60637 , n60639 );
buf ( n407717 , n60640 );
buf ( n407718 , n407280 );
buf ( n407719 , n407287 );
nand ( n60644 , n407718 , n407719 );
buf ( n407721 , n60644 );
buf ( n407722 , n407721 );
not ( n60647 , n407722 );
buf ( n407724 , n407120 );
not ( n60649 , n407724 );
buf ( n407726 , n60649 );
buf ( n407727 , n407726 );
not ( n60652 , n407727 );
or ( n60653 , n60647 , n60652 );
buf ( n407730 , n407721 );
not ( n60655 , n407730 );
buf ( n407732 , n60655 );
buf ( n407733 , n407732 );
buf ( n407734 , n407120 );
nand ( n60659 , n407733 , n407734 );
buf ( n407736 , n60659 );
buf ( n407737 , n407736 );
nand ( n60662 , n60653 , n407737 );
buf ( n407739 , n60662 );
not ( n60664 , n59898 );
and ( n60665 , n407739 , n60664 );
not ( n60666 , n407739 );
and ( n60667 , n60666 , n59898 );
nor ( n60668 , n60665 , n60667 );
buf ( n407745 , n60668 );
not ( n60670 , n407745 );
xor ( n60671 , n407160 , n60072 );
or ( n60672 , n407273 , n60671 );
nand ( n60673 , n60671 , n407273 );
nand ( n60674 , n60672 , n60673 );
buf ( n407751 , n60674 );
buf ( n407752 , n406145 );
buf ( n407753 , n406182 );
xor ( n60678 , n407752 , n407753 );
buf ( n407755 , n60678 );
xnor ( n60680 , n406170 , n407755 );
buf ( n407757 , n60680 );
not ( n60682 , n407757 );
buf ( n407759 , n60682 );
buf ( n407760 , n407759 );
nand ( n60685 , n407751 , n407760 );
buf ( n407762 , n60685 );
xor ( n60687 , n407230 , n407246 );
xor ( n60688 , n60687 , n407269 );
buf ( n407765 , n60688 );
buf ( n407766 , n407765 );
buf ( n407767 , n45260 );
not ( n60692 , n407767 );
buf ( n407769 , n392244 );
not ( n60694 , n407769 );
buf ( n407771 , n390178 );
not ( n60696 , n407771 );
or ( n60697 , n60694 , n60696 );
buf ( n407774 , n58545 );
not ( n60699 , n407774 );
buf ( n407776 , n399986 );
nand ( n60701 , n60699 , n407776 );
buf ( n407778 , n60701 );
buf ( n407779 , n407778 );
nand ( n60704 , n60697 , n407779 );
buf ( n407781 , n60704 );
buf ( n407782 , n407781 );
not ( n60707 , n407782 );
or ( n60708 , n60692 , n60707 );
buf ( n407785 , n407549 );
buf ( n407786 , n392740 );
nand ( n60711 , n407785 , n407786 );
buf ( n407788 , n60711 );
buf ( n407789 , n407788 );
nand ( n60714 , n60708 , n407789 );
buf ( n407791 , n60714 );
buf ( n407792 , n407791 );
xor ( n60717 , n407766 , n407792 );
buf ( n407794 , n390362 );
not ( n60719 , n407794 );
buf ( n407796 , n407423 );
not ( n60721 , n407796 );
or ( n60722 , n60719 , n60721 );
buf ( n407799 , n388102 );
not ( n60724 , n407799 );
buf ( n407801 , n388919 );
not ( n60726 , n407801 );
or ( n60727 , n60724 , n60726 );
buf ( n407804 , n396537 );
buf ( n407805 , n388105 );
nand ( n60730 , n407804 , n407805 );
buf ( n407807 , n60730 );
buf ( n407808 , n407807 );
nand ( n60733 , n60727 , n407808 );
buf ( n407810 , n60733 );
buf ( n407811 , n407810 );
buf ( n407812 , n43286 );
nand ( n60737 , n407811 , n407812 );
buf ( n407814 , n60737 );
buf ( n407815 , n407814 );
nand ( n60740 , n60722 , n407815 );
buf ( n407817 , n60740 );
buf ( n407818 , n407817 );
and ( n60743 , n358975 , n385975 );
not ( n60744 , n358975 );
and ( n60745 , n60744 , n379574 );
nor ( n60746 , n60743 , n60745 );
buf ( n407823 , n60746 );
not ( n60748 , n407823 );
buf ( n407825 , n389015 );
not ( n60750 , n407825 );
or ( n60751 , n60748 , n60750 );
buf ( n407828 , n389328 );
buf ( n407829 , n407373 );
nand ( n60754 , n407828 , n407829 );
buf ( n407831 , n60754 );
buf ( n407832 , n407831 );
nand ( n60757 , n60751 , n407832 );
buf ( n407834 , n60757 );
buf ( n407835 , n407834 );
xor ( n60760 , n407818 , n407835 );
buf ( n407837 , n389359 );
not ( n60762 , n407837 );
buf ( n407839 , n388965 );
not ( n60764 , n407839 );
or ( n60765 , n60762 , n60764 );
buf ( n407842 , n388962 );
buf ( n407843 , n389356 );
nand ( n60768 , n407842 , n407843 );
buf ( n407845 , n60768 );
buf ( n407846 , n407845 );
nand ( n60771 , n60765 , n407846 );
buf ( n407848 , n60771 );
buf ( n407849 , n407848 );
not ( n60774 , n407849 );
buf ( n407851 , n391553 );
not ( n60776 , n407851 );
or ( n60777 , n60774 , n60776 );
buf ( n407854 , n407208 );
buf ( n407855 , n49166 );
nand ( n60780 , n407854 , n407855 );
buf ( n407857 , n60780 );
buf ( n407858 , n407857 );
nand ( n60783 , n60777 , n407858 );
buf ( n407860 , n60783 );
buf ( n407861 , n407860 );
buf ( n407862 , n42073 );
not ( n60787 , n407862 );
buf ( n407864 , n51648 );
not ( n60789 , n407864 );
or ( n60790 , n60787 , n60789 );
buf ( n407867 , n49653 );
buf ( n407868 , n42074 );
nand ( n60793 , n407867 , n407868 );
buf ( n407870 , n60793 );
buf ( n407871 , n407870 );
nand ( n60796 , n60790 , n407871 );
buf ( n407873 , n60796 );
buf ( n407874 , n407873 );
not ( n60799 , n407874 );
buf ( n407876 , n397102 );
not ( n60801 , n407876 );
or ( n60802 , n60799 , n60801 );
buf ( n407879 , n407453 );
buf ( n407880 , n386477 );
nand ( n60805 , n407879 , n407880 );
buf ( n407882 , n60805 );
buf ( n407883 , n407882 );
nand ( n60808 , n60802 , n407883 );
buf ( n407885 , n60808 );
buf ( n407886 , n407885 );
not ( n60811 , n407886 );
buf ( n407888 , n388830 );
not ( n60813 , n407888 );
buf ( n407890 , n407499 );
not ( n60815 , n407890 );
or ( n60816 , n60813 , n60815 );
buf ( n407893 , n41342 );
not ( n60818 , n407893 );
buf ( n407895 , n46478 );
not ( n60820 , n407895 );
or ( n60821 , n60818 , n60820 );
buf ( n407898 , n49686 );
buf ( n407899 , n45897 );
nand ( n60824 , n407898 , n407899 );
buf ( n407901 , n60824 );
buf ( n407902 , n407901 );
nand ( n60827 , n60821 , n407902 );
buf ( n407904 , n60827 );
buf ( n407905 , n407904 );
buf ( n407906 , n388872 );
nand ( n60831 , n407905 , n407906 );
buf ( n407908 , n60831 );
buf ( n407909 , n407908 );
nand ( n60834 , n60816 , n407909 );
buf ( n407911 , n60834 );
buf ( n407912 , n407911 );
not ( n60837 , n407912 );
or ( n60838 , n60811 , n60837 );
buf ( n407915 , n407885 );
buf ( n407916 , n407911 );
or ( n60841 , n407915 , n407916 );
xor ( n60842 , n406466 , n406550 );
xor ( n60843 , n60842 , n406810 );
buf ( n407920 , n60843 );
not ( n60845 , n407920 );
buf ( n407922 , n47726 );
not ( n60847 , n407922 );
and ( n60848 , n28644 , n40653 );
not ( n60849 , n28644 );
buf ( n407926 , n40652 );
not ( n60851 , n407926 );
buf ( n407928 , n60851 );
and ( n60853 , n60849 , n407928 );
or ( n60854 , n60848 , n60853 );
buf ( n407931 , n60854 );
not ( n60856 , n407931 );
or ( n60857 , n60847 , n60856 );
buf ( n407934 , n40651 );
buf ( n60859 , n407934 );
buf ( n407936 , n60859 );
not ( n60861 , n407936 );
buf ( n407938 , n12471 );
not ( n60863 , n407938 );
buf ( n407940 , n60863 );
not ( n60865 , n407940 );
or ( n60866 , n60861 , n60865 );
buf ( n407943 , n12471 );
buf ( n407944 , n40653 );
nand ( n60869 , n407943 , n407944 );
buf ( n407946 , n60869 );
nand ( n60871 , n60866 , n407946 );
not ( n60872 , n50041 );
nand ( n60873 , n60871 , n60872 );
buf ( n407950 , n60873 );
nand ( n60875 , n60857 , n407950 );
buf ( n407952 , n60875 );
not ( n60877 , n407952 );
or ( n60878 , n60845 , n60877 );
or ( n60879 , n407952 , n407920 );
not ( n60880 , n41555 );
and ( n60881 , n388215 , n60880 );
not ( n60882 , n388215 );
and ( n60883 , n60882 , n53251 );
or ( n60884 , n60881 , n60883 );
buf ( n407961 , n60884 );
not ( n60886 , n407961 );
buf ( n407963 , n60886 );
not ( n60888 , n407963 );
not ( n60889 , n42951 );
and ( n60890 , n60888 , n60889 );
and ( n60891 , n59706 , n42924 );
nor ( n60892 , n60890 , n60891 );
not ( n60893 , n60892 );
nand ( n60894 , n60879 , n60893 );
nand ( n60895 , n60878 , n60894 );
buf ( n407972 , n60895 );
nand ( n60897 , n60841 , n407972 );
buf ( n407974 , n60897 );
buf ( n407975 , n407974 );
nand ( n60900 , n60838 , n407975 );
buf ( n407977 , n60900 );
buf ( n407978 , n407977 );
xor ( n60903 , n407861 , n407978 );
not ( n60904 , n390536 );
buf ( n407981 , n391443 );
buf ( n407982 , n37345 );
and ( n60907 , n407981 , n407982 );
not ( n60908 , n407981 );
buf ( n407985 , n388905 );
and ( n60910 , n60908 , n407985 );
or ( n60911 , n60907 , n60910 );
buf ( n407988 , n60911 );
not ( n60913 , n407988 );
not ( n60914 , n60913 );
or ( n60915 , n60904 , n60914 );
nand ( n60916 , n60437 , n37316 );
nand ( n60917 , n60915 , n60916 );
buf ( n407994 , n60917 );
and ( n60919 , n60903 , n407994 );
and ( n60920 , n407861 , n407978 );
or ( n60921 , n60919 , n60920 );
buf ( n407998 , n60921 );
buf ( n407999 , n407998 );
and ( n60924 , n60760 , n407999 );
and ( n60925 , n407818 , n407835 );
or ( n60926 , n60924 , n60925 );
buf ( n408003 , n60926 );
buf ( n408004 , n408003 );
and ( n60929 , n60717 , n408004 );
and ( n60930 , n407766 , n407792 );
or ( n60931 , n60929 , n60930 );
buf ( n408008 , n60931 );
and ( n60933 , n407762 , n408008 );
nor ( n60934 , n60674 , n407759 );
nor ( n60935 , n60933 , n60934 );
not ( n60936 , n60935 );
and ( n60937 , n407109 , C1 );
or ( n60940 , n60937 , C0 );
buf ( n408015 , n60940 );
buf ( n408016 , n407116 );
xnor ( n60943 , n408015 , n408016 );
buf ( n408018 , n60943 );
not ( n60945 , n408018 );
or ( n60946 , n60936 , n60945 );
or ( n60947 , n408018 , n60935 );
buf ( n408022 , n407034 );
buf ( n408023 , n51553 );
and ( n60950 , n408022 , n408023 );
buf ( n408025 , n47891 );
not ( n60952 , n408025 );
buf ( n408027 , n385774 );
not ( n60954 , n408027 );
or ( n60955 , n60952 , n60954 );
buf ( n408030 , n38227 );
buf ( n408031 , n50584 );
nand ( n60958 , n408030 , n408031 );
buf ( n408033 , n60958 );
buf ( n408034 , n408033 );
nand ( n60961 , n60955 , n408034 );
buf ( n408036 , n60961 );
buf ( n408037 , n408036 );
not ( n60964 , n408037 );
buf ( n408039 , n50580 );
nor ( n60966 , n60964 , n408039 );
buf ( n408041 , n60966 );
buf ( n408042 , n408041 );
nor ( n60969 , n60950 , n408042 );
buf ( n408044 , n60969 );
buf ( n408045 , n408044 );
buf ( n408046 , C1 );
buf ( n408047 , n408046 );
buf ( n408048 , C1 );
buf ( n408049 , n408048 );
buf ( n408050 , C1 );
nand ( n61007 , n60947 , n408050 );
nand ( n61008 , n60946 , n61007 );
buf ( n408053 , n61008 );
not ( n61010 , n408053 );
or ( n61011 , n60670 , n61010 );
xor ( n61012 , n406185 , n406210 );
xor ( n61013 , n61012 , n406215 );
buf ( n408058 , n61013 );
not ( n61015 , n408058 );
not ( n61016 , n58891 );
not ( n61017 , n61016 );
not ( n61018 , n58792 );
or ( n61019 , n61017 , n61018 );
nand ( n61020 , n58791 , n58891 );
nand ( n61021 , n61019 , n61020 );
not ( n61022 , n58796 );
not ( n61023 , n61022 );
and ( n61024 , n61021 , n61023 );
not ( n61025 , n61021 );
and ( n61026 , n61025 , n61022 );
nor ( n61027 , n61024 , n61026 );
not ( n61028 , n61027 );
nand ( n61029 , n61015 , n61028 );
not ( n61030 , n61029 );
xor ( n61031 , n60186 , n407277 );
xnor ( n61032 , n61031 , n60048 );
not ( n61033 , n61032 );
or ( n61034 , n61030 , n61033 );
nand ( n61035 , n408058 , n61027 );
nand ( n61036 , n61034 , n61035 );
buf ( n408081 , n61036 );
nand ( n61038 , n61011 , n408081 );
buf ( n408083 , n61038 );
not ( n61040 , n60668 );
not ( n61041 , n61008 );
nand ( n61042 , n61040 , n61041 );
nand ( n61043 , n408083 , n61042 );
buf ( n408088 , n61043 );
not ( n61045 , n408088 );
xor ( n61046 , n60195 , n407316 );
xor ( n61047 , n61046 , n60619 );
buf ( n408092 , n61047 );
not ( n61049 , n408092 );
or ( n61050 , n61045 , n61049 );
not ( n61051 , n61047 );
buf ( n408096 , n61051 );
not ( n61053 , n408096 );
not ( n61054 , n61043 );
buf ( n408099 , n61054 );
not ( n61056 , n408099 );
or ( n61057 , n61053 , n61056 );
xor ( n408102 , n407326 , n407322 );
xnor ( n61059 , n408102 , n60617 );
not ( n61060 , n61059 );
not ( n61061 , n61060 );
and ( n61062 , n407689 , n407335 );
or ( n61065 , n61062 , C0 );
and ( n61066 , n61065 , n407404 );
not ( n61067 , n61065 );
and ( n61068 , n61067 , n407401 );
nor ( n61069 , n61066 , n61068 );
not ( n61070 , n61069 );
buf ( n408113 , n406271 );
not ( n61072 , n408113 );
buf ( n408115 , n406946 );
not ( n61074 , n408115 );
or ( n61075 , n61072 , n61074 );
buf ( n408118 , n59156 );
buf ( n408119 , n406268 );
nand ( n61078 , n408118 , n408119 );
buf ( n408121 , n61078 );
buf ( n408122 , n408121 );
nand ( n61081 , n61075 , n408122 );
buf ( n408124 , n61081 );
buf ( n408125 , n408124 );
buf ( n408126 , n59812 );
not ( n61085 , n408126 );
buf ( n408128 , n61085 );
buf ( n408129 , n408128 );
and ( n61088 , n408125 , n408129 );
not ( n61089 , n408125 );
buf ( n408132 , n59812 );
and ( n61091 , n61089 , n408132 );
nor ( n61092 , n61088 , n61091 );
buf ( n408135 , n61092 );
not ( n61094 , n408135 );
and ( n61095 , n61070 , n61094 );
not ( n61096 , n384008 );
and ( n61097 , n394219 , n40824 );
not ( n61098 , n394219 );
and ( n61099 , n61098 , n40973 );
nor ( n61100 , n61097 , n61099 );
not ( n61101 , n61100 );
and ( n61102 , n61096 , n61101 );
buf ( n408145 , n407241 );
not ( n61104 , n408145 );
buf ( n408147 , n40969 );
nor ( n61106 , n61104 , n408147 );
buf ( n408149 , n61106 );
nor ( n61108 , n61102 , n408149 );
buf ( n408151 , n61108 );
not ( n61110 , n408151 );
buf ( n408153 , n49117 );
not ( n61112 , n408153 );
buf ( n408155 , n388419 );
not ( n61114 , n408155 );
or ( n61115 , n61112 , n61114 );
buf ( n408158 , n40943 );
buf ( n408159 , n49124 );
nand ( n61118 , n408158 , n408159 );
buf ( n408161 , n61118 );
buf ( n408162 , n408161 );
nand ( n61121 , n61115 , n408162 );
buf ( n408164 , n61121 );
buf ( n408165 , n408164 );
not ( n61124 , n408165 );
buf ( n408167 , n36801 );
not ( n61126 , n408167 );
or ( n61127 , n61124 , n61126 );
buf ( n408170 , n392111 );
buf ( n408171 , n407256 );
nand ( n61130 , n408170 , n408171 );
buf ( n408173 , n61130 );
buf ( n408174 , n408173 );
nand ( n61133 , n61127 , n408174 );
buf ( n408176 , n61133 );
buf ( n408177 , n408176 );
not ( n61136 , n408177 );
buf ( n408179 , n61136 );
buf ( n408180 , n408179 );
not ( n61139 , n408180 );
or ( n61140 , n61110 , n61139 );
xor ( n61141 , n407195 , n407213 );
xor ( n61142 , n61141 , n407225 );
buf ( n408185 , n61142 );
buf ( n408186 , n408185 );
nand ( n61145 , n61140 , n408186 );
buf ( n408188 , n61145 );
buf ( n408189 , n408188 );
buf ( n408190 , n61108 );
not ( n61149 , n408190 );
buf ( n408192 , n61149 );
buf ( n408193 , n408192 );
buf ( n408194 , n408176 );
nand ( n61153 , n408193 , n408194 );
buf ( n408196 , n61153 );
buf ( n408197 , n408196 );
nand ( n61156 , n408189 , n408197 );
buf ( n408199 , n61156 );
buf ( n408200 , n408199 );
buf ( n408201 , n393825 );
not ( n61160 , n408201 );
buf ( n408203 , n398116 );
not ( n61162 , n408203 );
buf ( n408205 , n385734 );
not ( n61164 , n408205 );
or ( n61165 , n61162 , n61164 );
buf ( n408208 , n390794 );
buf ( n408209 , n393369 );
or ( n61168 , n408208 , n408209 );
buf ( n408211 , n61168 );
buf ( n408212 , n408211 );
nand ( n61171 , n61165 , n408212 );
buf ( n408214 , n61171 );
buf ( n408215 , n408214 );
not ( n61174 , n408215 );
or ( n61175 , n61160 , n61174 );
buf ( n408218 , n406315 );
buf ( n408219 , n45954 );
nand ( n61178 , n408218 , n408219 );
buf ( n408221 , n61178 );
buf ( n408222 , n408221 );
nand ( n61181 , n61175 , n408222 );
buf ( n408224 , n61181 );
buf ( n408225 , n408224 );
xor ( n61184 , n408200 , n408225 );
xor ( n61185 , n407441 , n407511 );
xor ( n61186 , n61185 , n407523 );
buf ( n408229 , n61186 );
buf ( n408230 , n408229 );
buf ( n408231 , n383891 );
not ( n61190 , n408231 );
buf ( n408233 , n61190 );
buf ( n408234 , n408233 );
not ( n61193 , n408234 );
buf ( n408236 , n392887 );
buf ( n408237 , n40775 );
and ( n61196 , n408236 , n408237 );
not ( n61197 , n408236 );
buf ( n408240 , n389936 );
and ( n61199 , n61197 , n408240 );
nor ( n61200 , n61196 , n61199 );
buf ( n408243 , n61200 );
buf ( n408244 , n408243 );
not ( n61203 , n408244 );
and ( n61204 , n61193 , n61203 );
buf ( n408247 , n407632 );
not ( n61206 , n408247 );
buf ( n408249 , n383910 );
nor ( n61208 , n61206 , n408249 );
buf ( n408251 , n61208 );
buf ( n408252 , n408251 );
nor ( n61211 , n61204 , n408252 );
buf ( n408254 , n61211 );
buf ( n408255 , n408254 );
not ( n61214 , n408255 );
buf ( n408257 , n61214 );
not ( n61216 , n408257 );
not ( n61217 , n43286 );
not ( n61218 , n388102 );
buf ( n408261 , n375784 );
not ( n61220 , n408261 );
buf ( n408263 , n61220 );
not ( n61222 , n408263 );
or ( n61223 , n61218 , n61222 );
buf ( n408266 , n386147 );
buf ( n408267 , n388105 );
nand ( n61226 , n408266 , n408267 );
buf ( n408269 , n61226 );
nand ( n61228 , n61223 , n408269 );
not ( n61229 , n61228 );
or ( n61230 , n61217 , n61229 );
nand ( n61231 , n407810 , n390362 );
nand ( n61232 , n61230 , n61231 );
not ( n61233 , n61232 );
or ( n61234 , n61216 , n61233 );
not ( n61235 , n61232 );
not ( n61236 , n61235 );
not ( n61237 , n408254 );
or ( n61238 , n61236 , n61237 );
not ( n61239 , n60427 );
not ( n61240 , n407465 );
not ( n61241 , n60405 );
and ( n61242 , n61240 , n61241 );
and ( n61243 , n407465 , n60405 );
nor ( n61244 , n61242 , n61243 );
not ( n61245 , n61244 );
or ( n61246 , n61239 , n61245 );
or ( n61247 , n60427 , n61244 );
nand ( n61248 , n61246 , n61247 );
buf ( n61249 , n61248 );
nand ( n61250 , n61238 , n61249 );
nand ( n61251 , n61234 , n61250 );
buf ( n408294 , n61251 );
xor ( n61253 , n408230 , n408294 );
buf ( n408296 , n400440 );
not ( n61255 , n408296 );
buf ( n408298 , n384562 );
not ( n61257 , n408298 );
or ( n61258 , n61255 , n61257 );
buf ( n408301 , n395885 );
buf ( n408302 , n51185 );
nand ( n61261 , n408301 , n408302 );
buf ( n408304 , n61261 );
buf ( n408305 , n408304 );
nand ( n61264 , n61258 , n408305 );
buf ( n408307 , n61264 );
buf ( n408308 , n408307 );
not ( n61267 , n408308 );
buf ( n408310 , n384624 );
not ( n61269 , n408310 );
or ( n61270 , n61267 , n61269 );
buf ( n408313 , n60483 );
buf ( n408314 , n384554 );
nand ( n61273 , n408313 , n408314 );
buf ( n408316 , n61273 );
buf ( n408317 , n408316 );
nand ( n61276 , n61270 , n408317 );
buf ( n408319 , n61276 );
buf ( n408320 , n408319 );
and ( n61279 , n61253 , n408320 );
and ( n61280 , n408230 , n408294 );
or ( n61281 , n61279 , n61280 );
buf ( n408324 , n61281 );
buf ( n408325 , n408324 );
and ( n61284 , n61184 , n408325 );
and ( n61285 , n408200 , n408225 );
or ( n61286 , n61284 , n61285 );
buf ( n408329 , n61286 );
buf ( n408330 , n408329 );
xor ( n61289 , n407532 , n407557 );
xor ( n61290 , n61289 , n407685 );
buf ( n408333 , n61290 );
buf ( n408334 , n408333 );
xor ( n61293 , n408330 , n408334 );
buf ( n408336 , n51553 );
not ( n61295 , n408336 );
buf ( n408338 , n408036 );
not ( n61297 , n408338 );
or ( n61298 , n61295 , n61297 );
not ( n61299 , n47891 );
buf ( n408342 , n61299 );
buf ( n61301 , n408342 );
buf ( n408344 , n61301 );
buf ( n408345 , n408344 );
not ( n61304 , n408345 );
buf ( n408347 , n61304 );
buf ( n408348 , n408347 );
not ( n61307 , n408348 );
buf ( n408350 , n37147 );
not ( n61309 , n408350 );
or ( n61310 , n61307 , n61309 );
buf ( n408353 , n394463 );
buf ( n408354 , n408344 );
nand ( n61313 , n408353 , n408354 );
buf ( n408356 , n61313 );
buf ( n408357 , n408356 );
nand ( n61316 , n61310 , n408357 );
buf ( n408359 , n61316 );
buf ( n408360 , n408359 );
buf ( n408361 , n50579 );
nand ( n61320 , n408360 , n408361 );
buf ( n408363 , n61320 );
buf ( n408364 , n408363 );
nand ( n61323 , n61298 , n408364 );
buf ( n408366 , n61323 );
xor ( n61325 , n407359 , n407384 );
xor ( n61326 , n61325 , n407392 );
buf ( n408369 , n61326 );
xor ( n61328 , n408366 , n408369 );
buf ( n408371 , n43515 );
not ( n61330 , n408371 );
buf ( n408373 , n60505 );
not ( n61332 , n408373 );
or ( n61333 , n61330 , n61332 );
buf ( n408376 , n391027 );
not ( n61335 , n408376 );
buf ( n408378 , n388955 );
not ( n61337 , n408378 );
or ( n61338 , n61335 , n61337 );
nand ( n61339 , n37763 , n391024 );
buf ( n408382 , n61339 );
nand ( n61341 , n61338 , n408382 );
buf ( n408384 , n61341 );
buf ( n408385 , n408384 );
buf ( n408386 , n43727 );
nand ( n61345 , n408385 , n408386 );
buf ( n408388 , n61345 );
buf ( n408389 , n408388 );
nand ( n61348 , n61333 , n408389 );
buf ( n408391 , n61348 );
buf ( n408392 , n408391 );
buf ( n408393 , n400033 );
not ( n61352 , n408393 );
buf ( n408395 , n389598 );
not ( n61354 , n408395 );
or ( n61355 , n61352 , n61354 );
buf ( n408398 , n389589 );
buf ( n408399 , n400042 );
nand ( n61358 , n408398 , n408399 );
buf ( n408401 , n61358 );
buf ( n408402 , n408401 );
nand ( n61361 , n61355 , n408402 );
buf ( n408404 , n61361 );
buf ( n408405 , n408404 );
not ( n61364 , n408405 );
buf ( n408407 , n391917 );
not ( n61366 , n408407 );
or ( n61367 , n61364 , n61366 );
buf ( n408410 , n391173 );
buf ( n408411 , n59786 );
nand ( n61370 , n408410 , n408411 );
buf ( n408413 , n61370 );
buf ( n408414 , n408413 );
nand ( n61373 , n61367 , n408414 );
buf ( n408416 , n61373 );
buf ( n408417 , n408416 );
xor ( n61376 , n408392 , n408417 );
buf ( n408419 , n47726 );
not ( n61378 , n408419 );
buf ( n408421 , n59291 );
not ( n61380 , n408421 );
or ( n61381 , n61378 , n61380 );
buf ( n408424 , n60854 );
buf ( n408425 , n397476 );
nand ( n61384 , n408424 , n408425 );
buf ( n408427 , n61384 );
buf ( n408428 , n408427 );
nand ( n61387 , n61381 , n408428 );
buf ( n408430 , n61387 );
buf ( n408431 , n408430 );
buf ( n408432 , n388502 );
not ( n61391 , n408432 );
buf ( n408434 , n399164 );
not ( n61393 , n408434 );
or ( n61394 , n61391 , n61393 );
buf ( n408437 , n399167 );
buf ( n408438 , n54922 );
nand ( n61397 , n408437 , n408438 );
buf ( n408440 , n61397 );
buf ( n408441 , n408440 );
nand ( n61400 , n61394 , n408441 );
buf ( n408443 , n61400 );
buf ( n408444 , n408443 );
not ( n61403 , n408444 );
buf ( n408446 , n389122 );
not ( n61405 , n408446 );
or ( n61406 , n61403 , n61405 );
buf ( n408449 , n407479 );
buf ( n408450 , n46921 );
nand ( n61409 , n408449 , n408450 );
buf ( n408452 , n61409 );
buf ( n408453 , n408452 );
nand ( n61412 , n61406 , n408453 );
buf ( n408455 , n61412 );
buf ( n408456 , n408455 );
xor ( n61415 , n408431 , n408456 );
xor ( n61416 , n406447 , n406815 );
xor ( n61417 , n61416 , n406846 );
buf ( n408460 , n61417 );
buf ( n408461 , n408460 );
and ( n61420 , n61415 , n408461 );
and ( n61421 , n408431 , n408456 );
or ( n61422 , n61420 , n61421 );
buf ( n408465 , n61422 );
buf ( n408466 , n408465 );
not ( n61425 , n388746 );
and ( n61426 , n41118 , n405736 );
not ( n61427 , n41118 );
and ( n61428 , n61427 , n388757 );
or ( n61429 , n61426 , n61428 );
not ( n61430 , n61429 );
or ( n61431 , n61425 , n61430 );
buf ( n408474 , n407662 );
buf ( n408475 , n388809 );
nand ( n61434 , n408474 , n408475 );
buf ( n408477 , n61434 );
nand ( n61436 , n61431 , n408477 );
buf ( n408479 , n61436 );
xor ( n61438 , n408466 , n408479 );
buf ( n408481 , n386209 );
buf ( n408482 , n358975 );
and ( n61441 , n408481 , n408482 );
buf ( n408484 , n61441 );
buf ( n408485 , n408484 );
and ( n61444 , n61438 , n408485 );
and ( n61445 , n408466 , n408479 );
or ( n61446 , n61444 , n61445 );
buf ( n408489 , n61446 );
buf ( n408490 , n408489 );
and ( n61449 , n61376 , n408490 );
and ( n61450 , n408392 , n408417 );
or ( n61451 , n61449 , n61450 );
buf ( n408494 , n61451 );
and ( n61453 , n61328 , n408494 );
and ( n61454 , n408366 , n408369 );
or ( n61455 , n61453 , n61454 );
buf ( n408498 , n61455 );
and ( n61457 , n61293 , n408498 );
and ( n61458 , n408330 , n408334 );
or ( n61459 , n61457 , n61458 );
buf ( n408502 , n61459 );
buf ( n408503 , n61069 );
buf ( n408504 , n408135 );
nand ( n61463 , n408503 , n408504 );
buf ( n408506 , n61463 );
and ( n61465 , n408502 , n408506 );
nor ( n61466 , n61095 , n61465 );
not ( n61467 , n61466 );
not ( n61468 , n61467 );
or ( n61469 , n61061 , n61468 );
buf ( n408512 , n61059 );
not ( n61471 , n408512 );
buf ( n408514 , n61466 );
not ( n61473 , n408514 );
or ( n61474 , n61471 , n61473 );
xor ( n61475 , n406255 , n406953 );
xor ( n61476 , n61475 , n406960 );
buf ( n408519 , n61476 );
nand ( n61478 , n61474 , n408519 );
buf ( n408521 , n61478 );
nand ( n61480 , n61469 , n408521 );
buf ( n408523 , n61480 );
nand ( n61482 , n61057 , n408523 );
buf ( n408525 , n61482 );
buf ( n408526 , n408525 );
nand ( n61485 , n61050 , n408526 );
buf ( n408528 , n61485 );
buf ( n408529 , n408528 );
xor ( n61488 , n407717 , n408529 );
xor ( n61489 , n405651 , n406117 );
xor ( n61490 , n61489 , n406975 );
buf ( n408533 , n61490 );
buf ( n408534 , n408533 );
and ( n61493 , n61488 , n408534 );
and ( n61494 , n407717 , n408529 );
or ( n61495 , n61493 , n61494 );
buf ( n408538 , n61495 );
buf ( n408539 , n408538 );
not ( n408540 , n408539 );
buf ( n408541 , n408540 );
nand ( n61500 , n60627 , n408541 );
buf ( n408543 , n61500 );
xor ( n61502 , n407717 , n408529 );
xor ( n61503 , n61502 , n408534 );
buf ( n408546 , n61503 );
buf ( n408547 , n408546 );
not ( n61506 , n408547 );
buf ( n408549 , n61506 );
not ( n61508 , n61480 );
not ( n61509 , n61043 );
not ( n61510 , n61051 );
or ( n61511 , n61509 , n61510 );
or ( n61512 , n61051 , n61043 );
nand ( n61513 , n61511 , n61512 );
not ( n61514 , n61513 );
or ( n61515 , n61508 , n61514 );
not ( n61516 , n61043 );
not ( n61517 , n61051 );
or ( n61518 , n61516 , n61517 );
or ( n61519 , n61051 , n61043 );
nand ( n61520 , n61518 , n61519 );
or ( n61521 , n61520 , n61480 );
nand ( n61522 , n61515 , n61521 );
buf ( n408565 , n61522 );
not ( n61524 , n408565 );
buf ( n408567 , n61524 );
not ( n61526 , n408567 );
buf ( n408569 , n59123 );
buf ( n408570 , n406121 );
and ( n61529 , n408569 , n408570 );
not ( n61530 , n408569 );
buf ( n408573 , n406121 );
not ( n61532 , n408573 );
buf ( n408575 , n61532 );
buf ( n408576 , n408575 );
and ( n61535 , n61530 , n408576 );
nor ( n61536 , n61529 , n61535 );
buf ( n408579 , n61536 );
buf ( n408580 , n408579 );
buf ( n408581 , n59836 );
and ( n61540 , n408580 , n408581 );
not ( n61541 , n408580 );
buf ( n408584 , n59836 );
not ( n61543 , n408584 );
buf ( n408586 , n61543 );
buf ( n408587 , n408586 );
and ( n61546 , n61541 , n408587 );
nor ( n61547 , n61540 , n61546 );
buf ( n408590 , n61547 );
not ( n61549 , n408590 );
or ( n61550 , n61526 , n61549 );
buf ( n408593 , n408590 );
not ( n61552 , n408593 );
buf ( n408595 , n61552 );
not ( n61554 , n408595 );
not ( n61555 , n61522 );
or ( n61556 , n61554 , n61555 );
xor ( n61557 , n61036 , n60668 );
xnor ( n61558 , n61557 , n61041 );
buf ( n408601 , n61558 );
not ( n61560 , n408601 );
buf ( n408603 , n61560 );
buf ( n408604 , n408603 );
not ( n61563 , n408604 );
xor ( n61564 , n408330 , n408334 );
xor ( n61565 , n61564 , n408498 );
buf ( n408608 , n61565 );
not ( n61567 , n408608 );
buf ( n408610 , n60680 );
buf ( n408611 , n408008 );
xor ( n61570 , n408610 , n408611 );
buf ( n408613 , n60674 );
xnor ( n61572 , n61570 , n408613 );
buf ( n408615 , n61572 );
buf ( n408616 , n408615 );
not ( n61575 , n408616 );
buf ( n408618 , n408359 );
not ( n61577 , n50564 );
buf ( n408620 , n61577 );
and ( n61579 , n408618 , n408620 );
and ( n61580 , n37173 , n50584 );
not ( n61581 , n37173 );
and ( n61582 , n61581 , n47891 );
or ( n61583 , n61580 , n61582 );
buf ( n408626 , n61583 );
buf ( n408627 , n50579 );
and ( n61586 , n408626 , n408627 );
buf ( n408629 , n61586 );
buf ( n408630 , n408629 );
nor ( n61589 , n61579 , n408630 );
buf ( n408632 , n61589 );
buf ( n408633 , n408632 );
not ( n61592 , n408633 );
buf ( n408635 , n61592 );
buf ( n408636 , n408635 );
not ( n61595 , n408636 );
buf ( n408638 , n395362 );
not ( n61597 , n408638 );
and ( n61598 , n47863 , n390373 );
not ( n61599 , n47863 );
and ( n61600 , n61599 , n36188 );
or ( n61601 , n61598 , n61600 );
buf ( n408644 , n61601 );
not ( n61603 , n408644 );
or ( n61604 , n61597 , n61603 );
buf ( n408647 , n395315 );
not ( n61606 , n408647 );
buf ( n408649 , n61606 );
buf ( n408650 , n408649 );
not ( n61609 , n408650 );
buf ( n408652 , n42234 );
not ( n61611 , n408652 );
or ( n61612 , n61609 , n61611 );
buf ( n408655 , n36216 );
buf ( n408656 , n395315 );
nand ( n61615 , n408655 , n408656 );
buf ( n408658 , n61615 );
buf ( n408659 , n408658 );
nand ( n61618 , n61612 , n408659 );
buf ( n408661 , n61618 );
buf ( n408662 , n408661 );
buf ( n408663 , n395349 );
nand ( n61622 , n408662 , n408663 );
buf ( n408665 , n61622 );
buf ( n408666 , n408665 );
nand ( n61625 , n61604 , n408666 );
buf ( n408668 , n61625 );
buf ( n408669 , n408668 );
not ( n61628 , n408669 );
or ( n61629 , n61595 , n61628 );
buf ( n408672 , n408668 );
not ( n61631 , n408672 );
buf ( n408674 , n61631 );
buf ( n408675 , n408674 );
not ( n61634 , n408675 );
buf ( n408677 , n408632 );
not ( n61636 , n408677 );
or ( n61637 , n61634 , n61636 );
buf ( n408680 , n399274 );
not ( n61639 , n408680 );
buf ( n408682 , n384562 );
not ( n61641 , n408682 );
or ( n61642 , n61639 , n61641 );
buf ( n408685 , n395885 );
buf ( n408686 , n399283 );
nand ( n61645 , n408685 , n408686 );
buf ( n408688 , n61645 );
buf ( n408689 , n408688 );
nand ( n61648 , n61642 , n408689 );
buf ( n408691 , n61648 );
buf ( n408692 , n408691 );
not ( n61651 , n408692 );
buf ( n408694 , n392659 );
not ( n61653 , n408694 );
or ( n61654 , n61651 , n61653 );
buf ( n408697 , n408307 );
buf ( n408698 , n393602 );
nand ( n61657 , n408697 , n408698 );
buf ( n408700 , n61657 );
buf ( n408701 , n408700 );
nand ( n61660 , n61654 , n408701 );
buf ( n408703 , n61660 );
buf ( n408704 , n408703 );
buf ( n408705 , n45260 );
not ( n61664 , n408705 );
buf ( n408707 , n399986 );
not ( n61666 , n408707 );
buf ( n408709 , n38660 );
not ( n61668 , n408709 );
or ( n61669 , n61666 , n61668 );
not ( n61670 , n38153 );
not ( n61671 , n36562 );
or ( n61672 , n61670 , n61671 );
nand ( n61673 , n61672 , n44776 );
buf ( n408716 , n61673 );
nand ( n61675 , n61669 , n408716 );
buf ( n408718 , n61675 );
buf ( n408719 , n408718 );
not ( n61678 , n408719 );
or ( n61679 , n61664 , n61678 );
buf ( n408722 , n399986 );
not ( n61681 , n408722 );
buf ( n408724 , n384083 );
not ( n61683 , n408724 );
or ( n61684 , n61681 , n61683 );
buf ( n408727 , n385983 );
buf ( n408728 , n44776 );
nand ( n61687 , n408727 , n408728 );
buf ( n408730 , n61687 );
buf ( n408731 , n408730 );
nand ( n61690 , n61684 , n408731 );
buf ( n408733 , n61690 );
buf ( n408734 , n408733 );
buf ( n408735 , n392740 );
nand ( n61694 , n408734 , n408735 );
buf ( n408737 , n61694 );
buf ( n408738 , n408737 );
nand ( n61697 , n61679 , n408738 );
buf ( n408740 , n61697 );
buf ( n408741 , n408740 );
xor ( n61700 , n408704 , n408741 );
buf ( n408743 , n55055 );
not ( n61702 , n408743 );
buf ( n408745 , n391183 );
not ( n61704 , n408745 );
or ( n61705 , n61702 , n61704 );
buf ( n408748 , n385630 );
buf ( n408749 , n404855 );
nand ( n61708 , n408748 , n408749 );
buf ( n408751 , n61708 );
buf ( n408752 , n408751 );
nand ( n61711 , n61705 , n408752 );
buf ( n408754 , n61711 );
buf ( n408755 , n408754 );
not ( n61714 , n408755 );
buf ( n408757 , n391917 );
not ( n61716 , n408757 );
or ( n61717 , n61714 , n61716 );
buf ( n408760 , n391173 );
buf ( n408761 , n408404 );
nand ( n61720 , n408760 , n408761 );
buf ( n408763 , n61720 );
buf ( n408764 , n408763 );
nand ( n61723 , n61717 , n408764 );
buf ( n408766 , n61723 );
buf ( n408767 , n408766 );
and ( n61726 , n61700 , n408767 );
and ( n61727 , n408704 , n408741 );
or ( n61728 , n61726 , n61727 );
buf ( n408771 , n61728 );
buf ( n408772 , n408771 );
nand ( n61731 , n61637 , n408772 );
buf ( n408774 , n61731 );
buf ( n408775 , n408774 );
nand ( n61734 , n61629 , n408775 );
buf ( n408777 , n61734 );
buf ( n408778 , n408777 );
xor ( n61737 , n407766 , n407792 );
xor ( n61738 , n61737 , n408004 );
buf ( n408781 , n61738 );
buf ( n408782 , n408781 );
xor ( n61741 , n408778 , n408782 );
xor ( n61742 , n408200 , n408225 );
xor ( n61743 , n61742 , n408325 );
buf ( n408786 , n61743 );
buf ( n408787 , n408786 );
and ( n61746 , n61741 , n408787 );
and ( n61747 , n408778 , n408782 );
or ( n61748 , n61746 , n61747 );
buf ( n408791 , n61748 );
buf ( n408792 , n408791 );
not ( n61751 , n408792 );
buf ( n408794 , n61751 );
buf ( n408795 , n408794 );
nand ( n61754 , n61575 , n408795 );
buf ( n408797 , n61754 );
not ( n61756 , n408797 );
or ( n61757 , n61567 , n61756 );
buf ( n408800 , n408615 );
not ( n61759 , n408800 );
buf ( n408802 , n408794 );
nor ( n61761 , n61759 , n408802 );
buf ( n408804 , n61761 );
not ( n61763 , n408804 );
nand ( n61764 , n61757 , n61763 );
not ( n61765 , n61764 );
and ( n61767 , n407762 , n408008 );
nor ( n61768 , n61767 , n60934 );
not ( n61769 , n61768 );
not ( n61770 , n61769 );
or ( n61771 , C0 , n61770 );
nand ( n61773 , C0 , n61768 );
nand ( n61774 , n61771 , n61773 );
and ( n61775 , n61774 , n408018 );
not ( n61776 , n61774 );
not ( n61777 , n408018 );
and ( n61778 , n61776 , n61777 );
nor ( n61779 , n61775 , n61778 );
not ( n61780 , n61779 );
not ( n61781 , n61780 );
or ( n61782 , n61765 , n61781 );
not ( n61783 , n408608 );
not ( n61784 , n408797 );
or ( n61785 , n61783 , n61784 );
nand ( n61786 , n61785 , n61763 );
not ( n61787 , n61779 );
or ( n61788 , n61786 , n61787 );
not ( n61789 , n408502 );
not ( n61790 , n61789 );
not ( n61791 , n61069 );
or ( n61792 , n61790 , n61791 );
not ( n61793 , n61069 );
nand ( n61794 , n61793 , n408502 );
nand ( n61795 , n61792 , n61794 );
buf ( n61796 , n408135 );
and ( n61797 , n61795 , n61796 );
not ( n61798 , n61795 );
not ( n61799 , n61796 );
and ( n61800 , n61798 , n61799 );
nor ( n61801 , n61797 , n61800 );
nand ( n61802 , n61788 , n61801 );
nand ( n61803 , n61782 , n61802 );
not ( n61804 , n61803 );
buf ( n408845 , n61804 );
not ( n61806 , n408845 );
or ( n61807 , n61563 , n61806 );
xor ( n61808 , n406322 , n59204 );
xor ( n61809 , n61808 , n406936 );
buf ( n408850 , n408185 );
buf ( n408851 , n408176 );
xor ( n61829 , n408850 , n408851 );
buf ( n408853 , n408192 );
xnor ( n61831 , n61829 , n408853 );
buf ( n408855 , n61831 );
buf ( n408856 , n408855 );
not ( n61834 , n408856 );
or ( n61835 , n390810 , n393384 );
or ( n61836 , n41595 , n398116 );
nand ( n61837 , n61835 , n61836 );
buf ( n408861 , n61837 );
not ( n61839 , n408861 );
buf ( n408863 , n393404 );
not ( n61841 , n408863 );
and ( n61842 , n61839 , n61841 );
buf ( n408866 , n408214 );
buf ( n408867 , n45954 );
and ( n61845 , n408866 , n408867 );
nor ( n61846 , n61842 , n61845 );
buf ( n408870 , n61846 );
buf ( n408871 , n408870 );
not ( n61849 , n408871 );
or ( n61850 , n61834 , n61849 );
not ( n61851 , n390292 );
buf ( n408875 , n397495 );
buf ( n408876 , n395722 );
and ( n61854 , n408875 , n408876 );
not ( n61855 , n408875 );
buf ( n408879 , n396373 );
and ( n61857 , n61855 , n408879 );
nor ( n61858 , n61854 , n61857 );
buf ( n408882 , n61858 );
not ( n61860 , n408882 );
and ( n61861 , n61851 , n61860 );
and ( n61862 , n392111 , n408164 );
nor ( n61863 , n61861 , n61862 );
not ( n61864 , n61863 );
buf ( n408888 , n384008 );
not ( n61866 , n408888 );
buf ( n408890 , n394814 );
buf ( n408891 , n36397 );
and ( n61869 , n408890 , n408891 );
not ( n61870 , n408890 );
buf ( n408894 , n40835 );
and ( n61872 , n61870 , n408894 );
nor ( n61873 , n61869 , n61872 );
buf ( n408897 , n61873 );
buf ( n408898 , n408897 );
not ( n61876 , n408898 );
and ( n61877 , n61866 , n61876 );
buf ( n408901 , n394219 );
buf ( n408902 , n40835 );
and ( n61880 , n408901 , n408902 );
not ( n61881 , n408901 );
buf ( n408905 , n40974 );
and ( n61883 , n61881 , n408905 );
or ( n61884 , n61880 , n61883 );
buf ( n408908 , n61884 );
buf ( n408909 , n408908 );
buf ( n408910 , n383943 );
nor ( n61888 , n408909 , n408910 );
buf ( n408912 , n61888 );
buf ( n408913 , n408912 );
nor ( n61891 , n61877 , n408913 );
buf ( n408915 , n61891 );
not ( n61893 , n408915 );
or ( n61894 , n61864 , n61893 );
xor ( n61895 , n59724 , n406431 );
xnor ( n61896 , n61895 , n406889 );
nand ( n61897 , n61894 , n61896 );
buf ( n408921 , n61897 );
buf ( n408922 , n408915 );
not ( n61900 , n408922 );
buf ( n408924 , n61863 );
not ( n61902 , n408924 );
buf ( n408926 , n61902 );
buf ( n408927 , n408926 );
nand ( n61905 , n61900 , n408927 );
buf ( n408929 , n61905 );
buf ( n408930 , n408929 );
nand ( n61908 , n408921 , n408930 );
buf ( n408932 , n61908 );
buf ( n408933 , n408932 );
nand ( n61911 , n61850 , n408933 );
buf ( n408935 , n61911 );
buf ( n408936 , n408935 );
buf ( n408937 , n408870 );
not ( n61915 , n408937 );
buf ( n408939 , n408855 );
not ( n61917 , n408939 );
buf ( n408941 , n61917 );
buf ( n408942 , n408941 );
nand ( n61920 , n61915 , n408942 );
buf ( n408944 , n61920 );
buf ( n408945 , n408944 );
nand ( n61923 , n408936 , n408945 );
buf ( n408947 , n61923 );
buf ( n408948 , n408947 );
buf ( n408949 , C0 );
or ( n61929 , n408948 , n408949 );
buf ( n408951 , n407781 );
buf ( n408952 , n392740 );
and ( n408953 , n408951 , n408952 );
buf ( n408954 , n408733 );
not ( n61934 , n408954 );
buf ( n408956 , n44771 );
nor ( n61936 , n61934 , n408956 );
buf ( n408958 , n61936 );
buf ( n408959 , n408958 );
nor ( n61939 , n408953 , n408959 );
buf ( n408961 , n61939 );
not ( n61941 , n408961 );
not ( n61942 , n61941 );
xor ( n61943 , n407620 , n407669 );
xnor ( n61944 , n61943 , n407644 );
not ( n61945 , n61944 );
not ( n61946 , n61945 );
or ( n61947 , n61942 , n61946 );
not ( n61948 , n408961 );
not ( n61949 , n61944 );
or ( n61950 , n61948 , n61949 );
not ( n61951 , n406358 );
not ( n61952 , n406354 );
not ( n61953 , n61952 );
or ( n61954 , n61951 , n61953 );
not ( n61955 , n406358 );
nand ( n61956 , n61955 , n406354 );
nand ( n61957 , n61954 , n61956 );
xor ( n61958 , n61957 , n59766 );
not ( n61959 , n61958 );
nand ( n61960 , n61950 , n61959 );
nand ( n61961 , n61947 , n61960 );
buf ( n408983 , n61961 );
nand ( n61963 , n61929 , n408983 );
buf ( n408985 , n61963 );
nand ( n61965 , C1 , n408985 );
xor ( n61966 , n61809 , n61965 );
xor ( n61967 , n406904 , n406907 );
xor ( n61968 , n61967 , n406932 );
buf ( n408990 , n61968 );
buf ( n408991 , C0 );
buf ( n408992 , n408990 );
buf ( n408993 , n408991 );
or ( n61996 , n408992 , n408993 );
buf ( n408995 , n406867 );
buf ( n408996 , n389162 );
and ( n61999 , n408995 , n408996 );
buf ( n408998 , n46114 );
not ( n62001 , n408998 );
buf ( n409000 , n24116 );
not ( n62003 , n409000 );
or ( n62004 , n62001 , n62003 );
buf ( n409003 , n397069 );
not ( n62006 , n24116 );
buf ( n409005 , n62006 );
nand ( n62008 , n409003 , n409005 );
buf ( n409007 , n62008 );
buf ( n409008 , n409007 );
nand ( n62011 , n62004 , n409008 );
buf ( n409010 , n62011 );
buf ( n409011 , n409010 );
not ( n62014 , n409011 );
buf ( n409013 , n41710 );
nor ( n62016 , n62014 , n409013 );
buf ( n409015 , n62016 );
buf ( n409016 , n409015 );
nor ( n62019 , n61999 , n409016 );
buf ( n409018 , n62019 );
buf ( n409019 , n409018 );
not ( n62022 , n409019 );
buf ( n409021 , n389341 );
not ( n62024 , n409021 );
buf ( n409023 , n385488 );
not ( n62026 , n409023 );
or ( n62027 , n62024 , n62026 );
buf ( n409026 , n388962 );
buf ( n409027 , n393185 );
nand ( n62030 , n409026 , n409027 );
buf ( n409029 , n62030 );
buf ( n409030 , n409029 );
nand ( n62033 , n62027 , n409030 );
buf ( n409032 , n62033 );
buf ( n409033 , n409032 );
not ( n62036 , n409033 );
buf ( n409035 , n393544 );
not ( n62038 , n409035 );
or ( n62039 , n62036 , n62038 );
buf ( n409038 , n407848 );
buf ( n409039 , n51692 );
nand ( n62042 , n409038 , n409039 );
buf ( n409041 , n62042 );
buf ( n409042 , n409041 );
nand ( n62045 , n62039 , n409042 );
buf ( n409044 , n62045 );
buf ( n409045 , n409044 );
not ( n62048 , n409045 );
buf ( n409047 , n62048 );
buf ( n409048 , n409047 );
not ( n62051 , n409048 );
or ( n62052 , n62022 , n62051 );
buf ( n409051 , n388830 );
not ( n62054 , n409051 );
buf ( n409053 , n407904 );
not ( n62056 , n409053 );
or ( n62057 , n62054 , n62056 );
and ( n62058 , n27258 , n45897 );
not ( n62059 , n27258 );
and ( n62060 , n62059 , n41342 );
or ( n62061 , n62058 , n62060 );
buf ( n409060 , n62061 );
buf ( n409061 , n388872 );
nand ( n62064 , n409060 , n409061 );
buf ( n409063 , n62064 );
buf ( n409064 , n409063 );
nand ( n62067 , n62057 , n409064 );
buf ( n409066 , n62067 );
buf ( n409067 , n409066 );
xor ( n62070 , n406522 , n406542 );
xor ( n62071 , n62070 , n406546 );
xor ( n62072 , n406695 , n59677 );
xor ( n62073 , n62071 , n62072 );
buf ( n409072 , n62073 );
not ( n62075 , n40638 );
buf ( n409074 , n62075 );
not ( n62077 , n409074 );
buf ( n409076 , n62077 );
not ( n62079 , n409076 );
not ( n62080 , n60871 );
or ( n62081 , n62079 , n62080 );
buf ( n409080 , n50041 );
not ( n62083 , n409080 );
buf ( n409082 , n62083 );
buf ( n409083 , n409082 );
buf ( n409084 , n407936 );
not ( n62087 , n409084 );
buf ( n409086 , n406824 );
not ( n62089 , n409086 );
or ( n62090 , n62087 , n62089 );
buf ( n409089 , n388230 );
buf ( n409090 , n407936 );
not ( n62093 , n409090 );
buf ( n409092 , n62093 );
buf ( n409093 , n409092 );
nand ( n62096 , n409089 , n409093 );
buf ( n409095 , n62096 );
buf ( n409096 , n409095 );
nand ( n62099 , n62090 , n409096 );
buf ( n409098 , n62099 );
buf ( n409099 , n409098 );
nand ( n62102 , n409083 , n409099 );
buf ( n409101 , n62102 );
nand ( n62104 , n62081 , n409101 );
buf ( n409103 , n62104 );
or ( n62106 , n409072 , n409103 );
buf ( n409105 , n406720 );
buf ( n409106 , n406731 );
or ( n62109 , n409105 , n409106 );
buf ( n409108 , n406734 );
nand ( n62111 , n62109 , n409108 );
buf ( n409110 , n62111 );
buf ( n409111 , n409110 );
buf ( n409112 , n58166 );
buf ( n409113 , n55905 );
and ( n62116 , n409112 , n409113 );
buf ( n409115 , n58205 );
buf ( n409116 , n55895 );
and ( n62119 , n409115 , n409116 );
nor ( n62120 , n62116 , n62119 );
buf ( n409119 , n62120 );
buf ( n409120 , n409119 );
buf ( n409121 , n403120 );
or ( n62124 , n409120 , n409121 );
buf ( n409123 , n406642 );
buf ( n409124 , n403133 );
or ( n62127 , n409123 , n409124 );
nand ( n62128 , n62124 , n62127 );
buf ( n409127 , n62128 );
buf ( n409128 , n409127 );
xor ( n62131 , n409111 , n409128 );
not ( n62132 , n53758 );
not ( n62133 , n54252 );
or ( n62134 , n62132 , n62133 );
not ( n62135 , n54255 );
nand ( n62136 , n62134 , n62135 );
not ( n62137 , n54257 );
nand ( n62138 , n62137 , n53710 );
xnor ( n62139 , n62136 , n62138 );
buf ( n409138 , n62139 );
not ( n62141 , n409138 );
buf ( n409140 , n62141 );
buf ( n409141 , n409140 );
buf ( n409142 , n403083 );
or ( n62145 , n409141 , n409142 );
buf ( n409144 , n59596 );
not ( n62147 , n409144 );
buf ( n409146 , n62147 );
buf ( n409147 , n409146 );
buf ( n409148 , n403092 );
or ( n62151 , n409147 , n409148 );
nand ( n62152 , n62145 , n62151 );
buf ( n409151 , n62152 );
buf ( n409152 , n409151 );
buf ( n62155 , n9071 );
buf ( n409154 , n62155 );
not ( n62157 , n409154 );
buf ( n409156 , n62157 );
not ( n62159 , n59463 );
or ( n62160 , n409156 , n62159 );
or ( n62161 , n62155 , n59463 );
nand ( n62162 , n62160 , n62161 );
buf ( n409161 , n62162 );
buf ( n62164 , n1856 );
buf ( n409163 , n62164 );
buf ( n409164 , n409156 );
and ( n62167 , n409163 , n409164 );
not ( n62168 , n409163 );
buf ( n409167 , n62155 );
and ( n62170 , n62168 , n409167 );
or ( n62171 , n62167 , n62170 );
buf ( n409170 , n62171 );
buf ( n409171 , n409170 );
and ( n62174 , n409161 , n409171 );
buf ( n409173 , n62174 );
buf ( n409174 , n409173 );
buf ( n62177 , n59463 );
buf ( n409176 , n62177 );
not ( n62179 , n409176 );
buf ( n409178 , n62179 );
buf ( n409179 , n409178 );
nand ( n62182 , n409174 , n409179 );
buf ( n409181 , n62182 );
buf ( n409182 , n409181 );
buf ( n409183 , n409170 );
not ( n62186 , n409183 );
buf ( n409185 , n62186 );
buf ( n409186 , n409185 );
buf ( n409187 , n62159 );
nand ( n62190 , n409186 , n409187 );
buf ( n409189 , n62190 );
buf ( n409190 , n409189 );
and ( n62193 , n409182 , n409190 );
buf ( n409192 , n62193 );
buf ( n409193 , n409192 );
xor ( n62196 , n409152 , n409193 );
buf ( n409195 , n59435 );
buf ( n409196 , n403146 );
and ( n62199 , n409195 , n409196 );
buf ( n409198 , n406565 );
buf ( n409199 , n401695 );
and ( n62202 , n409198 , n409199 );
nor ( n62203 , n62199 , n62202 );
buf ( n409202 , n62203 );
buf ( n409203 , n409202 );
buf ( n409204 , n403158 );
or ( n62207 , n409203 , n409204 );
buf ( n409206 , n406706 );
buf ( n409207 , n403167 );
or ( n62210 , n409206 , n409207 );
nand ( n62211 , n62207 , n62210 );
buf ( n409210 , n62211 );
buf ( n409211 , n409210 );
and ( n62214 , n62196 , n409211 );
and ( n62215 , n409152 , n409193 );
or ( n62216 , n62214 , n62215 );
buf ( n409215 , n62216 );
buf ( n409216 , n409215 );
and ( n62219 , n62131 , n409216 );
and ( n62220 , n409111 , n409128 );
or ( n62221 , n62219 , n62220 );
buf ( n409220 , n62221 );
xor ( n62223 , n406651 , n406668 );
xor ( n62224 , n62223 , n406686 );
buf ( n409223 , n62224 );
xor ( n62226 , n409220 , n409223 );
xor ( n62227 , n406576 , n406605 );
xor ( n62228 , n62227 , n406622 );
xor ( n62229 , n406734 , n59662 );
xor ( n62230 , n62228 , n62229 );
and ( n62231 , n62226 , n62230 );
and ( n62232 , n409220 , n409223 );
or ( n62233 , n62231 , n62232 );
xor ( n62234 , n59667 , n406797 );
xor ( n62235 , n62234 , n406801 );
and ( n62236 , n62233 , n62235 );
buf ( n409235 , n54297 );
buf ( n409236 , n59628 );
and ( n62239 , n409235 , n409236 );
buf ( n409238 , n55919 );
buf ( n409239 , n59457 );
and ( n62242 , n409238 , n409239 );
nor ( n62243 , n62239 , n62242 );
buf ( n409242 , n62243 );
buf ( n409243 , n409242 );
buf ( n409244 , n59637 );
or ( n62247 , n409243 , n409244 );
buf ( n409246 , n406762 );
buf ( n409247 , n59467 );
or ( n62250 , n409246 , n409247 );
nand ( n62251 , n62247 , n62250 );
buf ( n409250 , n62251 );
buf ( n409251 , n409250 );
buf ( n409252 , n59596 );
buf ( n409253 , n403146 );
and ( n62256 , n409252 , n409253 );
buf ( n409255 , n409146 );
buf ( n409256 , n401695 );
and ( n62259 , n409255 , n409256 );
nor ( n62260 , n62256 , n62259 );
buf ( n409259 , n62260 );
buf ( n409260 , n409259 );
not ( n62263 , n409260 );
buf ( n409262 , n62263 );
buf ( n409263 , n409262 );
buf ( n409264 , n401674 );
and ( n62267 , n409263 , n409264 );
buf ( n409266 , n409202 );
not ( n62269 , n409266 );
buf ( n409268 , n62269 );
buf ( n409269 , n409268 );
buf ( n409270 , n403164 );
and ( n62273 , n409269 , n409270 );
nor ( n62274 , n62267 , n62273 );
buf ( n409273 , n62274 );
buf ( n409274 , n409273 );
nand ( n62277 , n62135 , n53758 );
xnor ( n62278 , n54252 , n62277 );
buf ( n409277 , n62278 );
buf ( n409278 , n401626 );
and ( n62281 , n409277 , n409278 );
buf ( n409280 , n62139 );
buf ( n409281 , n401650 );
and ( n62284 , n409280 , n409281 );
nor ( n62285 , n62281 , n62284 );
buf ( n409284 , n62285 );
buf ( n409285 , n409284 );
nand ( n62288 , n409274 , n409285 );
buf ( n409287 , n62288 );
buf ( n409288 , n409287 );
xor ( n62291 , n409251 , n409288 );
buf ( n409290 , n55846 );
buf ( n409291 , n405391 );
and ( n62294 , n409290 , n409291 );
buf ( n409293 , n403079 );
buf ( n409294 , n405388 );
and ( n62297 , n409293 , n409294 );
nor ( n62298 , n62294 , n62297 );
buf ( n409297 , n62298 );
buf ( n409298 , n409297 );
buf ( n409299 , n405407 );
or ( n62302 , n409298 , n409299 );
buf ( n409301 , n406745 );
buf ( n409302 , n405384 );
or ( n62305 , n409301 , n409302 );
nand ( n62306 , n62302 , n62305 );
buf ( n409305 , n62306 );
buf ( n409306 , n409305 );
and ( n62309 , n62291 , n409306 );
and ( n62310 , n409251 , n409288 );
or ( n62311 , n62309 , n62310 );
buf ( n409310 , n62311 );
xor ( n62313 , n406753 , n406769 );
xor ( n62314 , n62313 , n406786 );
and ( n62315 , n409310 , n62314 );
buf ( n409314 , n55895 );
buf ( n409315 , n58201 );
and ( n62318 , n409314 , n409315 );
not ( n62319 , n409314 );
buf ( n409318 , n58200 );
and ( n62321 , n62319 , n409318 );
nor ( n62322 , n62318 , n62321 );
buf ( n409321 , n62322 );
buf ( n409322 , n409321 );
buf ( n409323 , n403120 );
or ( n62326 , n409322 , n409323 );
buf ( n409325 , n409119 );
buf ( n409326 , n403133 );
or ( n62329 , n409325 , n409326 );
nand ( n62330 , n62326 , n62329 );
buf ( n409329 , n62330 );
buf ( n409330 , n409329 );
buf ( n409331 , n58090 );
buf ( n409332 , n405215 );
and ( n62335 , n409331 , n409332 );
buf ( n409334 , n405335 );
buf ( n409335 , n58061 );
and ( n62338 , n409334 , n409335 );
nor ( n62339 , n62335 , n62338 );
buf ( n409338 , n62339 );
buf ( n409339 , n409338 );
buf ( n409340 , n403293 );
or ( n62343 , n409339 , n409340 );
buf ( n409342 , n406778 );
buf ( n409343 , n405476 );
or ( n62346 , n409342 , n409343 );
nand ( n62347 , n62343 , n62346 );
buf ( n409346 , n62347 );
buf ( n409347 , n409346 );
xor ( n62350 , n409330 , n409347 );
xor ( n62351 , n409152 , n409193 );
xor ( n62352 , n62351 , n409211 );
buf ( n409351 , n62352 );
buf ( n409352 , n409351 );
and ( n62355 , n62350 , n409352 );
and ( n62356 , n409330 , n409347 );
or ( n62357 , n62355 , n62356 );
buf ( n409356 , n62357 );
xor ( n62359 , n406753 , n406769 );
xor ( n409358 , n62359 , n406786 );
and ( n62361 , n409356 , n409358 );
and ( n62362 , n409310 , n409356 );
or ( n62363 , n62315 , n62361 , n62362 );
xor ( n62364 , n409220 , n409223 );
xor ( n62365 , n62364 , n62230 );
and ( n62366 , n62363 , n62365 );
buf ( n409365 , n55984 );
buf ( n409366 , n405391 );
and ( n62369 , n409365 , n409366 );
buf ( n409368 , n58135 );
buf ( n409369 , n405388 );
and ( n62372 , n409368 , n409369 );
nor ( n62373 , n62369 , n62372 );
buf ( n409372 , n62373 );
buf ( n409373 , n409372 );
buf ( n409374 , n405407 );
or ( n62377 , n409373 , n409374 );
buf ( n409376 , n409297 );
buf ( n409377 , n405384 );
or ( n62380 , n409376 , n409377 );
nand ( n62381 , n62377 , n62380 );
buf ( n409380 , n62381 );
buf ( n409381 , n54433 );
buf ( n409382 , n59628 );
and ( n62385 , n409381 , n409382 );
buf ( n409384 , n403088 );
buf ( n409385 , n59457 );
and ( n62388 , n409384 , n409385 );
nor ( n62389 , n62385 , n62388 );
buf ( n409388 , n62389 );
buf ( n409389 , n409388 );
buf ( n409390 , n59637 );
or ( n62393 , n409389 , n409390 );
buf ( n409392 , n409242 );
buf ( n409393 , n59467 );
or ( n62396 , n409392 , n409393 );
nand ( n62397 , n62393 , n62396 );
buf ( n409396 , n62397 );
xor ( n62399 , n409380 , n409396 );
buf ( n409398 , n58166 );
buf ( n409399 , n405215 );
and ( n62402 , n409398 , n409399 );
buf ( n409401 , n58205 );
buf ( n409402 , n58061 );
and ( n62405 , n409401 , n409402 );
nor ( n62406 , n62402 , n62405 );
buf ( n409405 , n62406 );
buf ( n409406 , n409405 );
buf ( n409407 , n403293 );
or ( n62410 , n409406 , n409407 );
buf ( n409409 , n409338 );
buf ( n409410 , n405476 );
or ( n62413 , n409409 , n409410 );
nand ( n62414 , n62410 , n62413 );
buf ( n409413 , n62414 );
and ( n62416 , n62399 , n409413 );
and ( n62417 , n409380 , n409396 );
or ( n62418 , n62416 , n62417 );
buf ( n409417 , n62418 );
buf ( n409418 , n54336 );
buf ( n409419 , n62177 );
and ( n62422 , n409418 , n409419 );
buf ( n409421 , n401699 );
buf ( n409422 , n62159 );
and ( n62425 , n409421 , n409422 );
nor ( n62426 , n62422 , n62425 );
buf ( n409425 , n62426 );
buf ( n409426 , n409425 );
buf ( n409427 , n409173 );
not ( n62430 , n409427 );
buf ( n409429 , n62430 );
buf ( n409430 , n409429 );
or ( n62433 , n409426 , n409430 );
buf ( n409432 , n409189 );
nand ( n62435 , n62433 , n409432 );
buf ( n409434 , n62435 );
buf ( n409435 , n409434 );
buf ( n409436 , n58352 );
buf ( n409437 , n55905 );
and ( n62440 , n409436 , n409437 );
buf ( n409439 , n406571 );
buf ( n409440 , n55895 );
and ( n62443 , n409439 , n409440 );
nor ( n62444 , n62440 , n62443 );
buf ( n409443 , n62444 );
buf ( n409444 , n409443 );
buf ( n409445 , n403120 );
or ( n62448 , n409444 , n409445 );
buf ( n409447 , n409321 );
buf ( n409448 , n403133 );
or ( n62451 , n409447 , n409448 );
nand ( n62452 , n62448 , n62451 );
buf ( n409451 , n62452 );
buf ( n409452 , n409451 );
xor ( n62455 , n409435 , n409452 );
not ( n62456 , n54250 );
nand ( n62457 , n62456 , n53917 );
not ( n62458 , n62457 );
nand ( n62459 , n54240 , n53895 );
not ( n62460 , n53910 );
or ( n62461 , n62459 , n62460 );
not ( n62462 , n54248 );
nand ( n62463 , n62461 , n62462 );
not ( n62464 , n62463 );
or ( n62465 , n62458 , n62464 );
or ( n62466 , n62457 , n62463 );
nand ( n62467 , n62465 , n62466 );
buf ( n409466 , n62467 );
not ( n62469 , n409466 );
buf ( n409468 , n62469 );
buf ( n409469 , n409468 );
buf ( n409470 , n403083 );
or ( n62473 , n409469 , n409470 );
buf ( n409472 , n62278 );
not ( n62475 , n409472 );
buf ( n409474 , n62475 );
buf ( n409475 , n409474 );
buf ( n409476 , n403092 );
or ( n62479 , n409475 , n409476 );
nand ( n62480 , n62473 , n62479 );
buf ( n409479 , n62480 );
buf ( n409480 , n409479 );
buf ( n409481 , n62164 );
buf ( n409482 , n5744 );
not ( n62485 , n409482 );
buf ( n409484 , n62485 );
buf ( n409485 , n409484 );
and ( n62488 , n409481 , n409485 );
not ( n62489 , n409481 );
buf ( n409488 , n5744 );
and ( n62491 , n62489 , n409488 );
nor ( n62492 , n62488 , n62491 );
buf ( n409491 , n62492 );
buf ( n409492 , n409491 );
not ( n62495 , n348348 );
not ( n62496 , n62495 );
nand ( n62497 , n409484 , n62496 );
buf ( n409496 , n62497 );
buf ( n62499 , n62495 );
buf ( n409498 , n62499 );
buf ( n409499 , n5744 );
nand ( n62502 , n409498 , n409499 );
buf ( n409501 , n62502 );
buf ( n409502 , n409501 );
and ( n62505 , n409496 , n409502 );
buf ( n409504 , n62505 );
buf ( n409505 , n409504 );
and ( n62508 , n409492 , n409505 );
buf ( n409507 , n62508 );
buf ( n409508 , n409507 );
not ( n62511 , n62164 );
buf ( n409510 , n62511 );
nand ( n62513 , n409508 , n409510 );
buf ( n409512 , n62513 );
buf ( n409513 , n409512 );
buf ( n409514 , n409504 );
not ( n62517 , n409514 );
buf ( n409516 , n62517 );
buf ( n409517 , n409516 );
buf ( n409518 , n62511 );
nand ( n62521 , n409517 , n409518 );
buf ( n409520 , n62521 );
buf ( n409521 , n409520 );
and ( n62524 , n409513 , n409521 );
buf ( n409523 , n62524 );
buf ( n409524 , n409523 );
xor ( n62527 , n409480 , n409524 );
buf ( n409526 , n62139 );
buf ( n409527 , n403146 );
and ( n62530 , n409526 , n409527 );
buf ( n409529 , n409140 );
buf ( n409530 , n401695 );
and ( n62533 , n409529 , n409530 );
nor ( n62534 , n62530 , n62533 );
buf ( n409533 , n62534 );
buf ( n409534 , n409533 );
buf ( n409535 , n403158 );
or ( n62538 , n409534 , n409535 );
buf ( n409537 , n409259 );
buf ( n409538 , n403167 );
or ( n62541 , n409537 , n409538 );
nand ( n62542 , n62538 , n62541 );
buf ( n409541 , n62542 );
buf ( n409542 , n409541 );
and ( n62545 , n62527 , n409542 );
and ( n62546 , n409480 , n409524 );
or ( n62547 , n62545 , n62546 );
buf ( n409546 , n62547 );
buf ( n409547 , n409546 );
and ( n62550 , n62455 , n409547 );
and ( n62551 , n409435 , n409452 );
or ( n62552 , n62550 , n62551 );
buf ( n409551 , n62552 );
buf ( n409552 , n409551 );
xor ( n62555 , n409417 , n409552 );
xor ( n62556 , n409251 , n409288 );
xor ( n62557 , n62556 , n409306 );
buf ( n409556 , n62557 );
buf ( n409557 , n409556 );
and ( n62560 , n62555 , n409557 );
and ( n62561 , n409417 , n409552 );
or ( n62562 , n62560 , n62561 );
buf ( n409561 , n62562 );
xor ( n62564 , n409111 , n409128 );
xor ( n62565 , n62564 , n409216 );
buf ( n409564 , n62565 );
xor ( n62567 , n409561 , n409564 );
xor ( n62568 , n406753 , n406769 );
xor ( n62569 , n62568 , n406786 );
xor ( n62570 , n409310 , n409356 );
xor ( n62571 , n62569 , n62570 );
and ( n62572 , n62567 , n62571 );
and ( n62573 , n409561 , n409564 );
or ( n62574 , n62572 , n62573 );
xor ( n62575 , n409220 , n409223 );
xor ( n62576 , n62575 , n62230 );
and ( n62577 , n62574 , n62576 );
and ( n62578 , n62363 , n62574 );
or ( n62579 , n62366 , n62577 , n62578 );
xor ( n62580 , n59667 , n406797 );
xor ( n62581 , n62580 , n406801 );
and ( n62582 , n62579 , n62581 );
and ( n62583 , n62233 , n62579 );
or ( n62584 , n62236 , n62582 , n62583 );
buf ( n409583 , n62584 );
nand ( n62586 , n62106 , n409583 );
buf ( n409585 , n62586 );
buf ( n409586 , n409585 );
buf ( n409587 , n62104 );
buf ( n409588 , n62073 );
nand ( n62591 , n409587 , n409588 );
buf ( n409590 , n62591 );
buf ( n409591 , n409590 );
nand ( n62594 , n409586 , n409591 );
buf ( n409593 , n62594 );
buf ( n409594 , n409593 );
xor ( n62597 , n409067 , n409594 );
xor ( n62598 , n407920 , n60892 );
xnor ( n62599 , n62598 , n407952 );
buf ( n409598 , n62599 );
and ( n62601 , n62597 , n409598 );
and ( n62602 , n409067 , n409594 );
or ( n62603 , n62601 , n62602 );
buf ( n409602 , n62603 );
buf ( n409603 , n409602 );
nand ( n62606 , n62052 , n409603 );
buf ( n409605 , n62606 );
buf ( n409606 , n409605 );
buf ( n409607 , n409044 );
buf ( n409608 , n409018 );
not ( n62611 , n409608 );
buf ( n409610 , n62611 );
buf ( n409611 , n409610 );
nand ( n62614 , n409607 , n409611 );
buf ( n409613 , n62614 );
buf ( n409614 , n409613 );
nand ( n62617 , n409606 , n409614 );
buf ( n409616 , n62617 );
buf ( n409617 , n409616 );
buf ( n409618 , n43536 );
not ( n62621 , n409618 );
buf ( n409620 , n391027 );
not ( n62623 , n409620 );
buf ( n409622 , n389805 );
not ( n62625 , n409622 );
or ( n62626 , n62623 , n62625 );
buf ( n409625 , n385342 );
buf ( n409626 , n391024 );
nand ( n62629 , n409625 , n409626 );
buf ( n409628 , n62629 );
buf ( n409629 , n409628 );
nand ( n62632 , n62626 , n409629 );
buf ( n409631 , n62632 );
buf ( n409632 , n409631 );
not ( n62635 , n409632 );
or ( n62636 , n62621 , n62635 );
buf ( n409635 , n408384 );
buf ( n409636 , n43515 );
nand ( n62639 , n409635 , n409636 );
buf ( n409638 , n62639 );
buf ( n409639 , n409638 );
nand ( n62642 , n62636 , n409639 );
buf ( n409641 , n62642 );
buf ( n409642 , n409641 );
xor ( n62645 , n409617 , n409642 );
buf ( n409644 , n61429 );
buf ( n409645 , n388809 );
and ( n62648 , n409644 , n409645 );
buf ( n409647 , n405736 );
not ( n62650 , n409647 );
buf ( n409649 , n28215 );
not ( n62652 , n409649 );
or ( n62653 , n62650 , n62652 );
buf ( n409652 , n375822 );
buf ( n409653 , n388754 );
nand ( n62656 , n409652 , n409653 );
buf ( n409655 , n62656 );
buf ( n409656 , n409655 );
nand ( n62659 , n62653 , n409656 );
buf ( n409658 , n62659 );
buf ( n409659 , n409658 );
not ( n62662 , n409659 );
buf ( n409661 , n388743 );
nor ( n62664 , n62662 , n409661 );
buf ( n409663 , n62664 );
buf ( n409664 , n409663 );
nor ( n62667 , n62648 , n409664 );
buf ( n409666 , n62667 );
buf ( n409667 , n409666 );
not ( n62670 , n409667 );
buf ( n409669 , n43058 );
not ( n62672 , n409669 );
buf ( n409671 , n393562 );
not ( n62674 , n409671 );
buf ( n409673 , n392620 );
not ( n62676 , n409673 );
and ( n62677 , n62674 , n62676 );
buf ( n409676 , n393117 );
buf ( n409677 , n392620 );
and ( n62680 , n409676 , n409677 );
nor ( n62681 , n62677 , n62680 );
buf ( n409680 , n62681 );
buf ( n409681 , n409680 );
not ( n62684 , n409681 );
and ( n62685 , n62672 , n62684 );
buf ( n409684 , n407988 );
buf ( n409685 , n398665 );
nor ( n62688 , n409684 , n409685 );
buf ( n409687 , n62688 );
buf ( n409688 , n409687 );
nor ( n62691 , n62685 , n409688 );
buf ( n409690 , n62691 );
buf ( n409691 , n409690 );
not ( n62694 , n409691 );
or ( n62695 , n62670 , n62694 );
buf ( n409694 , n40990 );
not ( n62697 , n409694 );
buf ( n409696 , n399164 );
not ( n62699 , n409696 );
or ( n62700 , n62697 , n62699 );
buf ( n409699 , n24049 );
buf ( n409700 , n390460 );
nand ( n62703 , n409699 , n409700 );
buf ( n409702 , n62703 );
buf ( n409703 , n409702 );
nand ( n62706 , n62700 , n409703 );
buf ( n409705 , n62706 );
buf ( n409706 , n409705 );
not ( n62709 , n409706 );
buf ( n409708 , n396622 );
not ( n62711 , n409708 );
or ( n62712 , n62709 , n62711 );
buf ( n409711 , n408443 );
buf ( n409712 , n55831 );
nand ( n62715 , n409711 , n409712 );
buf ( n409714 , n62715 );
buf ( n409715 , n409714 );
nand ( n62718 , n62712 , n409715 );
buf ( n409717 , n62718 );
buf ( n409718 , n409717 );
not ( n62721 , n409718 );
buf ( n409720 , n389359 );
not ( n62723 , n409720 );
buf ( n409722 , n45102 );
not ( n62725 , n409722 );
or ( n62726 , n62723 , n62725 );
buf ( n409725 , n22982 );
buf ( n409726 , n389356 );
nand ( n62729 , n409725 , n409726 );
buf ( n409728 , n62729 );
buf ( n409729 , n409728 );
nand ( n62732 , n62726 , n409729 );
buf ( n409731 , n62732 );
buf ( n409732 , n409731 );
not ( n62735 , n409732 );
buf ( n409734 , n399031 );
not ( n62737 , n409734 );
or ( n62738 , n62735 , n62737 );
buf ( n409737 , n407873 );
buf ( n409738 , n395469 );
nand ( n62741 , n409737 , n409738 );
buf ( n409740 , n62741 );
buf ( n409741 , n409740 );
nand ( n62744 , n62738 , n409741 );
buf ( n409743 , n62744 );
buf ( n409744 , n409743 );
not ( n62747 , n409744 );
or ( n62748 , n62721 , n62747 );
buf ( n409747 , n409743 );
buf ( n409748 , n409717 );
or ( n62751 , n409747 , n409748 );
buf ( n409750 , n57569 );
not ( n62753 , n409750 );
buf ( n409752 , n24116 );
not ( n62755 , n409752 );
buf ( n409754 , n45699 );
not ( n62757 , n409754 );
or ( n62758 , n62755 , n62757 );
buf ( n409757 , n388643 );
buf ( n409758 , n62006 );
nand ( n62761 , n409757 , n409758 );
buf ( n409760 , n62761 );
buf ( n409761 , n409760 );
nand ( n62764 , n62758 , n409761 );
buf ( n409763 , n62764 );
buf ( n409764 , n409763 );
not ( n62767 , n409764 );
or ( n62768 , n62753 , n62767 );
buf ( n409767 , n389162 );
buf ( n409768 , n409010 );
nand ( n62771 , n409767 , n409768 );
buf ( n409770 , n62771 );
buf ( n409771 , n409770 );
nand ( n62774 , n62768 , n409771 );
buf ( n409773 , n62774 );
buf ( n409774 , n409773 );
nand ( n62777 , n62751 , n409774 );
buf ( n409776 , n62777 );
buf ( n409777 , n409776 );
nand ( n62780 , n62748 , n409777 );
buf ( n409779 , n62780 );
buf ( n409780 , n409779 );
nand ( n62783 , n62695 , n409780 );
buf ( n409782 , n62783 );
buf ( n409783 , n409782 );
or ( n62786 , n409690 , n409666 );
buf ( n409785 , n62786 );
nand ( n62788 , n409783 , n409785 );
buf ( n409787 , n62788 );
buf ( n409788 , n409787 );
and ( n62791 , n62645 , n409788 );
and ( n62792 , n409617 , n409642 );
or ( n62793 , n62791 , n62792 );
buf ( n409792 , n62793 );
buf ( n409793 , n409792 );
xor ( n62796 , n407818 , n407835 );
xor ( n62797 , n62796 , n407999 );
buf ( n409796 , n62797 );
buf ( n409797 , n409796 );
xor ( n62800 , n409793 , n409797 );
xor ( n62801 , n407861 , n407978 );
xor ( n62802 , n62801 , n407994 );
buf ( n409801 , n62802 );
buf ( n409802 , n409801 );
xor ( n62805 , n408431 , n408456 );
xor ( n62806 , n62805 , n408461 );
buf ( n409805 , n62806 );
buf ( n409806 , n409805 );
xor ( n62809 , n60895 , n407885 );
xor ( n62810 , n62809 , n407911 );
buf ( n409809 , n62810 );
xor ( n62812 , n409806 , n409809 );
buf ( n409811 , n394210 );
not ( n62814 , n409811 );
buf ( n409813 , n388299 );
not ( n62816 , n409813 );
or ( n62817 , n62814 , n62816 );
buf ( n409816 , n400355 );
buf ( n409817 , n394219 );
nand ( n62820 , n409816 , n409817 );
buf ( n409819 , n62820 );
buf ( n409820 , n409819 );
nand ( n62823 , n62817 , n409820 );
buf ( n409822 , n62823 );
buf ( n409823 , n409822 );
not ( n62826 , n409823 );
buf ( n409825 , n383891 );
not ( n62828 , n409825 );
or ( n62829 , n62826 , n62828 );
buf ( n409828 , n408243 );
not ( n62831 , n409828 );
buf ( n409830 , n388629 );
nand ( n62833 , n62831 , n409830 );
buf ( n409832 , n62833 );
buf ( n409833 , n409832 );
nand ( n62836 , n62829 , n409833 );
buf ( n409835 , n62836 );
buf ( n409836 , n409835 );
and ( n62839 , n62812 , n409836 );
and ( n62840 , n409806 , n409809 );
or ( n62841 , n62839 , n62840 );
buf ( n409840 , n62841 );
buf ( n409841 , n409840 );
xor ( n62844 , n409802 , n409841 );
xor ( n62845 , n408466 , n408479 );
xor ( n62846 , n62845 , n408485 );
buf ( n409845 , n62846 );
buf ( n409846 , n409845 );
and ( n62849 , n62844 , n409846 );
and ( n62850 , n409802 , n409841 );
or ( n62851 , n62849 , n62850 );
buf ( n409850 , n62851 );
buf ( n409851 , n409850 );
and ( n62854 , n62800 , n409851 );
and ( n62855 , n409793 , n409797 );
or ( n62856 , n62854 , n62855 );
buf ( n409855 , n62856 );
buf ( n409856 , n409855 );
nand ( n62859 , n61996 , n409856 );
buf ( n409858 , n62859 );
nand ( n62861 , C1 , n409858 );
and ( n62862 , n61966 , n62861 );
and ( n62863 , n61809 , n61965 );
or ( n62864 , n62862 , n62863 );
buf ( n409863 , n62864 );
not ( n62866 , n409863 );
buf ( n409865 , n407069 );
buf ( n409866 , n407092 );
and ( n62869 , n409865 , n409866 );
not ( n62870 , n409865 );
buf ( n409869 , n407103 );
and ( n62872 , n62870 , n409869 );
nor ( n62873 , n62869 , n62872 );
buf ( n409872 , n62873 );
and ( n62875 , n409872 , n59995 );
not ( n62876 , n409872 );
not ( n62877 , n59995 );
and ( n62878 , n62876 , n62877 );
nor ( n62879 , n62875 , n62878 );
buf ( n409878 , n62879 );
xor ( n62881 , n407352 , n407355 );
xor ( n62882 , n62881 , n407397 );
buf ( n409881 , n62882 );
buf ( n409882 , n409881 );
xor ( n62885 , n409878 , n409882 );
buf ( n409884 , n395349 );
not ( n62887 , n409884 );
buf ( n409886 , n61601 );
not ( n62889 , n409886 );
or ( n62890 , n62887 , n62889 );
nand ( n62891 , n60266 , n395362 );
buf ( n409890 , n62891 );
nand ( n62893 , n62890 , n409890 );
buf ( n409892 , n62893 );
buf ( n409893 , n409892 );
not ( n62896 , n407428 );
xor ( n62897 , n60350 , n62896 );
xnor ( n62898 , n62897 , n407527 );
buf ( n409897 , n62898 );
xor ( n62900 , n409893 , n409897 );
buf ( n409899 , n407574 );
not ( n62902 , n409899 );
buf ( n409901 , n407605 );
not ( n62904 , n409901 );
or ( n62905 , n62902 , n62904 );
buf ( n409904 , n407594 );
buf ( n409905 , n407600 );
nand ( n62908 , n409904 , n409905 );
buf ( n409907 , n62908 );
buf ( n409908 , n409907 );
nand ( n62911 , n62905 , n409908 );
buf ( n409910 , n62911 );
buf ( n409911 , n409910 );
buf ( n409912 , n407678 );
and ( n62915 , n409911 , n409912 );
not ( n62916 , n409911 );
buf ( n409915 , n407678 );
not ( n62918 , n409915 );
buf ( n409917 , n62918 );
buf ( n409918 , n409917 );
and ( n62921 , n62916 , n409918 );
nor ( n62922 , n62915 , n62921 );
buf ( n409921 , n62922 );
buf ( n409922 , n409921 );
and ( n62925 , n62900 , n409922 );
and ( n62926 , n409893 , n409897 );
or ( n62927 , n62925 , n62926 );
buf ( n409926 , n62927 );
buf ( n409927 , n409926 );
and ( n62930 , n62885 , n409927 );
and ( n62931 , n409878 , n409882 );
or ( n62932 , n62930 , n62931 );
buf ( n409931 , n62932 );
buf ( n409932 , n409931 );
not ( n62935 , n409932 );
and ( n62936 , n408058 , n61027 );
not ( n62937 , n408058 );
and ( n62938 , n62937 , n61028 );
nor ( n62939 , n62936 , n62938 );
and ( n62940 , n62939 , n61032 );
not ( n62941 , n62939 );
not ( n62942 , n61032 );
and ( n62943 , n62941 , n62942 );
nor ( n62944 , n62940 , n62943 );
buf ( n409943 , n62944 );
not ( n62946 , n409943 );
buf ( n409945 , n62946 );
buf ( n409946 , n409945 );
nand ( n62949 , n62935 , n409946 );
buf ( n409948 , n62949 );
buf ( n409949 , n409948 );
not ( n62952 , n409949 );
or ( n62953 , n62866 , n62952 );
buf ( n409952 , n409931 );
buf ( n409953 , n62944 );
nand ( n62956 , n409952 , n409953 );
buf ( n409955 , n62956 );
buf ( n409956 , n409955 );
nand ( n62959 , n62953 , n409956 );
buf ( n409958 , n62959 );
buf ( n409959 , n409958 );
nand ( n62962 , n61807 , n409959 );
buf ( n409961 , n62962 );
nand ( n62964 , n61803 , n61558 );
nand ( n62965 , n409961 , n62964 );
nand ( n62966 , n61556 , n62965 );
nand ( n62967 , n61550 , n62966 );
not ( n62968 , n62967 );
nand ( n62969 , n408549 , n62968 );
buf ( n409968 , n62969 );
and ( n62971 , n408543 , n409968 );
buf ( n409970 , n62971 );
xor ( n62973 , n56735 , n57214 );
xnor ( n62974 , n62973 , n57219 );
buf ( n409973 , n62974 );
xor ( n62976 , n406985 , n406988 );
and ( n62977 , n62976 , n60624 );
and ( n62978 , n406985 , n406988 );
or ( n62979 , n62977 , n62978 );
buf ( n409978 , n62979 );
xor ( n62981 , n409973 , n409978 );
xor ( n62982 , n404890 , n404894 );
xor ( n62983 , n62982 , n405592 );
buf ( n409982 , n62983 );
buf ( n409983 , n409982 );
xor ( n62986 , n62981 , n409983 );
buf ( n409985 , n62986 );
buf ( n409986 , n409985 );
not ( n62989 , n409986 );
buf ( n409988 , n62989 );
xor ( n62991 , n58490 , n406979 );
and ( n62992 , n62991 , n60625 );
and ( n62993 , n58490 , n406979 );
or ( n62994 , n62992 , n62993 );
buf ( n409993 , n62994 );
not ( n62996 , n409993 );
buf ( n409995 , n62996 );
nand ( n62998 , n409988 , n409995 );
buf ( n409997 , n62998 );
buf ( n63000 , n409997 );
buf ( n409999 , n63000 );
xor ( n63002 , n58450 , n405596 );
xnor ( n63003 , n63002 , n58460 );
buf ( n410002 , n63003 );
not ( n63005 , n410002 );
buf ( n410004 , n63005 );
buf ( n410005 , n410004 );
xor ( n63008 , n409973 , n409978 );
and ( n63009 , n63008 , n409983 );
and ( n63010 , n409973 , n409978 );
or ( n63011 , n63009 , n63010 );
buf ( n410010 , n63011 );
buf ( n410011 , n410010 );
not ( n63014 , n410011 );
buf ( n410013 , n63014 );
buf ( n410014 , n410013 );
nand ( n63017 , n410005 , n410014 );
buf ( n410016 , n63017 );
and ( n63019 , n409970 , n409999 , n410016 );
xor ( n63020 , n409893 , n409897 );
xor ( n63021 , n63020 , n409922 );
buf ( n410020 , n63021 );
xor ( n63023 , n408392 , n408417 );
xor ( n63024 , n63023 , n408490 );
buf ( n410023 , n63024 );
not ( n63026 , n410023 );
xor ( n63027 , n408230 , n408294 );
xor ( n63028 , n63027 , n408320 );
buf ( n410027 , n63028 );
not ( n63030 , n410027 );
or ( n63031 , n63026 , n63030 );
buf ( n410030 , n410023 );
buf ( n410031 , n410027 );
or ( n63034 , n410030 , n410031 );
buf ( n410033 , n61248 );
buf ( n410034 , n61232 );
xor ( n63037 , n410033 , n410034 );
buf ( n410036 , n408257 );
xor ( n63039 , n63037 , n410036 );
buf ( n410038 , n63039 );
buf ( n410039 , n410038 );
buf ( n410040 , n393825 );
not ( n63043 , n410040 );
buf ( n410042 , n393369 );
not ( n63045 , n410042 );
buf ( n410044 , n389467 );
not ( n63047 , n410044 );
or ( n63048 , n63045 , n63047 );
buf ( n410047 , n384974 );
buf ( n410048 , n393384 );
nand ( n63051 , n410047 , n410048 );
buf ( n410050 , n63051 );
buf ( n410051 , n410050 );
nand ( n63054 , n63048 , n410051 );
buf ( n410053 , n63054 );
buf ( n410054 , n410053 );
not ( n63057 , n410054 );
or ( n63058 , n63043 , n63057 );
buf ( n410057 , n61837 );
not ( n63060 , n410057 );
buf ( n410059 , n45954 );
nand ( n63062 , n63060 , n410059 );
buf ( n410061 , n63062 );
buf ( n410062 , n410061 );
nand ( n63065 , n63058 , n410062 );
buf ( n410064 , n63065 );
buf ( n410065 , n410064 );
xor ( n63068 , n410039 , n410065 );
buf ( n410067 , n61228 );
not ( n63070 , n410067 );
buf ( n410069 , n390362 );
not ( n63072 , n410069 );
or ( n63073 , n63070 , n63072 );
buf ( n410072 , n388102 );
not ( n63075 , n410072 );
buf ( n410074 , n40777 );
not ( n63077 , n410074 );
or ( n63078 , n63075 , n63077 );
buf ( n410077 , n40758 );
buf ( n410078 , n40600 );
nand ( n63081 , n410077 , n410078 );
buf ( n410080 , n63081 );
buf ( n410081 , n410080 );
nand ( n63084 , n63078 , n410081 );
buf ( n410083 , n63084 );
buf ( n410084 , n410083 );
buf ( n410085 , n43286 );
nand ( n63088 , n410084 , n410085 );
buf ( n410087 , n63088 );
buf ( n410088 , n410087 );
nand ( n63091 , n63073 , n410088 );
buf ( n410090 , n63091 );
not ( n63093 , n410090 );
buf ( n410092 , n63093 );
not ( n63095 , n410092 );
buf ( n410094 , n384008 );
not ( n63097 , n410094 );
buf ( n410096 , n40839 );
not ( n63099 , n410096 );
buf ( n410098 , n49124 );
not ( n63101 , n410098 );
and ( n63102 , n63099 , n63101 );
buf ( n410101 , n40840 );
buf ( n410102 , n49124 );
and ( n63105 , n410101 , n410102 );
nor ( n63106 , n63102 , n63105 );
buf ( n410105 , n63106 );
buf ( n410106 , n410105 );
not ( n63109 , n410106 );
and ( n63110 , n63097 , n63109 );
buf ( n410109 , n408897 );
buf ( n410110 , n383943 );
nor ( n63113 , n410109 , n410110 );
buf ( n410112 , n63113 );
buf ( n410113 , n410112 );
nor ( n63116 , n63110 , n410113 );
buf ( n410115 , n63116 );
buf ( n410116 , n410115 );
not ( n63119 , n410116 );
or ( n63120 , n63095 , n63119 );
buf ( n410119 , n388502 );
not ( n63122 , n410119 );
buf ( n410121 , n51822 );
not ( n63124 , n410121 );
or ( n63125 , n63122 , n63124 );
buf ( n410124 , n24070 );
buf ( n410125 , n388502 );
not ( n63128 , n410125 );
buf ( n410127 , n63128 );
buf ( n410128 , n410127 );
nand ( n63131 , n410124 , n410128 );
buf ( n410130 , n63131 );
buf ( n410131 , n410130 );
nand ( n63134 , n63125 , n410131 );
buf ( n410133 , n63134 );
buf ( n410134 , n410133 );
not ( n63137 , n410134 );
buf ( n410136 , n52812 );
not ( n63139 , n410136 );
or ( n63140 , n63137 , n63139 );
buf ( n410139 , n60884 );
buf ( n410140 , n400143 );
nand ( n63143 , n410139 , n410140 );
buf ( n410142 , n63143 );
buf ( n410143 , n410142 );
nand ( n63146 , n63140 , n410143 );
buf ( n410145 , n63146 );
buf ( n410146 , n410145 );
buf ( n410147 , n388830 );
not ( n63150 , n410147 );
buf ( n410149 , n62061 );
not ( n63152 , n410149 );
or ( n63153 , n63150 , n63152 );
and ( n63154 , n28644 , n45897 );
not ( n63155 , n28644 );
and ( n63156 , n63155 , n41342 );
or ( n63157 , n63154 , n63156 );
buf ( n410156 , n63157 );
buf ( n410157 , n388872 );
nand ( n63160 , n410156 , n410157 );
buf ( n410159 , n63160 );
buf ( n410160 , n410159 );
nand ( n63163 , n63153 , n410160 );
buf ( n410162 , n63163 );
buf ( n410163 , n410162 );
xor ( n63166 , n410146 , n410163 );
buf ( n410165 , n62584 );
buf ( n410166 , n62073 );
xnor ( n63169 , n410165 , n410166 );
buf ( n410168 , n63169 );
buf ( n410169 , n410168 );
not ( n63172 , n410169 );
buf ( n410171 , n62104 );
not ( n63174 , n410171 );
or ( n63175 , n63172 , n63174 );
buf ( n410174 , n62104 );
buf ( n410175 , n410168 );
or ( n63178 , n410174 , n410175 );
nand ( n63179 , n63175 , n63178 );
buf ( n410178 , n63179 );
buf ( n410179 , n410178 );
and ( n63182 , n63166 , n410179 );
and ( n63183 , n410146 , n410163 );
or ( n63184 , n63182 , n63183 );
buf ( n410183 , n63184 );
buf ( n410184 , n410183 );
buf ( n410185 , n388809 );
not ( n63188 , n410185 );
buf ( n410187 , n409658 );
not ( n63190 , n410187 );
or ( n63191 , n63188 , n63190 );
buf ( n410190 , n405736 );
not ( n63193 , n410190 );
buf ( n410192 , n388409 );
not ( n63195 , n410192 );
or ( n63196 , n63193 , n63195 );
buf ( n410195 , n388406 );
buf ( n410196 , n388754 );
nand ( n63199 , n410195 , n410196 );
buf ( n410198 , n63199 );
buf ( n410199 , n410198 );
nand ( n63202 , n63196 , n410199 );
buf ( n410201 , n63202 );
buf ( n410202 , n410201 );
buf ( n410203 , n388746 );
nand ( n63206 , n410202 , n410203 );
buf ( n410205 , n63206 );
buf ( n410206 , n410205 );
nand ( n63209 , n63191 , n410206 );
buf ( n410208 , n63209 );
buf ( n410209 , n410208 );
xor ( n63212 , n410184 , n410209 );
buf ( n410211 , n385473 );
not ( n63214 , n410211 );
buf ( n410213 , n391443 );
not ( n63216 , n410213 );
and ( n63217 , n63214 , n63216 );
buf ( n410216 , n385473 );
buf ( n410217 , n391443 );
and ( n63220 , n410216 , n410217 );
nor ( n63221 , n63217 , n63220 );
buf ( n410220 , n63221 );
buf ( n410221 , n410220 );
not ( n63224 , n410221 );
buf ( n410223 , n63224 );
buf ( n410224 , n410223 );
not ( n63227 , n410224 );
buf ( n410226 , n393544 );
not ( n63229 , n410226 );
or ( n63230 , n63227 , n63229 );
buf ( n410229 , n409032 );
buf ( n410230 , n49166 );
nand ( n63233 , n410229 , n410230 );
buf ( n410232 , n63233 );
buf ( n410233 , n410232 );
nand ( n63236 , n63230 , n410233 );
buf ( n410235 , n63236 );
buf ( n410236 , n410235 );
and ( n63239 , n63212 , n410236 );
and ( n63240 , n410184 , n410209 );
or ( n63241 , n63239 , n63240 );
buf ( n410240 , n63241 );
buf ( n410241 , n410240 );
nand ( n63244 , n63120 , n410241 );
buf ( n410243 , n63244 );
buf ( n410244 , n410243 );
buf ( n410245 , n410115 );
not ( n63248 , n410245 );
buf ( n410247 , n410090 );
nand ( n63250 , n63248 , n410247 );
buf ( n410249 , n63250 );
buf ( n410250 , n410249 );
nand ( n63253 , n410244 , n410250 );
buf ( n410252 , n63253 );
buf ( n410253 , n410252 );
and ( n63256 , n63068 , n410253 );
and ( n63257 , n410039 , n410065 );
or ( n63258 , n63256 , n63257 );
buf ( n410257 , n63258 );
buf ( n410258 , n410257 );
nand ( n63261 , n63034 , n410258 );
buf ( n410260 , n63261 );
nand ( n63263 , n63031 , n410260 );
xor ( n63264 , n410020 , n63263 );
xor ( n63265 , n408366 , n408369 );
xor ( n63266 , n63265 , n408494 );
xor ( n63267 , n63264 , n63266 );
buf ( n410266 , n63267 );
xor ( n63269 , n409802 , n409841 );
xor ( n63270 , n63269 , n409846 );
buf ( n410269 , n63270 );
buf ( n410270 , n410269 );
xor ( n63273 , n409806 , n409809 );
xor ( n63274 , n63273 , n409836 );
buf ( n410273 , n63274 );
buf ( n410274 , n410273 );
buf ( n410275 , n358975 );
buf ( n410276 , n385729 );
and ( n63279 , n410275 , n410276 );
not ( n63280 , n410275 );
buf ( n410279 , n383426 );
and ( n63282 , n63280 , n410279 );
nor ( n63283 , n63279 , n63282 );
buf ( n410282 , n63283 );
buf ( n410283 , n410282 );
not ( n63286 , n410283 );
buf ( n410285 , n391917 );
not ( n63288 , n410285 );
or ( n63289 , n63286 , n63288 );
buf ( n410288 , n393903 );
buf ( n410289 , n408754 );
nand ( n63292 , n410288 , n410289 );
buf ( n410291 , n63292 );
buf ( n410292 , n410291 );
nand ( n63295 , n63289 , n410292 );
buf ( n410294 , n63295 );
buf ( n410295 , n410294 );
xor ( n63298 , n410274 , n410295 );
buf ( n410297 , n394817 );
not ( n63300 , n410297 );
buf ( n410299 , n388299 );
not ( n63302 , n410299 );
or ( n63303 , n63300 , n63302 );
buf ( n410302 , n388608 );
buf ( n410303 , n394814 );
nand ( n63306 , n410302 , n410303 );
buf ( n410305 , n63306 );
buf ( n410306 , n410305 );
nand ( n63309 , n63303 , n410306 );
buf ( n410308 , n63309 );
buf ( n410309 , n410308 );
not ( n63312 , n410309 );
buf ( n410311 , n383894 );
not ( n63314 , n410311 );
or ( n63315 , n63312 , n63314 );
buf ( n410314 , n409822 );
buf ( n410315 , n383907 );
nand ( n63318 , n410314 , n410315 );
buf ( n410317 , n63318 );
buf ( n410318 , n410317 );
nand ( n63321 , n63315 , n410318 );
buf ( n410320 , n63321 );
buf ( n410321 , n410320 );
not ( n63324 , n389162 );
not ( n63325 , n409763 );
or ( n63326 , n63324 , n63325 );
not ( n63327 , n41710 );
buf ( n410326 , n389856 );
not ( n63329 , n410326 );
buf ( n410328 , n24116 );
not ( n63331 , n410328 );
or ( n63332 , n63329 , n63331 );
buf ( n410331 , n49686 );
buf ( n410332 , n62006 );
nand ( n63335 , n410331 , n410332 );
buf ( n410334 , n63335 );
buf ( n410335 , n410334 );
nand ( n63338 , n63332 , n410335 );
buf ( n410337 , n63338 );
nand ( n63340 , n63327 , n410337 );
nand ( n63341 , n63326 , n63340 );
not ( n63342 , n63341 );
buf ( n410341 , n63342 );
not ( n63344 , n410341 );
not ( n63345 , n46062 );
not ( n63346 , n410220 );
and ( n63347 , n63345 , n63346 );
buf ( n410346 , n392611 );
not ( n63349 , n410346 );
buf ( n410348 , n388965 );
not ( n63351 , n410348 );
or ( n63352 , n63349 , n63351 );
buf ( n410351 , n385473 );
buf ( n410352 , n392620 );
nand ( n63355 , n410351 , n410352 );
buf ( n410354 , n63355 );
buf ( n410355 , n410354 );
nand ( n63358 , n63352 , n410355 );
buf ( n410357 , n63358 );
not ( n63360 , n410357 );
nor ( n63361 , n63360 , n391550 );
nor ( n63362 , n63347 , n63361 );
buf ( n410361 , n63362 );
not ( n63364 , n410361 );
or ( n63365 , n63344 , n63364 );
xor ( n63366 , n59667 , n406797 );
xor ( n63367 , n63366 , n406801 );
xor ( n63368 , n62233 , n62579 );
xor ( n63369 , n63367 , n63368 );
buf ( n410368 , n63369 );
buf ( n410369 , n12480 );
buf ( n410370 , n388192 );
and ( n63373 , n410369 , n410370 );
not ( n63374 , n410369 );
buf ( n410373 , n409092 );
and ( n63376 , n63374 , n410373 );
nor ( n63377 , n63373 , n63376 );
buf ( n410376 , n63377 );
buf ( n410377 , n410376 );
not ( n63380 , n410377 );
buf ( n410379 , n60872 );
not ( n63382 , n410379 );
or ( n63383 , n63380 , n63382 );
buf ( n410382 , n409098 );
buf ( n410383 , n47726 );
nand ( n63386 , n410382 , n410383 );
buf ( n410385 , n63386 );
buf ( n410386 , n410385 );
nand ( n63389 , n63383 , n410386 );
buf ( n410388 , n63389 );
buf ( n410389 , n410388 );
xor ( n63392 , n410368 , n410389 );
buf ( n410391 , n388830 );
not ( n63394 , n410391 );
buf ( n410393 , n63157 );
not ( n63396 , n410393 );
or ( n63397 , n63394 , n63396 );
buf ( n410396 , n41342 );
not ( n63399 , n410396 );
buf ( n410398 , n12471 );
not ( n63401 , n410398 );
buf ( n410400 , n63401 );
buf ( n410401 , n410400 );
not ( n63404 , n410401 );
or ( n63405 , n63399 , n63404 );
buf ( n410404 , n12471 );
buf ( n410405 , n23840 );
buf ( n63408 , n410405 );
buf ( n410407 , n63408 );
buf ( n410408 , n410407 );
nand ( n63411 , n410404 , n410408 );
buf ( n410410 , n63411 );
buf ( n410411 , n410410 );
nand ( n63414 , n63405 , n410411 );
buf ( n410413 , n63414 );
nand ( n63416 , n410413 , n41373 );
buf ( n410415 , n63416 );
nand ( n63418 , n63397 , n410415 );
buf ( n410417 , n63418 );
buf ( n410418 , n410417 );
xor ( n63421 , n63392 , n410418 );
buf ( n410420 , n63421 );
not ( n63423 , n410420 );
buf ( n410422 , n40990 );
not ( n63425 , n410422 );
buf ( n410424 , n51822 );
not ( n63427 , n410424 );
or ( n63428 , n63425 , n63427 );
buf ( n410427 , n41559 );
buf ( n410428 , n390460 );
nand ( n63431 , n410427 , n410428 );
buf ( n410430 , n63431 );
buf ( n410431 , n410430 );
nand ( n63434 , n63428 , n410431 );
buf ( n410433 , n63434 );
buf ( n410434 , n410433 );
not ( n63437 , n410434 );
buf ( n410436 , n390429 );
not ( n63439 , n410436 );
or ( n63440 , n63437 , n63439 );
buf ( n410439 , n410133 );
buf ( n410440 , n400143 );
nand ( n63443 , n410439 , n410440 );
buf ( n410442 , n63443 );
buf ( n410443 , n410442 );
nand ( n63446 , n63440 , n410443 );
buf ( n410445 , n63446 );
buf ( n410446 , n410445 );
not ( n63449 , n410446 );
xor ( n63450 , n409220 , n409223 );
xor ( n63451 , n63450 , n62230 );
xor ( n63452 , n62363 , n62574 );
xor ( n63453 , n63451 , n63452 );
buf ( n410452 , n63453 );
buf ( n410453 , n58200 );
buf ( n410454 , n405215 );
and ( n63457 , n410453 , n410454 );
buf ( n410456 , n58201 );
buf ( n410457 , n58061 );
and ( n63460 , n410456 , n410457 );
nor ( n63461 , n63457 , n63460 );
buf ( n410460 , n63461 );
buf ( n410461 , n410460 );
buf ( n410462 , n403293 );
or ( n63465 , n410461 , n410462 );
buf ( n410464 , n409405 );
buf ( n410465 , n405476 );
or ( n63468 , n410464 , n410465 );
nand ( n63469 , n63465 , n63468 );
buf ( n410468 , n63469 );
buf ( n410469 , n54297 );
buf ( n410470 , n62177 );
and ( n63473 , n410469 , n410470 );
buf ( n410472 , n55919 );
buf ( n410473 , n62159 );
and ( n63476 , n410472 , n410473 );
nor ( n63477 , n63473 , n63476 );
buf ( n410476 , n63477 );
buf ( n410477 , n410476 );
buf ( n410478 , n409429 );
or ( n63481 , n410477 , n410478 );
buf ( n410480 , n409425 );
buf ( n410481 , n409170 );
or ( n63484 , n410480 , n410481 );
nand ( n63485 , n63481 , n63484 );
buf ( n410484 , n63485 );
xor ( n63487 , n410468 , n410484 );
buf ( n410486 , n55846 );
buf ( n410487 , n59628 );
and ( n63490 , n410486 , n410487 );
buf ( n410489 , n403079 );
buf ( n410490 , n59457 );
and ( n63493 , n410489 , n410490 );
nor ( n63494 , n63490 , n63493 );
buf ( n410493 , n63494 );
buf ( n410494 , n410493 );
buf ( n410495 , n59637 );
or ( n63498 , n410494 , n410495 );
buf ( n410497 , n409388 );
buf ( n410498 , n59467 );
or ( n63501 , n410497 , n410498 );
nand ( n63502 , n63498 , n63501 );
buf ( n410501 , n63502 );
and ( n63504 , n63487 , n410501 );
and ( n63505 , n410468 , n410484 );
or ( n63506 , n63504 , n63505 );
buf ( n410505 , n63506 );
buf ( n410506 , n409273 );
buf ( n410507 , n409284 );
or ( n63510 , n410506 , n410507 );
buf ( n410509 , n409287 );
nand ( n63512 , n63510 , n410509 );
buf ( n410511 , n63512 );
buf ( n410512 , n410511 );
xor ( n63515 , n410505 , n410512 );
buf ( n410514 , n59435 );
buf ( n410515 , n55905 );
and ( n63518 , n410514 , n410515 );
buf ( n410517 , n406565 );
buf ( n410518 , n55895 );
and ( n63521 , n410517 , n410518 );
nor ( n63522 , n63518 , n63521 );
buf ( n410521 , n63522 );
buf ( n410522 , n410521 );
buf ( n410523 , n403120 );
or ( n63526 , n410522 , n410523 );
buf ( n410525 , n409443 );
buf ( n410526 , n403133 );
or ( n63529 , n410525 , n410526 );
nand ( n63530 , n63526 , n63529 );
buf ( n410529 , n63530 );
buf ( n410530 , n410529 );
buf ( n410531 , n62278 );
buf ( n410532 , n403146 );
and ( n63535 , n410531 , n410532 );
buf ( n410534 , n409474 );
buf ( n410535 , n401695 );
and ( n63538 , n410534 , n410535 );
nor ( n63539 , n63535 , n63538 );
buf ( n410538 , n63539 );
buf ( n410539 , n410538 );
not ( n63542 , n410539 );
buf ( n410541 , n63542 );
buf ( n410542 , n410541 );
buf ( n410543 , n401674 );
and ( n63546 , n410542 , n410543 );
buf ( n410545 , n409533 );
not ( n63548 , n410545 );
buf ( n410547 , n63548 );
buf ( n410548 , n410547 );
buf ( n410549 , n403164 );
and ( n63552 , n410548 , n410549 );
nor ( n63553 , n63546 , n63552 );
buf ( n410552 , n63553 );
buf ( n410553 , n410552 );
nand ( n63556 , n54247 , n53910 );
not ( n63557 , n63556 );
not ( n63558 , n54244 );
nand ( n63559 , n62459 , n63558 );
not ( n63560 , n63559 );
or ( n63561 , n63557 , n63560 );
not ( n63562 , n63556 );
nand ( n63563 , n63562 , n62459 , n63558 );
nand ( n63564 , n63561 , n63563 );
buf ( n410563 , n63564 );
buf ( n410564 , n401626 );
and ( n63567 , n410563 , n410564 );
buf ( n63568 , n62467 );
buf ( n410567 , n63568 );
buf ( n410568 , n401650 );
and ( n63571 , n410567 , n410568 );
nor ( n63572 , n63567 , n63571 );
buf ( n410571 , n63572 );
buf ( n410572 , n410571 );
nand ( n63575 , n410553 , n410572 );
buf ( n410574 , n63575 );
buf ( n410575 , n410574 );
xor ( n63578 , n410530 , n410575 );
buf ( n410577 , n58178 );
buf ( n410578 , n405391 );
and ( n63581 , n410577 , n410578 );
buf ( n410580 , n405335 );
buf ( n410581 , n405388 );
and ( n63584 , n410580 , n410581 );
nor ( n63585 , n63581 , n63584 );
buf ( n410584 , n63585 );
buf ( n410585 , n410584 );
buf ( n410586 , n405407 );
or ( n63589 , n410585 , n410586 );
buf ( n410588 , n409372 );
buf ( n410589 , n405384 );
or ( n63592 , n410588 , n410589 );
nand ( n63593 , n63589 , n63592 );
buf ( n410592 , n63593 );
buf ( n410593 , n410592 );
and ( n63596 , n63578 , n410593 );
and ( n63597 , n410530 , n410575 );
or ( n63598 , n63596 , n63597 );
buf ( n410597 , n63598 );
buf ( n410598 , n410597 );
and ( n63601 , n63515 , n410598 );
and ( n63602 , n410505 , n410512 );
or ( n63603 , n63601 , n63602 );
buf ( n410602 , n63603 );
xor ( n63605 , n409330 , n409347 );
xor ( n63606 , n63605 , n409352 );
buf ( n410605 , n63606 );
xor ( n410606 , n410602 , n410605 );
xor ( n63609 , n409417 , n409552 );
xor ( n63610 , n63609 , n409557 );
buf ( n410609 , n63610 );
and ( n63612 , n410606 , n410609 );
and ( n63613 , n410602 , n410605 );
or ( n63614 , n63612 , n63613 );
xor ( n63615 , n409561 , n409564 );
xor ( n63616 , n63615 , n62571 );
and ( n63617 , n63614 , n63616 );
xor ( n63618 , n409435 , n409452 );
xor ( n63619 , n63618 , n409547 );
buf ( n410618 , n63619 );
xor ( n63621 , n409380 , n409396 );
xor ( n63622 , n63621 , n409413 );
and ( n63623 , n410618 , n63622 );
buf ( n410622 , n54336 );
not ( n63625 , n62511 );
buf ( n410624 , n63625 );
and ( n63627 , n410622 , n410624 );
buf ( n410626 , n401699 );
not ( n63629 , n63625 );
buf ( n410628 , n63629 );
and ( n63631 , n410626 , n410628 );
nor ( n63632 , n63627 , n63631 );
buf ( n410631 , n63632 );
buf ( n410632 , n410631 );
buf ( n410633 , n409507 );
not ( n63636 , n410633 );
buf ( n410635 , n63636 );
buf ( n410636 , n410635 );
or ( n63639 , n410632 , n410636 );
buf ( n410638 , n409520 );
nand ( n63641 , n63639 , n410638 );
buf ( n410640 , n63641 );
buf ( n410641 , n410640 );
buf ( n410642 , n59596 );
buf ( n410643 , n55905 );
and ( n63646 , n410642 , n410643 );
buf ( n410645 , n409146 );
buf ( n410646 , n55895 );
and ( n63649 , n410645 , n410646 );
nor ( n63650 , n63646 , n63649 );
buf ( n410649 , n63650 );
buf ( n410650 , n410649 );
buf ( n410651 , n403120 );
or ( n63654 , n410650 , n410651 );
buf ( n410653 , n410521 );
buf ( n410654 , n403133 );
or ( n63657 , n410653 , n410654 );
nand ( n63658 , n63654 , n63657 );
buf ( n410657 , n63658 );
buf ( n410658 , n410657 );
xor ( n63661 , n410641 , n410658 );
buf ( n410660 , n58352 );
buf ( n410661 , n405215 );
and ( n63664 , n410660 , n410661 );
buf ( n410663 , n406571 );
buf ( n410664 , n58061 );
and ( n63667 , n410663 , n410664 );
nor ( n63668 , n63664 , n63667 );
buf ( n410667 , n63668 );
buf ( n410668 , n410667 );
buf ( n410669 , n403293 );
or ( n63672 , n410668 , n410669 );
buf ( n410671 , n410460 );
buf ( n410672 , n405476 );
or ( n63675 , n410671 , n410672 );
nand ( n63676 , n63672 , n63675 );
buf ( n410675 , n63676 );
buf ( n410676 , n410675 );
and ( n63679 , n63661 , n410676 );
and ( n63680 , n410641 , n410658 );
or ( n63681 , n63679 , n63680 );
buf ( n410680 , n63681 );
buf ( n410681 , n410680 );
xor ( n63684 , n409480 , n409524 );
xor ( n63685 , n63684 , n409542 );
buf ( n410684 , n63685 );
buf ( n410685 , n410684 );
xor ( n63688 , n410681 , n410685 );
buf ( n410687 , n58042 );
buf ( n410688 , n62177 );
and ( n63691 , n410687 , n410688 );
buf ( n410690 , n403088 );
buf ( n410691 , n62159 );
and ( n63694 , n410690 , n410691 );
nor ( n63695 , n63691 , n63694 );
buf ( n410694 , n63695 );
buf ( n410695 , n410694 );
buf ( n410696 , n409429 );
or ( n63699 , n410695 , n410696 );
buf ( n410698 , n410476 );
buf ( n410699 , n409170 );
or ( n63702 , n410698 , n410699 );
nand ( n63703 , n63699 , n63702 );
buf ( n410702 , n63703 );
buf ( n410703 , n410702 );
nand ( n63706 , n63558 , n53895 );
xnor ( n63707 , n54240 , n63706 );
buf ( n410706 , n63707 );
buf ( n410707 , n401626 );
and ( n63710 , n410706 , n410707 );
buf ( n410709 , n63564 );
buf ( n410710 , n401650 );
and ( n63713 , n410709 , n410710 );
nor ( n63714 , n63710 , n63713 );
buf ( n410713 , n63714 );
buf ( n410714 , n410713 );
buf ( n410715 , n62495 );
not ( n63718 , n410715 );
buf ( n410717 , n63718 );
buf ( n410718 , n410717 );
buf ( n410719 , n348158 );
not ( n63722 , n410719 );
buf ( n410721 , n63722 );
buf ( n410722 , n410721 );
nand ( n63725 , n410718 , n410722 );
buf ( n410724 , n63725 );
buf ( n410725 , n410724 );
buf ( n410726 , n410717 );
buf ( n410727 , n348158 );
nand ( n63730 , n410726 , n410727 );
buf ( n410729 , n63730 );
buf ( n410730 , n410729 );
nand ( n63733 , n410725 , n410730 );
buf ( n410732 , n63733 );
buf ( n410733 , n410732 );
nand ( n63736 , n410714 , n410733 );
buf ( n410735 , n63736 );
buf ( n410736 , n410735 );
xor ( n63739 , n410703 , n410736 );
buf ( n410738 , n405388 );
buf ( n410739 , n58205 );
and ( n63742 , n410738 , n410739 );
not ( n63743 , n410738 );
buf ( n410742 , n58166 );
and ( n63745 , n63743 , n410742 );
nor ( n63746 , n63742 , n63745 );
buf ( n410745 , n63746 );
buf ( n410746 , n410745 );
buf ( n410747 , n405407 );
or ( n63750 , n410746 , n410747 );
buf ( n410749 , n410584 );
buf ( n410750 , n405384 );
or ( n63753 , n410749 , n410750 );
nand ( n63754 , n63750 , n63753 );
buf ( n410753 , n63754 );
buf ( n410754 , n410753 );
and ( n63757 , n63739 , n410754 );
and ( n63758 , n410703 , n410736 );
or ( n63759 , n63757 , n63758 );
buf ( n410758 , n63759 );
buf ( n410759 , n410758 );
and ( n63762 , n63688 , n410759 );
and ( n63763 , n410681 , n410685 );
or ( n63764 , n63762 , n63763 );
buf ( n410763 , n63764 );
xor ( n63766 , n409380 , n409396 );
xor ( n63767 , n63766 , n409413 );
and ( n63768 , n410763 , n63767 );
and ( n63769 , n410618 , n410763 );
or ( n63770 , n63623 , n63768 , n63769 );
xor ( n63771 , n410602 , n410605 );
xor ( n63772 , n63771 , n410609 );
and ( n63773 , n63770 , n63772 );
xor ( n63774 , n410530 , n410575 );
xor ( n63775 , n63774 , n410593 );
buf ( n410774 , n63775 );
xor ( n63777 , n410468 , n410484 );
xor ( n63778 , n63777 , n410501 );
and ( n63779 , n410774 , n63778 );
buf ( n410778 , n55984 );
buf ( n410779 , n59628 );
and ( n63782 , n410778 , n410779 );
buf ( n410781 , n58135 );
buf ( n410782 , n59457 );
and ( n63785 , n410781 , n410782 );
nor ( n63786 , n63782 , n63785 );
buf ( n410785 , n63786 );
buf ( n410786 , n410785 );
buf ( n410787 , n59637 );
or ( n63790 , n410786 , n410787 );
buf ( n410789 , n410493 );
buf ( n410790 , n59467 );
or ( n63793 , n410789 , n410790 );
nand ( n63794 , n63790 , n63793 );
buf ( n410793 , n63794 );
buf ( n410794 , n410552 );
buf ( n410795 , n410571 );
or ( n63798 , n410794 , n410795 );
buf ( n410797 , n410574 );
nand ( n63800 , n63798 , n410797 );
buf ( n410799 , n63800 );
xor ( n63802 , n410793 , n410799 );
buf ( n410801 , n55895 );
buf ( n410802 , n409140 );
and ( n63805 , n410801 , n410802 );
not ( n63806 , n410801 );
buf ( n410805 , n62139 );
and ( n63808 , n63806 , n410805 );
nor ( n63809 , n63805 , n63808 );
buf ( n410808 , n63809 );
buf ( n410809 , n410808 );
buf ( n410810 , n403120 );
or ( n63813 , n410809 , n410810 );
buf ( n410812 , n410649 );
buf ( n410813 , n403133 );
or ( n63816 , n410812 , n410813 );
nand ( n63817 , n63813 , n63816 );
buf ( n410816 , n63817 );
buf ( n410817 , n410816 );
buf ( n410818 , n62467 );
buf ( n410819 , n403146 );
and ( n63822 , n410818 , n410819 );
buf ( n410821 , n409468 );
buf ( n410822 , n401695 );
and ( n63825 , n410821 , n410822 );
nor ( n63826 , n63822 , n63825 );
buf ( n410825 , n63826 );
buf ( n410826 , n410825 );
buf ( n410827 , n403158 );
or ( n63830 , n410826 , n410827 );
buf ( n410829 , n410538 );
buf ( n410830 , n403167 );
or ( n63833 , n410829 , n410830 );
nand ( n63834 , n63830 , n63833 );
buf ( n410833 , n63834 );
buf ( n410834 , n410833 );
xor ( n63837 , n410817 , n410834 );
buf ( n410836 , n59435 );
buf ( n410837 , n405215 );
and ( n63840 , n410836 , n410837 );
buf ( n410839 , n406565 );
buf ( n410840 , n58061 );
and ( n63843 , n410839 , n410840 );
nor ( n63844 , n63840 , n63843 );
buf ( n410843 , n63844 );
buf ( n410844 , n410843 );
buf ( n410845 , n403293 );
or ( n63848 , n410844 , n410845 );
buf ( n410847 , n410667 );
buf ( n410848 , n405476 );
or ( n63851 , n410847 , n410848 );
nand ( n63852 , n63848 , n63851 );
buf ( n410851 , n63852 );
buf ( n410852 , n410851 );
and ( n63855 , n63837 , n410852 );
and ( n63856 , n410817 , n410834 );
or ( n63857 , n63855 , n63856 );
buf ( n410856 , n63857 );
and ( n63859 , n63802 , n410856 );
and ( n63860 , n410793 , n410799 );
or ( n63861 , n63859 , n63860 );
xor ( n63862 , n410468 , n410484 );
xor ( n63863 , n63862 , n410501 );
and ( n63864 , n63861 , n63863 );
and ( n63865 , n410774 , n63861 );
or ( n63866 , n63779 , n63864 , n63865 );
xor ( n63867 , n410505 , n410512 );
xor ( n63868 , n63867 , n410598 );
buf ( n410867 , n63868 );
or ( n63870 , n63866 , n410867 );
not ( n63871 , n63870 );
xor ( n63872 , n409380 , n409396 );
xor ( n63873 , n63872 , n409413 );
xor ( n63874 , n410618 , n410763 );
xor ( n63875 , n63873 , n63874 );
not ( n63876 , n63875 );
or ( n63877 , n63871 , n63876 );
nand ( n63878 , n410867 , n63866 );
nand ( n63879 , n63877 , n63878 );
xor ( n63880 , n410602 , n410605 );
xor ( n63881 , n63880 , n410609 );
and ( n63882 , n63879 , n63881 );
and ( n63883 , n63770 , n63879 );
or ( n63884 , n63773 , n63882 , n63883 );
xor ( n63885 , n409561 , n409564 );
xor ( n63886 , n63885 , n62571 );
and ( n63887 , n63884 , n63886 );
and ( n63888 , n63614 , n63884 );
or ( n63889 , n63617 , n63887 , n63888 );
buf ( n410888 , n63889 );
xor ( n63891 , n410452 , n410888 );
buf ( n410890 , n388502 );
not ( n63893 , n410890 );
buf ( n410892 , n40653 );
not ( n63895 , n410892 );
or ( n63896 , n63893 , n63895 );
buf ( n410895 , n407928 );
buf ( n410896 , n410127 );
nand ( n63899 , n410895 , n410896 );
buf ( n410898 , n63899 );
buf ( n410899 , n410898 );
nand ( n63902 , n63896 , n410899 );
buf ( n410901 , n63902 );
buf ( n410902 , n410901 );
not ( n63905 , n410902 );
nand ( n63906 , n62075 , n40695 , n40698 );
buf ( n410905 , n63906 );
not ( n63908 , n410905 );
buf ( n410907 , n63908 );
buf ( n410908 , n410907 );
not ( n63911 , n410908 );
or ( n63912 , n63905 , n63911 );
buf ( n410911 , n410376 );
buf ( n410912 , n409076 );
nand ( n63915 , n410911 , n410912 );
buf ( n410914 , n63915 );
buf ( n410915 , n410914 );
nand ( n63918 , n63912 , n410915 );
buf ( n410917 , n63918 );
buf ( n410918 , n410917 );
and ( n63921 , n63891 , n410918 );
and ( n63922 , n410452 , n410888 );
or ( n63923 , n63921 , n63922 );
buf ( n410922 , n63923 );
buf ( n410923 , n410922 );
not ( n63926 , n410923 );
buf ( n410925 , n63926 );
buf ( n410926 , n410925 );
nand ( n63929 , n63449 , n410926 );
buf ( n410928 , n63929 );
not ( n63931 , n410928 );
or ( n63932 , n63423 , n63931 );
buf ( n410931 , n410922 );
buf ( n410932 , n410445 );
nand ( n63935 , n410931 , n410932 );
buf ( n410934 , n63935 );
nand ( n63937 , n63932 , n410934 );
buf ( n410936 , n63937 );
nand ( n63939 , n63365 , n410936 );
buf ( n410938 , n63939 );
buf ( n410939 , n410938 );
buf ( n410940 , n63362 );
not ( n63943 , n410940 );
buf ( n410942 , n63341 );
nand ( n63945 , n63943 , n410942 );
buf ( n410944 , n63945 );
buf ( n410945 , n410944 );
nand ( n63948 , n410939 , n410945 );
buf ( n410947 , n63948 );
buf ( n410948 , n410947 );
xor ( n63951 , n410321 , n410948 );
buf ( n410950 , n40943 );
not ( n63953 , n410950 );
buf ( n410952 , n399283 );
not ( n63955 , n410952 );
and ( n63956 , n63953 , n63955 );
buf ( n410955 , n40943 );
buf ( n410956 , n399283 );
and ( n63959 , n410955 , n410956 );
nor ( n63960 , n63956 , n63959 );
buf ( n410959 , n63960 );
buf ( n410960 , n410959 );
not ( n63963 , n410960 );
buf ( n410962 , n63963 );
buf ( n410963 , n410962 );
not ( n63966 , n410963 );
buf ( n410965 , n36801 );
not ( n63968 , n410965 );
or ( n63969 , n63966 , n63968 );
buf ( n410968 , n388669 );
buf ( n410969 , n400440 );
not ( n63972 , n410969 );
buf ( n410971 , n388419 );
not ( n63974 , n410971 );
or ( n63975 , n63972 , n63974 );
buf ( n410974 , n390307 );
buf ( n410975 , n51185 );
nand ( n63978 , n410974 , n410975 );
buf ( n410977 , n63978 );
buf ( n410978 , n410977 );
nand ( n63981 , n63975 , n410978 );
buf ( n410980 , n63981 );
buf ( n410981 , n410980 );
nand ( n63984 , n410968 , n410981 );
buf ( n410983 , n63984 );
buf ( n410984 , n410983 );
nand ( n63987 , n63969 , n410984 );
buf ( n410986 , n63987 );
buf ( n410987 , n410986 );
and ( n63990 , n63951 , n410987 );
and ( n63991 , n410321 , n410948 );
or ( n63992 , n63990 , n63991 );
buf ( n410991 , n63992 );
buf ( n410992 , n410991 );
and ( n63995 , n63298 , n410992 );
and ( n63996 , n410274 , n410295 );
or ( n63997 , n63995 , n63996 );
buf ( n410996 , n63997 );
buf ( n410997 , n410996 );
xor ( n64000 , n410270 , n410997 );
not ( n64001 , n42390 );
buf ( n411000 , n35820 );
buf ( n64003 , n411000 );
buf ( n411002 , n64003 );
nor ( n64005 , n64001 , n411002 );
not ( n64006 , n64005 );
not ( n64007 , n402819 );
and ( n64008 , n64006 , n64007 );
buf ( n411007 , n411002 );
not ( n64010 , n411007 );
buf ( n411009 , n395885 );
not ( n411010 , n411009 );
or ( n64013 , n64010 , n411010 );
buf ( n411012 , n389589 );
nand ( n64015 , n64013 , n411012 );
buf ( n411014 , n64015 );
nor ( n64017 , n64008 , n411014 );
not ( n64018 , n410980 );
not ( n64019 , n36801 );
or ( n64020 , n64018 , n64019 );
buf ( n411019 , n408882 );
not ( n64022 , n411019 );
buf ( n411021 , n384413 );
nand ( n64024 , n64022 , n411021 );
buf ( n411023 , n64024 );
nand ( n64026 , n64020 , n411023 );
xor ( n64027 , n64017 , n64026 );
not ( n64028 , n409602 );
not ( n64029 , n64028 );
buf ( n411028 , n409610 );
not ( n64031 , n411028 );
buf ( n411030 , n409047 );
not ( n64033 , n411030 );
or ( n64034 , n64031 , n64033 );
buf ( n411033 , n409047 );
buf ( n411034 , n409610 );
or ( n64037 , n411033 , n411034 );
nand ( n64038 , n64034 , n64037 );
buf ( n411037 , n64038 );
not ( n64040 , n411037 );
or ( n64041 , n64029 , n64040 );
or ( n64042 , n411037 , n64028 );
nand ( n64043 , n64041 , n64042 );
xor ( n64044 , n64027 , n64043 );
buf ( n411043 , n64044 );
not ( n64046 , n411043 );
not ( n64047 , n395362 );
not ( n64048 , n47863 );
not ( n64049 , n384211 );
or ( n64050 , n64048 , n64049 );
not ( n64051 , n389067 );
nand ( n64052 , n64051 , n395315 );
nand ( n64053 , n64050 , n64052 );
not ( n64054 , n64053 );
or ( n64055 , n64047 , n64054 );
not ( n64056 , n395312 );
not ( n64057 , n389692 );
or ( n64058 , n64056 , n64057 );
or ( n64059 , n38472 , n395315 );
nand ( n64060 , n64058 , n64059 );
buf ( n411059 , n64060 );
buf ( n411060 , n395349 );
nand ( n64063 , n411059 , n411060 );
buf ( n411062 , n64063 );
nand ( n64065 , n64055 , n411062 );
buf ( n411064 , n64065 );
not ( n64067 , n411064 );
or ( n64068 , n64046 , n64067 );
buf ( n411067 , n64044 );
buf ( n411068 , n64065 );
or ( n64071 , n411067 , n411068 );
xor ( n64072 , n410184 , n410209 );
xor ( n64073 , n64072 , n410236 );
buf ( n411072 , n64073 );
buf ( n411073 , n411072 );
not ( n64076 , n43272 );
not ( n64077 , n410105 );
not ( n64078 , n64077 );
or ( n64079 , n64076 , n64078 );
or ( n64080 , n40824 , n397498 );
nand ( n64081 , n40977 , n397498 );
nand ( n64082 , n64080 , n64081 );
not ( n64083 , n64082 );
nand ( n64084 , n64083 , n388460 );
nand ( n64085 , n64079 , n64084 );
buf ( n411084 , n64085 );
xor ( n64087 , n411073 , n411084 );
buf ( n411086 , n391173 );
buf ( n411087 , n358975 );
and ( n64090 , n411086 , n411087 );
buf ( n411089 , n64090 );
buf ( n411090 , n411089 );
and ( n64093 , n64087 , n411090 );
and ( n64094 , n411073 , n411084 );
or ( n64095 , n64093 , n64094 );
buf ( n411094 , n64095 );
buf ( n411095 , n411094 );
nand ( n64098 , n64071 , n411095 );
buf ( n411097 , n64098 );
buf ( n411098 , n411097 );
nand ( n64101 , n64068 , n411098 );
buf ( n411100 , n64101 );
buf ( n411101 , n411100 );
and ( n64104 , n64000 , n411101 );
and ( n64105 , n410270 , n410997 );
or ( n64106 , n64104 , n64105 );
buf ( n411105 , n64106 );
buf ( n411106 , n411105 );
buf ( n411107 , C0 );
buf ( n411108 , n411107 );
not ( n64135 , n392740 );
not ( n64136 , n44776 );
buf ( n411111 , n64136 );
not ( n64138 , n411111 );
buf ( n411113 , n388955 );
not ( n64140 , n411113 );
or ( n64141 , n64138 , n64140 );
buf ( n411116 , n37763 );
buf ( n411117 , n44776 );
nand ( n64144 , n411116 , n411117 );
buf ( n411119 , n64144 );
buf ( n411120 , n411119 );
nand ( n64147 , n64141 , n411120 );
buf ( n411122 , n64147 );
not ( n64149 , n411122 );
or ( n64150 , n64135 , n64149 );
and ( n64151 , n64136 , n391483 );
not ( n64152 , n64136 );
and ( n64153 , n64152 , n385342 );
or ( n64154 , n64151 , n64153 );
nand ( n64155 , n64154 , n45260 );
nand ( n64156 , n64150 , n64155 );
not ( n64157 , n64156 );
buf ( n411132 , n64157 );
not ( n64159 , n411132 );
buf ( n411134 , n390362 );
not ( n64161 , n411134 );
buf ( n411136 , n388102 );
not ( n64163 , n411136 );
buf ( n411138 , n43044 );
not ( n64165 , n411138 );
or ( n64166 , n64163 , n64165 );
buf ( n411141 , n27196 );
buf ( n411142 , n40600 );
nand ( n64169 , n411141 , n411142 );
buf ( n411144 , n64169 );
buf ( n411145 , n411144 );
nand ( n64172 , n64166 , n411145 );
buf ( n411147 , n64172 );
buf ( n411148 , n411147 );
not ( n64175 , n411148 );
or ( n64176 , n64161 , n64175 );
buf ( n411151 , n388102 );
not ( n64178 , n411151 );
buf ( n411153 , n391569 );
not ( n64180 , n411153 );
or ( n64181 , n64178 , n64180 );
buf ( n411156 , n40818 );
buf ( n411157 , n40600 );
nand ( n64184 , n411156 , n411157 );
buf ( n411159 , n64184 );
buf ( n411160 , n411159 );
nand ( n64187 , n64181 , n411160 );
buf ( n411162 , n64187 );
buf ( n411163 , n411162 );
buf ( n411164 , n43286 );
nand ( n64191 , n411163 , n411164 );
buf ( n411166 , n64191 );
buf ( n411167 , n411166 );
nand ( n64194 , n64176 , n411167 );
buf ( n411169 , n64194 );
buf ( n411170 , n411169 );
not ( n64197 , n391563 );
not ( n64198 , n394219 );
and ( n64199 , n64197 , n64198 );
not ( n64200 , n393562 );
and ( n64201 , n64200 , n394219 );
nor ( n64202 , n64199 , n64201 );
not ( n64203 , n64202 );
not ( n64204 , n45662 );
or ( n64205 , n64203 , n64204 );
buf ( n411180 , n392884 );
not ( n64207 , n411180 );
buf ( n411182 , n388897 );
not ( n64209 , n411182 );
or ( n64210 , n64207 , n64209 );
buf ( n411185 , n393117 );
buf ( n411186 , n392887 );
nand ( n64213 , n411185 , n411186 );
buf ( n411188 , n64213 );
buf ( n411189 , n411188 );
nand ( n64216 , n64210 , n411189 );
buf ( n411191 , n64216 );
buf ( n411192 , n411191 );
buf ( n411193 , n37314 );
nand ( n64220 , n411192 , n411193 );
buf ( n411195 , n64220 );
nand ( n64222 , n64205 , n411195 );
buf ( n411197 , n64222 );
or ( n64224 , n411170 , n411197 );
buf ( n411199 , n64224 );
buf ( n411200 , n389359 );
not ( n64227 , n411200 );
buf ( n411202 , n399164 );
not ( n64229 , n411202 );
or ( n64230 , n64227 , n64229 );
buf ( n411205 , n24049 );
buf ( n411206 , n389356 );
nand ( n64233 , n411205 , n411206 );
buf ( n411208 , n64233 );
buf ( n411209 , n411208 );
nand ( n64236 , n64230 , n411209 );
buf ( n411211 , n64236 );
buf ( n411212 , n411211 );
not ( n64239 , n411212 );
buf ( n411214 , n396622 );
not ( n64241 , n411214 );
or ( n64242 , n64239 , n64241 );
buf ( n411217 , n46921 );
buf ( n411218 , n42073 );
not ( n64245 , n411218 );
buf ( n411220 , n399164 );
not ( n64247 , n411220 );
or ( n64248 , n64245 , n64247 );
buf ( n411223 , n24049 );
buf ( n411224 , n42074 );
nand ( n64251 , n411223 , n411224 );
buf ( n411226 , n64251 );
buf ( n411227 , n411226 );
nand ( n64254 , n64248 , n411227 );
buf ( n411229 , n64254 );
buf ( n411230 , n411229 );
nand ( n64257 , n411217 , n411230 );
buf ( n411232 , n64257 );
buf ( n411233 , n411232 );
nand ( n64260 , n64242 , n411233 );
buf ( n411235 , n64260 );
not ( n64262 , n411235 );
buf ( n411237 , n389162 );
not ( n64264 , n411237 );
buf ( n411239 , n410337 );
not ( n64266 , n411239 );
or ( n64267 , n64264 , n64266 );
buf ( n64268 , n24116 );
not ( n64269 , n64268 );
not ( n64270 , n394663 );
or ( n64271 , n64269 , n64270 );
buf ( n411246 , n27258 );
not ( n64273 , n64268 );
buf ( n411248 , n64273 );
nand ( n64275 , n411246 , n411248 );
buf ( n411250 , n64275 );
nand ( n64277 , n64271 , n411250 );
nand ( n64278 , n64277 , n57569 );
buf ( n411253 , n64278 );
nand ( n64280 , n64267 , n411253 );
buf ( n411255 , n64280 );
not ( n64282 , n411255 );
or ( n64283 , n64262 , n64282 );
not ( n64284 , n411235 );
not ( n64285 , n64284 );
not ( n64286 , n411255 );
not ( n64287 , n64286 );
or ( n64288 , n64285 , n64287 );
not ( n64289 , n22982 );
not ( n64290 , n391443 );
or ( n64291 , n64289 , n64290 );
nand ( n64292 , n46906 , n391446 );
nand ( n64293 , n64291 , n64292 );
not ( n64294 , n64293 );
buf ( n411269 , n48025 );
not ( n64296 , n411269 );
buf ( n411271 , n64296 );
not ( n64298 , n411271 );
or ( n64299 , n64294 , n64298 );
buf ( n411274 , n389341 );
buf ( n411275 , n54957 );
and ( n64302 , n411274 , n411275 );
not ( n64303 , n411274 );
buf ( n411278 , n22982 );
and ( n64305 , n64303 , n411278 );
nor ( n64306 , n64302 , n64305 );
buf ( n411281 , n64306 );
or ( n64308 , n386474 , n411281 );
nand ( n64309 , n64299 , n64308 );
nand ( n64310 , n64288 , n64309 );
nand ( n64311 , n64283 , n64310 );
and ( n64312 , n411199 , n64311 );
buf ( n411287 , n411169 );
buf ( n411288 , n64222 );
and ( n64315 , n411287 , n411288 );
buf ( n411290 , n64315 );
nor ( n64317 , n64312 , n411290 );
buf ( n411292 , n64317 );
not ( n64319 , n411292 );
or ( n64320 , n64159 , n64319 );
xor ( n64321 , n410146 , n410163 );
xor ( n64322 , n64321 , n410179 );
buf ( n411297 , n64322 );
not ( n64324 , n411297 );
buf ( n411299 , n388809 );
not ( n64326 , n411299 );
buf ( n411301 , n410201 );
not ( n64328 , n411301 );
or ( n64329 , n64326 , n64328 );
nand ( n64330 , n405736 , n388367 );
not ( n64331 , n64330 );
buf ( n411306 , n397069 );
buf ( n411307 , n388754 );
nand ( n64334 , n411306 , n411307 );
buf ( n411309 , n64334 );
not ( n64336 , n411309 );
or ( n64337 , n64331 , n64336 );
nand ( n64338 , n64337 , n388746 );
buf ( n411313 , n64338 );
nand ( n64340 , n64329 , n411313 );
buf ( n411315 , n64340 );
not ( n64342 , n411315 );
nand ( n64343 , n64324 , n64342 );
not ( n64344 , n64343 );
buf ( n411319 , n391870 );
buf ( n411320 , n36809 );
buf ( n411321 , n384614 );
nand ( n64348 , n411320 , n411321 );
buf ( n411323 , n64348 );
buf ( n411324 , n411323 );
buf ( n411325 , n358975 );
and ( n64352 , n411324 , n411325 );
buf ( n411327 , n36810 );
buf ( n411328 , n384606 );
and ( n64355 , n411327 , n411328 );
nor ( n64356 , n64352 , n64355 );
buf ( n411331 , n64356 );
buf ( n411332 , n411331 );
and ( n64359 , n411319 , n411332 );
buf ( n411334 , n64359 );
not ( n64361 , n411334 );
or ( n64362 , n64344 , n64361 );
nand ( n64363 , n411315 , n411297 );
nand ( n64364 , n64362 , n64363 );
buf ( n411339 , n64364 );
nand ( n64366 , n64320 , n411339 );
buf ( n411341 , n64366 );
buf ( n411342 , n64317 );
not ( n64369 , n411342 );
buf ( n411344 , n64369 );
buf ( n411345 , n411344 );
buf ( n411346 , n64156 );
nand ( n64373 , n411345 , n411346 );
buf ( n411348 , n64373 );
nand ( n64375 , n411341 , n411348 );
buf ( n411350 , n64375 );
not ( n64377 , n411350 );
buf ( n411352 , n45954 );
not ( n64379 , n411352 );
buf ( n411354 , n410053 );
not ( n64381 , n411354 );
or ( n64382 , n64379 , n64381 );
and ( n64383 , n390651 , n393369 );
not ( n64384 , n390651 );
and ( n64385 , n64384 , n393381 );
or ( n64386 , n64383 , n64385 );
buf ( n411361 , n64386 );
buf ( n411362 , n393825 );
nand ( n64389 , n411361 , n411362 );
buf ( n411364 , n64389 );
buf ( n411365 , n411364 );
nand ( n64392 , n64382 , n411365 );
buf ( n411367 , n64392 );
buf ( n411368 , n411367 );
not ( n64395 , n411368 );
or ( n64396 , n64377 , n64395 );
buf ( n411371 , n410240 );
not ( n64398 , n411371 );
buf ( n411373 , n64398 );
and ( n64400 , n63093 , n411373 );
not ( n64401 , n63093 );
and ( n64402 , n64401 , n410240 );
nor ( n64403 , n64400 , n64402 );
not ( n64404 , n410115 );
and ( n64405 , n64403 , n64404 );
not ( n64406 , n64403 );
and ( n64407 , n64406 , n410115 );
nor ( n64408 , n64405 , n64407 );
not ( n64409 , n411367 );
nand ( n411384 , n64409 , n411341 , n411348 );
nand ( n64411 , n64408 , n411384 );
buf ( n411386 , n64411 );
nand ( n64413 , n64396 , n411386 );
buf ( n411388 , n64413 );
buf ( n411389 , n411388 );
xor ( n64416 , n411108 , n411389 );
xor ( n64417 , n410039 , n410065 );
xor ( n64418 , n64417 , n410253 );
buf ( n411393 , n64418 );
buf ( n411394 , n411393 );
and ( n64421 , n64416 , n411394 );
or ( n64423 , n64421 , C0 );
buf ( n411397 , n64423 );
buf ( n411398 , n411397 );
xor ( n64426 , n411106 , n411398 );
buf ( n411400 , n410027 );
buf ( n411401 , n410023 );
xor ( n64429 , n411400 , n411401 );
buf ( n411403 , n410257 );
xor ( n64431 , n64429 , n411403 );
buf ( n411405 , n64431 );
buf ( n411406 , n411405 );
and ( n64434 , n64426 , n411406 );
and ( n64435 , n411106 , n411398 );
or ( n64436 , n64434 , n64435 );
buf ( n411410 , n64436 );
buf ( n411411 , n411410 );
xor ( n64439 , n410266 , n411411 );
and ( n64440 , n61958 , n61944 );
not ( n64441 , n61958 );
and ( n64442 , n64441 , n61945 );
nor ( n64443 , n64440 , n64442 );
and ( n64444 , n64443 , n61941 );
not ( n64445 , n64443 );
and ( n64446 , n64445 , n408961 );
nor ( n64447 , n64444 , n64446 );
buf ( n411421 , n64447 );
buf ( n411422 , C0 );
buf ( n411423 , n411422 );
xor ( n64474 , n411421 , n411423 );
xor ( n64475 , n64017 , n64026 );
and ( n64476 , n64475 , n64043 );
and ( n64477 , n64017 , n64026 );
or ( n64478 , n64476 , n64477 );
buf ( n411429 , n64478 );
not ( n64480 , n408915 );
xor ( n64481 , n61896 , n64480 );
xor ( n64482 , n64481 , n408926 );
buf ( n411433 , n64482 );
xor ( n64484 , n411429 , n411433 );
buf ( n411435 , n395349 );
not ( n64486 , n411435 );
buf ( n411437 , n64053 );
not ( n64488 , n411437 );
or ( n64489 , n64486 , n64488 );
buf ( n411440 , n408661 );
buf ( n411441 , n395362 );
nand ( n64492 , n411440 , n411441 );
buf ( n411443 , n64492 );
buf ( n411444 , n411443 );
nand ( n64495 , n64489 , n411444 );
buf ( n411446 , n64495 );
buf ( n411447 , n411446 );
and ( n64498 , n64484 , n411447 );
and ( n64499 , n411429 , n411433 );
or ( n64500 , n64498 , n64499 );
buf ( n411451 , n64500 );
buf ( n411452 , n411451 );
xor ( n64503 , n64474 , n411452 );
buf ( n411454 , n64503 );
buf ( n411455 , n411454 );
not ( n64506 , n390485 );
buf ( n411457 , n400033 );
not ( n64508 , n411457 );
buf ( n411459 , n391129 );
not ( n64510 , n411459 );
or ( n64511 , n64508 , n64510 );
buf ( n411462 , n389897 );
buf ( n411463 , n400042 );
nand ( n64514 , n411462 , n411463 );
buf ( n411465 , n64514 );
buf ( n411466 , n411465 );
nand ( n64517 , n64511 , n411466 );
buf ( n411468 , n64517 );
not ( n64519 , n411468 );
or ( n64520 , n64506 , n64519 );
buf ( n411471 , n408691 );
buf ( n411472 , n391638 );
nand ( n64523 , n411471 , n411472 );
buf ( n411474 , n64523 );
nand ( n64525 , n64520 , n411474 );
buf ( n411476 , n409717 );
buf ( n411477 , n409773 );
xor ( n64528 , n411476 , n411477 );
buf ( n411479 , n409743 );
xnor ( n64530 , n64528 , n411479 );
buf ( n411481 , n64530 );
buf ( n411482 , n411481 );
not ( n64533 , n411482 );
buf ( n411484 , n64533 );
not ( n64535 , n411484 );
buf ( n411486 , n43286 );
not ( n64537 , n411486 );
buf ( n411488 , n411147 );
not ( n64539 , n411488 );
or ( n64540 , n64537 , n64539 );
buf ( n411491 , n390362 );
buf ( n411492 , n410083 );
nand ( n64543 , n411491 , n411492 );
buf ( n411494 , n64543 );
buf ( n411495 , n411494 );
nand ( n64546 , n64540 , n411495 );
buf ( n411497 , n64546 );
buf ( n411498 , n411497 );
not ( n64549 , n411498 );
buf ( n411500 , n43536 );
not ( n64551 , n411500 );
buf ( n411502 , n391024 );
not ( n64553 , n411502 );
buf ( n411504 , n64553 );
buf ( n411505 , n411504 );
not ( n64556 , n411505 );
buf ( n411507 , n386150 );
not ( n64558 , n411507 );
or ( n64559 , n64556 , n64558 );
buf ( n411510 , n386147 );
buf ( n411511 , n391024 );
nand ( n64562 , n411510 , n411511 );
buf ( n411513 , n64562 );
buf ( n411514 , n411513 );
nand ( n64565 , n64559 , n411514 );
buf ( n411516 , n64565 );
buf ( n411517 , n411516 );
not ( n64568 , n411517 );
or ( n64569 , n64551 , n64568 );
buf ( n411520 , n411504 );
not ( n64571 , n411520 );
buf ( n411522 , n388919 );
not ( n64573 , n411522 );
or ( n64574 , n64571 , n64573 );
buf ( n411525 , n396537 );
buf ( n411526 , n391024 );
nand ( n64577 , n411525 , n411526 );
buf ( n411528 , n64577 );
buf ( n411529 , n411528 );
nand ( n64580 , n64574 , n411529 );
buf ( n411531 , n64580 );
buf ( n411532 , n411531 );
buf ( n411533 , n43515 );
nand ( n64584 , n411532 , n411533 );
buf ( n411535 , n64584 );
buf ( n411536 , n411535 );
nand ( n64587 , n64569 , n411536 );
buf ( n411538 , n64587 );
buf ( n411539 , n411538 );
not ( n64590 , n411539 );
buf ( n411541 , n64590 );
buf ( n411542 , n411541 );
nand ( n64593 , n64549 , n411542 );
buf ( n411544 , n64593 );
not ( n64595 , n411544 );
or ( n64596 , n64535 , n64595 );
nand ( n64597 , n411538 , n411497 );
nand ( n64598 , n64596 , n64597 );
xor ( n64599 , n64525 , n64598 );
xor ( n64600 , n409779 , n409666 );
xnor ( n64601 , n64600 , n409690 );
not ( n64602 , n64601 );
xnor ( n64603 , n64599 , n64602 );
buf ( n411554 , n64603 );
not ( n64605 , n411554 );
not ( n64606 , n47891 );
not ( n64607 , n42153 );
or ( n64608 , n64606 , n64607 );
buf ( n411559 , n49525 );
buf ( n411560 , n50584 );
nand ( n64611 , n411559 , n411560 );
buf ( n411562 , n64611 );
nand ( n64613 , n64608 , n411562 );
buf ( n411564 , n64613 );
buf ( n411565 , n51553 );
and ( n64616 , n411564 , n411565 );
and ( n64617 , n36216 , n397990 );
not ( n64618 , n36216 );
and ( n64619 , n64618 , n50584 );
nor ( n64620 , n64617 , n64619 );
not ( n64621 , n64620 );
nor ( n64622 , n64621 , n50580 );
buf ( n411573 , n64622 );
nor ( n64624 , n64616 , n411573 );
buf ( n411575 , n64624 );
buf ( n411576 , n411575 );
not ( n64627 , n411576 );
or ( n64628 , n64605 , n64627 );
buf ( n411579 , n411497 );
not ( n64630 , n411579 );
buf ( n411581 , n411481 );
not ( n64632 , n411581 );
or ( n64633 , n64630 , n64632 );
buf ( n411584 , n411497 );
buf ( n411585 , n411481 );
or ( n64636 , n411584 , n411585 );
nand ( n64637 , n64633 , n64636 );
buf ( n411588 , n64637 );
buf ( n411589 , n411588 );
buf ( n411590 , n411538 );
and ( n64641 , n411589 , n411590 );
not ( n64642 , n411589 );
buf ( n411593 , n411541 );
and ( n64644 , n64642 , n411593 );
nor ( n64645 , n64641 , n64644 );
buf ( n411596 , n64645 );
buf ( n411597 , n411596 );
not ( n64648 , n411597 );
buf ( n411599 , n64648 );
buf ( n411600 , n411599 );
not ( n64651 , n43515 );
not ( n64652 , n411516 );
or ( n64653 , n64651 , n64652 );
buf ( n411604 , n411504 );
not ( n64655 , n411604 );
buf ( n411606 , n40971 );
not ( n64657 , n411606 );
or ( n64658 , n64655 , n64657 );
buf ( n411609 , n27613 );
buf ( n411610 , n391024 );
nand ( n64661 , n411609 , n411610 );
buf ( n411612 , n64661 );
buf ( n411613 , n411612 );
nand ( n64664 , n64658 , n411613 );
buf ( n411615 , n64664 );
buf ( n411616 , n411615 );
buf ( n411617 , n43536 );
nand ( n64668 , n411616 , n411617 );
buf ( n411619 , n64668 );
nand ( n64670 , n64653 , n411619 );
buf ( n411621 , n64670 );
not ( n64672 , n411621 );
buf ( n411623 , n49117 );
not ( n64674 , n411623 );
buf ( n411625 , n391764 );
not ( n64676 , n411625 );
or ( n64677 , n64674 , n64676 );
buf ( n411628 , n388263 );
buf ( n411629 , n49124 );
nand ( n64680 , n411628 , n411629 );
buf ( n411631 , n64680 );
buf ( n411632 , n411631 );
nand ( n64683 , n64677 , n411632 );
buf ( n411634 , n64683 );
not ( n64685 , n411634 );
not ( n64686 , n383894 );
or ( n64687 , n64685 , n64686 );
buf ( n411638 , n410308 );
buf ( n411639 , n388629 );
nand ( n64690 , n411638 , n411639 );
buf ( n411641 , n64690 );
nand ( n64692 , n64687 , n411641 );
buf ( n411643 , n64692 );
not ( n64694 , n411643 );
or ( n64695 , n64672 , n64694 );
buf ( n411646 , n64670 );
buf ( n411647 , n64692 );
or ( n64698 , n411646 , n411647 );
buf ( n411649 , n389122 );
buf ( n411650 , n411229 );
and ( n64701 , n411649 , n411650 );
buf ( n411652 , n409705 );
not ( n64703 , n411652 );
buf ( n411654 , n41562 );
nor ( n64705 , n64703 , n411654 );
buf ( n411656 , n64705 );
buf ( n411657 , n411656 );
nor ( n64708 , n64701 , n411657 );
buf ( n411659 , n64708 );
not ( n64710 , n411659 );
xor ( n64711 , n410368 , n410389 );
and ( n64712 , n64711 , n410418 );
and ( n64713 , n410368 , n410389 );
or ( n64714 , n64712 , n64713 );
buf ( n411665 , n64714 );
not ( n64716 , n411665 );
or ( n64717 , n64710 , n64716 );
not ( n64718 , n411659 );
buf ( n411669 , n411665 );
not ( n64720 , n411669 );
buf ( n411671 , n64720 );
nand ( n64722 , n64718 , n411671 );
nand ( n64723 , n64717 , n64722 );
buf ( n411674 , n38960 );
not ( n64725 , n411674 );
buf ( n411676 , n411281 );
not ( n64727 , n411676 );
and ( n64728 , n64725 , n64727 );
buf ( n411679 , n409731 );
not ( n64730 , n411679 );
buf ( n411681 , n386474 );
nor ( n64732 , n64730 , n411681 );
buf ( n411683 , n64732 );
buf ( n411684 , n411683 );
nor ( n64735 , n64728 , n411684 );
buf ( n411686 , n64735 );
xnor ( n64737 , n64723 , n411686 );
buf ( n411688 , n64737 );
nand ( n64739 , n64698 , n411688 );
buf ( n411690 , n64739 );
buf ( n411691 , n411690 );
nand ( n64742 , n64695 , n411691 );
buf ( n411693 , n64742 );
buf ( n411694 , n411693 );
not ( n64745 , n411694 );
buf ( n411696 , n64745 );
buf ( n411697 , n411696 );
nand ( n64748 , n411600 , n411697 );
buf ( n411699 , n64748 );
buf ( n411700 , n411699 );
not ( n64751 , n411700 );
buf ( n411702 , n388746 );
not ( n64753 , n411702 );
buf ( n411704 , n405736 );
not ( n64755 , n411704 );
buf ( n411706 , n394330 );
not ( n64757 , n411706 );
or ( n64758 , n64755 , n64757 );
buf ( n411709 , n27301 );
buf ( n411710 , n388754 );
nand ( n64761 , n411709 , n411710 );
buf ( n411712 , n64761 );
buf ( n411713 , n411712 );
nand ( n64764 , n64758 , n411713 );
buf ( n411715 , n64764 );
buf ( n411716 , n411715 );
not ( n64767 , n411716 );
or ( n64768 , n64753 , n64767 );
not ( n64769 , n64330 );
not ( n64770 , n411309 );
or ( n64771 , n64769 , n64770 );
nand ( n64772 , n64771 , n388809 );
buf ( n411723 , n64772 );
nand ( n64774 , n64768 , n411723 );
buf ( n411725 , n64774 );
buf ( n411726 , n411725 );
not ( n64777 , n41373 );
and ( n64778 , n406821 , n410407 );
not ( n64779 , n406821 );
not ( n64780 , n41341 );
and ( n64781 , n64779 , n64780 );
or ( n64782 , n64778 , n64781 );
not ( n64783 , n64782 );
or ( n64784 , n64777 , n64783 );
nand ( n64785 , n410413 , n388830 );
nand ( n64786 , n64784 , n64785 );
buf ( n411737 , n64786 );
and ( n64788 , n28390 , n41555 );
not ( n64789 , n28390 );
and ( n64790 , n64789 , n41559 );
or ( n64791 , n64788 , n64790 );
buf ( n411742 , n64791 );
not ( n64793 , n411742 );
buf ( n411744 , n390429 );
not ( n64795 , n411744 );
or ( n64796 , n64793 , n64795 );
buf ( n411747 , n410433 );
buf ( n411748 , n42924 );
nand ( n64799 , n411747 , n411748 );
buf ( n411750 , n64799 );
buf ( n411751 , n411750 );
nand ( n411752 , n64796 , n411751 );
buf ( n411753 , n411752 );
buf ( n411754 , n411753 );
xor ( n64805 , n411737 , n411754 );
not ( n64806 , n389162 );
not ( n64807 , n64277 );
or ( n64808 , n64806 , n64807 );
and ( n64809 , n28644 , n64273 );
not ( n64810 , n28644 );
and ( n64811 , n64810 , n64268 );
or ( n64812 , n64809 , n64811 );
buf ( n411763 , n64812 );
buf ( n411764 , n57569 );
nand ( n64815 , n411763 , n411764 );
buf ( n411766 , n64815 );
nand ( n64817 , n64808 , n411766 );
buf ( n411768 , n64817 );
and ( n64819 , n64805 , n411768 );
and ( n64820 , n411737 , n411754 );
or ( n64821 , n64819 , n64820 );
buf ( n411772 , n64821 );
buf ( n411773 , n411772 );
or ( n64824 , n411726 , n411773 );
xor ( n64825 , n410445 , n410925 );
xnor ( n64826 , n64825 , n410420 );
buf ( n411777 , n64826 );
nand ( n64828 , n64824 , n411777 );
buf ( n411779 , n64828 );
buf ( n411780 , n411779 );
buf ( n411781 , n411725 );
buf ( n411782 , n411772 );
nand ( n64833 , n411781 , n411782 );
buf ( n411784 , n64833 );
buf ( n411785 , n411784 );
nand ( n64836 , n411780 , n411785 );
buf ( n411787 , n64836 );
buf ( n411788 , n411787 );
buf ( n411789 , n50992 );
not ( n64840 , n411789 );
buf ( n411791 , n51185 );
not ( n64842 , n411791 );
and ( n64843 , n64840 , n64842 );
buf ( n411794 , n50992 );
buf ( n411795 , n51185 );
and ( n64846 , n411794 , n411795 );
nor ( n64847 , n64843 , n64846 );
buf ( n411798 , n64847 );
not ( n64849 , n411798 );
not ( n64850 , n64849 );
not ( n64851 , n36434 );
not ( n64852 , n64851 );
or ( n64853 , n64850 , n64852 );
or ( n64854 , n64082 , n40969 );
nand ( n64855 , n64853 , n64854 );
buf ( n411806 , n64855 );
xor ( n64857 , n411788 , n411806 );
buf ( n411808 , n390292 );
buf ( n411809 , n400042 );
buf ( n411810 , n40943 );
and ( n64861 , n411809 , n411810 );
not ( n64862 , n411809 );
buf ( n411813 , n396373 );
and ( n64864 , n64862 , n411813 );
nor ( n64865 , n64861 , n64864 );
buf ( n411816 , n64865 );
buf ( n411817 , n411816 );
or ( n64868 , n411808 , n411817 );
buf ( n411819 , n36845 );
buf ( n411820 , n410959 );
or ( n64871 , n411819 , n411820 );
nand ( n64872 , n64868 , n64871 );
buf ( n411823 , n64872 );
buf ( n411824 , n411823 );
and ( n64875 , n64857 , n411824 );
and ( n64876 , n411788 , n411806 );
or ( n64877 , n64875 , n64876 );
buf ( n411828 , n64877 );
buf ( n411829 , n411828 );
not ( n64880 , n411829 );
or ( n64881 , n64751 , n64880 );
buf ( n411832 , n411596 );
buf ( n411833 , n411693 );
nand ( n64884 , n411832 , n411833 );
buf ( n411835 , n64884 );
buf ( n411836 , n411835 );
nand ( n64887 , n64881 , n411836 );
buf ( n411838 , n64887 );
buf ( n411839 , n411838 );
nand ( n64890 , n64628 , n411839 );
buf ( n411841 , n64890 );
buf ( n411842 , n411575 );
not ( n64893 , n411842 );
buf ( n411844 , n64603 );
not ( n64895 , n411844 );
buf ( n411846 , n64895 );
buf ( n411847 , n411846 );
nand ( n64898 , n64893 , n411847 );
buf ( n411849 , n64898 );
nand ( n64900 , n411841 , n411849 );
buf ( n411851 , n64900 );
not ( n64902 , n411851 );
xor ( n64903 , n411429 , n411433 );
xor ( n64904 , n64903 , n411447 );
buf ( n411855 , n64904 );
buf ( n411856 , n411855 );
not ( n64907 , n411856 );
or ( n64908 , n64902 , n64907 );
not ( n64909 , n411855 );
nand ( n64910 , n64909 , n411841 , n411849 );
buf ( n411861 , C1 );
buf ( n411862 , n43515 );
not ( n64948 , n411862 );
buf ( n411864 , n409631 );
not ( n64950 , n411864 );
or ( n64951 , n64948 , n64950 );
buf ( n411867 , n411531 );
buf ( n411868 , n43536 );
nand ( n64954 , n411867 , n411868 );
buf ( n411870 , n64954 );
buf ( n411871 , n411870 );
nand ( n64957 , n64951 , n411871 );
buf ( n411873 , n64957 );
not ( n64959 , n411659 );
not ( n64960 , n411671 );
or ( n64961 , n64959 , n64960 );
not ( n64962 , n64718 );
not ( n64963 , n411665 );
or ( n64964 , n64962 , n64963 );
nand ( n64965 , n64964 , n411686 );
nand ( n64966 , n64961 , n64965 );
buf ( n411882 , n64966 );
not ( n64968 , n411882 );
buf ( n411884 , n64968 );
buf ( n411885 , n411884 );
not ( n64971 , n411885 );
buf ( n411887 , n43058 );
not ( n64973 , n411887 );
buf ( n411889 , n411191 );
not ( n64975 , n411889 );
buf ( n411891 , n64975 );
buf ( n411892 , n411891 );
not ( n64978 , n411892 );
and ( n64979 , n64973 , n64978 );
buf ( n411895 , n409680 );
buf ( n411896 , n37315 );
nor ( n64982 , n411895 , n411896 );
buf ( n411898 , n64982 );
buf ( n411899 , n411898 );
nor ( n64985 , n64979 , n411899 );
buf ( n411901 , n64985 );
buf ( n411902 , n411901 );
not ( n64988 , n411902 );
buf ( n411904 , n64988 );
buf ( n411905 , n411904 );
not ( n64991 , n411905 );
or ( n64992 , n64971 , n64991 );
buf ( n411908 , n64966 );
not ( n64994 , n411908 );
buf ( n411910 , n411901 );
not ( n64996 , n411910 );
or ( n64997 , n64994 , n64996 );
xor ( n64998 , n409067 , n409594 );
xor ( n64999 , n64998 , n409598 );
buf ( n411915 , n64999 );
buf ( n411916 , n411915 );
nand ( n65002 , n64997 , n411916 );
buf ( n411918 , n65002 );
buf ( n411919 , n411918 );
nand ( n65005 , n64992 , n411919 );
buf ( n411921 , n65005 );
xor ( n65007 , n411873 , n411921 );
buf ( n411923 , n411122 );
not ( n65009 , n411923 );
buf ( n411925 , n44771 );
nor ( n65011 , n65009 , n411925 );
buf ( n411927 , n65011 );
not ( n65013 , n411927 );
nand ( n65014 , n408718 , n392740 );
nand ( n65015 , n65013 , n65014 );
xnor ( n65016 , n65007 , n65015 );
not ( n65022 , n65016 );
or ( n65024 , n65022 , C0 );
buf ( n411934 , n45954 );
not ( n65026 , n411934 );
buf ( n411936 , n64386 );
not ( n65028 , n411936 );
or ( n65029 , n65026 , n65028 );
buf ( n411939 , n398116 );
not ( n65031 , n411939 );
buf ( n411941 , n46161 );
not ( n65033 , n411941 );
or ( n65034 , n65031 , n65033 );
buf ( n411944 , n38155 );
buf ( n411945 , n393384 );
nand ( n65037 , n411944 , n411945 );
buf ( n411947 , n65037 );
buf ( n411948 , n411947 );
nand ( n65040 , n65034 , n411948 );
buf ( n411950 , n65040 );
buf ( n411951 , n411950 );
buf ( n411952 , n393825 );
nand ( n65044 , n411951 , n411952 );
buf ( n411954 , n65044 );
buf ( n411955 , n411954 );
nand ( n65047 , n65029 , n411955 );
buf ( n411957 , n65047 );
buf ( n411958 , n411957 );
buf ( n411959 , n55055 );
not ( n65051 , n411959 );
buf ( n411961 , n384562 );
not ( n65053 , n411961 );
or ( n65054 , n65051 , n65053 );
buf ( n411964 , n395885 );
buf ( n411965 , n404855 );
nand ( n65057 , n411964 , n411965 );
buf ( n411967 , n65057 );
buf ( n411968 , n411967 );
nand ( n65060 , n65054 , n411968 );
buf ( n411970 , n65060 );
buf ( n411971 , n411970 );
not ( n65063 , n411971 );
buf ( n411973 , n392659 );
not ( n65065 , n411973 );
or ( n65066 , n65063 , n65065 );
buf ( n411976 , n411468 );
buf ( n411977 , n389908 );
nand ( n65069 , n411976 , n411977 );
buf ( n411979 , n65069 );
buf ( n411980 , n411979 );
nand ( n65072 , n65066 , n411980 );
buf ( n411982 , n65072 );
buf ( n411983 , n411982 );
or ( n65075 , n411958 , n411983 );
buf ( n411985 , n411915 );
buf ( n411986 , n411884 );
xor ( n65078 , n411985 , n411986 );
buf ( n411988 , n411904 );
xor ( n65080 , n65078 , n411988 );
buf ( n411990 , n65080 );
buf ( n411991 , n411990 );
nand ( n65083 , n65075 , n411991 );
buf ( n411993 , n65083 );
buf ( n411994 , n411993 );
buf ( n411995 , n411957 );
buf ( n411996 , n411982 );
nand ( n65088 , n411995 , n411996 );
buf ( n411998 , n65088 );
buf ( n411999 , n411998 );
nand ( n65091 , n411994 , n411999 );
buf ( n412001 , n65091 );
nand ( n65093 , n65024 , n412001 );
nand ( n65094 , C1 , n65093 );
nand ( n65095 , n64910 , n65094 );
buf ( n412005 , n65095 );
nand ( n65097 , n64908 , n412005 );
buf ( n412007 , n65097 );
buf ( n412008 , n412007 );
xor ( n65100 , n411455 , n412008 );
xor ( n65101 , n409617 , n409642 );
xor ( n65102 , n65101 , n409788 );
buf ( n412012 , n65102 );
buf ( n412013 , n412012 );
not ( n65105 , n411873 );
not ( n65106 , n411921 );
or ( n65107 , n65105 , n65106 );
nor ( n65108 , n411921 , n411873 );
not ( n65109 , n65015 );
or ( n65110 , n65108 , n65109 );
nand ( n65111 , n65107 , n65110 );
buf ( n412021 , n65111 );
xor ( n65113 , n412013 , n412021 );
not ( n65114 , n64525 );
buf ( n412024 , n65114 );
not ( n65116 , n412024 );
buf ( n412026 , n64601 );
not ( n65118 , n412026 );
or ( n65119 , n65116 , n65118 );
not ( n65120 , n411484 );
not ( n65121 , n411544 );
or ( n65122 , n65120 , n65121 );
nand ( n65123 , n65122 , n64597 );
buf ( n412033 , n65123 );
nand ( n65125 , n65119 , n412033 );
buf ( n412035 , n65125 );
buf ( n412036 , n412035 );
buf ( n412037 , n64602 );
buf ( n412038 , n64525 );
nand ( n65130 , n412037 , n412038 );
buf ( n412040 , n65130 );
buf ( n412041 , n412040 );
nand ( n65133 , n412036 , n412041 );
buf ( n412043 , n65133 );
buf ( n412044 , n412043 );
and ( n65136 , n65113 , n412044 );
and ( n65137 , n412013 , n412021 );
or ( n65138 , n65136 , n65137 );
buf ( n412048 , n65138 );
buf ( n412049 , n412048 );
not ( n65141 , n412049 );
buf ( n412051 , C1 );
or ( n65167 , n65141 , C0 );
nand ( n65171 , n65167 , C1 );
buf ( n412054 , n65171 );
buf ( n412055 , n412054 );
xor ( n65174 , n408870 , n408932 );
and ( n65175 , n65174 , n408941 );
not ( n65176 , n65174 );
and ( n65177 , n65176 , n408855 );
nor ( n65178 , n65175 , n65177 );
buf ( n412061 , n65178 );
not ( n65180 , n412061 );
buf ( n412063 , n65180 );
buf ( n412064 , n412063 );
and ( n65183 , n412055 , n412064 );
not ( n65184 , n412055 );
buf ( n412067 , n65178 );
and ( n65186 , n65184 , n412067 );
nor ( n65187 , n65183 , n65186 );
buf ( n412070 , n65187 );
buf ( n412071 , n412070 );
and ( n65190 , n65100 , n412071 );
and ( n65191 , n411455 , n412008 );
or ( n65192 , n65190 , n65191 );
buf ( n412075 , n65192 );
buf ( n412076 , n412075 );
xor ( n65195 , n64439 , n412076 );
buf ( n412078 , n65195 );
buf ( n412079 , n412078 );
xor ( n65198 , n411106 , n411398 );
xor ( n65199 , n65198 , n411406 );
buf ( n412082 , n65199 );
buf ( n412083 , n412082 );
xor ( n65202 , n411455 , n412008 );
xor ( n65203 , n65202 , n412071 );
buf ( n412086 , n65203 );
buf ( n412087 , n412086 );
xor ( n65206 , n412083 , n412087 );
buf ( n412089 , n408668 );
buf ( n412090 , n408635 );
xor ( n65209 , n412089 , n412090 );
buf ( n412092 , n408771 );
xor ( n65211 , n65209 , n412092 );
buf ( n412094 , n65211 );
buf ( n412095 , n412094 );
buf ( n412096 , C0 );
buf ( n412097 , n50579 );
not ( n65229 , n412097 );
buf ( n412099 , n64613 );
not ( n65231 , n412099 );
or ( n65232 , n65229 , n65231 );
buf ( n412102 , n61583 );
buf ( n412103 , n61577 );
nand ( n65235 , n412102 , n412103 );
buf ( n412105 , n65235 );
buf ( n412106 , n412105 );
nand ( n65238 , n65232 , n412106 );
buf ( n412108 , n65238 );
buf ( n412109 , n412108 );
buf ( n412110 , n412096 );
or ( n65245 , n412109 , n412110 );
xor ( n65246 , n408704 , n408741 );
xor ( n65247 , n65246 , n408767 );
buf ( n412114 , n65247 );
buf ( n412115 , n412114 );
nand ( n65250 , n65245 , n412115 );
buf ( n412117 , n65250 );
buf ( n412118 , n412117 );
nand ( n65253 , C1 , n412118 );
buf ( n412120 , n65253 );
buf ( n412121 , n412120 );
xor ( n65256 , n412095 , n412121 );
buf ( n412123 , n65256 );
buf ( n412124 , n412123 );
xor ( n65259 , n409793 , n409797 );
xor ( n65260 , n65259 , n409851 );
buf ( n412127 , n65260 );
buf ( n412128 , n412127 );
xor ( n65263 , n412124 , n412128 );
buf ( n412130 , n65263 );
buf ( n412131 , n412130 );
xor ( n65266 , n412013 , n412021 );
xor ( n65267 , n65266 , n412044 );
buf ( n412134 , n65267 );
buf ( n412135 , n412134 );
buf ( n412136 , n50579 );
not ( n65271 , n412136 );
buf ( n412138 , n50584 );
buf ( n412139 , n384202 );
and ( n65274 , n412138 , n412139 );
not ( n65275 , n412138 );
buf ( n412142 , n384205 );
and ( n65277 , n65275 , n412142 );
nor ( n65278 , n65274 , n65277 );
buf ( n412145 , n65278 );
buf ( n412146 , n412145 );
not ( n65281 , n412146 );
or ( n65282 , n65271 , n65281 );
nand ( n65283 , n64620 , n51553 );
buf ( n412150 , n65283 );
nand ( n65285 , n65282 , n412150 );
buf ( n412152 , n65285 );
not ( n65287 , n412152 );
buf ( n412154 , n408649 );
buf ( n412155 , n384280 );
and ( n65290 , n412154 , n412155 );
not ( n65291 , n412154 );
buf ( n412158 , n58546 );
and ( n65293 , n65291 , n412158 );
nor ( n65294 , n65290 , n65293 );
buf ( n412161 , n65294 );
not ( n65296 , n412161 );
not ( n65297 , n395352 );
and ( n65298 , n65296 , n65297 );
and ( n65299 , n64060 , n395362 );
nor ( n65300 , n65298 , n65299 );
buf ( n412167 , n65300 );
not ( n65302 , n412167 );
buf ( n412169 , n65302 );
not ( n65304 , n412169 );
or ( n65305 , n65287 , n65304 );
buf ( n412172 , n412152 );
buf ( n412173 , n412169 );
nor ( n65308 , n412172 , n412173 );
buf ( n412175 , n65308 );
buf ( n412176 , n392740 );
not ( n65311 , n412176 );
buf ( n412178 , n64154 );
not ( n65313 , n412178 );
or ( n65314 , n65311 , n65313 );
buf ( n412181 , n64136 );
not ( n65316 , n412181 );
buf ( n412183 , n396534 );
not ( n65318 , n412183 );
or ( n65319 , n65316 , n65318 );
buf ( n412186 , n396537 );
buf ( n412187 , n44776 );
nand ( n65322 , n412186 , n412187 );
buf ( n412189 , n65322 );
buf ( n412190 , n412189 );
nand ( n65325 , n65319 , n412190 );
buf ( n412192 , n65325 );
buf ( n412193 , n412192 );
buf ( n412194 , n45260 );
nand ( n65329 , n412193 , n412194 );
buf ( n412196 , n65329 );
buf ( n412197 , n412196 );
nand ( n65332 , n65314 , n412197 );
buf ( n412199 , n65332 );
buf ( n412200 , n412199 );
not ( n65335 , n412200 );
buf ( n412202 , n65335 );
not ( n65337 , n412202 );
and ( n65338 , n63937 , n63342 );
not ( n65339 , n63937 );
and ( n65340 , n65339 , n63341 );
or ( n65341 , n65338 , n65340 );
xor ( n65342 , n63362 , n65341 );
not ( n65343 , n65342 );
and ( n65344 , n65337 , n65343 );
xor ( n65345 , n411297 , n64342 );
xnor ( n65346 , n65345 , n411334 );
buf ( n412213 , n412202 );
buf ( n412214 , n65342 );
nand ( n65349 , n412213 , n412214 );
buf ( n412216 , n65349 );
and ( n65351 , n65346 , n412216 );
nor ( n65352 , n65344 , n65351 );
or ( n65353 , n412175 , n65352 );
nand ( n65354 , n65305 , n65353 );
buf ( n412221 , n65354 );
xor ( n65356 , n410274 , n410295 );
xor ( n65357 , n65356 , n410992 );
buf ( n412224 , n65357 );
buf ( n412225 , n412224 );
buf ( n412226 , C0 );
buf ( n412227 , n412226 );
and ( n65382 , n412221 , n412225 );
or ( n65383 , C0 , n65382 );
buf ( n412230 , n65383 );
buf ( n412231 , n412230 );
xor ( n65386 , n412135 , n412231 );
xor ( n65387 , n410270 , n410997 );
xor ( n65388 , n65387 , n411101 );
buf ( n412235 , n65388 );
buf ( n412236 , n412235 );
and ( n65391 , n65386 , n412236 );
and ( n65392 , n412135 , n412231 );
or ( n65393 , n65391 , n65392 );
buf ( n412240 , n65393 );
buf ( n412241 , n412240 );
xor ( n65396 , n412131 , n412241 );
buf ( n412243 , n412114 );
not ( n65398 , n412243 );
buf ( n412245 , n65398 );
buf ( n412246 , n412245 );
not ( n65401 , n412246 );
xor ( n65402 , n412096 , n412108 );
buf ( n412249 , n65402 );
not ( n65404 , n412249 );
or ( n65405 , n65401 , n65404 );
buf ( n412252 , n65402 );
buf ( n412253 , n412245 );
or ( n65408 , n412252 , n412253 );
nand ( n65409 , n65405 , n65408 );
buf ( n412256 , n65409 );
buf ( n412257 , n412256 );
xor ( n65412 , n411108 , n411389 );
xor ( n65413 , n65412 , n411394 );
buf ( n412260 , n65413 );
buf ( n412261 , n412260 );
xor ( n65416 , n412257 , n412261 );
xor ( n65417 , n410321 , n410948 );
xor ( n65418 , n65417 , n410987 );
buf ( n412265 , n65418 );
not ( n65420 , n412265 );
buf ( n412267 , C0 );
xor ( n65435 , n411073 , n411084 );
xor ( n65436 , n65435 , n411090 );
buf ( n412270 , n65436 );
buf ( n412271 , n412270 );
or ( n65439 , n412267 , n412271 );
buf ( n412273 , n65439 );
not ( n65441 , n412273 );
or ( n65442 , n65420 , n65441 );
buf ( n412276 , C0 );
nand ( n65448 , n65442 , C1 );
not ( n65449 , n65448 );
or ( n65450 , n64065 , n64044 );
nand ( n65451 , n64044 , n64065 );
nand ( n65452 , n65450 , n65451 );
and ( n65453 , n65452 , n411094 );
not ( n65454 , n65452 );
not ( n65455 , n411094 );
and ( n65456 , n65454 , n65455 );
nor ( n65457 , n65453 , n65456 );
not ( n65458 , n65457 );
not ( n65459 , n65458 );
or ( n65460 , n65449 , n65459 );
not ( n65461 , n65457 );
and ( n65462 , n412273 , n412265 );
nor ( n65463 , n65462 , n412276 );
not ( n65464 , n65463 );
or ( n65465 , n65461 , n65464 );
not ( n65466 , n411367 );
not ( n65467 , n65466 );
and ( n65468 , n64408 , n65467 );
not ( n65469 , n64408 );
and ( n65470 , n65469 , n65466 );
nor ( n65471 , n65468 , n65470 );
buf ( n412301 , n64375 );
buf ( n65473 , n412301 );
buf ( n412303 , n65473 );
and ( n65475 , n65471 , n412303 );
not ( n65476 , n65471 );
not ( n65477 , n412303 );
and ( n65478 , n65476 , n65477 );
nor ( n65479 , n65475 , n65478 );
nand ( n65480 , n65465 , n65479 );
nand ( n65481 , n65460 , n65480 );
buf ( n412311 , n65481 );
and ( n65483 , n65416 , n412311 );
and ( n65484 , n412257 , n412261 );
or ( n65485 , n65483 , n65484 );
buf ( n412315 , n65485 );
buf ( n412316 , n412315 );
xor ( n65488 , n65396 , n412316 );
buf ( n412318 , n65488 );
buf ( n412319 , n412318 );
and ( n65491 , n65206 , n412319 );
and ( n65492 , n412083 , n412087 );
or ( n65493 , n65491 , n65492 );
buf ( n412323 , n65493 );
buf ( n412324 , n412323 );
xor ( n65496 , n412079 , n412324 );
buf ( n412326 , n61961 );
buf ( n412327 , C0 );
xor ( n65499 , n412326 , n412327 );
buf ( n412329 , n408947 );
xnor ( n65501 , n65499 , n412329 );
buf ( n412331 , n65501 );
buf ( n412332 , n412331 );
not ( n65504 , n412332 );
buf ( n412334 , n65504 );
not ( n65506 , n412334 );
xor ( n65507 , n411421 , n411423 );
and ( n65508 , n65507 , n411452 );
or ( n65510 , n65508 , C0 );
buf ( n412339 , n65510 );
not ( n65512 , n412339 );
not ( n65513 , n65512 );
or ( n65514 , n65506 , n65513 );
nand ( n65515 , n412339 , n412331 );
nand ( n65516 , n65514 , n65515 );
buf ( n412345 , n412051 );
buf ( n412346 , n65178 );
nand ( n65522 , n412345 , n412346 );
buf ( n412348 , n65522 );
and ( n65524 , n412348 , n412048 );
nor ( n65525 , C0 , n65524 );
buf ( n412351 , n65525 );
buf ( n65527 , n412351 );
buf ( n412353 , n65527 );
buf ( n412354 , n412353 );
not ( n65530 , n412354 );
buf ( n412356 , n65530 );
and ( n65532 , n65516 , n412356 );
not ( n65533 , n65516 );
and ( n65534 , n65533 , n412353 );
nor ( n65535 , n65532 , n65534 );
or ( n65536 , n412120 , n412094 );
and ( n65537 , n65536 , n412127 );
and ( n65538 , n412095 , n412121 );
buf ( n412364 , n65538 );
nor ( n65540 , n65537 , n412364 );
buf ( n65541 , n65540 );
not ( n65542 , n65541 );
xor ( n65543 , n408778 , n408782 );
xor ( n65544 , n65543 , n408787 );
buf ( n412370 , n65544 );
not ( n65546 , n412370 );
not ( n65547 , n65546 );
buf ( n412373 , n408990 );
buf ( n412374 , n408991 );
xor ( n65550 , n412373 , n412374 );
buf ( n412376 , n409855 );
xnor ( n65552 , n65550 , n412376 );
buf ( n412378 , n65552 );
buf ( n412379 , n412378 );
not ( n65555 , n412379 );
buf ( n412381 , n65555 );
not ( n65557 , n412381 );
or ( n65558 , n65547 , n65557 );
buf ( n412384 , n412370 );
buf ( n412385 , n412378 );
nand ( n65561 , n412384 , n412385 );
buf ( n412387 , n65561 );
nand ( n65563 , n65558 , n412387 );
not ( n65564 , n65563 );
or ( n65565 , n65542 , n65564 );
or ( n65566 , n65541 , n65563 );
nand ( n65567 , n65565 , n65566 );
xor ( n412393 , n65535 , n65567 );
xor ( n65569 , n412131 , n412241 );
and ( n65570 , n65569 , n412316 );
and ( n65571 , n412131 , n412241 );
or ( n65572 , n65570 , n65571 );
buf ( n412398 , n65572 );
xor ( n65574 , n412393 , n412398 );
buf ( n412400 , n65574 );
and ( n65576 , n65496 , n412400 );
and ( n65577 , n412079 , n412324 );
or ( n65578 , n65576 , n65577 );
buf ( n412404 , n65578 );
not ( n65580 , n412404 );
not ( n65581 , n65580 );
xor ( n65582 , n410266 , n411411 );
and ( n65583 , n65582 , n412076 );
and ( n65584 , n410266 , n411411 );
or ( n65585 , n65583 , n65584 );
buf ( n412411 , n65585 );
buf ( n412412 , n412411 );
xor ( n65588 , n65535 , n65567 );
and ( n65589 , n65588 , n412398 );
and ( n65590 , n65535 , n65567 );
or ( n65591 , n65589 , n65590 );
buf ( n412417 , n65591 );
xor ( n65593 , n412412 , n412417 );
xor ( n65594 , n61809 , n61965 );
xor ( n65595 , n65594 , n62861 );
buf ( n412421 , n65595 );
not ( n65597 , n65525 );
not ( n65598 , n65597 );
not ( n65599 , n412334 );
or ( n65600 , n65598 , n65599 );
not ( n65601 , n412331 );
not ( n65602 , n65525 );
or ( n65603 , n65601 , n65602 );
nand ( n65604 , n65603 , n412339 );
nand ( n65605 , n65600 , n65604 );
buf ( n412431 , n65605 );
and ( n65607 , n412421 , n412431 );
not ( n65608 , n412421 );
buf ( n412434 , n65605 );
not ( n65610 , n412434 );
buf ( n412436 , n65610 );
buf ( n412437 , n412436 );
and ( n65613 , n65608 , n412437 );
nor ( n65614 , n65607 , n65613 );
buf ( n412440 , n65614 );
buf ( n412441 , n65546 );
not ( n65617 , n412441 );
buf ( n412443 , n65540 );
not ( n65619 , n412443 );
or ( n65620 , n65617 , n65619 );
buf ( n412446 , n412381 );
nand ( n65622 , n65620 , n412446 );
buf ( n412448 , n65622 );
buf ( n412449 , n65540 );
not ( n65625 , n412449 );
not ( n65626 , n65546 );
buf ( n412452 , n65626 );
nand ( n65628 , n65625 , n412452 );
buf ( n412454 , n65628 );
nand ( n65630 , n412448 , n412454 );
xor ( n65631 , n412440 , n65630 );
buf ( n412457 , n408615 );
buf ( n412458 , n408794 );
xor ( n65634 , n412457 , n412458 );
buf ( n412460 , n408608 );
xnor ( n65636 , n65634 , n412460 );
buf ( n412462 , n65636 );
xor ( n65638 , n408045 , n408047 );
xor ( n65639 , n65638 , n408049 );
buf ( n412465 , n65639 );
buf ( n412466 , n412465 );
buf ( n412467 , n410020 );
not ( n65643 , n412467 );
buf ( n412469 , n63266 );
not ( n65645 , n412469 );
or ( n65646 , n65643 , n65645 );
buf ( n412472 , n63266 );
buf ( n412473 , n410020 );
or ( n65649 , n412472 , n412473 );
buf ( n412475 , n63263 );
nand ( n65651 , n65649 , n412475 );
buf ( n412477 , n65651 );
buf ( n412478 , n412477 );
nand ( n65654 , n65646 , n412478 );
buf ( n412480 , n65654 );
buf ( n412481 , n412480 );
xor ( n65657 , n412466 , n412481 );
xor ( n65658 , n409878 , n409882 );
xor ( n65659 , n65658 , n409927 );
buf ( n412485 , n65659 );
buf ( n412486 , n412485 );
xnor ( n65662 , n65657 , n412486 );
buf ( n412488 , n65662 );
buf ( n412489 , n412488 );
not ( n65665 , n412489 );
buf ( n412491 , n65665 );
and ( n65667 , n412462 , n412491 );
not ( n65668 , n412462 );
and ( n65669 , n65668 , n412488 );
or ( n65670 , n65667 , n65669 );
xor ( n65671 , n65631 , n65670 );
buf ( n412497 , n65671 );
xor ( n65673 , n65593 , n412497 );
buf ( n412499 , n65673 );
not ( n65675 , n412499 );
not ( n65676 , n65675 );
and ( n65677 , n65581 , n65676 );
not ( n65678 , n61780 );
not ( n65679 , n61786 );
not ( n65680 , n65679 );
or ( n65681 , n65678 , n65680 );
nand ( n65682 , n61764 , n61779 );
nand ( n65683 , n65681 , n65682 );
buf ( n412509 , n65683 );
buf ( n412510 , n61801 );
not ( n65686 , n412510 );
buf ( n412512 , n65686 );
buf ( n412513 , n412512 );
and ( n65689 , n412509 , n412513 );
not ( n65690 , n412509 );
buf ( n65691 , n61801 );
buf ( n412517 , n65691 );
and ( n65693 , n65690 , n412517 );
nor ( n65694 , n65689 , n65693 );
buf ( n412520 , n65694 );
buf ( n412521 , n412520 );
not ( n65697 , n412491 );
xor ( n65698 , n408615 , n408794 );
xor ( n65699 , n65698 , n408608 );
not ( n65700 , n65699 );
and ( n65701 , n65697 , n65700 );
buf ( n412527 , n412491 );
buf ( n412528 , n65699 );
nand ( n65704 , n412527 , n412528 );
buf ( n412530 , n65704 );
and ( n65706 , n412530 , n65631 );
nor ( n65707 , n65701 , n65706 );
buf ( n412533 , n65707 );
xor ( n65709 , n412521 , n412533 );
buf ( n412535 , n412465 );
not ( n65711 , n412535 );
buf ( n412537 , n412485 );
not ( n65713 , n412537 );
buf ( n412539 , n65713 );
buf ( n412540 , n412539 );
not ( n65716 , n412540 );
or ( n65717 , n65711 , n65716 );
buf ( n412543 , n412480 );
nand ( n65719 , n65717 , n412543 );
buf ( n412545 , n65719 );
buf ( n412546 , n412545 );
buf ( n412547 , n412465 );
not ( n65723 , n412547 );
buf ( n412549 , n412485 );
nand ( n65725 , n65723 , n412549 );
buf ( n412551 , n65725 );
buf ( n412552 , n412551 );
and ( n65728 , n412546 , n412552 );
buf ( n412554 , n65728 );
buf ( n412555 , n412554 );
and ( n65731 , n409931 , n409945 );
not ( n65732 , n409931 );
and ( n65733 , n65732 , n62944 );
nor ( n65734 , n65731 , n65733 );
xor ( n65735 , n62864 , n65734 );
buf ( n412561 , n65735 );
xor ( n65737 , n412555 , n412561 );
not ( n65738 , n65630 );
not ( n65739 , n65738 );
buf ( n412565 , n412436 );
buf ( n65741 , n412565 );
buf ( n412567 , n65741 );
not ( n65743 , n412567 );
and ( n65744 , n65739 , n65743 );
nand ( n65745 , n412567 , n65738 );
buf ( n412571 , n65595 );
buf ( n65747 , n412571 );
buf ( n412573 , n65747 );
and ( n65749 , n65745 , n412573 );
nor ( n65750 , n65744 , n65749 );
buf ( n412576 , n65750 );
xor ( n65752 , n65737 , n412576 );
buf ( n412578 , n65752 );
buf ( n412579 , n412578 );
xor ( n65755 , n65709 , n412579 );
buf ( n412581 , n65755 );
not ( n65757 , n412581 );
xor ( n65758 , n412412 , n412417 );
and ( n65759 , n65758 , n412497 );
and ( n65760 , n412412 , n412417 );
or ( n65761 , n65759 , n65760 );
buf ( n412587 , n65761 );
and ( n65763 , n65757 , n412587 );
nor ( n65764 , n65677 , n65763 );
not ( n65765 , n61467 );
not ( n65766 , n61476 );
not ( n65767 , n65766 );
or ( n65768 , n65765 , n65767 );
nand ( n65769 , n61476 , n61466 );
nand ( n65770 , n65768 , n65769 );
and ( n65771 , n65770 , n61059 );
not ( n65772 , n65770 );
and ( n65773 , n65772 , n61060 );
nor ( n65774 , n65771 , n65773 );
buf ( n412600 , n65774 );
xor ( n65776 , n412555 , n412561 );
and ( n65777 , n65776 , n412576 );
and ( n65778 , n412555 , n412561 );
or ( n65779 , n65777 , n65778 );
buf ( n412605 , n65779 );
buf ( n412606 , n412605 );
xor ( n65782 , n412600 , n412606 );
xor ( n65783 , n409958 , n61558 );
xnor ( n65784 , n65783 , n61803 );
buf ( n412610 , n65784 );
xor ( n65786 , n65782 , n412610 );
buf ( n412612 , n65786 );
buf ( n412613 , n412612 );
not ( n65789 , n412613 );
buf ( n412615 , n65789 );
xor ( n65791 , n412521 , n412533 );
and ( n65792 , n65791 , n412579 );
and ( n65793 , n412521 , n412533 );
or ( n65794 , n65792 , n65793 );
buf ( n412620 , n65794 );
buf ( n412621 , n412620 );
not ( n65797 , n412621 );
buf ( n412623 , n65797 );
nand ( n65799 , n412615 , n412623 );
xor ( n65800 , n412079 , n412324 );
xor ( n65801 , n65800 , n412400 );
buf ( n412627 , n65801 );
not ( n65803 , n41407 );
not ( n65804 , n394814 );
or ( n65805 , n65803 , n65804 );
nand ( n65806 , n388897 , n394817 );
nand ( n65807 , n65805 , n65806 );
not ( n65808 , n65807 );
and ( n65809 , n37336 , n37334 );
not ( n65810 , n65809 );
or ( n65811 , n65808 , n65810 );
not ( n65812 , n37336 );
nand ( n65813 , n65812 , n64202 );
nand ( n65814 , n65811 , n65813 );
buf ( n412640 , n65814 );
buf ( n412641 , n384545 );
buf ( n412642 , n402819 );
nor ( n65818 , n412641 , n412642 );
buf ( n412644 , n65818 );
buf ( n412645 , n412644 );
xor ( n65821 , n412640 , n412645 );
not ( n65822 , n43536 );
buf ( n412648 , n411504 );
not ( n65824 , n412648 );
buf ( n412650 , n41118 );
not ( n65826 , n412650 );
or ( n65827 , n65824 , n65826 );
buf ( n412653 , n27195 );
buf ( n412654 , n391024 );
nand ( n65830 , n412653 , n412654 );
buf ( n412656 , n65830 );
buf ( n412657 , n412656 );
nand ( n65833 , n65827 , n412657 );
buf ( n412659 , n65833 );
not ( n65835 , n412659 );
or ( n65836 , n65822 , n65835 );
nand ( n65837 , n411615 , n43515 );
nand ( n65838 , n65836 , n65837 );
buf ( n412664 , n65838 );
and ( n65840 , n65821 , n412664 );
and ( n65841 , n412640 , n412645 );
or ( n65842 , n65840 , n65841 );
buf ( n412668 , n65842 );
buf ( n412669 , n412668 );
buf ( n412670 , n392884 );
not ( n65846 , n412670 );
buf ( n412672 , n393525 );
not ( n65848 , n412672 );
or ( n65849 , n65846 , n65848 );
buf ( n412675 , n385473 );
buf ( n412676 , n392887 );
nand ( n65852 , n412675 , n412676 );
buf ( n412678 , n65852 );
buf ( n412679 , n412678 );
nand ( n65855 , n65849 , n412679 );
buf ( n412681 , n65855 );
buf ( n412682 , n412681 );
not ( n65858 , n412682 );
buf ( n412684 , n393544 );
not ( n65860 , n412684 );
or ( n65861 , n65858 , n65860 );
buf ( n412687 , n410357 );
buf ( n412688 , n41447 );
nand ( n65864 , n412687 , n412688 );
buf ( n412690 , n65864 );
buf ( n412691 , n412690 );
nand ( n65867 , n65861 , n412691 );
buf ( n412693 , n65867 );
buf ( n412694 , n412693 );
buf ( n412695 , n43286 );
not ( n65871 , n412695 );
buf ( n412697 , n40601 );
not ( n65873 , n412697 );
buf ( n412699 , n388409 );
not ( n65875 , n412699 );
or ( n65876 , n65873 , n65875 );
buf ( n412702 , n398292 );
not ( n65878 , n412702 );
buf ( n412704 , n40600 );
nand ( n65880 , n65878 , n412704 );
buf ( n412706 , n65880 );
buf ( n412707 , n412706 );
nand ( n65883 , n65876 , n412707 );
buf ( n412709 , n65883 );
buf ( n412710 , n412709 );
not ( n65886 , n412710 );
or ( n65887 , n65871 , n65886 );
buf ( n412713 , n411162 );
buf ( n412714 , n390362 );
nand ( n65890 , n412713 , n412714 );
buf ( n412716 , n65890 );
buf ( n412717 , n412716 );
nand ( n65893 , n65887 , n412717 );
buf ( n412719 , n65893 );
buf ( n412720 , n412719 );
xor ( n65896 , n412694 , n412720 );
buf ( n412722 , n389341 );
not ( n65898 , n412722 );
buf ( n412724 , n399164 );
not ( n65900 , n412724 );
or ( n65901 , n65898 , n65900 );
buf ( n412727 , n24049 );
buf ( n412728 , n393185 );
nand ( n65904 , n412727 , n412728 );
buf ( n412730 , n65904 );
buf ( n412731 , n412730 );
nand ( n65907 , n65901 , n412731 );
buf ( n412733 , n65907 );
buf ( n412734 , n412733 );
not ( n65910 , n412734 );
buf ( n412736 , n396622 );
not ( n65912 , n412736 );
or ( n65913 , n65910 , n65912 );
buf ( n412739 , n411211 );
buf ( n412740 , n41563 );
nand ( n65916 , n412739 , n412740 );
buf ( n412742 , n65916 );
buf ( n412743 , n412742 );
nand ( n65919 , n65913 , n412743 );
buf ( n412745 , n65919 );
buf ( n412746 , n412745 );
buf ( n412747 , n392611 );
not ( n65923 , n412747 );
buf ( n412749 , n49661 );
not ( n65925 , n412749 );
or ( n65926 , n65923 , n65925 );
buf ( n412752 , n49653 );
buf ( n412753 , n392620 );
nand ( n65929 , n412752 , n412753 );
buf ( n412755 , n65929 );
buf ( n412756 , n412755 );
nand ( n65932 , n65926 , n412756 );
buf ( n412758 , n65932 );
buf ( n412759 , n412758 );
not ( n65935 , n412759 );
buf ( n412761 , n399031 );
not ( n65937 , n412761 );
or ( n65938 , n65935 , n65937 );
nand ( n65939 , n64293 , n395469 );
buf ( n412765 , n65939 );
nand ( n65941 , n65938 , n412765 );
buf ( n412767 , n65941 );
buf ( n412768 , n412767 );
xor ( n65944 , n412746 , n412768 );
buf ( n412770 , n411715 );
not ( n65946 , n412770 );
buf ( n412772 , n65946 );
buf ( n412773 , n412772 );
buf ( n412774 , n388806 );
or ( n65950 , n412773 , n412774 );
buf ( n412776 , n405736 );
not ( n65952 , n412776 );
buf ( n412778 , n389856 );
not ( n65954 , n412778 );
or ( n65955 , n65952 , n65954 );
buf ( n412781 , n28297 );
buf ( n412782 , n388754 );
nand ( n65958 , n412781 , n412782 );
buf ( n412784 , n65958 );
buf ( n412785 , n412784 );
nand ( n65961 , n65955 , n412785 );
buf ( n412787 , n65961 );
buf ( n412788 , n412787 );
buf ( n412789 , n388746 );
nand ( n65965 , n412788 , n412789 );
buf ( n412791 , n65965 );
buf ( n412792 , n412791 );
nand ( n65968 , n65950 , n412792 );
buf ( n412794 , n65968 );
buf ( n412795 , n412794 );
and ( n65971 , n65944 , n412795 );
and ( n65972 , n412746 , n412768 );
or ( n65973 , n65971 , n65972 );
buf ( n412799 , n65973 );
buf ( n412800 , n412799 );
and ( n65976 , n65896 , n412800 );
and ( n65977 , n412694 , n412720 );
or ( n65978 , n65976 , n65977 );
buf ( n412804 , n65978 );
buf ( n412805 , n412804 );
xor ( n65981 , n412669 , n412805 );
buf ( n412807 , n45954 );
not ( n65983 , n412807 );
buf ( n412809 , n411950 );
not ( n65985 , n412809 );
or ( n65986 , n65983 , n65985 );
buf ( n412812 , n393369 );
not ( n65988 , n412812 );
buf ( n412814 , n41904 );
not ( n65990 , n412814 );
or ( n65991 , n65988 , n65990 );
buf ( n412817 , n388952 );
buf ( n412818 , n393381 );
nand ( n65994 , n412817 , n412818 );
buf ( n412820 , n65994 );
buf ( n412821 , n412820 );
nand ( n65997 , n65991 , n412821 );
buf ( n412823 , n65997 );
buf ( n412824 , n412823 );
buf ( n412825 , n393825 );
nand ( n66001 , n412824 , n412825 );
buf ( n412827 , n66001 );
buf ( n412828 , n412827 );
nand ( n66004 , n65986 , n412828 );
buf ( n412830 , n66004 );
buf ( n412831 , n412830 );
and ( n66007 , n65981 , n412831 );
and ( n66008 , n412669 , n412805 );
or ( n66009 , n66007 , n66008 );
buf ( n412835 , n66009 );
not ( n66011 , n64156 );
not ( n66012 , n64364 );
or ( n66013 , n66011 , n66012 );
or ( n66014 , n64364 , n64156 );
nand ( n66015 , n66013 , n66014 );
and ( n66016 , n66015 , n411344 );
not ( n66017 , n66015 );
and ( n66018 , n66017 , n64317 );
or ( n66019 , n66016 , n66018 );
xor ( n66020 , n412835 , n66019 );
buf ( n412846 , n358975 );
not ( n66022 , n412846 );
buf ( n412848 , n394392 );
not ( n66024 , n412848 );
or ( n66025 , n66022 , n66024 );
buf ( n412851 , n395885 );
buf ( n412852 , n402819 );
nand ( n66028 , n412851 , n412852 );
buf ( n412854 , n66028 );
buf ( n412855 , n412854 );
nand ( n66031 , n66025 , n412855 );
buf ( n412857 , n66031 );
buf ( n412858 , n412857 );
not ( n66034 , n412858 );
buf ( n412860 , n392659 );
not ( n66036 , n412860 );
or ( n66037 , n66034 , n66036 );
buf ( n412863 , n393602 );
buf ( n412864 , n411970 );
nand ( n66040 , n412863 , n412864 );
buf ( n412866 , n66040 );
buf ( n412867 , n412866 );
nand ( n66043 , n66037 , n412867 );
buf ( n412869 , n66043 );
buf ( n412870 , n412869 );
buf ( n412871 , n64222 );
buf ( n412872 , n64311 );
xor ( n66048 , n412871 , n412872 );
buf ( n412874 , n411169 );
xor ( n66050 , n66048 , n412874 );
buf ( n412876 , n66050 );
buf ( n412877 , n412876 );
xor ( n66053 , n412870 , n412877 );
xor ( n66054 , n410452 , n410888 );
xor ( n66055 , n66054 , n410918 );
buf ( n412881 , n66055 );
buf ( n412882 , n412881 );
not ( n66058 , n412882 );
xor ( n66059 , n409561 , n409564 );
xor ( n66060 , n66059 , n62571 );
xor ( n66061 , n63614 , n63884 );
xor ( n66062 , n66060 , n66061 );
not ( n66063 , n66062 );
buf ( n412889 , n66063 );
buf ( n412890 , n27320 );
not ( n66066 , n412890 );
buf ( n412892 , n66066 );
not ( n66068 , n412892 );
not ( n66069 , n407928 );
or ( n66070 , n66068 , n66069 );
nand ( n66071 , n40652 , n27320 );
nand ( n66072 , n66070 , n66071 );
buf ( n412898 , n66072 );
not ( n66074 , n412898 );
buf ( n412900 , n410907 );
not ( n66076 , n412900 );
or ( n66077 , n66074 , n66076 );
buf ( n412903 , n410901 );
buf ( n412904 , n409076 );
nand ( n66080 , n412903 , n412904 );
buf ( n412906 , n66080 );
buf ( n412907 , n412906 );
nand ( n66083 , n66077 , n412907 );
buf ( n412909 , n66083 );
buf ( n412910 , n412909 );
not ( n66086 , n412910 );
buf ( n412912 , n66086 );
buf ( n412913 , n412912 );
xor ( n66089 , n412889 , n412913 );
and ( n66090 , n388830 , n64782 );
buf ( n412916 , n41365 );
not ( n66092 , n412916 );
buf ( n412918 , n12480 );
not ( n66094 , n412918 );
buf ( n412920 , n66094 );
buf ( n412921 , n412920 );
not ( n66097 , n412921 );
or ( n66098 , n66092 , n66097 );
buf ( n412924 , n12480 );
buf ( n412925 , n410407 );
nand ( n66101 , n412924 , n412925 );
buf ( n412927 , n66101 );
buf ( n412928 , n412927 );
nand ( n66104 , n66098 , n412928 );
buf ( n412930 , n66104 );
buf ( n412931 , n412930 );
not ( n66107 , n412931 );
buf ( n412933 , n41374 );
nor ( n66109 , n66107 , n412933 );
buf ( n412935 , n66109 );
nor ( n66111 , n66090 , n412935 );
buf ( n412937 , n66111 );
and ( n66113 , n66089 , n412937 );
and ( n66114 , n412889 , n412913 );
or ( n66115 , n66113 , n66114 );
buf ( n412941 , n66115 );
buf ( n412942 , n412941 );
nand ( n66118 , n66058 , n412942 );
buf ( n412944 , n66118 );
buf ( n412945 , n412944 );
not ( n66121 , n412945 );
xor ( n66122 , n410602 , n410605 );
xor ( n66123 , n66122 , n410609 );
xor ( n66124 , n63770 , n63879 );
xor ( n66125 , n66123 , n66124 );
buf ( n412951 , n66125 );
not ( n66127 , n412951 );
not ( n66128 , n41371 );
buf ( n412954 , n66128 );
buf ( n412955 , n28353 );
not ( n66131 , n412955 );
not ( n66132 , n23841 );
buf ( n412958 , n66132 );
not ( n66134 , n412958 );
or ( n66135 , n66131 , n66134 );
buf ( n412961 , n41365 );
buf ( n412962 , n28353 );
not ( n66138 , n412962 );
buf ( n412964 , n66138 );
buf ( n412965 , n412964 );
nand ( n66141 , n412961 , n412965 );
buf ( n412967 , n66141 );
buf ( n412968 , n412967 );
nand ( n66144 , n66135 , n412968 );
buf ( n412970 , n66144 );
buf ( n412971 , n412970 );
and ( n66147 , n412954 , n412971 );
buf ( n412973 , n412930 );
buf ( n412974 , n41332 );
not ( n66150 , n412974 );
buf ( n412976 , n66150 );
buf ( n412977 , n412976 );
and ( n66153 , n412973 , n412977 );
nor ( n66154 , n66147 , n66153 );
buf ( n412980 , n66154 );
buf ( n412981 , n412980 );
nand ( n66157 , n66127 , n412981 );
buf ( n412983 , n66157 );
buf ( n412984 , n412983 );
buf ( n412985 , n58200 );
buf ( n412986 , n405391 );
and ( n66162 , n412985 , n412986 );
buf ( n412988 , n58201 );
buf ( n412989 , n405388 );
and ( n66165 , n412988 , n412989 );
nor ( n66166 , n66162 , n66165 );
buf ( n412992 , n66166 );
buf ( n412993 , n412992 );
buf ( n412994 , n405407 );
or ( n66170 , n412993 , n412994 );
buf ( n412996 , n410745 );
buf ( n412997 , n405384 );
or ( n66173 , n412996 , n412997 );
nand ( n66174 , n66170 , n66173 );
buf ( n413000 , n66174 );
buf ( n413001 , n410713 );
buf ( n413002 , n410732 );
or ( n66178 , n413001 , n413002 );
buf ( n413004 , n410735 );
nand ( n66180 , n66178 , n413004 );
buf ( n413006 , n66180 );
xor ( n66182 , n413000 , n413006 );
buf ( n413008 , n58090 );
buf ( n413009 , n59628 );
and ( n66185 , n413008 , n413009 );
buf ( n413011 , n405335 );
buf ( n413012 , n59457 );
and ( n66188 , n413011 , n413012 );
nor ( n66189 , n66185 , n66188 );
buf ( n413015 , n66189 );
buf ( n413016 , n413015 );
buf ( n413017 , n59637 );
or ( n66193 , n413016 , n413017 );
buf ( n413019 , n410785 );
buf ( n413020 , n59467 );
or ( n66196 , n413019 , n413020 );
nand ( n66197 , n66193 , n66196 );
buf ( n413023 , n66197 );
and ( n66199 , n66182 , n413023 );
and ( n66200 , n413000 , n413006 );
or ( n66201 , n66199 , n66200 );
buf ( n413027 , n66201 );
xor ( n66203 , n410641 , n410658 );
xor ( n66204 , n66203 , n410676 );
buf ( n413030 , n66204 );
buf ( n413031 , n413030 );
xor ( n66207 , n413027 , n413031 );
buf ( n413033 , n55846 );
buf ( n413034 , n62177 );
and ( n66210 , n413033 , n413034 );
buf ( n413036 , n403079 );
buf ( n413037 , n62159 );
and ( n66213 , n413036 , n413037 );
nor ( n66214 , n66210 , n66213 );
buf ( n413040 , n66214 );
buf ( n413041 , n413040 );
buf ( n413042 , n409429 );
or ( n66218 , n413041 , n413042 );
buf ( n413044 , n410694 );
buf ( n413045 , n409170 );
or ( n66221 , n413044 , n413045 );
nand ( n66222 , n66218 , n66221 );
buf ( n413048 , n66222 );
buf ( n413049 , n413048 );
buf ( n413050 , n54297 );
buf ( n413051 , n63625 );
and ( n66227 , n413050 , n413051 );
buf ( n413053 , n55919 );
buf ( n413054 , n63629 );
and ( n66230 , n413053 , n413054 );
nor ( n66231 , n66227 , n66230 );
buf ( n413057 , n66231 );
buf ( n413058 , n413057 );
buf ( n413059 , n410635 );
or ( n66235 , n413058 , n413059 );
buf ( n413061 , n410631 );
buf ( n413062 , n409504 );
or ( n66238 , n413061 , n413062 );
nand ( n66239 , n66235 , n66238 );
buf ( n413065 , n66239 );
buf ( n413066 , n413065 );
xor ( n66242 , n413049 , n413066 );
buf ( n413068 , n63564 );
buf ( n413069 , n403146 );
and ( n66245 , n413068 , n413069 );
buf ( n413071 , n63564 );
not ( n66247 , n413071 );
buf ( n413073 , n66247 );
buf ( n413074 , n413073 );
buf ( n413075 , n401695 );
and ( n66251 , n413074 , n413075 );
nor ( n66252 , n66245 , n66251 );
buf ( n413078 , n66252 );
buf ( n413079 , n413078 );
buf ( n413080 , n403158 );
or ( n66256 , n413079 , n413080 );
buf ( n413082 , n410825 );
buf ( n413083 , n403167 );
or ( n66259 , n413082 , n413083 );
nand ( n66260 , n66256 , n66259 );
buf ( n413086 , n66260 );
buf ( n413087 , n413086 );
not ( n66263 , n54000 );
not ( n66264 , n66263 );
not ( n66265 , n54233 );
or ( n66266 , n66264 , n66265 );
not ( n66267 , n54236 );
nand ( n66268 , n66266 , n66267 );
nand ( n66269 , n53968 , n54238 );
xnor ( n66270 , n66268 , n66269 );
buf ( n413096 , n66270 );
not ( n66272 , n413096 );
buf ( n413098 , n66272 );
buf ( n413099 , n413098 );
buf ( n413100 , n403083 );
or ( n66276 , n413099 , n413100 );
buf ( n413102 , n63707 );
not ( n66278 , n413102 );
buf ( n413104 , n66278 );
buf ( n413105 , n413104 );
buf ( n413106 , n403092 );
or ( n66282 , n413105 , n413106 );
nand ( n66283 , n66276 , n66282 );
buf ( n413109 , n66283 );
buf ( n413110 , n413109 );
xor ( n66286 , n413087 , n413110 );
buf ( n413112 , n56064 );
not ( n66288 , n413112 );
buf ( n413114 , n59596 );
buf ( n413115 , n405215 );
and ( n66291 , n413114 , n413115 );
buf ( n413117 , n409146 );
buf ( n413118 , n58061 );
and ( n66294 , n413117 , n413118 );
nor ( n66295 , n66291 , n66294 );
buf ( n413121 , n66295 );
buf ( n413122 , n413121 );
not ( n66298 , n413122 );
buf ( n413124 , n66298 );
buf ( n413125 , n413124 );
not ( n66301 , n413125 );
or ( n66302 , n66288 , n66301 );
buf ( n413128 , n410843 );
buf ( n413129 , n405476 );
or ( n66305 , n413128 , n413129 );
nand ( n66306 , n66302 , n66305 );
buf ( n413132 , n66306 );
buf ( n413133 , n413132 );
and ( n66309 , n66286 , n413133 );
and ( n413135 , n413087 , n413110 );
or ( n66311 , n66309 , n413135 );
buf ( n413137 , n66311 );
buf ( n413138 , n413137 );
and ( n66314 , n66242 , n413138 );
and ( n66315 , n413049 , n413066 );
or ( n66316 , n66314 , n66315 );
buf ( n413142 , n66316 );
buf ( n413143 , n413142 );
and ( n66319 , n66207 , n413143 );
and ( n66320 , n413027 , n413031 );
or ( n66321 , n66319 , n66320 );
buf ( n413147 , n66321 );
xor ( n66323 , n410681 , n410685 );
xor ( n66324 , n66323 , n410759 );
buf ( n413150 , n66324 );
xor ( n66326 , n413147 , n413150 );
xor ( n66327 , n410468 , n410484 );
xor ( n66328 , n66327 , n410501 );
xor ( n66329 , n410774 , n63861 );
xor ( n66330 , n66328 , n66329 );
and ( n66331 , n66326 , n66330 );
and ( n66332 , n413147 , n413150 );
or ( n66333 , n66331 , n66332 );
not ( n66334 , n66333 );
not ( n66335 , n63870 );
and ( n66336 , n63875 , n66335 );
not ( n66337 , n63878 );
and ( n66338 , n63875 , n66337 );
nor ( n66339 , n66336 , n66338 );
not ( n66340 , n63866 );
not ( n66341 , n63875 );
nand ( n66342 , n66340 , n66341 , n410867 );
not ( n66343 , n63866 );
nor ( n66344 , n66343 , n410867 );
nand ( n66345 , n66341 , n66344 );
and ( n66346 , n66339 , n66342 , n66345 );
nand ( n66347 , n66334 , n66346 );
not ( n66348 , n66347 );
xor ( n66349 , n410703 , n410736 );
xor ( n66350 , n66349 , n410754 );
buf ( n413176 , n66350 );
xor ( n66352 , n410793 , n410799 );
xor ( n66353 , n66352 , n410856 );
and ( n66354 , n413176 , n66353 );
xor ( n66355 , n410817 , n410834 );
xor ( n66356 , n66355 , n410852 );
buf ( n413182 , n66356 );
and ( n66358 , n66267 , n66263 );
xor ( n66359 , n66358 , n54233 );
buf ( n413185 , n66359 );
not ( n66361 , n413185 );
buf ( n413187 , n66361 );
buf ( n413188 , n413187 );
buf ( n413189 , n403083 );
or ( n66365 , n413188 , n413189 );
buf ( n413191 , n413098 );
buf ( n413192 , n403092 );
or ( n66368 , n413191 , n413192 );
nand ( n66369 , n66365 , n66368 );
buf ( n413195 , n66369 );
buf ( n413196 , n413195 );
buf ( n413197 , n63707 );
buf ( n413198 , n403146 );
and ( n66374 , n413197 , n413198 );
buf ( n413200 , n413104 );
buf ( n413201 , n401695 );
and ( n66377 , n413200 , n413201 );
nor ( n66378 , n66374 , n66377 );
buf ( n413204 , n66378 );
buf ( n413205 , n413204 );
buf ( n413206 , n403158 );
or ( n66382 , n413205 , n413206 );
buf ( n413208 , n413078 );
buf ( n413209 , n403167 );
or ( n66385 , n413208 , n413209 );
nand ( n66386 , n66382 , n66385 );
buf ( n413212 , n66386 );
buf ( n413213 , n413212 );
and ( n66389 , n413196 , n413213 );
buf ( n413215 , n66389 );
buf ( n413216 , n413215 );
buf ( n413217 , n62278 );
buf ( n413218 , n55905 );
and ( n66394 , n413217 , n413218 );
buf ( n413220 , n409474 );
buf ( n413221 , n55895 );
and ( n66397 , n413220 , n413221 );
nor ( n66398 , n66394 , n66397 );
buf ( n413224 , n66398 );
buf ( n413225 , n413224 );
buf ( n413226 , n403120 );
or ( n66402 , n413225 , n413226 );
buf ( n413228 , n410808 );
buf ( n413229 , n403133 );
or ( n66405 , n413228 , n413229 );
nand ( n66406 , n66402 , n66405 );
buf ( n413232 , n66406 );
buf ( n413233 , n413232 );
xor ( n66409 , n413216 , n413233 );
buf ( n413235 , n54336 );
buf ( n66411 , n62495 );
buf ( n413237 , n66411 );
and ( n66413 , n413235 , n413237 );
buf ( n413239 , n401699 );
buf ( n413240 , n62496 );
and ( n66416 , n413239 , n413240 );
nor ( n66417 , n66413 , n66416 );
buf ( n413243 , n66417 );
buf ( n413244 , n413243 );
buf ( n413245 , n410724 );
or ( n66421 , n413244 , n413245 );
buf ( n413247 , n410729 );
nand ( n66423 , n66421 , n413247 );
buf ( n413249 , n66423 );
buf ( n413250 , n413249 );
and ( n66426 , n66409 , n413250 );
and ( n66427 , n413216 , n413233 );
or ( n66428 , n66426 , n66427 );
buf ( n413254 , n66428 );
xor ( n66430 , n413182 , n413254 );
buf ( n413256 , n58042 );
buf ( n413257 , n63625 );
and ( n66433 , n413256 , n413257 );
buf ( n413259 , n403088 );
buf ( n413260 , n63629 );
and ( n66436 , n413259 , n413260 );
nor ( n66437 , n66433 , n66436 );
buf ( n413263 , n66437 );
buf ( n413264 , n413263 );
buf ( n413265 , n410635 );
or ( n66441 , n413264 , n413265 );
buf ( n413267 , n413057 );
buf ( n413268 , n409504 );
or ( n66444 , n413267 , n413268 );
nand ( n66445 , n66441 , n66444 );
buf ( n413271 , n66445 );
buf ( n413272 , n413271 );
buf ( n413273 , n58352 );
buf ( n413274 , n405391 );
and ( n66450 , n413273 , n413274 );
buf ( n413276 , n406571 );
buf ( n413277 , n405388 );
and ( n66453 , n413276 , n413277 );
nor ( n66454 , n66450 , n66453 );
buf ( n413280 , n66454 );
buf ( n413281 , n413280 );
buf ( n413282 , n405407 );
or ( n66458 , n413281 , n413282 );
buf ( n413284 , n412992 );
buf ( n413285 , n405384 );
or ( n66461 , n413284 , n413285 );
nand ( n66462 , n66458 , n66461 );
buf ( n413288 , n66462 );
buf ( n413289 , n413288 );
xor ( n66465 , n413272 , n413289 );
buf ( n413291 , n59468 );
not ( n66467 , n413291 );
buf ( n413293 , n58166 );
buf ( n413294 , n59628 );
and ( n66470 , n413293 , n413294 );
buf ( n413296 , n58205 );
buf ( n413297 , n59457 );
and ( n66473 , n413296 , n413297 );
nor ( n66474 , n66470 , n66473 );
buf ( n413300 , n66474 );
buf ( n413301 , n413300 );
not ( n66477 , n413301 );
buf ( n413303 , n66477 );
buf ( n413304 , n413303 );
not ( n66480 , n413304 );
or ( n66481 , n66467 , n66480 );
buf ( n413307 , n413015 );
buf ( n413308 , n59467 );
or ( n66484 , n413307 , n413308 );
nand ( n66485 , n66481 , n66484 );
buf ( n413311 , n66485 );
buf ( n413312 , n413311 );
and ( n66488 , n66465 , n413312 );
and ( n66489 , n413272 , n413289 );
or ( n66490 , n66488 , n66489 );
buf ( n413316 , n66490 );
and ( n66492 , n66430 , n413316 );
and ( n66493 , n413182 , n413254 );
or ( n66494 , n66492 , n66493 );
xor ( n66495 , n410793 , n410799 );
xor ( n66496 , n66495 , n410856 );
and ( n66497 , n66494 , n66496 );
and ( n66498 , n413176 , n66494 );
or ( n66499 , n66354 , n66497 , n66498 );
xor ( n66500 , n413147 , n413150 );
xor ( n66501 , n66500 , n66330 );
xor ( n66502 , n66499 , n66501 );
xor ( n66503 , n413027 , n413031 );
xor ( n66504 , n66503 , n413143 );
buf ( n413330 , n66504 );
buf ( n413331 , n413330 );
xor ( n66507 , n413087 , n413110 );
xor ( n66508 , n66507 , n413133 );
buf ( n413334 , n66508 );
buf ( n413335 , n55984 );
buf ( n413336 , n62177 );
and ( n66512 , n413335 , n413336 );
buf ( n413338 , n58135 );
buf ( n413339 , n62159 );
and ( n66515 , n413338 , n413339 );
nor ( n66516 , n66512 , n66515 );
buf ( n413342 , n66516 );
buf ( n413343 , n413342 );
buf ( n413344 , n409429 );
or ( n66520 , n413343 , n413344 );
buf ( n413346 , n413040 );
buf ( n413347 , n409170 );
or ( n66523 , n413346 , n413347 );
nand ( n66524 , n66520 , n66523 );
buf ( n413350 , n66524 );
xor ( n66526 , n413334 , n413350 );
buf ( n413352 , n62139 );
buf ( n413353 , n405215 );
and ( n66529 , n413352 , n413353 );
buf ( n413355 , n409140 );
buf ( n413356 , n58061 );
and ( n66532 , n413355 , n413356 );
nor ( n66533 , n66529 , n66532 );
buf ( n413359 , n66533 );
buf ( n413360 , n413359 );
buf ( n413361 , n403293 );
or ( n66537 , n413360 , n413361 );
buf ( n413363 , n413121 );
buf ( n413364 , n405476 );
or ( n66540 , n413363 , n413364 );
nand ( n66541 , n66537 , n66540 );
buf ( n413367 , n66541 );
buf ( n413368 , n62467 );
buf ( n413369 , n55905 );
and ( n66545 , n413368 , n413369 );
buf ( n413371 , n409468 );
buf ( n413372 , n55895 );
and ( n66548 , n413371 , n413372 );
nor ( n66549 , n66545 , n66548 );
buf ( n413375 , n66549 );
buf ( n413376 , n413375 );
buf ( n413377 , n403120 );
or ( n66553 , n413376 , n413377 );
buf ( n413379 , n413224 );
buf ( n413380 , n403133 );
or ( n66556 , n413379 , n413380 );
nand ( n66557 , n66553 , n66556 );
buf ( n413383 , n66557 );
xor ( n66559 , n413367 , n413383 );
xor ( n66560 , n413196 , n413213 );
buf ( n413386 , n66560 );
and ( n66562 , n66559 , n413386 );
and ( n66563 , n413367 , n413383 );
or ( n66564 , n66562 , n66563 );
and ( n66565 , n66526 , n66564 );
and ( n66566 , n413334 , n413350 );
or ( n66567 , n66565 , n66566 );
xor ( n66568 , n413000 , n413006 );
xor ( n66569 , n66568 , n413023 );
and ( n66570 , n66567 , n66569 );
xor ( n66571 , n413049 , n413066 );
xor ( n66572 , n66571 , n413138 );
buf ( n413398 , n66572 );
xor ( n66574 , n413000 , n413006 );
xor ( n66575 , n66574 , n413023 );
and ( n66576 , n413398 , n66575 );
and ( n66577 , n66567 , n413398 );
or ( n66578 , n66570 , n66576 , n66577 );
buf ( n413404 , n66578 );
xor ( n66580 , n413331 , n413404 );
xor ( n66581 , n410793 , n410799 );
xor ( n66582 , n66581 , n410856 );
xor ( n66583 , n413176 , n66494 );
xor ( n66584 , n66582 , n66583 );
buf ( n413410 , n66584 );
and ( n66586 , n66580 , n413410 );
and ( n66587 , n413331 , n413404 );
or ( n66588 , n66586 , n66587 );
buf ( n413414 , n66588 );
and ( n66590 , n66502 , n413414 );
and ( n66591 , n66499 , n66501 );
or ( n66592 , n66590 , n66591 );
not ( n66593 , n66592 );
or ( n66594 , n66348 , n66593 );
not ( n66595 , n66346 );
nand ( n66596 , n66595 , n66333 );
nand ( n66597 , n66594 , n66596 );
buf ( n413423 , n66597 );
and ( n66599 , n412984 , n413423 );
buf ( n413425 , n66125 );
not ( n66601 , n413425 );
buf ( n413427 , n412980 );
nor ( n66603 , n66601 , n413427 );
buf ( n413429 , n66603 );
buf ( n413430 , n413429 );
nor ( n66606 , n66599 , n413430 );
buf ( n413432 , n66606 );
buf ( n413433 , n413432 );
and ( n66609 , n64812 , n389162 );
not ( n66610 , n64268 );
not ( n66611 , n407940 );
or ( n66612 , n66610 , n66611 );
buf ( n413438 , n12471 );
buf ( n413439 , n64273 );
nand ( n66615 , n413438 , n413439 );
buf ( n413441 , n66615 );
nand ( n66617 , n66612 , n413441 );
not ( n66618 , n66617 );
nor ( n66619 , n66618 , n41710 );
nor ( n66620 , n66609 , n66619 );
buf ( n413446 , n66620 );
xor ( n66622 , n413433 , n413446 );
buf ( n413448 , n389359 );
not ( n66624 , n413448 );
buf ( n413450 , n24071 );
not ( n66626 , n413450 );
or ( n66627 , n66624 , n66626 );
buf ( n413453 , n60880 );
buf ( n413454 , n389356 );
nand ( n66630 , n413453 , n413454 );
buf ( n413456 , n66630 );
buf ( n413457 , n413456 );
nand ( n66633 , n66627 , n413457 );
buf ( n413459 , n66633 );
buf ( n413460 , n413459 );
not ( n66636 , n413460 );
buf ( n413462 , n66636 );
not ( n66638 , n413462 );
not ( n66639 , n42951 );
and ( n66640 , n66638 , n66639 );
and ( n66641 , n42924 , n64791 );
nor ( n66642 , n66640 , n66641 );
buf ( n413468 , n66642 );
and ( n66644 , n66622 , n413468 );
and ( n66645 , n413433 , n413446 );
or ( n66646 , n66644 , n66645 );
buf ( n413472 , n66646 );
buf ( n413473 , n413472 );
not ( n66649 , n413473 );
buf ( n413475 , n66649 );
buf ( n413476 , n413475 );
not ( n66652 , n413476 );
or ( n66653 , n66121 , n66652 );
buf ( n413479 , n412941 );
not ( n66655 , n413479 );
buf ( n413481 , n412881 );
nand ( n66657 , n66655 , n413481 );
buf ( n413483 , n66657 );
buf ( n413484 , n413483 );
nand ( n66660 , n66653 , n413484 );
buf ( n413486 , n66660 );
buf ( n413487 , n413486 );
xor ( n66663 , n411235 , n64286 );
xnor ( n66664 , n66663 , n64309 );
buf ( n413490 , n66664 );
xor ( n66666 , n413487 , n413490 );
buf ( n413492 , n397498 );
not ( n66668 , n413492 );
buf ( n413494 , n388299 );
not ( n66670 , n413494 );
or ( n66671 , n66668 , n66670 );
buf ( n413497 , n400355 );
buf ( n413498 , n397495 );
nand ( n66674 , n413497 , n413498 );
buf ( n413500 , n66674 );
buf ( n413501 , n413500 );
nand ( n66677 , n66671 , n413501 );
buf ( n413503 , n66677 );
buf ( n413504 , n413503 );
not ( n66680 , n413504 );
buf ( n413506 , n383894 );
not ( n66682 , n413506 );
or ( n66683 , n66680 , n66682 );
buf ( n413509 , n411634 );
buf ( n413510 , n383907 );
nand ( n66686 , n413509 , n413510 );
buf ( n413512 , n66686 );
buf ( n413513 , n413512 );
nand ( n66689 , n66683 , n413513 );
buf ( n413515 , n66689 );
buf ( n413516 , n413515 );
and ( n66692 , n66666 , n413516 );
and ( n66693 , n413487 , n413490 );
or ( n66694 , n66692 , n66693 );
buf ( n413520 , n66694 );
buf ( n413521 , n413520 );
and ( n66697 , n66053 , n413521 );
and ( n66698 , n412870 , n412877 );
or ( n66699 , n66697 , n66698 );
buf ( n413525 , n66699 );
and ( n66701 , n66020 , n413525 );
and ( n66702 , n412835 , n66019 );
or ( n66703 , n66701 , n66702 );
buf ( n413529 , n412001 );
buf ( n413530 , n65016 );
xor ( n66706 , n413529 , n413530 );
buf ( n413532 , n411861 );
xor ( n66708 , n66706 , n413532 );
buf ( n413534 , n66708 );
or ( n66710 , n66703 , n413534 );
buf ( n413536 , n411575 );
not ( n66712 , n413536 );
buf ( n413538 , n411838 );
not ( n66714 , n413538 );
and ( n66715 , n66712 , n66714 );
buf ( n413541 , n411838 );
buf ( n413542 , n411575 );
and ( n66718 , n413541 , n413542 );
nor ( n66719 , n66715 , n66718 );
buf ( n413545 , n66719 );
buf ( n413546 , n413545 );
buf ( n413547 , n64603 );
and ( n66723 , n413546 , n413547 );
not ( n66724 , n413546 );
buf ( n413550 , n411846 );
and ( n66726 , n66724 , n413550 );
nor ( n66727 , n66723 , n66726 );
buf ( n413553 , n66727 );
nand ( n66729 , n66710 , n413553 );
buf ( n413555 , n66729 );
buf ( n413556 , n413534 );
buf ( n413557 , n66703 );
nand ( n66733 , n413556 , n413557 );
buf ( n413559 , n66733 );
buf ( n413560 , n413559 );
nand ( n66736 , n413555 , n413560 );
buf ( n413562 , n66736 );
not ( n66738 , n413562 );
xor ( n66739 , n412135 , n412231 );
xor ( n66740 , n66739 , n412236 );
buf ( n413566 , n66740 );
buf ( n413567 , n413566 );
not ( n66743 , n413567 );
buf ( n413569 , n66743 );
buf ( n413570 , n413569 );
xor ( n66746 , n65094 , n411855 );
buf ( n413572 , n66746 );
buf ( n413573 , n64900 );
and ( n66749 , n413572 , n413573 );
not ( n66750 , n413572 );
buf ( n413576 , n64900 );
not ( n66752 , n413576 );
buf ( n413578 , n66752 );
buf ( n413579 , n413578 );
and ( n66755 , n66750 , n413579 );
nor ( n66756 , n66749 , n66755 );
buf ( n413582 , n66756 );
buf ( n413583 , n413582 );
not ( n66759 , n413583 );
buf ( n413585 , n66759 );
buf ( n413586 , n413585 );
nand ( n66762 , n413570 , n413586 );
buf ( n413588 , n66762 );
not ( n66764 , n413588 );
or ( n66765 , n66738 , n66764 );
nand ( n66766 , n413566 , n413582 );
nand ( n66767 , n66765 , n66766 );
buf ( n66768 , n66767 );
not ( n66769 , n66768 );
not ( n66770 , n66769 );
xor ( n66771 , n412083 , n412087 );
xor ( n66772 , n66771 , n412319 );
buf ( n413598 , n66772 );
buf ( n413599 , n413598 );
not ( n66775 , n413599 );
buf ( n413601 , n66775 );
not ( n66777 , n413601 );
or ( n66778 , n66770 , n66777 );
xor ( n66779 , n412257 , n412261 );
xor ( n66780 , n66779 , n412311 );
buf ( n413606 , n66780 );
not ( n66782 , n413606 );
xor ( n66783 , n412221 , n412225 );
xor ( n66784 , n66783 , n412227 );
buf ( n413610 , n66784 );
not ( n66786 , n413610 );
xor ( n66805 , n412640 , n412645 );
xor ( n66806 , n66805 , n412664 );
buf ( n413614 , n66806 );
buf ( n413615 , n413614 );
buf ( n413616 , n55543 );
not ( n66810 , n413616 );
buf ( n413618 , n388299 );
not ( n66812 , n413618 );
or ( n66813 , n66810 , n66812 );
buf ( n413621 , n388263 );
buf ( n413622 , n51185 );
nand ( n66816 , n413621 , n413622 );
buf ( n413624 , n66816 );
buf ( n413625 , n413624 );
nand ( n66819 , n66813 , n413625 );
buf ( n413627 , n66819 );
buf ( n413628 , n413627 );
not ( n66822 , n413628 );
buf ( n413630 , n383891 );
not ( n66824 , n413630 );
or ( n66825 , n66822 , n66824 );
buf ( n413633 , n413503 );
buf ( n413634 , n383904 );
nand ( n66828 , n413633 , n413634 );
buf ( n413636 , n66828 );
buf ( n413637 , n413636 );
nand ( n66831 , n66825 , n413637 );
buf ( n413639 , n66831 );
buf ( n413640 , n413639 );
buf ( n413641 , n392224 );
not ( n66835 , n413641 );
buf ( n413643 , n66835 );
not ( n66837 , n413643 );
buf ( n413645 , n399986 );
not ( n66839 , n413645 );
buf ( n413647 , n390704 );
not ( n66841 , n413647 );
or ( n66842 , n66839 , n66841 );
buf ( n413650 , n397277 );
buf ( n413651 , n44776 );
nand ( n66845 , n413650 , n413651 );
buf ( n413653 , n66845 );
buf ( n413654 , n413653 );
nand ( n66848 , n66842 , n413654 );
buf ( n413656 , n66848 );
not ( n66850 , n413656 );
or ( n66851 , n66837 , n66850 );
not ( n66852 , n64136 );
not ( n66853 , n40759 );
or ( n66854 , n66852 , n66853 );
buf ( n413662 , n40760 );
buf ( n413663 , n44776 );
nand ( n66857 , n413662 , n413663 );
buf ( n413665 , n66857 );
nand ( n66859 , n66854 , n413665 );
nand ( n66860 , n66859 , n45260 );
nand ( n66861 , n66851 , n66860 );
buf ( n413669 , n66861 );
xor ( n66863 , n413640 , n413669 );
xor ( n66864 , n412746 , n412768 );
xor ( n66865 , n66864 , n412795 );
buf ( n413673 , n66865 );
buf ( n413674 , n413673 );
and ( n66868 , n66863 , n413674 );
and ( n66869 , n413640 , n413669 );
or ( n66870 , n66868 , n66869 );
buf ( n413678 , n66870 );
buf ( n413679 , n413678 );
xor ( n66873 , n413615 , n413679 );
buf ( n413681 , n395349 );
not ( n66875 , n413681 );
buf ( n413683 , n47863 );
not ( n66877 , n413683 );
buf ( n413685 , n46161 );
not ( n66879 , n413685 );
or ( n66880 , n66877 , n66879 );
buf ( n413688 , n38155 );
buf ( n413689 , n395312 );
nand ( n66883 , n413688 , n413689 );
buf ( n413691 , n66883 );
buf ( n413692 , n413691 );
nand ( n66886 , n66880 , n413692 );
buf ( n413694 , n66886 );
buf ( n413695 , n413694 );
not ( n66889 , n413695 );
or ( n66890 , n66875 , n66889 );
buf ( n413698 , n47863 );
not ( n66892 , n413698 );
buf ( n413700 , n390651 );
not ( n66894 , n413700 );
or ( n66895 , n66892 , n66894 );
buf ( n413703 , n36509 );
buf ( n413704 , n395315 );
nand ( n66898 , n413703 , n413704 );
buf ( n413706 , n66898 );
buf ( n413707 , n413706 );
nand ( n66901 , n66895 , n413707 );
buf ( n413709 , n66901 );
buf ( n413710 , n413709 );
buf ( n413711 , n395362 );
nand ( n66905 , n413710 , n413711 );
buf ( n413713 , n66905 );
buf ( n413714 , n413713 );
nand ( n66908 , n66890 , n413714 );
buf ( n413716 , n66908 );
buf ( n413717 , n413716 );
and ( n66911 , n66873 , n413717 );
and ( n66912 , n413615 , n413679 );
or ( n66913 , n66911 , n66912 );
buf ( n413721 , n66913 );
buf ( n413722 , n413721 );
not ( n66916 , n413722 );
buf ( n413724 , n66916 );
not ( n66918 , n413724 );
or ( n66919 , C0 , n66918 );
xor ( n66920 , n411788 , n411806 );
xor ( n66921 , n66920 , n411824 );
buf ( n413729 , n66921 );
nand ( n66923 , n66919 , n413729 );
nand ( n66925 , n66923 , C1 );
not ( n66926 , n66925 );
not ( n66927 , n66926 );
buf ( n413734 , n411693 );
not ( n66929 , n413734 );
buf ( n413736 , n411599 );
not ( n66931 , n413736 );
or ( n66932 , n66929 , n66931 );
buf ( n413739 , n411596 );
buf ( n413740 , n411696 );
nand ( n66935 , n413739 , n413740 );
buf ( n413742 , n66935 );
buf ( n413743 , n413742 );
nand ( n66938 , n66932 , n413743 );
buf ( n413745 , n66938 );
buf ( n413746 , n413745 );
buf ( n413747 , n411828 );
not ( n66942 , n413747 );
buf ( n413749 , n66942 );
buf ( n413750 , n413749 );
and ( n66945 , n413746 , n413750 );
not ( n66946 , n413746 );
buf ( n413753 , n411828 );
and ( n66948 , n66946 , n413753 );
nor ( n66949 , n66945 , n66948 );
buf ( n413756 , n66949 );
buf ( n413757 , n413756 );
buf ( n66952 , n413757 );
buf ( n413759 , n66952 );
not ( n66954 , n413759 );
and ( n66955 , n66927 , n66954 );
buf ( n413762 , n66926 );
buf ( n413763 , n413759 );
nand ( n66958 , n413762 , n413763 );
buf ( n413765 , n66958 );
not ( n66960 , n413709 );
not ( n66961 , n395349 );
or ( n66962 , n66960 , n66961 );
not ( n66963 , n412161 );
nand ( n66964 , n66963 , n395362 );
nand ( n66965 , n66962 , n66964 );
buf ( n413772 , n66965 );
not ( n66967 , n413772 );
buf ( n413774 , n66967 );
buf ( n413775 , n413774 );
not ( n66970 , n413775 );
buf ( n413777 , n36434 );
not ( n66972 , n413777 );
buf ( n413779 , n36396 );
not ( n66974 , n413779 );
buf ( n413781 , n399283 );
not ( n66976 , n413781 );
and ( n66977 , n66974 , n66976 );
buf ( n413784 , n40839 );
buf ( n413785 , n399283 );
and ( n66980 , n413784 , n413785 );
nor ( n66981 , n66977 , n66980 );
buf ( n413788 , n66981 );
buf ( n413789 , n413788 );
not ( n66984 , n413789 );
and ( n66985 , n66972 , n66984 );
buf ( n413792 , n388349 );
buf ( n413793 , n411798 );
nor ( n66988 , n413792 , n413793 );
buf ( n413795 , n66988 );
buf ( n413796 , n413795 );
nor ( n66991 , n66985 , n413796 );
buf ( n413798 , n66991 );
buf ( n413799 , n413798 );
not ( n66994 , n413799 );
buf ( n413801 , n66994 );
buf ( n413802 , n413801 );
not ( n66997 , n413802 );
buf ( n413804 , n390292 );
not ( n66999 , n413804 );
or ( n67000 , n40885 , n55055 );
nand ( n67001 , n36821 , n55055 );
nand ( n67002 , n67000 , n67001 );
buf ( n413809 , n67002 );
not ( n67004 , n413809 );
and ( n67005 , n66999 , n67004 );
buf ( n413812 , n388402 );
buf ( n413813 , n411816 );
nor ( n67008 , n413812 , n413813 );
buf ( n413815 , n67008 );
buf ( n413816 , n413815 );
nor ( n67011 , n67005 , n413816 );
buf ( n413818 , n67011 );
buf ( n413819 , n413818 );
not ( n67014 , n413819 );
buf ( n413821 , n67014 );
buf ( n413822 , n413821 );
not ( n67017 , n413822 );
or ( n67018 , n66997 , n67017 );
buf ( n413825 , n413798 );
not ( n67020 , n413825 );
buf ( n413827 , n413818 );
not ( n67022 , n413827 );
or ( n67023 , n67020 , n67022 );
buf ( n413830 , n390362 );
not ( n67025 , n413830 );
buf ( n413832 , n412709 );
not ( n67027 , n413832 );
or ( n413834 , n67025 , n67027 );
buf ( n413835 , n40601 );
not ( n67030 , n413835 );
buf ( n413837 , n397072 );
not ( n67032 , n413837 );
or ( n67033 , n67030 , n67032 );
buf ( n413840 , n393557 );
buf ( n413841 , n40600 );
nand ( n67036 , n413840 , n413841 );
buf ( n413843 , n67036 );
buf ( n413844 , n413843 );
nand ( n67039 , n67033 , n413844 );
buf ( n413846 , n67039 );
buf ( n413847 , n413846 );
not ( n67042 , n40590 );
buf ( n413849 , n67042 );
nand ( n67044 , n413847 , n413849 );
buf ( n413851 , n67044 );
buf ( n413852 , n413851 );
nand ( n67047 , n413834 , n413852 );
buf ( n413854 , n67047 );
buf ( n413855 , n413854 );
xor ( n67050 , n412881 , n412941 );
xor ( n67051 , n67050 , n413472 );
buf ( n413858 , n67051 );
xor ( n67053 , n413855 , n413858 );
buf ( n413860 , n411504 );
not ( n67055 , n413860 );
buf ( n413862 , n50317 );
not ( n67057 , n413862 );
or ( n67058 , n67055 , n67057 );
buf ( n413865 , n40818 );
buf ( n413866 , n391024 );
nand ( n67061 , n413865 , n413866 );
buf ( n413868 , n67061 );
buf ( n413869 , n413868 );
nand ( n67064 , n67058 , n413869 );
buf ( n413871 , n67064 );
not ( n67066 , n413871 );
not ( n67067 , n43536 );
or ( n67068 , n67066 , n67067 );
buf ( n413875 , n412659 );
not ( n67070 , n413875 );
buf ( n413877 , n67070 );
or ( n67072 , n413877 , n43516 );
nand ( n67073 , n67068 , n67072 );
buf ( n413880 , n67073 );
and ( n67075 , n67053 , n413880 );
and ( n67076 , n413855 , n413858 );
or ( n67077 , n67075 , n67076 );
buf ( n413884 , n67077 );
buf ( n413885 , n413884 );
nand ( n67080 , n67023 , n413885 );
buf ( n413887 , n67080 );
buf ( n413888 , n413887 );
nand ( n67083 , n67018 , n413888 );
buf ( n413890 , n67083 );
buf ( n413891 , n413890 );
not ( n67086 , n413891 );
buf ( n413893 , n67086 );
buf ( n413894 , n413893 );
not ( n67089 , n413894 );
or ( n67090 , n66970 , n67089 );
buf ( n413897 , n45949 );
not ( n67092 , n413897 );
buf ( n413899 , n393369 );
not ( n67094 , n413899 );
buf ( n413901 , n44007 );
not ( n67096 , n413901 );
or ( n67097 , n67094 , n67096 );
buf ( n413904 , n385342 );
buf ( n413905 , n393381 );
nand ( n67100 , n413904 , n413905 );
buf ( n413907 , n67100 );
buf ( n413908 , n413907 );
nand ( n67103 , n67097 , n413908 );
buf ( n413910 , n67103 );
buf ( n413911 , n413910 );
not ( n67106 , n413911 );
or ( n67107 , n67092 , n67106 );
buf ( n413914 , n412823 );
buf ( n413915 , n45954 );
nand ( n67110 , n413914 , n413915 );
buf ( n413917 , n67110 );
buf ( n413918 , n413917 );
nand ( n67113 , n67107 , n413918 );
buf ( n413920 , n67113 );
buf ( n413921 , n413920 );
not ( n67116 , n36757 );
not ( n67117 , n36395 );
or ( n67118 , n67116 , n67117 );
nand ( n67119 , n67118 , n358975 );
nand ( n67120 , n40839 , n36758 );
nand ( n67121 , n67119 , n395722 , n67120 );
buf ( n413928 , n67121 );
not ( n67123 , n413928 );
buf ( n413930 , n45661 );
not ( n67125 , n413930 );
buf ( n67126 , n49116 );
buf ( n413933 , n67126 );
buf ( n413934 , n388905 );
and ( n67129 , n413933 , n413934 );
not ( n67130 , n413933 );
buf ( n413937 , n388908 );
and ( n67132 , n67130 , n413937 );
nor ( n67133 , n67129 , n67132 );
buf ( n413940 , n67133 );
buf ( n413941 , n413940 );
not ( n67136 , n413941 );
and ( n67137 , n67125 , n67136 );
buf ( n413944 , n65807 );
not ( n67139 , n413944 );
buf ( n413946 , n37313 );
nor ( n67141 , n67139 , n413946 );
buf ( n413948 , n67141 );
buf ( n413949 , n413948 );
nor ( n67144 , n67137 , n413949 );
buf ( n413951 , n67144 );
buf ( n413952 , n413951 );
not ( n67147 , n413952 );
or ( n67148 , n67123 , n67147 );
not ( n67149 , n389119 );
buf ( n413956 , n391446 );
not ( n67151 , n413956 );
buf ( n413958 , n399164 );
not ( n67153 , n413958 );
or ( n67154 , n67151 , n67153 );
buf ( n413961 , n24049 );
buf ( n413962 , n391443 );
nand ( n67157 , n413961 , n413962 );
buf ( n413964 , n67157 );
buf ( n413965 , n413964 );
nand ( n67160 , n67154 , n413965 );
buf ( n413967 , n67160 );
buf ( n413968 , n413967 );
not ( n67163 , n413968 );
buf ( n413970 , n67163 );
not ( n67165 , n413970 );
and ( n67166 , n67149 , n67165 );
and ( n67167 , n412733 , n46921 );
nor ( n67168 , n67166 , n67167 );
buf ( n413975 , n67168 );
not ( n67170 , n413975 );
buf ( n413977 , n40592 );
not ( n67172 , n413977 );
buf ( n413979 , n40601 );
not ( n67174 , n413979 );
buf ( n413981 , n52763 );
not ( n67176 , n413981 );
or ( n67177 , n67174 , n67176 );
buf ( n413984 , n388643 );
buf ( n413985 , n40600 );
nand ( n67180 , n413984 , n413985 );
buf ( n413987 , n67180 );
buf ( n413988 , n413987 );
nand ( n67183 , n67177 , n413988 );
buf ( n413990 , n67183 );
buf ( n413991 , n413990 );
not ( n67186 , n413991 );
or ( n67187 , n67172 , n67186 );
buf ( n413994 , n413846 );
buf ( n413995 , n390362 );
nand ( n67190 , n413994 , n413995 );
buf ( n413997 , n67190 );
buf ( n413998 , n413997 );
nand ( n67193 , n67187 , n413998 );
buf ( n414000 , n67193 );
not ( n67195 , n414000 );
buf ( n414002 , n67195 );
not ( n67197 , n414002 );
or ( n67198 , n67170 , n67197 );
xor ( n67199 , n413433 , n413446 );
xor ( n67200 , n67199 , n413468 );
buf ( n414007 , n67200 );
buf ( n414008 , n414007 );
not ( n67203 , n414008 );
buf ( n414010 , n67203 );
buf ( n414011 , n414010 );
nand ( n67206 , n67198 , n414011 );
buf ( n414013 , n67206 );
buf ( n414014 , n414013 );
buf ( n414015 , n67168 );
not ( n67210 , n414015 );
buf ( n414017 , n414000 );
nand ( n67212 , n67210 , n414017 );
buf ( n414019 , n67212 );
buf ( n414020 , n414019 );
nand ( n67215 , n414014 , n414020 );
buf ( n414022 , n67215 );
buf ( n414023 , n414022 );
nand ( n67218 , n67148 , n414023 );
buf ( n414025 , n67218 );
buf ( n414026 , n414025 );
buf ( n414027 , n413951 );
not ( n67222 , n414027 );
buf ( n414029 , n67121 );
not ( n67224 , n414029 );
buf ( n414031 , n67224 );
buf ( n414032 , n414031 );
nand ( n67227 , n67222 , n414032 );
buf ( n414034 , n67227 );
buf ( n414035 , n414034 );
nand ( n67230 , n414026 , n414035 );
buf ( n414037 , n67230 );
buf ( n414038 , n414037 );
xor ( n67233 , n413921 , n414038 );
xor ( n67234 , n412694 , n412720 );
xor ( n67235 , n67234 , n412800 );
buf ( n414042 , n67235 );
buf ( n414043 , n414042 );
and ( n67238 , n67233 , n414043 );
and ( n67239 , n413921 , n414038 );
or ( n67240 , n67238 , n67239 );
buf ( n414047 , n67240 );
buf ( n414048 , n414047 );
nand ( n67243 , n67090 , n414048 );
buf ( n414050 , n67243 );
buf ( n414051 , n414050 );
buf ( n414052 , n413890 );
buf ( n414053 , n66965 );
nand ( n67248 , n414052 , n414053 );
buf ( n414055 , n67248 );
buf ( n414056 , n414055 );
nand ( n67251 , n414051 , n414056 );
buf ( n414058 , n67251 );
and ( n67253 , n413765 , n414058 );
nor ( n67254 , n66955 , n67253 );
buf ( n414061 , n67254 );
not ( n67256 , n414061 );
buf ( n414063 , n67256 );
not ( n67258 , n414063 );
or ( n67259 , n66786 , n67258 );
buf ( n414066 , n413610 );
not ( n67261 , n414066 );
buf ( n414068 , n67261 );
buf ( n414069 , n414068 );
not ( n67264 , n414069 );
buf ( n414071 , n67254 );
not ( n67266 , n414071 );
or ( n67267 , n67264 , n67266 );
buf ( n414074 , C0 );
buf ( n67283 , n64692 );
not ( n67284 , n64737 );
not ( n67285 , n64670 );
or ( n67286 , n67284 , n67285 );
or ( n67287 , n64670 , n64737 );
nand ( n67288 , n67286 , n67287 );
xor ( n67289 , n67283 , n67288 );
nand ( n67290 , n61577 , n412145 );
buf ( n414083 , n408347 );
not ( n67292 , n414083 );
buf ( n414085 , n384239 );
not ( n67294 , n414085 );
or ( n67295 , n67292 , n67294 );
buf ( n414088 , n389692 );
buf ( n414089 , n408344 );
nand ( n67298 , n414088 , n414089 );
buf ( n414091 , n67298 );
buf ( n414092 , n414091 );
nand ( n67301 , n67295 , n414092 );
buf ( n414094 , n67301 );
buf ( n414095 , n414094 );
buf ( n414096 , n50579 );
nand ( n67305 , n414095 , n414096 );
buf ( n414098 , n67305 );
nand ( n67307 , n67289 , n67290 , n414098 );
not ( n67308 , n67307 );
not ( n67309 , n45260 );
not ( n67310 , n413656 );
or ( n67311 , n67309 , n67310 );
nand ( n67312 , n412192 , n392740 );
nand ( n67313 , n67311 , n67312 );
not ( n67314 , n67313 );
xor ( n67315 , n411725 , n411772 );
buf ( n414108 , n67315 );
buf ( n414109 , n64826 );
xnor ( n67318 , n414108 , n414109 );
buf ( n414111 , n67318 );
not ( n67320 , n414111 );
not ( n67321 , n67320 );
or ( n67322 , n67314 , n67321 );
buf ( n414115 , n67313 );
not ( n67324 , n414115 );
buf ( n414117 , n67324 );
not ( n67326 , n414117 );
not ( n67327 , n414111 );
or ( n67328 , n67326 , n67327 );
xor ( n67329 , n411737 , n411754 );
xor ( n67330 , n67329 , n411768 );
buf ( n414123 , n67330 );
buf ( n414124 , n414123 );
not ( n67333 , n414124 );
buf ( n414126 , n67333 );
buf ( n414127 , n414126 );
not ( n67336 , n414127 );
not ( n67337 , n41447 );
not ( n67338 , n412681 );
or ( n67339 , n67337 , n67338 );
not ( n67340 , n394210 );
not ( n67341 , n393525 );
or ( n67342 , n67340 , n67341 );
nand ( n67343 , n394219 , n388962 );
nand ( n67344 , n67342 , n67343 );
nand ( n67345 , n393544 , n67344 );
nand ( n67346 , n67339 , n67345 );
buf ( n414139 , n67346 );
not ( n67348 , n414139 );
buf ( n414141 , n67348 );
buf ( n414142 , n414141 );
not ( n67351 , n414142 );
or ( n67352 , n67336 , n67351 );
buf ( n414145 , n388809 );
not ( n67354 , n414145 );
buf ( n414147 , n412787 );
not ( n67356 , n414147 );
or ( n67357 , n67354 , n67356 );
and ( n67358 , n27258 , n388754 );
not ( n67359 , n27258 );
and ( n67360 , n67359 , n405736 );
or ( n67361 , n67358 , n67360 );
buf ( n414154 , n67361 );
buf ( n414155 , n388746 );
nand ( n67364 , n414154 , n414155 );
buf ( n414157 , n67364 );
buf ( n414158 , n414157 );
nand ( n67367 , n67357 , n414158 );
buf ( n414160 , n67367 );
buf ( n414161 , n414160 );
not ( n67370 , n414161 );
buf ( n414163 , n67370 );
not ( n67372 , n414163 );
xor ( n67373 , n412889 , n412913 );
xor ( n67374 , n67373 , n412937 );
buf ( n414167 , n67374 );
not ( n67376 , n414167 );
or ( n67377 , n67372 , n67376 );
buf ( n414170 , n42066 );
not ( n67379 , n414170 );
buf ( n414172 , n404601 );
not ( n67381 , n414172 );
or ( n67382 , n67379 , n67381 );
buf ( n414175 , n407928 );
buf ( n414176 , n42065 );
nand ( n67385 , n414175 , n414176 );
buf ( n414178 , n67385 );
buf ( n414179 , n414178 );
nand ( n67388 , n67382 , n414179 );
buf ( n414181 , n67388 );
buf ( n414182 , n414181 );
not ( n67391 , n414182 );
buf ( n414184 , n409082 );
not ( n67393 , n414184 );
or ( n67394 , n67391 , n67393 );
buf ( n414187 , n66072 );
buf ( n414188 , n394134 );
nand ( n67397 , n414187 , n414188 );
buf ( n414190 , n67397 );
buf ( n414191 , n414190 );
nand ( n67400 , n67394 , n414191 );
buf ( n414193 , n67400 );
not ( n67402 , n414193 );
not ( n67403 , n389162 );
not ( n67404 , n66617 );
or ( n67405 , n67403 , n67404 );
not ( n67406 , n64268 );
not ( n67407 , n388227 );
or ( n67408 , n67406 , n67407 );
buf ( n414201 , n27234 );
buf ( n414202 , n64273 );
nand ( n67411 , n414201 , n414202 );
buf ( n414204 , n67411 );
nand ( n67413 , n67408 , n414204 );
buf ( n414206 , n67413 );
buf ( n414207 , n45076 );
nand ( n67416 , n414206 , n414207 );
buf ( n414209 , n67416 );
nand ( n67418 , n67405 , n414209 );
not ( n67419 , n67418 );
or ( n67420 , n67402 , n67419 );
or ( n67421 , n414193 , n67418 );
xor ( n67422 , n66597 , n66125 );
xnor ( n67423 , n67422 , n412980 );
nand ( n67424 , n67421 , n67423 );
nand ( n67425 , n67420 , n67424 );
nand ( n67426 , n67377 , n67425 );
buf ( n414219 , n67426 );
buf ( n414220 , n414167 );
not ( n67429 , n414220 );
buf ( n414222 , n414160 );
nand ( n67431 , n67429 , n414222 );
buf ( n414224 , n67431 );
buf ( n414225 , n414224 );
nand ( n67434 , n414219 , n414225 );
buf ( n414227 , n67434 );
buf ( n414228 , n414227 );
nand ( n67437 , n67352 , n414228 );
buf ( n414230 , n67437 );
buf ( n414231 , n414230 );
buf ( n414232 , n67346 );
buf ( n414233 , n414123 );
nand ( n67442 , n414232 , n414233 );
buf ( n414235 , n67442 );
buf ( n414236 , n414235 );
nand ( n67445 , n414231 , n414236 );
buf ( n414238 , n67445 );
nand ( n67447 , n67328 , n414238 );
nand ( n67448 , n67322 , n67447 );
not ( n67449 , n67448 );
or ( n67450 , n67308 , n67449 );
not ( n67451 , n67289 );
nand ( n67452 , n67290 , n414098 );
nand ( n67453 , n67451 , n67452 );
nand ( n67454 , n67450 , n67453 );
xor ( n67455 , n414074 , n67454 );
xor ( n67456 , n411982 , n411957 );
xor ( n67457 , n67456 , n411990 );
and ( n67458 , n67455 , n67457 );
or ( n67460 , n67458 , C0 );
buf ( n414252 , n67460 );
nand ( n67462 , n67267 , n414252 );
buf ( n414254 , n67462 );
nand ( n67464 , n67259 , n414254 );
not ( n67465 , n67464 );
or ( n67466 , n66782 , n67465 );
xor ( n67467 , n65479 , n65448 );
xor ( n67468 , n67467 , n65457 );
not ( n67469 , n67468 );
xor ( n67470 , n412835 , n66019 );
xor ( n67471 , n67470 , n413525 );
not ( n67472 , n67471 );
xor ( n67473 , n65300 , n412152 );
xor ( n67474 , n67473 , n65352 );
not ( n67475 , n67474 );
not ( n67476 , n412270 );
xor ( n67477 , n412265 , n67476 );
xor ( n67478 , n67477 , C0 );
nand ( n67479 , n67475 , n67478 );
not ( n67480 , n67479 );
or ( n67481 , n67472 , n67480 );
not ( n67482 , n67478 );
nand ( n67483 , n67482 , n67474 );
nand ( n67484 , n67481 , n67483 );
not ( n67485 , n67484 );
not ( n67486 , n67485 );
and ( n67487 , n67469 , n67486 );
nand ( n67488 , n67468 , n67485 );
xor ( n67489 , n412669 , n412805 );
xor ( n67490 , n67489 , n412831 );
buf ( n414282 , n67490 );
buf ( n414283 , n414282 );
buf ( n414284 , n412199 );
buf ( n414285 , n65342 );
xor ( n67495 , n414284 , n414285 );
buf ( n414287 , n65346 );
xnor ( n67497 , n67495 , n414287 );
buf ( n414289 , n67497 );
buf ( n414290 , n414289 );
xor ( n67500 , n414283 , n414290 );
xor ( n67501 , n412870 , n412877 );
xor ( n67502 , n67501 , n413521 );
buf ( n414294 , n67502 );
buf ( n414295 , n414294 );
and ( n67505 , n67500 , n414295 );
and ( n67506 , n414283 , n414290 );
or ( n67507 , n67505 , n67506 );
buf ( n414299 , n67507 );
buf ( n414300 , n414299 );
xor ( n67535 , n67448 , n67452 );
xor ( n67536 , n67535 , n67289 );
not ( n67540 , n67536 );
or ( n67541 , C0 , n67540 );
buf ( n414305 , C0 );
buf ( n414306 , n414305 );
xor ( n67563 , n414238 , n414117 );
xnor ( n67564 , n67563 , n67320 );
buf ( n414309 , n67564 );
xor ( n67566 , n414306 , n414309 );
buf ( n414311 , n50579 );
not ( n67568 , n414311 );
buf ( n414313 , n408347 );
not ( n67570 , n414313 );
buf ( n414315 , n384280 );
not ( n67572 , n414315 );
or ( n67573 , n67570 , n67572 );
buf ( n414318 , n384974 );
buf ( n414319 , n50584 );
nand ( n67576 , n414318 , n414319 );
buf ( n414321 , n67576 );
buf ( n414322 , n414321 );
nand ( n67579 , n67573 , n414322 );
buf ( n414324 , n67579 );
buf ( n414325 , n414324 );
not ( n67582 , n414325 );
or ( n67583 , n67568 , n67582 );
buf ( n414328 , n414094 );
buf ( n414329 , n51553 );
nand ( n67586 , n414328 , n414329 );
buf ( n414331 , n67586 );
buf ( n414332 , n414331 );
nand ( n67589 , n67583 , n414332 );
buf ( n414334 , n67589 );
buf ( n414335 , n414334 );
and ( n67592 , n67566 , n414335 );
or ( n67594 , n67592 , C0 );
buf ( n414338 , n67594 );
nand ( n67596 , n67541 , n414338 );
nand ( n67597 , C1 , n67596 );
buf ( n414341 , n67597 );
xor ( n67599 , n414300 , n414341 );
xor ( n67600 , n414074 , n67454 );
xor ( n67601 , n67600 , n67457 );
buf ( n414345 , n67601 );
and ( n67603 , n67599 , n414345 );
and ( n67604 , n414300 , n414341 );
or ( n67605 , n67603 , n67604 );
buf ( n414349 , n67605 );
and ( n67607 , n67488 , n414349 );
nor ( n67608 , n67487 , n67607 );
nor ( n67609 , n413606 , n67464 );
or ( n67610 , n67608 , n67609 );
nand ( n67611 , n67466 , n67610 );
buf ( n67612 , n67611 );
nand ( n67613 , n66778 , n67612 );
nand ( n67614 , n66768 , n413598 );
nand ( n67615 , n67613 , n67614 );
nand ( n67616 , n412627 , n67615 );
not ( n67617 , n67616 );
nand ( n67618 , n65675 , n65580 );
nand ( n67619 , n67617 , n67618 );
nand ( n67620 , n65764 , n65799 , n67619 );
not ( n67621 , n412587 );
nand ( n67622 , n67621 , n412581 );
not ( n67623 , n67622 );
buf ( n414367 , n412612 );
buf ( n414368 , n412620 );
nand ( n67626 , n414367 , n414368 );
buf ( n414370 , n67626 );
not ( n67628 , n414370 );
or ( n67629 , n67623 , n67628 );
nand ( n67630 , n67629 , n65799 );
buf ( n414374 , n408590 );
buf ( n414375 , n62965 );
xor ( n67633 , n414374 , n414375 );
buf ( n414377 , n408567 );
xnor ( n67635 , n67633 , n414377 );
buf ( n414379 , n67635 );
xor ( n67637 , n412600 , n412606 );
and ( n67638 , n67637 , n412610 );
and ( n67639 , n412600 , n412606 );
or ( n67640 , n67638 , n67639 );
buf ( n414384 , n67640 );
nand ( n67642 , n414379 , n414384 );
nand ( n67643 , n67620 , n67630 , n67642 );
buf ( n414387 , n413598 );
not ( n67645 , n414387 );
not ( n67646 , n66767 );
not ( n67647 , n67611 );
or ( n67648 , n67646 , n67647 );
or ( n67649 , n67611 , n66767 );
nand ( n67650 , n67648 , n67649 );
buf ( n414394 , n67650 );
not ( n67652 , n414394 );
and ( n67653 , n67645 , n67652 );
buf ( n414397 , n413598 );
buf ( n414398 , n67650 );
and ( n67656 , n414397 , n414398 );
nor ( n67657 , n67653 , n67656 );
buf ( n414401 , n67657 );
buf ( n414402 , n413562 );
not ( n67660 , n414402 );
buf ( n414404 , n413585 );
not ( n67662 , n414404 );
or ( n67663 , n67660 , n67662 );
buf ( n414407 , n413562 );
not ( n67665 , n414407 );
buf ( n414409 , n413582 );
nand ( n67667 , n67665 , n414409 );
buf ( n414411 , n67667 );
buf ( n414412 , n414411 );
nand ( n67670 , n67663 , n414412 );
buf ( n414414 , n67670 );
buf ( n414415 , n414414 );
buf ( n414416 , n413569 );
and ( n67674 , n414415 , n414416 );
not ( n67675 , n414415 );
buf ( n414419 , n413566 );
and ( n67677 , n67675 , n414419 );
nor ( n67678 , n67674 , n67677 );
buf ( n414422 , n67678 );
buf ( n414423 , n414422 );
buf ( n414424 , n66703 );
buf ( n414425 , n413534 );
xor ( n67683 , n414424 , n414425 );
buf ( n414427 , n413553 );
xnor ( n67685 , n67683 , n414427 );
buf ( n414429 , n67685 );
buf ( n414430 , n414429 );
buf ( n414431 , n67460 );
buf ( n414432 , n413610 );
xor ( n67690 , n414431 , n414432 );
buf ( n414434 , n414063 );
xnor ( n67692 , n67690 , n414434 );
buf ( n414436 , n67692 );
buf ( n414437 , n414436 );
xor ( n67695 , n414430 , n414437 );
xor ( n67696 , n414283 , n414290 );
xor ( n67697 , n67696 , n414295 );
buf ( n414441 , n67697 );
buf ( n414442 , n414441 );
xor ( n67700 , n413615 , n413679 );
xor ( n67701 , n67700 , n413717 );
buf ( n414445 , n67701 );
not ( n67703 , n414445 );
buf ( n414447 , C1 );
nand ( n67724 , n67703 , n414447 );
not ( n67725 , n67724 );
xor ( n67726 , n413855 , n413858 );
xor ( n67727 , n67726 , n413880 );
buf ( n414452 , n67727 );
buf ( n414453 , n414452 );
xor ( n67730 , n414031 , n414022 );
xnor ( n67731 , n67730 , n413951 );
buf ( n414456 , n67731 );
xor ( n67733 , n414453 , n414456 );
buf ( n414458 , n399274 );
not ( n67735 , n414458 );
buf ( n414460 , n391764 );
not ( n67737 , n414460 );
or ( n67738 , n67735 , n67737 );
buf ( n414463 , n388263 );
buf ( n414464 , n399283 );
nand ( n67741 , n414463 , n414464 );
buf ( n414466 , n67741 );
buf ( n414467 , n414466 );
nand ( n67744 , n67738 , n414467 );
buf ( n414469 , n67744 );
buf ( n414470 , n414469 );
not ( n67747 , n414470 );
buf ( n414472 , n383894 );
not ( n67749 , n414472 );
or ( n67750 , n67747 , n67749 );
buf ( n414475 , n413627 );
buf ( n414476 , n383907 );
nand ( n67753 , n414475 , n414476 );
buf ( n414478 , n67753 );
buf ( n414479 , n414478 );
nand ( n67756 , n67750 , n414479 );
buf ( n414481 , n67756 );
not ( n67758 , n414481 );
buf ( n414483 , n392884 );
not ( n67760 , n414483 );
buf ( n414485 , n46906 );
not ( n67762 , n414485 );
or ( n67763 , n67760 , n67762 );
buf ( n414488 , n49660 );
buf ( n414489 , n392887 );
nand ( n67766 , n414488 , n414489 );
buf ( n414491 , n67766 );
buf ( n414492 , n414491 );
nand ( n67769 , n67763 , n414492 );
buf ( n414494 , n67769 );
buf ( n414495 , n414494 );
not ( n67772 , n414495 );
buf ( n414497 , n411271 );
not ( n67774 , n414497 );
or ( n67775 , n67772 , n67774 );
buf ( n414500 , n412758 );
buf ( n414501 , n395469 );
nand ( n67778 , n414500 , n414501 );
buf ( n414503 , n67778 );
buf ( n414504 , n414503 );
nand ( n67781 , n67775 , n414504 );
buf ( n414506 , n67781 );
buf ( n414507 , n389341 );
not ( n67784 , n414507 );
buf ( n414509 , n24071 );
not ( n67786 , n414509 );
or ( n67787 , n67784 , n67786 );
buf ( n414512 , n51821 );
buf ( n414513 , n393185 );
nand ( n67790 , n414512 , n414513 );
buf ( n414515 , n67790 );
buf ( n414516 , n414515 );
nand ( n67793 , n67787 , n414516 );
buf ( n414518 , n67793 );
not ( n67795 , n414518 );
not ( n67796 , n52812 );
or ( n67797 , n67795 , n67796 );
buf ( n414522 , n413459 );
buf ( n414523 , n42924 );
nand ( n67800 , n414522 , n414523 );
buf ( n414525 , n67800 );
nand ( n67802 , n67797 , n414525 );
not ( n67803 , n67802 );
buf ( n414528 , n388809 );
not ( n67805 , n414528 );
buf ( n414530 , n67361 );
not ( n67807 , n414530 );
or ( n67808 , n67805 , n67807 );
xor ( n67809 , n405736 , n28644 );
buf ( n414534 , n67809 );
buf ( n414535 , n388746 );
nand ( n67812 , n414534 , n414535 );
buf ( n414537 , n67812 );
buf ( n414538 , n414537 );
nand ( n67815 , n67808 , n414538 );
buf ( n414540 , n67815 );
buf ( n414541 , n414540 );
not ( n67818 , n414541 );
buf ( n414543 , n67818 );
nand ( n67820 , n67803 , n414543 );
not ( n67821 , n67820 );
not ( n67822 , n45076 );
and ( n67823 , n12480 , n64273 );
not ( n67824 , n12480 );
and ( n67825 , n67824 , n64268 );
or ( n67826 , n67823 , n67825 );
not ( n67827 , n67826 );
or ( n67828 , n67822 , n67827 );
nand ( n67829 , n67413 , n41664 );
nand ( n67830 , n67828 , n67829 );
not ( n67831 , n66128 );
buf ( n67832 , n23841 );
not ( n67833 , n67832 );
not ( n67834 , n412892 );
or ( n67835 , n67833 , n67834 );
nand ( n67836 , n410407 , n27320 );
nand ( n67837 , n67835 , n67836 );
not ( n67838 , n67837 );
or ( n67839 , n67831 , n67838 );
nand ( n67840 , n412970 , n412976 );
nand ( n67841 , n67839 , n67840 );
or ( n67842 , n67830 , n67841 );
buf ( n414567 , n67842 );
xor ( n67844 , n66333 , n66346 );
xnor ( n67845 , n67844 , n66592 );
buf ( n414570 , n67845 );
and ( n67847 , n414567 , n414570 );
and ( n67848 , n67830 , n67841 );
buf ( n414573 , n67848 );
nor ( n67850 , n67847 , n414573 );
buf ( n414575 , n67850 );
buf ( n414576 , n414575 );
not ( n67853 , n414576 );
buf ( n414578 , n67853 );
not ( n67855 , n414578 );
or ( n67856 , n67821 , n67855 );
buf ( n414581 , n414540 );
buf ( n414582 , n67802 );
nand ( n67859 , n414581 , n414582 );
buf ( n414584 , n67859 );
nand ( n67861 , n67856 , n414584 );
xor ( n67862 , n414506 , n67861 );
buf ( n414587 , n394817 );
not ( n67864 , n414587 );
buf ( n414589 , n388965 );
not ( n67866 , n414589 );
or ( n67867 , n67864 , n67866 );
buf ( n414592 , n385473 );
buf ( n414593 , n394814 );
nand ( n67870 , n414592 , n414593 );
buf ( n414595 , n67870 );
buf ( n414596 , n414595 );
nand ( n67873 , n67867 , n414596 );
buf ( n414598 , n67873 );
buf ( n414599 , n414598 );
not ( n67876 , n414599 );
buf ( n414601 , n393544 );
not ( n67878 , n414601 );
or ( n67879 , n67876 , n67878 );
buf ( n414604 , n67344 );
buf ( n414605 , n51692 );
nand ( n67882 , n414604 , n414605 );
buf ( n414607 , n67882 );
buf ( n414608 , n414607 );
nand ( n67885 , n67879 , n414608 );
buf ( n414610 , n67885 );
buf ( n414611 , n414610 );
not ( n67888 , n414611 );
buf ( n414613 , n67888 );
xor ( n67890 , n67862 , n414613 );
nand ( n67891 , n67758 , n67890 );
not ( n67892 , n67891 );
and ( n67893 , n51821 , n391443 );
not ( n67894 , n51821 );
and ( n67895 , n67894 , n391446 );
or ( n67896 , n67893 , n67895 );
buf ( n414621 , n67896 );
not ( n67898 , n414621 );
buf ( n414623 , n52812 );
not ( n67900 , n414623 );
or ( n67901 , n67898 , n67900 );
buf ( n414626 , n42923 );
not ( n67903 , n414626 );
buf ( n414628 , n414518 );
nand ( n67905 , n67903 , n414628 );
buf ( n414630 , n67905 );
buf ( n414631 , n414630 );
nand ( n67908 , n67901 , n414631 );
buf ( n414633 , n67908 );
buf ( n414634 , n414633 );
not ( n67911 , n414634 );
buf ( n414636 , n67911 );
not ( n67913 , n414636 );
xor ( n67914 , n67845 , n67841 );
xor ( n67915 , n67914 , n67830 );
not ( n67916 , n67915 );
not ( n67917 , n67916 );
or ( n67918 , n67913 , n67917 );
not ( n67919 , n41373 );
not ( n67920 , n66132 );
not ( n67921 , n42066 );
or ( n67922 , n67920 , n67921 );
buf ( n414647 , n41365 );
buf ( n414648 , n42065 );
nand ( n67925 , n414647 , n414648 );
buf ( n414650 , n67925 );
nand ( n67927 , n67922 , n414650 );
not ( n67928 , n67927 );
or ( n67929 , n67919 , n67928 );
nand ( n67930 , n412976 , n67837 );
nand ( n67931 , n67929 , n67930 );
xor ( n67932 , n413182 , n413254 );
xor ( n67933 , n67932 , n413316 );
buf ( n414658 , n59435 );
buf ( n414659 , n405391 );
and ( n67936 , n414658 , n414659 );
buf ( n414661 , n406565 );
buf ( n414662 , n405391 );
not ( n67939 , n414662 );
buf ( n414664 , n67939 );
buf ( n414665 , n414664 );
and ( n67942 , n414661 , n414665 );
nor ( n67943 , n67936 , n67942 );
buf ( n414668 , n67943 );
buf ( n414669 , n414668 );
buf ( n414670 , n405407 );
or ( n67947 , n414669 , n414670 );
buf ( n414672 , n413280 );
buf ( n414673 , n405384 );
or ( n67950 , n414672 , n414673 );
nand ( n67951 , n67947 , n67950 );
buf ( n414676 , n67951 );
buf ( n414677 , n414676 );
buf ( n414678 , n401695 );
buf ( n414679 , n66270 );
and ( n67956 , n414678 , n414679 );
not ( n67957 , n414678 );
buf ( n414682 , n413098 );
and ( n67959 , n67957 , n414682 );
nor ( n67960 , n67956 , n67959 );
buf ( n414685 , n67960 );
buf ( n414686 , n414685 );
not ( n67963 , n414686 );
buf ( n414688 , n67963 );
buf ( n414689 , n414688 );
buf ( n414690 , n403158 );
or ( n67967 , n414689 , n414690 );
buf ( n414692 , n413204 );
buf ( n414693 , n403167 );
or ( n67970 , n414692 , n414693 );
nand ( n67971 , n67967 , n67970 );
buf ( n414696 , n67971 );
buf ( n414697 , n414696 );
not ( n67974 , n54229 );
not ( n67975 , n67974 );
not ( n67976 , n54068 );
nand ( n67977 , n67976 , n54226 );
not ( n67978 , n67977 );
or ( n67979 , n67975 , n67978 );
nand ( n67980 , n54231 , n54034 );
nand ( n67981 , n67979 , n67980 );
not ( n67982 , n67976 );
not ( n67983 , n54226 );
or ( n67984 , n67982 , n67983 );
nor ( n67985 , n54229 , n67980 );
nand ( n67986 , n67984 , n67985 );
nand ( n67987 , n67981 , n67986 );
buf ( n414712 , n67987 );
not ( n67989 , n414712 );
buf ( n414714 , n67989 );
buf ( n414715 , n414714 );
buf ( n414716 , n403083 );
or ( n67993 , n414715 , n414716 );
buf ( n414718 , n413187 );
buf ( n414719 , n403092 );
or ( n67996 , n414718 , n414719 );
nand ( n67997 , n67993 , n67996 );
buf ( n414722 , n67997 );
buf ( n414723 , n414722 );
xor ( n68000 , n414697 , n414723 );
nand ( n68001 , n67976 , n67974 );
xnor ( n68002 , n54226 , n68001 );
buf ( n414727 , n68002 );
not ( n68004 , n414727 );
buf ( n414729 , n68004 );
buf ( n414730 , n414729 );
buf ( n414731 , n401623 );
or ( n68008 , n414730 , n414731 );
buf ( n414733 , n403092 );
buf ( n414734 , n414714 );
or ( n68011 , n414733 , n414734 );
nand ( n68012 , n68008 , n68011 );
buf ( n414737 , n68012 );
buf ( n414738 , n414737 );
buf ( n414739 , n403164 );
not ( n68016 , n414739 );
buf ( n414741 , n414685 );
not ( n68018 , n414741 );
or ( n68019 , n68016 , n68018 );
buf ( n414744 , n401695 );
buf ( n414745 , n413187 );
and ( n68022 , n414744 , n414745 );
not ( n68023 , n414744 );
buf ( n414748 , n66359 );
and ( n68025 , n68023 , n414748 );
nor ( n68026 , n68022 , n68025 );
buf ( n414751 , n68026 );
buf ( n414752 , n414751 );
buf ( n414753 , n403158 );
or ( n68030 , n414752 , n414753 );
nand ( n68031 , n68019 , n68030 );
buf ( n414756 , n68031 );
buf ( n414757 , n414756 );
and ( n68034 , n414738 , n414757 );
buf ( n414759 , n68034 );
buf ( n414760 , n414759 );
and ( n68037 , n68000 , n414760 );
and ( n68038 , n414697 , n414723 );
or ( n68039 , n68037 , n68038 );
buf ( n414764 , n68039 );
buf ( n414765 , n414764 );
xor ( n68042 , n414677 , n414765 );
not ( n68043 , n409504 );
not ( n68044 , n68043 );
not ( n68045 , n413263 );
not ( n68046 , n68045 );
or ( n68047 , n68044 , n68046 );
and ( n68048 , n403079 , n63629 );
and ( n68049 , n63625 , n55846 );
nor ( n68050 , n68048 , n68049 );
not ( n68051 , n68050 );
nand ( n68052 , n68051 , n409507 );
nand ( n68053 , n68047 , n68052 );
buf ( n414778 , n68053 );
and ( n68055 , n68042 , n414778 );
and ( n68056 , n414677 , n414765 );
or ( n68057 , n68055 , n68056 );
buf ( n414782 , n68057 );
buf ( n414783 , n414782 );
xor ( n414784 , n413216 , n413233 );
xor ( n68061 , n414784 , n413250 );
buf ( n414786 , n68061 );
buf ( n414787 , n414786 );
xor ( n68064 , n414783 , n414787 );
buf ( n414789 , n58178 );
buf ( n414790 , n62177 );
and ( n68067 , n414789 , n414790 );
buf ( n414792 , n405335 );
buf ( n414793 , n62159 );
and ( n68070 , n414792 , n414793 );
nor ( n68071 , n68067 , n68070 );
buf ( n414796 , n68071 );
buf ( n414797 , n414796 );
buf ( n414798 , n409429 );
or ( n68075 , n414797 , n414798 );
buf ( n414800 , n413342 );
buf ( n414801 , n409170 );
or ( n68078 , n414800 , n414801 );
nand ( n68079 , n68075 , n68078 );
buf ( n414804 , n68079 );
buf ( n414805 , n414804 );
buf ( n414806 , n54297 );
buf ( n414807 , n66411 );
and ( n68084 , n414806 , n414807 );
buf ( n414809 , n55919 );
buf ( n414810 , n62496 );
and ( n68087 , n414809 , n414810 );
nor ( n68088 , n68084 , n68087 );
buf ( n414813 , n68088 );
buf ( n414814 , n414813 );
buf ( n414815 , n410724 );
or ( n68092 , n414814 , n414815 );
buf ( n414817 , n413243 );
buf ( n414818 , n410721 );
or ( n68095 , n414817 , n414818 );
nand ( n68096 , n68092 , n68095 );
buf ( n414821 , n68096 );
buf ( n414822 , n414821 );
xor ( n68099 , n414805 , n414822 );
buf ( n414824 , n62278 );
buf ( n414825 , n405215 );
and ( n68102 , n414824 , n414825 );
buf ( n414827 , n409474 );
buf ( n414828 , n58061 );
and ( n68105 , n414827 , n414828 );
nor ( n68106 , n68102 , n68105 );
buf ( n414831 , n68106 );
buf ( n414832 , n414831 );
buf ( n414833 , n403293 );
or ( n68110 , n414832 , n414833 );
buf ( n414835 , n413359 );
buf ( n414836 , n405476 );
or ( n68113 , n414835 , n414836 );
nand ( n68114 , n68110 , n68113 );
buf ( n414839 , n68114 );
buf ( n414840 , n414839 );
buf ( n414841 , n63564 );
buf ( n414842 , n55905 );
and ( n68119 , n414841 , n414842 );
buf ( n414844 , n413073 );
buf ( n414845 , n55895 );
and ( n68122 , n414844 , n414845 );
nor ( n68123 , n68119 , n68122 );
buf ( n414848 , n68123 );
buf ( n414849 , n414848 );
buf ( n414850 , n403120 );
or ( n68127 , n414849 , n414850 );
buf ( n414852 , n413375 );
buf ( n414853 , n403133 );
or ( n68130 , n414852 , n414853 );
nand ( n68131 , n68127 , n68130 );
buf ( n414856 , n68131 );
buf ( n414857 , n414856 );
xor ( n68134 , n414840 , n414857 );
buf ( n414859 , n405381 );
not ( n68136 , n414859 );
buf ( n414861 , n414668 );
not ( n68138 , n414861 );
buf ( n414863 , n68138 );
buf ( n414864 , n414863 );
not ( n68141 , n414864 );
or ( n68142 , n68136 , n68141 );
buf ( n414867 , n409146 );
buf ( n414868 , n414664 );
or ( n68145 , n414867 , n414868 );
buf ( n414870 , n59596 );
buf ( n414871 , n405391 );
or ( n68148 , n414870 , n414871 );
nand ( n68149 , n68145 , n68148 );
buf ( n414874 , n68149 );
buf ( n414875 , n414874 );
not ( n68152 , n414875 );
buf ( n414877 , n68152 );
buf ( n414878 , n414877 );
buf ( n414879 , n405407 );
or ( n68156 , n414878 , n414879 );
nand ( n68157 , n68142 , n68156 );
buf ( n414882 , n68157 );
buf ( n414883 , n414882 );
and ( n68160 , n68134 , n414883 );
and ( n68161 , n414840 , n414857 );
or ( n68162 , n68160 , n68161 );
buf ( n414887 , n68162 );
buf ( n414888 , n414887 );
and ( n68165 , n68099 , n414888 );
and ( n68166 , n414805 , n414822 );
or ( n68167 , n68165 , n68166 );
buf ( n414892 , n68167 );
buf ( n414893 , n414892 );
and ( n68170 , n68064 , n414893 );
and ( n68171 , n414783 , n414787 );
or ( n68172 , n68170 , n68171 );
buf ( n414897 , n68172 );
xor ( n68174 , n413000 , n413006 );
xor ( n68175 , n68174 , n413023 );
xor ( n68176 , n66567 , n413398 );
xor ( n68177 , n68175 , n68176 );
xor ( n68178 , n414897 , n68177 );
xor ( n68179 , n67933 , n68178 );
not ( n68180 , n68179 );
and ( n68181 , n406571 , n59457 );
and ( n68182 , n58352 , n59628 );
nor ( n68183 , n68181 , n68182 );
or ( n68184 , n68183 , n59637 );
and ( n68185 , n58201 , n59457 );
and ( n68186 , n58200 , n59628 );
nor ( n68187 , n68185 , n68186 );
or ( n68188 , n68187 , n59467 );
nand ( n68189 , n68184 , n68188 );
xor ( n68190 , n414697 , n414723 );
xor ( n68191 , n68190 , n414760 );
buf ( n414916 , n68191 );
xor ( n68193 , n68189 , n414916 );
not ( n68194 , n409507 );
buf ( n414919 , n55984 );
buf ( n414920 , n63625 );
and ( n68197 , n414919 , n414920 );
buf ( n414922 , n58135 );
buf ( n414923 , n63629 );
and ( n68200 , n414922 , n414923 );
nor ( n68201 , n68197 , n68200 );
buf ( n414926 , n68201 );
buf ( n414927 , n414926 );
not ( n68204 , n414927 );
buf ( n414929 , n68204 );
not ( n68206 , n414929 );
or ( n68207 , n68194 , n68206 );
or ( n68208 , n68050 , n409504 );
nand ( n68209 , n68207 , n68208 );
and ( n68210 , n68193 , n68209 );
and ( n68211 , n68189 , n414916 );
or ( n68212 , n68210 , n68211 );
buf ( n414937 , n68212 );
or ( n68214 , n414796 , n409170 );
not ( n68215 , n409429 );
and ( n68216 , n58205 , n59463 );
and ( n68217 , n58166 , n62159 );
nor ( n68218 , n68216 , n68217 );
nand ( n68219 , n68215 , n68218 );
nand ( n68220 , n68214 , n68219 );
buf ( n414945 , n68220 );
buf ( n414946 , n54433 );
buf ( n414947 , n66411 );
and ( n68224 , n414946 , n414947 );
buf ( n414949 , n403088 );
buf ( n414950 , n62496 );
and ( n68227 , n414949 , n414950 );
nor ( n68228 , n68224 , n68227 );
buf ( n414953 , n68228 );
or ( n68230 , n414953 , n410724 );
not ( n68231 , n414813 );
nand ( n68232 , n68231 , n348158 );
nand ( n68233 , n68230 , n68232 );
buf ( n414958 , n68233 );
xor ( n68235 , n414945 , n414958 );
xor ( n68236 , n414738 , n414757 );
buf ( n414961 , n68236 );
buf ( n414962 , n414961 );
buf ( n414963 , n63707 );
buf ( n414964 , n55905 );
and ( n68241 , n414963 , n414964 );
buf ( n414966 , n413104 );
buf ( n414967 , n55895 );
and ( n68244 , n414966 , n414967 );
nor ( n68245 , n68241 , n68244 );
buf ( n414970 , n68245 );
buf ( n414971 , n414970 );
buf ( n414972 , n403120 );
or ( n68249 , n414971 , n414972 );
buf ( n414974 , n414848 );
buf ( n414975 , n403133 );
or ( n68252 , n414974 , n414975 );
nand ( n68253 , n68249 , n68252 );
buf ( n414978 , n68253 );
buf ( n414979 , n414978 );
xor ( n68256 , n414962 , n414979 );
buf ( n414981 , n405381 );
not ( n68258 , n414981 );
buf ( n414983 , n414874 );
not ( n68260 , n414983 );
or ( n68261 , n68258 , n68260 );
buf ( n414986 , n62139 );
buf ( n414987 , n405391 );
and ( n68264 , n414986 , n414987 );
buf ( n414989 , n409140 );
buf ( n414990 , n405388 );
and ( n68267 , n414989 , n414990 );
nor ( n68268 , n68264 , n68267 );
buf ( n414993 , n68268 );
buf ( n414994 , n414993 );
buf ( n414995 , n405407 );
or ( n68272 , n414994 , n414995 );
nand ( n68273 , n68261 , n68272 );
buf ( n414998 , n68273 );
buf ( n414999 , n414998 );
and ( n68276 , n68256 , n414999 );
and ( n68277 , n414962 , n414979 );
or ( n68278 , n68276 , n68277 );
buf ( n415003 , n68278 );
buf ( n415004 , n415003 );
and ( n68281 , n68235 , n415004 );
and ( n68282 , n414945 , n414958 );
or ( n68283 , n68281 , n68282 );
buf ( n415008 , n68283 );
buf ( n415009 , n415008 );
xor ( n68286 , n414937 , n415009 );
xor ( n68287 , n414805 , n414822 );
xor ( n68288 , n68287 , n414888 );
buf ( n415013 , n68288 );
buf ( n415014 , n415013 );
and ( n68291 , n68286 , n415014 );
and ( n68292 , n414937 , n415009 );
or ( n68293 , n68291 , n68292 );
buf ( n415018 , n68293 );
buf ( n415019 , n415018 );
xor ( n68296 , n414783 , n414787 );
xor ( n68297 , n68296 , n414893 );
buf ( n415022 , n68297 );
buf ( n415023 , n415022 );
xor ( n68300 , n415019 , n415023 );
xor ( n68301 , n413334 , n413350 );
xor ( n68302 , n68301 , n66564 );
xor ( n68303 , n413272 , n413289 );
xor ( n68304 , n68303 , n413312 );
buf ( n415029 , n68304 );
or ( n68306 , n413300 , n59467 );
or ( n68307 , n68187 , n59637 );
nand ( n68308 , n68306 , n68307 );
xor ( n68309 , n413367 , n413383 );
xor ( n68310 , n68309 , n413386 );
and ( n68311 , n68308 , n68310 );
xor ( n68312 , n414677 , n414765 );
xor ( n68313 , n68312 , n414778 );
buf ( n415038 , n68313 );
xor ( n68315 , n413367 , n413383 );
xor ( n68316 , n68315 , n413386 );
and ( n68317 , n415038 , n68316 );
and ( n68318 , n68308 , n415038 );
or ( n68319 , n68311 , n68317 , n68318 );
xor ( n68320 , n415029 , n68319 );
xor ( n68321 , n68302 , n68320 );
buf ( n415046 , n68321 );
and ( n68323 , n68300 , n415046 );
and ( n68324 , n415019 , n415023 );
or ( n68325 , n68323 , n68324 );
buf ( n415050 , n68325 );
not ( n68327 , n415050 );
xor ( n68328 , n413334 , n413350 );
xor ( n68329 , n68328 , n66564 );
and ( n68330 , n415029 , n68329 );
xor ( n68331 , n413334 , n413350 );
xor ( n68332 , n68331 , n66564 );
and ( n68333 , n68319 , n68332 );
and ( n68334 , n415029 , n68319 );
or ( n68335 , n68330 , n68333 , n68334 );
not ( n68336 , n68335 );
nand ( n68337 , n68327 , n68336 );
not ( n68338 , n68337 );
or ( n68339 , n68180 , n68338 );
nand ( n68340 , n415050 , n68335 );
nand ( n68341 , n68339 , n68340 );
not ( n68342 , n68341 );
xor ( n68343 , n413331 , n413404 );
xor ( n68344 , n68343 , n413410 );
buf ( n415069 , n68344 );
not ( n68346 , n415069 );
xor ( n68347 , n413182 , n413254 );
xor ( n68348 , n68347 , n413316 );
and ( n68349 , n414897 , n68348 );
xor ( n68350 , n413182 , n413254 );
xor ( n68351 , n68350 , n413316 );
and ( n68352 , n68177 , n68351 );
and ( n68353 , n414897 , n68177 );
or ( n68354 , n68349 , n68352 , n68353 );
not ( n68355 , n68354 );
nand ( n68356 , n68346 , n68355 );
not ( n68357 , n68356 );
or ( n68358 , n68342 , n68357 );
nor ( n68359 , n68346 , n68355 );
not ( n68360 , n68359 );
nand ( n68361 , n68358 , n68360 );
buf ( n415086 , n68361 );
xor ( n68363 , n66499 , n66501 );
xor ( n68364 , n68363 , n413414 );
buf ( n415089 , n68364 );
xor ( n68366 , n415086 , n415089 );
buf ( n415091 , n68366 );
xor ( n68368 , n67931 , n415091 );
not ( n68369 , n68368 );
buf ( n415094 , n45076 );
buf ( n415095 , n64268 );
not ( n68372 , n415095 );
buf ( n415097 , n412964 );
not ( n68374 , n415097 );
or ( n68375 , n68372 , n68374 );
not ( n68376 , n24116 );
buf ( n415101 , n68376 );
buf ( n415102 , n28353 );
nand ( n68379 , n415101 , n415102 );
buf ( n415104 , n68379 );
buf ( n415105 , n415104 );
nand ( n68382 , n68375 , n415105 );
buf ( n415107 , n68382 );
buf ( n415108 , n415107 );
nand ( n68385 , n415094 , n415108 );
buf ( n415110 , n68385 );
nand ( n68387 , n67826 , n41664 );
nand ( n68388 , n415110 , n68387 );
not ( n68389 , n68388 );
not ( n68390 , n406422 );
buf ( n415115 , n407928 );
not ( n415116 , n415115 );
buf ( n415117 , n393185 );
not ( n68394 , n415117 );
and ( n68395 , n415116 , n68394 );
buf ( n415120 , n407936 );
buf ( n415121 , n393185 );
and ( n68398 , n415120 , n415121 );
nor ( n68399 , n68395 , n68398 );
buf ( n415124 , n68399 );
not ( n68401 , n415124 );
not ( n68402 , n68401 );
or ( n68403 , n68390 , n68402 );
buf ( n415128 , n389356 );
buf ( n415129 , n407928 );
and ( n68406 , n415128 , n415129 );
not ( n68407 , n415128 );
buf ( n415132 , n409092 );
and ( n68409 , n68407 , n415132 );
nor ( n68410 , n68406 , n68409 );
buf ( n415135 , n68410 );
or ( n68412 , n415135 , n62075 );
nand ( n68413 , n68403 , n68412 );
not ( n68414 , n68413 );
nand ( n68415 , n68389 , n68414 );
not ( n68416 , n68415 );
or ( n68417 , n68369 , n68416 );
nand ( n68418 , n68413 , n68388 );
nand ( n68419 , n68417 , n68418 );
nand ( n68420 , n67918 , n68419 );
buf ( n415145 , n68420 );
buf ( n415146 , n67916 );
not ( n68423 , n415146 );
buf ( n415148 , n414633 );
nand ( n68425 , n68423 , n415148 );
buf ( n415150 , n68425 );
buf ( n415151 , n415150 );
nand ( n68428 , n415145 , n415151 );
buf ( n415153 , n68428 );
buf ( n415154 , n415153 );
buf ( n415155 , n49117 );
not ( n68432 , n415155 );
buf ( n415157 , n385488 );
not ( n68434 , n415157 );
or ( n68435 , n68432 , n68434 );
buf ( n415160 , n388962 );
buf ( n415161 , n67126 );
nand ( n68438 , n415160 , n415161 );
buf ( n415163 , n68438 );
buf ( n415164 , n415163 );
nand ( n68441 , n68435 , n415164 );
buf ( n415166 , n68441 );
buf ( n415167 , n415166 );
not ( n68444 , n415167 );
buf ( n415169 , n393544 );
not ( n68446 , n415169 );
or ( n68447 , n68444 , n68446 );
buf ( n415172 , n414598 );
buf ( n415173 , n49166 );
nand ( n68450 , n415172 , n415173 );
buf ( n415175 , n68450 );
buf ( n415176 , n415175 );
nand ( n68453 , n68447 , n415176 );
buf ( n415178 , n68453 );
buf ( n415179 , n415178 );
xor ( n68456 , n415154 , n415179 );
buf ( n415181 , n43515 );
not ( n68458 , n415181 );
buf ( n415183 , n411504 );
not ( n68460 , n415183 );
buf ( n415185 , n388409 );
not ( n68462 , n415185 );
or ( n68463 , n68460 , n68462 );
buf ( n415188 , n405785 );
buf ( n415189 , n391024 );
nand ( n68466 , n415188 , n415189 );
buf ( n415191 , n68466 );
buf ( n415192 , n415191 );
nand ( n68469 , n68463 , n415192 );
buf ( n415194 , n68469 );
buf ( n415195 , n415194 );
not ( n68472 , n415195 );
or ( n68473 , n68458 , n68472 );
buf ( n415198 , n411504 );
not ( n68475 , n415198 );
buf ( n415200 , n388367 );
not ( n68477 , n415200 );
or ( n68478 , n68475 , n68477 );
buf ( n415203 , n397069 );
buf ( n415204 , n391024 );
nand ( n68481 , n415203 , n415204 );
buf ( n415206 , n68481 );
buf ( n415207 , n415206 );
nand ( n68484 , n68478 , n415207 );
buf ( n415209 , n68484 );
buf ( n415210 , n415209 );
buf ( n415211 , n43536 );
nand ( n68488 , n415210 , n415211 );
buf ( n415213 , n68488 );
buf ( n415214 , n415213 );
nand ( n68491 , n68473 , n415214 );
buf ( n415216 , n68491 );
buf ( n415217 , n415216 );
and ( n68494 , n68456 , n415217 );
and ( n68495 , n415154 , n415179 );
or ( n68496 , n68494 , n68495 );
buf ( n415221 , n68496 );
not ( n68498 , n415221 );
or ( n68499 , n67892 , n68498 );
buf ( n415224 , n414481 );
buf ( n415225 , n67890 );
not ( n68502 , n415225 );
buf ( n415227 , n68502 );
buf ( n415228 , n415227 );
nand ( n68505 , n415224 , n415228 );
buf ( n415230 , n68505 );
nand ( n68507 , n68499 , n415230 );
buf ( n415232 , n68507 );
and ( n68509 , n67733 , n415232 );
and ( n68510 , n414453 , n414456 );
or ( n68511 , n68509 , n68510 );
buf ( n415236 , n68511 );
not ( n68513 , n415236 );
or ( n68514 , n67725 , n68513 );
buf ( n415239 , C1 );
nand ( n68520 , n68514 , n415239 );
buf ( n415241 , n68520 );
xor ( n68522 , n414442 , n415241 );
not ( n68524 , n413721 );
and ( n68525 , n68524 , C1 );
nor ( n68526 , C0 , n68525 );
buf ( n415246 , n68526 );
buf ( n415247 , n413729 );
xor ( n68529 , n415246 , n415247 );
buf ( n415249 , n68529 );
buf ( n415250 , n415249 );
and ( n68532 , n68522 , n415250 );
and ( n68533 , n414442 , n415241 );
or ( n68534 , n68532 , n68533 );
buf ( n415254 , n68534 );
buf ( n415255 , n415254 );
not ( n68537 , n415255 );
buf ( n415257 , n68537 );
not ( n68539 , n415257 );
xor ( n68540 , n414058 , n413756 );
and ( n68541 , n68540 , n66926 );
not ( n68542 , n68540 );
and ( n68543 , n68542 , n66925 );
nor ( n68544 , n68541 , n68543 );
not ( n68545 , n68544 );
not ( n68546 , n68545 );
and ( n68547 , n68539 , n68546 );
buf ( n415267 , n415257 );
buf ( n415268 , n68545 );
nand ( n68550 , n415267 , n415268 );
buf ( n415270 , n68550 );
buf ( n415271 , n66965 );
not ( n68553 , n415271 );
buf ( n415273 , n413893 );
not ( n68555 , n415273 );
or ( n68556 , n68553 , n68555 );
buf ( n415276 , n413890 );
buf ( n415277 , n413774 );
nand ( n68559 , n415276 , n415277 );
buf ( n415279 , n68559 );
buf ( n415280 , n415279 );
nand ( n68562 , n68556 , n415280 );
buf ( n415282 , n68562 );
xnor ( n68564 , n415282 , n414047 );
buf ( n415284 , n68564 );
not ( n68566 , n415284 );
buf ( n415286 , n68566 );
buf ( n415287 , n415286 );
not ( n68569 , n415287 );
and ( n68570 , n413884 , n413798 );
not ( n68571 , n413884 );
and ( n68572 , n68571 , n413801 );
or ( n68573 , n68570 , n68572 );
xnor ( n68574 , n68573 , n413821 );
not ( n68575 , n68574 );
xor ( n68576 , n413921 , n414038 );
xor ( n68577 , n68576 , n414043 );
buf ( n415297 , n68577 );
buf ( n415298 , n415297 );
not ( n68580 , n415298 );
buf ( n415300 , n68580 );
not ( n68582 , n415300 );
and ( n68583 , n68575 , n68582 );
buf ( n415303 , n68574 );
buf ( n415304 , n415300 );
nand ( n68586 , n415303 , n415304 );
buf ( n415306 , n68586 );
not ( n68588 , n395362 );
not ( n68589 , n413694 );
or ( n68590 , n68588 , n68589 );
buf ( n415310 , n47863 );
not ( n68592 , n415310 );
buf ( n415312 , n388955 );
not ( n68594 , n415312 );
or ( n68595 , n68592 , n68594 );
buf ( n415315 , n37763 );
buf ( n415316 , n395312 );
nand ( n68598 , n415315 , n415316 );
buf ( n415318 , n68598 );
buf ( n415319 , n415318 );
nand ( n68601 , n68595 , n415319 );
buf ( n415321 , n68601 );
buf ( n415322 , n415321 );
buf ( n415323 , n395349 );
nand ( n68605 , n415322 , n415323 );
buf ( n415325 , n68605 );
nand ( n68607 , n68590 , n415325 );
not ( n68608 , n68607 );
not ( n68609 , n67195 );
not ( n68610 , n414010 );
or ( n68611 , n68609 , n68610 );
nand ( n68612 , n414007 , n414000 );
nand ( n68613 , n68611 , n68612 );
not ( n68614 , n67168 );
and ( n68615 , n68613 , n68614 );
not ( n68616 , n68613 );
and ( n68617 , n68616 , n67168 );
nor ( n68618 , n68615 , n68617 );
not ( n68619 , n397102 );
buf ( n415339 , n394210 );
not ( n68621 , n415339 );
buf ( n415341 , n46906 );
not ( n68623 , n415341 );
or ( n68624 , n68621 , n68623 );
buf ( n415344 , n22982 );
buf ( n415345 , n394207 );
nand ( n68627 , n415344 , n415345 );
buf ( n415347 , n68627 );
buf ( n415348 , n415347 );
nand ( n68630 , n68624 , n415348 );
buf ( n415350 , n68630 );
not ( n68632 , n415350 );
or ( n68633 , n68619 , n68632 );
buf ( n415353 , n414494 );
buf ( n415354 , n393127 );
nand ( n68636 , n415353 , n415354 );
buf ( n415356 , n68636 );
nand ( n68638 , n68633 , n415356 );
not ( n68639 , n68638 );
not ( n68640 , n390362 );
not ( n68641 , n413990 );
or ( n68642 , n68640 , n68641 );
and ( n68643 , n46476 , n46474 );
and ( n68644 , n40601 , n68643 );
not ( n68645 , n40601 );
and ( n68646 , n68645 , n49686 );
or ( n68647 , n68644 , n68646 );
nand ( n68648 , n68647 , n67042 );
nand ( n68649 , n68642 , n68648 );
not ( n68650 , n68649 );
or ( n68651 , n68639 , n68650 );
buf ( n415371 , n68638 );
not ( n68653 , n415371 );
buf ( n415373 , n68653 );
not ( n68655 , n415373 );
buf ( n415375 , n68649 );
not ( n68657 , n415375 );
buf ( n415377 , n68657 );
not ( n68659 , n415377 );
or ( n68660 , n68655 , n68659 );
not ( n68661 , n414578 );
not ( n68662 , n414543 );
or ( n68663 , n68661 , n68662 );
buf ( n415383 , n414540 );
buf ( n415384 , n414575 );
nand ( n68666 , n415383 , n415384 );
buf ( n415386 , n68666 );
nand ( n68668 , n68663 , n415386 );
buf ( n68669 , n67802 );
xor ( n68670 , n68668 , n68669 );
nand ( n68671 , n68660 , n68670 );
nand ( n68672 , n68651 , n68671 );
not ( n68673 , n68672 );
buf ( n415393 , n393369 );
not ( n68675 , n415393 );
buf ( n415395 , n38630 );
not ( n68677 , n415395 );
or ( n68678 , n68675 , n68677 );
buf ( n415398 , n388928 );
buf ( n415399 , n393381 );
nand ( n68681 , n415398 , n415399 );
buf ( n415401 , n68681 );
buf ( n415402 , n415401 );
nand ( n68684 , n68678 , n415402 );
buf ( n415404 , n68684 );
nand ( n68686 , n415404 , n45954 );
nand ( n68687 , n388293 , n393369 );
not ( n68688 , n68687 );
buf ( n415408 , n375784 );
buf ( n415409 , n393381 );
nand ( n68691 , n415408 , n415409 );
buf ( n415411 , n68691 );
not ( n68693 , n415411 );
or ( n68694 , n68688 , n68693 );
nand ( n68695 , n68694 , n45949 );
nand ( n68696 , n68673 , n68686 , n68695 );
and ( n68697 , n68618 , n68696 );
nand ( n68698 , n68686 , n68695 );
and ( n68699 , n68698 , n68672 );
nor ( n68700 , n68697 , n68699 );
nand ( n68701 , n68608 , n68700 );
not ( n68702 , n68701 );
not ( n68703 , n43515 );
not ( n68704 , n413871 );
or ( n68705 , n68703 , n68704 );
buf ( n415425 , n415194 );
buf ( n415426 , n43536 );
nand ( n68708 , n415425 , n415426 );
buf ( n415428 , n68708 );
nand ( n68710 , n68705 , n415428 );
not ( n68711 , n68710 );
not ( n68712 , n414163 );
not ( n68713 , n414167 );
not ( n68714 , n68713 );
or ( n68715 , n68712 , n68714 );
nand ( n68716 , n414167 , n414160 );
nand ( n68717 , n68715 , n68716 );
and ( n415437 , n68717 , n67425 );
not ( n68719 , n68717 );
not ( n68720 , n67425 );
and ( n68721 , n68719 , n68720 );
nor ( n68722 , n415437 , n68721 );
not ( n68723 , n68722 );
nand ( n68724 , n68711 , n68723 );
not ( n68725 , n68724 );
not ( n68726 , n398668 );
not ( n68727 , n413940 );
not ( n68728 , n68727 );
or ( n68729 , n68726 , n68728 );
buf ( n415449 , n397498 );
not ( n68731 , n415449 );
buf ( n415451 , n391563 );
not ( n68733 , n415451 );
or ( n68734 , n68731 , n68733 );
buf ( n415454 , n388905 );
buf ( n415455 , n397495 );
nand ( n68737 , n415454 , n415455 );
buf ( n415457 , n68737 );
buf ( n415458 , n415457 );
nand ( n68740 , n68734 , n415458 );
buf ( n415460 , n68740 );
nand ( n68742 , n415460 , n37338 );
nand ( n68743 , n68729 , n68742 );
not ( n68744 , n68743 );
or ( n68745 , n68725 , n68744 );
nand ( n68746 , n68722 , n68710 );
nand ( n68747 , n68745 , n68746 );
not ( n68748 , n68747 );
or ( n68749 , n68702 , n68748 );
not ( n68750 , n68700 );
nand ( n68751 , n68750 , n68607 );
nand ( n68752 , n68749 , n68751 );
buf ( n415472 , n68752 );
buf ( n68754 , n415472 );
buf ( n415474 , n68754 );
and ( n68756 , n415306 , n415474 );
nor ( n68757 , n68583 , n68756 );
buf ( n415477 , n68757 );
not ( n68759 , n415477 );
buf ( n415479 , n68759 );
buf ( n415480 , n415479 );
not ( n68762 , n415480 );
or ( n68763 , n68569 , n68762 );
buf ( n415483 , n68564 );
not ( n68765 , n415483 );
buf ( n415485 , n68757 );
not ( n68767 , n415485 );
or ( n68768 , n68765 , n68767 );
xor ( n68769 , n413487 , n413490 );
xor ( n68770 , n68769 , n413516 );
buf ( n415490 , n68770 );
buf ( n415491 , n415490 );
not ( n68773 , n415491 );
buf ( n415493 , n68773 );
buf ( n415494 , n415493 );
not ( n68776 , n415494 );
buf ( n415496 , n413788 );
not ( n68778 , n415496 );
buf ( n415498 , n40969 );
not ( n68780 , n415498 );
and ( n68781 , n68778 , n68780 );
buf ( n415501 , n390260 );
buf ( n415502 , n400033 );
not ( n68784 , n415502 );
buf ( n415504 , n36395 );
not ( n68786 , n415504 );
or ( n68787 , n68784 , n68786 );
buf ( n415507 , n40977 );
buf ( n415508 , n400042 );
nand ( n68790 , n415507 , n415508 );
buf ( n415510 , n68790 );
buf ( n415511 , n415510 );
nand ( n68793 , n68787 , n415511 );
buf ( n415513 , n68793 );
buf ( n415514 , n415513 );
and ( n68796 , n415501 , n415514 );
nor ( n68797 , n68781 , n68796 );
buf ( n415517 , n68797 );
not ( n68799 , n415517 );
buf ( n415519 , n358975 );
buf ( n415520 , n390307 );
and ( n68802 , n415519 , n415520 );
not ( n68803 , n415519 );
buf ( n415523 , n40886 );
and ( n68805 , n68803 , n415523 );
nor ( n68806 , n68802 , n68805 );
buf ( n415526 , n68806 );
buf ( n415527 , n415526 );
not ( n68809 , n415527 );
buf ( n415529 , n36801 );
not ( n68811 , n415529 );
or ( n68812 , n68809 , n68811 );
buf ( n415532 , n67002 );
not ( n68814 , n415532 );
buf ( n415534 , n388669 );
nand ( n68816 , n68814 , n415534 );
buf ( n415536 , n68816 );
buf ( n415537 , n415536 );
nand ( n68819 , n68812 , n415537 );
buf ( n415539 , n68819 );
buf ( n415540 , n415539 );
not ( n68822 , n415540 );
buf ( n415542 , n68822 );
not ( n68824 , n415542 );
and ( n68825 , n68799 , n68824 );
buf ( n415545 , n415517 );
buf ( n415546 , n415542 );
nand ( n68828 , n415545 , n415546 );
buf ( n415548 , n68828 );
not ( n68830 , n414506 );
nand ( n68831 , n68830 , n414613 );
not ( n68832 , n68831 );
not ( n68833 , n67861 );
or ( n68834 , n68832 , n68833 );
buf ( n415554 , n414610 );
buf ( n415555 , n414506 );
nand ( n68837 , n415554 , n415555 );
buf ( n415557 , n68837 );
nand ( n68839 , n68834 , n415557 );
and ( n68840 , n415548 , n68839 );
nor ( n68841 , n68825 , n68840 );
buf ( n415561 , n68841 );
not ( n68843 , n415561 );
or ( n68844 , n68776 , n68843 );
xor ( n68845 , n414126 , n414227 );
xnor ( n68846 , n68845 , n414141 );
buf ( n415566 , n68846 );
not ( n68848 , n415566 );
buf ( n415568 , n68848 );
buf ( n415569 , n415568 );
not ( n68851 , n415569 );
buf ( n415571 , n45954 );
not ( n68853 , n415571 );
buf ( n415573 , n413910 );
not ( n68855 , n415573 );
or ( n68856 , n68853 , n68855 );
buf ( n415576 , n415404 );
buf ( n415577 , n45949 );
nand ( n68859 , n415576 , n415577 );
buf ( n415579 , n68859 );
buf ( n415580 , n415579 );
nand ( n68862 , n68856 , n415580 );
buf ( n415582 , n68862 );
buf ( n415583 , n415582 );
not ( n68865 , n415583 );
or ( n68866 , n68851 , n68865 );
buf ( n415586 , n415582 );
not ( n68868 , n415586 );
buf ( n415588 , n68868 );
buf ( n415589 , n415588 );
not ( n68871 , n415589 );
buf ( n415591 , n68846 );
not ( n68873 , n415591 );
or ( n68874 , n68871 , n68873 );
buf ( n415594 , n392611 );
not ( n68876 , n415594 );
buf ( n415596 , n399164 );
not ( n68878 , n415596 );
or ( n68879 , n68876 , n68878 );
buf ( n415599 , n24049 );
buf ( n415600 , n392620 );
nand ( n68882 , n415599 , n415600 );
buf ( n415602 , n68882 );
buf ( n415603 , n415602 );
nand ( n68885 , n68879 , n415603 );
buf ( n415605 , n68885 );
buf ( n415606 , n415605 );
not ( n68888 , n415606 );
buf ( n415608 , n396622 );
not ( n68890 , n415608 );
or ( n68891 , n68888 , n68890 );
buf ( n415611 , n46921 );
buf ( n415612 , n413967 );
nand ( n68894 , n415611 , n415612 );
buf ( n415614 , n68894 );
buf ( n415615 , n415614 );
nand ( n68897 , n68891 , n415615 );
buf ( n415617 , n68897 );
not ( n68899 , n415617 );
buf ( n415619 , n415135 );
not ( n68901 , n415619 );
buf ( n415621 , n68901 );
buf ( n415622 , n415621 );
not ( n68904 , n415622 );
buf ( n415624 , n60872 );
not ( n68906 , n415624 );
or ( n68907 , n68904 , n68906 );
buf ( n415627 , n414181 );
buf ( n415628 , n409076 );
nand ( n68910 , n415627 , n415628 );
buf ( n415630 , n68910 );
buf ( n415631 , n415630 );
nand ( n68913 , n68907 , n415631 );
buf ( n415633 , n68913 );
or ( n68915 , n68361 , n68364 );
not ( n68916 , n68915 );
not ( n68917 , n67931 );
or ( n68918 , n68916 , n68917 );
nand ( n68919 , n68361 , n68364 );
nand ( n68920 , n68918 , n68919 );
xor ( n68921 , n415633 , n68920 );
buf ( n415641 , n388809 );
not ( n68923 , n415641 );
buf ( n415643 , n67809 );
not ( n68925 , n415643 );
or ( n68926 , n68923 , n68925 );
and ( n68927 , n12471 , n388754 );
not ( n68928 , n12471 );
and ( n68929 , n68928 , n405736 );
or ( n68930 , n68927 , n68929 );
buf ( n415650 , n68930 );
buf ( n415651 , n388746 );
nand ( n68933 , n415650 , n415651 );
buf ( n415653 , n68933 );
buf ( n415654 , n415653 );
nand ( n68936 , n68926 , n415654 );
buf ( n415656 , n68936 );
and ( n68938 , n68921 , n415656 );
and ( n68939 , n415633 , n68920 );
or ( n68940 , n68938 , n68939 );
not ( n68941 , n68940 );
or ( n68942 , n68899 , n68941 );
buf ( n415662 , n68940 );
not ( n68944 , n415662 );
buf ( n415664 , n68944 );
not ( n68946 , n415664 );
buf ( n415666 , n415617 );
not ( n68948 , n415666 );
buf ( n415668 , n68948 );
not ( n68950 , n415668 );
or ( n68951 , n68946 , n68950 );
xor ( n68952 , n67418 , n414193 );
xnor ( n68953 , n68952 , n67423 );
buf ( n415673 , n68953 );
not ( n68955 , n415673 );
buf ( n415675 , n68955 );
nand ( n68957 , n68951 , n415675 );
nand ( n68958 , n68942 , n68957 );
buf ( n415678 , n68958 );
buf ( n415679 , n45260 );
not ( n68961 , n415679 );
buf ( n415681 , n44776 );
buf ( n415682 , n43044 );
and ( n68964 , n415681 , n415682 );
not ( n68965 , n415681 );
buf ( n415685 , n27195 );
and ( n68967 , n68965 , n415685 );
nor ( n68968 , n68964 , n68967 );
buf ( n415688 , n68968 );
buf ( n415689 , n415688 );
not ( n68971 , n415689 );
or ( n68972 , n68961 , n68971 );
nand ( n68973 , n66859 , n413643 );
buf ( n415693 , n68973 );
nand ( n68975 , n68972 , n415693 );
buf ( n415695 , n68975 );
buf ( n415696 , n415695 );
xor ( n68978 , n415678 , n415696 );
buf ( n415698 , n388402 );
buf ( n415699 , n402819 );
nor ( n68981 , n415698 , n415699 );
buf ( n415701 , n68981 );
buf ( n415702 , n415701 );
and ( n68984 , n68978 , n415702 );
and ( n68985 , n415678 , n415696 );
or ( n68986 , n68984 , n68985 );
buf ( n415706 , n68986 );
buf ( n415707 , n415706 );
nand ( n68989 , n68874 , n415707 );
buf ( n415709 , n68989 );
buf ( n415710 , n415709 );
nand ( n68992 , n68866 , n415710 );
buf ( n415712 , n68992 );
buf ( n415713 , n415712 );
nand ( n68995 , n68844 , n415713 );
buf ( n415715 , n68995 );
buf ( n415716 , n415715 );
buf ( n415717 , n415493 );
not ( n68999 , n415717 );
buf ( n415719 , n68841 );
not ( n69001 , n415719 );
buf ( n415721 , n69001 );
buf ( n415722 , n415721 );
nand ( n69004 , n68999 , n415722 );
buf ( n415724 , n69004 );
buf ( n415725 , n415724 );
nand ( n69007 , n415716 , n415725 );
buf ( n415727 , n69007 );
buf ( n415728 , n415727 );
nand ( n69010 , n68768 , n415728 );
buf ( n415730 , n69010 );
buf ( n415731 , n415730 );
nand ( n69013 , n68763 , n415731 );
buf ( n415733 , n69013 );
buf ( n415734 , n415733 );
not ( n69016 , n415734 );
buf ( n415736 , n69016 );
buf ( n415737 , n415736 );
not ( n69019 , n415737 );
buf ( n415739 , n69019 );
and ( n69021 , n415270 , n415739 );
nor ( n69022 , n68547 , n69021 );
buf ( n415742 , n69022 );
and ( n69024 , n67695 , n415742 );
and ( n69025 , n414430 , n414437 );
or ( n69026 , n69024 , n69025 );
buf ( n415746 , n69026 );
buf ( n415747 , n415746 );
xor ( n69029 , n414423 , n415747 );
not ( n69030 , n67464 );
buf ( n415750 , n413606 );
not ( n69032 , n415750 );
buf ( n415752 , n69032 );
not ( n69034 , n415752 );
or ( n69035 , n69030 , n69034 );
not ( n69036 , n67464 );
nand ( n69037 , n69036 , n413606 );
nand ( n415757 , n69035 , n69037 );
xor ( n69039 , n415757 , n67608 );
buf ( n415759 , n69039 );
and ( n69041 , n69029 , n415759 );
and ( n69042 , n414423 , n415747 );
or ( n69043 , n69041 , n69042 );
buf ( n415763 , n69043 );
nand ( n69045 , n414401 , n415763 );
buf ( n415765 , n69045 );
xor ( n69047 , n414423 , n415747 );
xor ( n69048 , n69047 , n415759 );
buf ( n415768 , n69048 );
buf ( n415769 , n415768 );
not ( n69051 , n67485 );
buf ( n415771 , n67468 );
not ( n69053 , n415771 );
buf ( n415773 , n69053 );
not ( n69055 , n415773 );
or ( n69056 , n69051 , n69055 );
nand ( n69057 , n67468 , n67484 );
nand ( n69058 , n69056 , n69057 );
buf ( n415778 , n69058 );
buf ( n415779 , n414349 );
not ( n69061 , n415779 );
buf ( n415781 , n69061 );
buf ( n415782 , n415781 );
and ( n69064 , n415778 , n415782 );
not ( n69065 , n415778 );
buf ( n415785 , n414349 );
and ( n69067 , n69065 , n415785 );
nor ( n69068 , n69064 , n69067 );
buf ( n415788 , n69068 );
buf ( n415789 , n415788 );
buf ( n415790 , n68544 );
buf ( n415791 , n415733 );
and ( n69073 , n415790 , n415791 );
not ( n69074 , n415790 );
buf ( n415794 , n415736 );
and ( n69076 , n69074 , n415794 );
nor ( n69077 , n69073 , n69076 );
buf ( n415797 , n69077 );
buf ( n415798 , n415797 );
buf ( n415799 , n415254 );
and ( n69081 , n415798 , n415799 );
not ( n69082 , n415798 );
buf ( n415802 , n415257 );
and ( n69084 , n69082 , n415802 );
nor ( n69085 , n69081 , n69084 );
buf ( n415805 , n69085 );
buf ( n415806 , n415805 );
xor ( n69088 , n414300 , n414341 );
xor ( n69089 , n69088 , n414345 );
buf ( n415809 , n69089 );
not ( n69091 , n415809 );
buf ( n415811 , n69091 );
buf ( n415812 , n67474 );
buf ( n415813 , n67471 );
xor ( n69095 , n415812 , n415813 );
buf ( n415815 , n67482 );
xnor ( n69097 , n69095 , n415815 );
buf ( n415817 , n69097 );
buf ( n415818 , n415817 );
nand ( n69100 , n415811 , n415818 );
buf ( n415820 , n69100 );
buf ( n415821 , n415820 );
nand ( n69103 , n415806 , n415821 );
buf ( n415823 , n69103 );
buf ( n415824 , n415823 );
buf ( n415825 , n69091 );
buf ( n415826 , n415817 );
or ( n69108 , n415825 , n415826 );
buf ( n415828 , n69108 );
buf ( n415829 , n415828 );
and ( n69111 , n415824 , n415829 );
buf ( n415831 , n69111 );
buf ( n415832 , n415831 );
xor ( n69114 , n415789 , n415832 );
xor ( n69115 , n414430 , n414437 );
xor ( n69116 , n69115 , n415742 );
buf ( n415836 , n69116 );
buf ( n415837 , n415836 );
and ( n69119 , n69114 , n415837 );
and ( n69120 , n415789 , n415832 );
or ( n69121 , n69119 , n69120 );
buf ( n415841 , n69121 );
buf ( n415842 , n415841 );
nand ( n69124 , n415769 , n415842 );
buf ( n415844 , n69124 );
buf ( n415845 , n415844 );
xor ( n69127 , n415789 , n415832 );
xor ( n69128 , n69127 , n415837 );
buf ( n415848 , n69128 );
buf ( n415849 , n415848 );
xor ( n69131 , n415817 , n415809 );
xnor ( n69132 , n69131 , n415805 );
buf ( n415852 , n69132 );
buf ( n69134 , n415852 );
buf ( n415854 , n69134 );
buf ( n415855 , n415854 );
not ( n69137 , n67536 );
not ( n69138 , n414338 );
nand ( n69139 , n69137 , n69138 , C1 );
nand ( n69140 , n67536 , n414338 , C1 );
nand ( n69144 , n69139 , n69140 , C1 , C1 );
xor ( n69145 , n413640 , n413669 );
xor ( n69146 , n69145 , n413674 );
buf ( n415863 , n69146 );
buf ( n415864 , n415863 );
buf ( n415865 , C0 );
buf ( n415866 , n415865 );
xor ( n69174 , n415864 , n415866 );
buf ( n415868 , n55055 );
not ( n69176 , n415868 );
buf ( n415870 , n40978 );
not ( n69178 , n415870 );
or ( n69179 , n69176 , n69178 );
buf ( n415873 , n36396 );
buf ( n415874 , n55054 );
nand ( n69182 , n415873 , n415874 );
buf ( n415876 , n69182 );
buf ( n415877 , n415876 );
nand ( n69185 , n69179 , n415877 );
buf ( n415879 , n69185 );
buf ( n415880 , n415879 );
not ( n69188 , n415880 );
buf ( n415882 , n388460 );
not ( n69190 , n415882 );
or ( n69191 , n69188 , n69190 );
buf ( n415885 , n415513 );
buf ( n415886 , n43272 );
nand ( n69194 , n415885 , n415886 );
buf ( n415888 , n69194 );
buf ( n415889 , n415888 );
nand ( n69197 , n69191 , n415889 );
buf ( n415891 , n69197 );
buf ( n415892 , n415891 );
buf ( n415893 , n395349 );
not ( n69201 , n415893 );
and ( n69202 , n47863 , n391483 );
not ( n69203 , n47863 );
and ( n69204 , n69203 , n29077 );
or ( n69205 , n69202 , n69204 );
buf ( n415899 , n69205 );
not ( n69207 , n415899 );
or ( n69208 , n69201 , n69207 );
buf ( n415902 , n415321 );
buf ( n415903 , n395362 );
nand ( n69211 , n415902 , n415903 );
buf ( n415905 , n69211 );
buf ( n415906 , n415905 );
nand ( n69214 , n69208 , n415906 );
buf ( n415908 , n69214 );
buf ( n415909 , n415908 );
xor ( n69217 , n415892 , n415909 );
buf ( n415911 , n389936 );
not ( n69219 , n415911 );
buf ( n415913 , n36360 );
not ( n69221 , n415913 );
or ( n69222 , n69219 , n69221 );
buf ( n415916 , n358975 );
nand ( n69224 , n69222 , n415916 );
buf ( n415918 , n69224 );
buf ( n415919 , n415918 );
buf ( n415920 , n40839 );
buf ( n415921 , n36360 );
not ( n69229 , n415921 );
buf ( n415923 , n40775 );
nand ( n69231 , n69229 , n415923 );
buf ( n415925 , n69231 );
buf ( n415926 , n415925 );
nand ( n69234 , n415919 , n415920 , n415926 );
buf ( n415928 , n69234 );
buf ( n415929 , n415928 );
not ( n69237 , n415929 );
buf ( n415931 , n69237 );
buf ( n415932 , n415931 );
not ( n69240 , n415932 );
buf ( n415934 , n413643 );
not ( n69242 , n415934 );
buf ( n415936 , n415688 );
not ( n69244 , n415936 );
or ( n69245 , n69242 , n69244 );
not ( n69246 , n40813 );
not ( n69247 , n44776 );
and ( n69248 , n28213 , n69247 );
not ( n69249 , n28213 );
not ( n69250 , n399986 );
and ( n69251 , n69249 , n69250 );
or ( n69252 , n69248 , n69251 );
and ( n69253 , n69246 , n69252 );
not ( n69254 , n69246 );
not ( n69255 , n44776 );
and ( n69256 , n28203 , n69255 );
not ( n69257 , n28203 );
not ( n69258 , n399986 );
and ( n69259 , n69257 , n69258 );
or ( n69260 , n69256 , n69259 );
and ( n69261 , n69254 , n69260 );
or ( n69262 , n69253 , n69261 );
nand ( n69263 , n69262 , n45260 );
buf ( n415957 , n69263 );
nand ( n69265 , n69245 , n415957 );
buf ( n415959 , n69265 );
buf ( n415960 , n415959 );
not ( n69268 , n415960 );
or ( n69269 , n69240 , n69268 );
buf ( n415963 , n415928 );
not ( n69271 , n415963 );
buf ( n415965 , n415959 );
not ( n69273 , n415965 );
buf ( n415967 , n69273 );
buf ( n415968 , n415967 );
not ( n69276 , n415968 );
or ( n69277 , n69271 , n69276 );
not ( n69278 , n43515 );
not ( n69279 , n415209 );
or ( n69280 , n69278 , n69279 );
not ( n69281 , n45699 );
not ( n69282 , n411504 );
or ( n69283 , n69281 , n69282 );
or ( n69284 , n52763 , n411504 );
nand ( n69285 , n69283 , n69284 );
nand ( n69286 , n69285 , n43536 );
nand ( n69287 , n69280 , n69286 );
not ( n69288 , n390362 );
not ( n69289 , n68647 );
or ( n69290 , n69288 , n69289 );
buf ( n415984 , n40601 );
not ( n69292 , n415984 );
buf ( n415986 , n388566 );
not ( n69294 , n415986 );
or ( n69295 , n69292 , n69294 );
buf ( n415989 , n27258 );
buf ( n415990 , n40600 );
nand ( n69298 , n415989 , n415990 );
buf ( n415992 , n69298 );
buf ( n415993 , n415992 );
nand ( n69301 , n69295 , n415993 );
buf ( n415995 , n69301 );
buf ( n415996 , n415995 );
buf ( n415997 , n40592 );
nand ( n69305 , n415996 , n415997 );
buf ( n415999 , n69305 );
nand ( n69307 , n69290 , n415999 );
or ( n69308 , n69287 , n69307 );
xor ( n69309 , n415633 , n68920 );
xor ( n69310 , n69309 , n415656 );
nand ( n69311 , n69308 , n69310 );
buf ( n416005 , n69311 );
buf ( n416006 , n69287 );
buf ( n416007 , n69307 );
nand ( n69315 , n416006 , n416007 );
buf ( n416009 , n69315 );
buf ( n416010 , n416009 );
and ( n69318 , n416005 , n416010 );
buf ( n416012 , n69318 );
buf ( n416013 , n416012 );
not ( n69321 , n416013 );
buf ( n416015 , n69321 );
buf ( n416016 , n416015 );
nand ( n69324 , n69277 , n416016 );
buf ( n416018 , n69324 );
buf ( n416019 , n416018 );
nand ( n69327 , n69269 , n416019 );
buf ( n416021 , n69327 );
buf ( n416022 , n416021 );
and ( n69330 , n69217 , n416022 );
and ( n69331 , n415892 , n415909 );
or ( n69332 , n69330 , n69331 );
buf ( n416026 , n69332 );
buf ( n416027 , n416026 );
and ( n69335 , n69174 , n416027 );
or ( n69337 , n69335 , C0 );
buf ( n416030 , n69337 );
buf ( n416031 , n416030 );
not ( n69340 , n416031 );
xor ( n69341 , n414306 , n414309 );
xor ( n69342 , n69341 , n414335 );
buf ( n416035 , n69342 );
buf ( n416036 , n416035 );
buf ( n69345 , n416036 );
buf ( n416038 , n69345 );
buf ( n416039 , n416038 );
not ( n69348 , n416039 );
or ( n69349 , n69340 , n69348 );
buf ( n416042 , n416038 );
buf ( n416043 , n416030 );
or ( n416044 , n416042 , n416043 );
buf ( n416045 , n415490 );
buf ( n416046 , n415712 );
xor ( n69355 , n416045 , n416046 );
buf ( n416048 , n415721 );
xor ( n69357 , n69355 , n416048 );
buf ( n416050 , n69357 );
buf ( n416051 , n416050 );
nand ( n69360 , n416044 , n416051 );
buf ( n416053 , n69360 );
buf ( n416054 , n416053 );
nand ( n69363 , n69349 , n416054 );
buf ( n416056 , n69363 );
xor ( n69365 , n69144 , n416056 );
buf ( n416058 , n61577 );
not ( n69367 , n416058 );
buf ( n416060 , n414324 );
not ( n69369 , n416060 );
or ( n69370 , n69367 , n69369 );
not ( n69371 , n50584 );
not ( n69372 , n385983 );
or ( n69373 , n69371 , n69372 );
nand ( n69374 , n390651 , n47891 );
nand ( n69375 , n69373 , n69374 );
buf ( n416068 , n69375 );
buf ( n416069 , n50579 );
nand ( n69378 , n416068 , n416069 );
buf ( n416071 , n69378 );
buf ( n416072 , n416071 );
nand ( n69381 , n69370 , n416072 );
buf ( n416074 , n69381 );
buf ( n416075 , n416074 );
buf ( n416076 , n68839 );
buf ( n416077 , n415539 );
xor ( n69386 , n416076 , n416077 );
buf ( n416079 , n415517 );
xnor ( n69388 , n69386 , n416079 );
buf ( n416081 , n69388 );
buf ( n416082 , n416081 );
xor ( n69391 , n416075 , n416082 );
buf ( n416084 , n68638 );
not ( n69393 , n416084 );
buf ( n416086 , n415377 );
not ( n69395 , n416086 );
or ( n69396 , n69393 , n69395 );
buf ( n416089 , n68649 );
buf ( n416090 , n415373 );
nand ( n69399 , n416089 , n416090 );
buf ( n416092 , n69399 );
buf ( n416093 , n416092 );
nand ( n69402 , n69396 , n416093 );
buf ( n416095 , n69402 );
buf ( n416096 , n416095 );
buf ( n416097 , n68670 );
not ( n69406 , n416097 );
buf ( n416099 , n69406 );
buf ( n416100 , n416099 );
and ( n69409 , n416096 , n416100 );
not ( n69410 , n416096 );
buf ( n416103 , n68670 );
and ( n69412 , n69410 , n416103 );
nor ( n69413 , n69409 , n69412 );
buf ( n416106 , n69413 );
buf ( n416107 , n416106 );
not ( n69416 , n416107 );
buf ( n416109 , n69416 );
not ( n69418 , n416109 );
buf ( n416111 , n393369 );
buf ( n416112 , n40759 );
and ( n69421 , n416111 , n416112 );
not ( n69422 , n416111 );
buf ( n416115 , n40758 );
and ( n69424 , n69422 , n416115 );
nor ( n69425 , n69421 , n69424 );
buf ( n416118 , n69425 );
not ( n69427 , n416118 );
not ( n69428 , n393404 );
and ( n69429 , n69427 , n69428 );
nand ( n69430 , n415411 , n68687 );
and ( n69431 , n69430 , n45954 );
nor ( n69432 , n69429 , n69431 );
buf ( n416125 , n69432 );
not ( n69434 , n416125 );
buf ( n416127 , n69434 );
not ( n69436 , n416127 );
or ( n69437 , n69418 , n69436 );
not ( n69438 , n69432 );
not ( n69439 , n416106 );
or ( n69440 , n69438 , n69439 );
buf ( n416133 , n415664 );
not ( n69442 , n416133 );
buf ( n416135 , n415675 );
not ( n69444 , n416135 );
or ( n69445 , n69442 , n69444 );
buf ( n416138 , n68953 );
buf ( n416139 , n68940 );
nand ( n69448 , n416138 , n416139 );
buf ( n416141 , n69448 );
buf ( n416142 , n416141 );
nand ( n69451 , n69445 , n416142 );
buf ( n416144 , n69451 );
and ( n69453 , n416144 , n415668 );
not ( n69454 , n416144 );
and ( n69455 , n69454 , n415617 );
nor ( n69456 , n69453 , n69455 );
buf ( n416149 , n69456 );
not ( n69458 , n416149 );
buf ( n416151 , n69458 );
nand ( n69460 , n69440 , n416151 );
nand ( n69461 , n69437 , n69460 );
buf ( n416154 , n394817 );
not ( n69463 , n416154 );
buf ( n416156 , n54957 );
not ( n69465 , n416156 );
or ( n69466 , n69463 , n69465 );
buf ( n416159 , n49653 );
buf ( n416160 , n394814 );
nand ( n69469 , n416159 , n416160 );
buf ( n416162 , n69469 );
buf ( n416163 , n416162 );
nand ( n69472 , n69466 , n416163 );
buf ( n416165 , n69472 );
buf ( n416166 , n416165 );
not ( n69475 , n416166 );
buf ( n416168 , n399031 );
not ( n69477 , n416168 );
or ( n69478 , n69475 , n69477 );
buf ( n416171 , n415350 );
buf ( n416172 , n395469 );
nand ( n69481 , n416171 , n416172 );
buf ( n416174 , n69481 );
buf ( n416175 , n416174 );
nand ( n69484 , n69478 , n416175 );
buf ( n416177 , n69484 );
not ( n69486 , n416177 );
buf ( n416179 , n392884 );
not ( n69488 , n416179 );
buf ( n416181 , n399164 );
not ( n69490 , n416181 );
or ( n69491 , n69488 , n69490 );
buf ( n416184 , n24049 );
buf ( n416185 , n392887 );
nand ( n69494 , n416184 , n416185 );
buf ( n416187 , n69494 );
buf ( n416188 , n416187 );
nand ( n69497 , n69491 , n416188 );
buf ( n416190 , n69497 );
buf ( n416191 , n416190 );
not ( n69500 , n416191 );
buf ( n416193 , n389122 );
not ( n69502 , n416193 );
or ( n69503 , n69500 , n69502 );
buf ( n416196 , n415605 );
buf ( n416197 , n41563 );
nand ( n69506 , n416196 , n416197 );
buf ( n416199 , n69506 );
buf ( n416200 , n416199 );
nand ( n69509 , n69503 , n416200 );
buf ( n416202 , n69509 );
not ( n69511 , n416202 );
or ( n69512 , n69486 , n69511 );
buf ( n416205 , n416202 );
buf ( n416206 , n416177 );
nor ( n69515 , n416205 , n416206 );
buf ( n416208 , n69515 );
buf ( n416209 , n392611 );
not ( n69518 , n416209 );
buf ( n416211 , n51822 );
not ( n69520 , n416211 );
or ( n69521 , n69518 , n69520 );
buf ( n416214 , n24072 );
buf ( n416215 , n392620 );
nand ( n69524 , n416214 , n416215 );
buf ( n416217 , n69524 );
buf ( n416218 , n416217 );
nand ( n69527 , n69521 , n416218 );
buf ( n416220 , n69527 );
buf ( n416221 , n416220 );
not ( n69530 , n416221 );
buf ( n416223 , n390429 );
not ( n69532 , n416223 );
or ( n69533 , n69530 , n69532 );
buf ( n416226 , n67896 );
buf ( n416227 , n42924 );
nand ( n69536 , n416226 , n416227 );
buf ( n416229 , n69536 );
buf ( n416230 , n416229 );
nand ( n69539 , n69533 , n416230 );
buf ( n416232 , n69539 );
buf ( n416233 , n416232 );
buf ( n416234 , n68930 );
buf ( n416235 , n388803 );
and ( n69544 , n416234 , n416235 );
buf ( n416237 , n405736 );
not ( n69546 , n416237 );
buf ( n416239 , n406824 );
not ( n69548 , n416239 );
or ( n69549 , n69546 , n69548 );
buf ( n416242 , n406821 );
buf ( n416243 , n388754 );
nand ( n69552 , n416242 , n416243 );
buf ( n416245 , n69552 );
buf ( n416246 , n416245 );
nand ( n69555 , n69549 , n416246 );
buf ( n416248 , n69555 );
and ( n69557 , n416248 , n388740 );
buf ( n416250 , n69557 );
nor ( n69559 , n69544 , n416250 );
buf ( n416252 , n69559 );
buf ( n416253 , n416252 );
not ( n69562 , n416253 );
buf ( n416255 , n69562 );
buf ( n416256 , n416255 );
or ( n69565 , n416233 , n416256 );
and ( n69566 , n68341 , n68359 );
not ( n69567 , n68341 );
nor ( n69568 , n415069 , n68355 );
and ( n69569 , n69567 , n69568 );
nor ( n69570 , n69566 , n69569 );
and ( n69571 , n68341 , n68356 );
not ( n69572 , n68341 );
nand ( n69573 , n415069 , n68355 );
and ( n69574 , n69572 , n69573 );
or ( n69575 , n69571 , n69574 );
nand ( n69576 , n69570 , n69575 );
buf ( n416269 , n69576 );
and ( n69578 , n27320 , n62006 );
not ( n69579 , n27320 );
and ( n69580 , n69579 , n24116 );
or ( n69581 , n69578 , n69580 );
buf ( n416274 , n69581 );
not ( n69583 , n416274 );
buf ( n416276 , n45076 );
not ( n69585 , n416276 );
or ( n69586 , n69583 , n69585 );
buf ( n416279 , n415107 );
buf ( n416280 , n41664 );
nand ( n69589 , n416279 , n416280 );
buf ( n416282 , n69589 );
buf ( n416283 , n416282 );
nand ( n69592 , n69586 , n416283 );
buf ( n416285 , n69592 );
buf ( n416286 , n416285 );
xor ( n69595 , n416269 , n416286 );
buf ( n416288 , n41861 );
not ( n69597 , n416288 );
buf ( n416290 , n41365 );
not ( n69599 , n416290 );
buf ( n416292 , n69599 );
buf ( n416293 , n416292 );
not ( n69602 , n416293 );
or ( n69603 , n69597 , n69602 );
buf ( n416296 , n410407 );
not ( n69605 , n416296 );
buf ( n416298 , n69605 );
buf ( n416299 , n416298 );
buf ( n416300 , n389356 );
nand ( n69609 , n416299 , n416300 );
buf ( n416302 , n69609 );
buf ( n416303 , n416302 );
nand ( n69612 , n69603 , n416303 );
buf ( n416305 , n69612 );
buf ( n416306 , n416305 );
not ( n69615 , n416306 );
buf ( n416308 , n66128 );
not ( n69617 , n416308 );
or ( n69618 , n69615 , n69617 );
buf ( n416311 , n412976 );
buf ( n416312 , n67927 );
nand ( n69621 , n416311 , n416312 );
buf ( n416314 , n69621 );
buf ( n416315 , n416314 );
nand ( n69624 , n69618 , n416315 );
buf ( n416317 , n69624 );
buf ( n416318 , n416317 );
and ( n69627 , n69595 , n416318 );
and ( n69628 , n416269 , n416286 );
or ( n69629 , n69627 , n69628 );
buf ( n416322 , n69629 );
buf ( n416323 , n416322 );
nand ( n69632 , n69565 , n416323 );
buf ( n416325 , n69632 );
buf ( n416326 , n416325 );
buf ( n416327 , n416232 );
buf ( n416328 , n416255 );
nand ( n69637 , n416327 , n416328 );
buf ( n416330 , n69637 );
buf ( n416331 , n416330 );
and ( n69640 , n416326 , n416331 );
buf ( n416333 , n69640 );
or ( n69642 , n416208 , n416333 );
nand ( n69643 , n69512 , n69642 );
buf ( n416336 , n69643 );
buf ( n416337 , n55543 );
not ( n69646 , n416337 );
buf ( n416339 , n37346 );
not ( n69648 , n416339 );
or ( n69649 , n69646 , n69648 );
buf ( n416342 , n395478 );
buf ( n416343 , n51185 );
nand ( n69652 , n416342 , n416343 );
buf ( n416345 , n69652 );
buf ( n416346 , n416345 );
nand ( n69655 , n69649 , n416346 );
buf ( n416348 , n69655 );
buf ( n416349 , n416348 );
not ( n69658 , n416349 );
buf ( n416351 , n390536 );
not ( n416352 , n416351 );
or ( n69661 , n69658 , n416352 );
buf ( n416354 , n415460 );
buf ( n416355 , n37314 );
nand ( n69664 , n416354 , n416355 );
buf ( n416357 , n69664 );
buf ( n416358 , n416357 );
nand ( n69667 , n69661 , n416358 );
buf ( n416360 , n69667 );
buf ( n416361 , n416360 );
xor ( n69670 , n416336 , n416361 );
buf ( n416363 , n400033 );
not ( n69672 , n416363 );
buf ( n416365 , n36251 );
not ( n69674 , n416365 );
or ( n69675 , n69672 , n69674 );
buf ( n416368 , n389928 );
buf ( n416369 , n400042 );
nand ( n69678 , n416368 , n416369 );
buf ( n416371 , n69678 );
buf ( n416372 , n416371 );
nand ( n69681 , n69675 , n416372 );
buf ( n416374 , n69681 );
buf ( n416375 , n416374 );
not ( n69684 , n416375 );
buf ( n416377 , n383894 );
not ( n69686 , n416377 );
or ( n69687 , n69684 , n69686 );
buf ( n416380 , n414469 );
buf ( n416381 , n388629 );
nand ( n69690 , n416380 , n416381 );
buf ( n416383 , n69690 );
buf ( n416384 , n416383 );
nand ( n69693 , n69687 , n416384 );
buf ( n416386 , n69693 );
buf ( n416387 , n416386 );
and ( n69696 , n69670 , n416387 );
and ( n69697 , n416336 , n416361 );
or ( n69698 , n69696 , n69697 );
buf ( n416391 , n69698 );
xor ( n69700 , n69461 , n416391 );
xor ( n69701 , n415678 , n415696 );
xor ( n69702 , n69701 , n415702 );
buf ( n416395 , n69702 );
and ( n69704 , n69700 , n416395 );
and ( n69705 , n69461 , n416391 );
or ( n69706 , n69704 , n69705 );
buf ( n416399 , n69706 );
and ( n69708 , n69391 , n416399 );
and ( n69709 , n416075 , n416082 );
or ( n69710 , n69708 , n69709 );
buf ( n416403 , n69710 );
buf ( n416404 , n416403 );
xor ( n69713 , n415297 , n68752 );
xnor ( n69714 , n69713 , n68574 );
buf ( n416407 , n69714 );
xor ( n69716 , n416404 , n416407 );
xor ( n69717 , n415582 , n68846 );
xnor ( n69718 , n69717 , n415706 );
buf ( n416411 , n69718 );
not ( n69720 , n51553 );
not ( n69721 , n69375 );
or ( n69722 , n69720 , n69721 );
and ( n69723 , n38155 , n50584 );
not ( n69724 , n38155 );
and ( n69725 , n69724 , n408347 );
or ( n69726 , n69723 , n69725 );
nand ( n69727 , n69726 , n50579 );
nand ( n69728 , n69722 , n69727 );
not ( n69729 , n68743 );
and ( n69730 , n68723 , n68710 );
nand ( n69731 , n69729 , n69730 );
not ( n69732 , n68724 );
nand ( n69733 , n69732 , n68743 );
and ( n69734 , n68711 , n68722 );
nand ( n69735 , n69734 , n69729 );
nand ( n69736 , n68743 , n68722 , n68710 );
nand ( n69737 , n69731 , n69733 , n69735 , n69736 );
xor ( n69738 , n69728 , n69737 );
not ( n69739 , n68698 );
and ( n69740 , n68673 , n69739 );
not ( n69741 , n68673 );
and ( n69742 , n69741 , n68698 );
nor ( n69743 , n69740 , n69742 );
and ( n69744 , n69743 , n68618 );
not ( n69745 , n69743 );
not ( n69746 , n68618 );
and ( n69747 , n69745 , n69746 );
nor ( n69748 , n69744 , n69747 );
and ( n69749 , n69738 , n69748 );
and ( n69750 , n69728 , n69737 );
or ( n69751 , n69749 , n69750 );
buf ( n416444 , n69751 );
xor ( n69753 , n416411 , n416444 );
xor ( n69754 , n414453 , n414456 );
xor ( n69755 , n69754 , n415232 );
buf ( n416448 , n69755 );
buf ( n416449 , n416448 );
and ( n69758 , n69753 , n416449 );
and ( n69759 , n416411 , n416444 );
or ( n69760 , n69758 , n69759 );
buf ( n416453 , n69760 );
buf ( n416454 , n416453 );
and ( n69763 , n69716 , n416454 );
and ( n69764 , n416404 , n416407 );
or ( n69765 , n69763 , n69764 );
buf ( n416458 , n69765 );
and ( n69767 , n69365 , n416458 );
and ( n69768 , n69144 , n416056 );
or ( n69769 , n69767 , n69768 );
buf ( n416462 , n69769 );
buf ( n416463 , n415727 );
buf ( n416464 , n415286 );
xor ( n69773 , n416463 , n416464 );
buf ( n416466 , n415479 );
xor ( n69775 , n69773 , n416466 );
buf ( n416468 , n69775 );
buf ( n416469 , n416468 );
xor ( n69778 , n414442 , n415241 );
xor ( n69779 , n69778 , n415250 );
buf ( n416472 , n69779 );
buf ( n416473 , n416472 );
xor ( n69782 , n416469 , n416473 );
and ( n69783 , n68608 , n68747 );
not ( n69784 , n68608 );
not ( n69785 , n68747 );
and ( n69786 , n69784 , n69785 );
nor ( n69787 , n69783 , n69786 );
not ( n69788 , n68750 );
and ( n69789 , n69787 , n69788 );
not ( n69790 , n69787 );
and ( n69791 , n69790 , n68750 );
nor ( n69792 , n69789 , n69791 );
buf ( n416485 , n69792 );
not ( n69799 , n45893 );
buf ( n416487 , C0 );
buf ( n416488 , n416487 );
xor ( n69815 , n416485 , n416488 );
buf ( n416490 , n67890 );
not ( n69834 , n416490 );
buf ( n416492 , n414481 );
not ( n69836 , n416492 );
or ( n69837 , n69834 , n69836 );
buf ( n416495 , n414481 );
buf ( n416496 , n67890 );
or ( n69840 , n416495 , n416496 );
nand ( n69841 , n69837 , n69840 );
buf ( n416499 , n69841 );
xor ( n69843 , n415221 , n416499 );
nor ( n69844 , C0 , n69843 );
buf ( n416502 , n395362 );
not ( n69846 , n416502 );
buf ( n416504 , n69205 );
not ( n69848 , n416504 );
or ( n69849 , n69846 , n69848 );
and ( n69850 , n47863 , n388931 );
not ( n69851 , n47863 );
and ( n69852 , n69851 , n388922 );
or ( n69853 , n69850 , n69852 );
buf ( n416511 , n69853 );
buf ( n416512 , n395349 );
nand ( n69856 , n416511 , n416512 );
buf ( n416514 , n69856 );
buf ( n416515 , n416514 );
nand ( n69859 , n69849 , n416515 );
buf ( n416517 , n69859 );
buf ( n416518 , n416517 );
not ( n69862 , n416518 );
buf ( n416520 , n69862 );
buf ( n416521 , n416520 );
not ( n69865 , n416521 );
buf ( n416523 , n384008 );
not ( n69867 , n416523 );
buf ( n416525 , n402819 );
buf ( n416526 , n40824 );
and ( n69870 , n416525 , n416526 );
not ( n69871 , n416525 );
buf ( n416529 , n36398 );
and ( n69873 , n69871 , n416529 );
nor ( n69874 , n69870 , n69873 );
buf ( n416532 , n69874 );
buf ( n416533 , n416532 );
not ( n69877 , n416533 );
and ( n69878 , n69867 , n69877 );
not ( n69879 , n415879 );
nor ( n69880 , n69879 , n383943 );
buf ( n416538 , n69880 );
nor ( n69882 , n69878 , n416538 );
buf ( n416540 , n69882 );
buf ( n416541 , n416540 );
not ( n69885 , n416541 );
or ( n69886 , n69865 , n69885 );
buf ( n416544 , n36363 );
buf ( n416545 , n358975 );
nand ( n69889 , n416544 , n416545 );
buf ( n416547 , n69889 );
not ( n69891 , n416547 );
buf ( n416549 , n397489 );
not ( n69893 , n416549 );
buf ( n416551 , n388965 );
not ( n69895 , n416551 );
or ( n69896 , n69893 , n69895 );
buf ( n416554 , n388962 );
buf ( n416555 , n397492 );
nand ( n69899 , n416554 , n416555 );
buf ( n416557 , n69899 );
buf ( n416558 , n416557 );
nand ( n69902 , n69896 , n416558 );
buf ( n416560 , n69902 );
buf ( n416561 , n416560 );
not ( n69905 , n416561 );
buf ( n416563 , n46056 );
not ( n69907 , n416563 );
or ( n69908 , n69905 , n69907 );
buf ( n416566 , n415166 );
buf ( n416567 , n51692 );
nand ( n69911 , n416566 , n416567 );
buf ( n416569 , n69911 );
buf ( n416570 , n416569 );
nand ( n69914 , n69908 , n416570 );
buf ( n416572 , n69914 );
nor ( n69916 , n69891 , n416572 );
not ( n69917 , n68419 );
not ( n69918 , n67916 );
not ( n69919 , n414633 );
or ( n69920 , n69918 , n69919 );
nand ( n69921 , n67915 , n414636 );
nand ( n69922 , n69920 , n69921 );
not ( n69923 , n69922 );
or ( n69924 , n69917 , n69923 );
not ( n69925 , n67916 );
not ( n69926 , n414633 );
or ( n69927 , n69925 , n69926 );
nand ( n69928 , n69927 , n69921 );
or ( n69929 , n68419 , n69928 );
nand ( n69930 , n69924 , n69929 );
or ( n69931 , n69916 , n69930 );
not ( n69932 , n416547 );
nand ( n69933 , n69932 , n416572 );
nand ( n69934 , n69931 , n69933 );
buf ( n416592 , n69934 );
nand ( n69936 , n69886 , n416592 );
buf ( n416594 , n69936 );
buf ( n416595 , n416594 );
buf ( n416596 , n416540 );
not ( n69940 , n416596 );
buf ( n416598 , n69940 );
buf ( n416599 , n416598 );
buf ( n416600 , n416517 );
nand ( n69944 , n416599 , n416600 );
buf ( n416602 , n69944 );
buf ( n416603 , n416602 );
nand ( n69947 , n416595 , n416603 );
buf ( n416605 , n69947 );
not ( n69949 , n416605 );
or ( n69950 , n69844 , n69949 );
nand ( n69952 , n69950 , C1 );
buf ( n416609 , n69952 );
and ( n69954 , n69815 , n416609 );
or ( n69956 , n69954 , C0 );
buf ( n416612 , n69956 );
buf ( n416613 , n416612 );
xor ( n69959 , n414445 , n414447 );
not ( n69960 , n415236 );
xor ( n69961 , n69959 , n69960 );
buf ( n416617 , n69961 );
xor ( n69963 , n416613 , n416617 );
xor ( n69964 , n415864 , n415866 );
xor ( n69965 , n69964 , n416027 );
buf ( n416621 , n69965 );
buf ( n416622 , n416621 );
buf ( n416623 , C0 );
buf ( n416624 , n416623 );
xor ( n69993 , n415892 , n415909 );
xor ( n69994 , n69993 , n416022 );
buf ( n416627 , n69994 );
buf ( n416628 , n416627 );
xor ( n69997 , n416624 , n416628 );
xor ( n69998 , n415154 , n415179 );
xor ( n69999 , n69998 , n415217 );
buf ( n416632 , n69999 );
buf ( n416633 , n416632 );
not ( n70002 , n416633 );
buf ( n416635 , n49117 );
not ( n70004 , n416635 );
buf ( n416637 , n49661 );
not ( n70006 , n416637 );
or ( n70007 , n70004 , n70006 );
buf ( n416640 , n49653 );
buf ( n416641 , n67126 );
nand ( n70010 , n416640 , n416641 );
buf ( n416643 , n70010 );
buf ( n416644 , n416643 );
nand ( n70013 , n70007 , n416644 );
buf ( n416646 , n70013 );
buf ( n416647 , n416646 );
not ( n70016 , n416647 );
buf ( n416649 , n397102 );
not ( n70018 , n416649 );
or ( n70019 , n70016 , n70018 );
buf ( n416652 , n416165 );
buf ( n416653 , n386477 );
nand ( n70022 , n416652 , n416653 );
buf ( n416655 , n70022 );
buf ( n416656 , n416655 );
nand ( n70025 , n70019 , n416656 );
buf ( n416658 , n70025 );
buf ( n416659 , n416658 );
not ( n70028 , n416659 );
buf ( n416661 , n70028 );
buf ( n416662 , n416661 );
not ( n70031 , n416662 );
buf ( n416664 , n41407 );
not ( n70033 , n416664 );
buf ( n416666 , n383863 );
nand ( n70035 , n70033 , n416666 );
buf ( n416668 , n70035 );
and ( n70037 , n416668 , n358975 );
and ( n70038 , n393117 , n36312 );
nor ( n70039 , n70037 , n70038 );
nand ( n70040 , n388608 , n70039 );
buf ( n416673 , n70040 );
not ( n70042 , n416673 );
or ( n70043 , n70031 , n70042 );
buf ( n416676 , n43515 );
not ( n70045 , n416676 );
buf ( n416678 , n69285 );
not ( n70047 , n416678 );
or ( n70048 , n70045 , n70047 );
buf ( n416681 , n411504 );
not ( n70050 , n416681 );
buf ( n416683 , n389856 );
not ( n70052 , n416683 );
or ( n70053 , n70050 , n70052 );
buf ( n416686 , n49686 );
buf ( n416687 , n391024 );
nand ( n70056 , n416686 , n416687 );
buf ( n416689 , n70056 );
buf ( n416690 , n416689 );
nand ( n70059 , n70053 , n416690 );
buf ( n416692 , n70059 );
buf ( n416693 , n416692 );
buf ( n416694 , n43536 );
nand ( n70063 , n416693 , n416694 );
buf ( n416696 , n70063 );
buf ( n416697 , n416696 );
nand ( n70066 , n70048 , n416697 );
buf ( n416699 , n70066 );
buf ( n416700 , n416699 );
nand ( n70069 , n70043 , n416700 );
buf ( n416702 , n70069 );
buf ( n416703 , n416702 );
buf ( n416704 , n70040 );
not ( n70073 , n416704 );
buf ( n416706 , n416658 );
nand ( n70075 , n70073 , n416706 );
buf ( n416708 , n70075 );
buf ( n416709 , n416708 );
nand ( n70078 , n416703 , n416709 );
buf ( n416711 , n70078 );
buf ( n416712 , n416711 );
buf ( n416713 , n69307 );
buf ( n416714 , n69310 );
xor ( n70083 , n416713 , n416714 );
buf ( n416716 , n69287 );
xor ( n70085 , n70083 , n416716 );
buf ( n416718 , n70085 );
buf ( n416719 , n416718 );
xor ( n70088 , n416712 , n416719 );
not ( n70089 , n395349 );
and ( n70090 , n47863 , n390271 );
not ( n70091 , n47863 );
and ( n70092 , n70091 , n386147 );
or ( n70093 , n70090 , n70092 );
not ( n70094 , n70093 );
or ( n70095 , n70089 , n70094 );
buf ( n416728 , n69853 );
buf ( n416729 , n395362 );
nand ( n70098 , n416728 , n416729 );
buf ( n416731 , n70098 );
nand ( n70100 , n70095 , n416731 );
buf ( n416733 , n70100 );
and ( n70102 , n70088 , n416733 );
and ( n70103 , n416712 , n416719 );
or ( n70104 , n70102 , n70103 );
buf ( n416737 , n70104 );
buf ( n416738 , n416737 );
not ( n70107 , n416738 );
or ( n70108 , n70002 , n70107 );
buf ( n416741 , n416737 );
buf ( n416742 , n416632 );
or ( n70111 , n416741 , n416742 );
xor ( n70112 , n68336 , n415050 );
xnor ( n70113 , n70112 , n68179 );
not ( n70114 , n70113 );
buf ( n416747 , n42066 );
not ( n70116 , n416747 );
buf ( n416749 , n68376 );
not ( n70118 , n416749 );
or ( n70119 , n70116 , n70118 );
buf ( n416752 , n24116 );
buf ( n416753 , n43144 );
nand ( n70122 , n416752 , n416753 );
buf ( n416755 , n70122 );
buf ( n416756 , n416755 );
nand ( n70125 , n70119 , n416756 );
buf ( n416758 , n70125 );
not ( n70127 , n416758 );
buf ( n416760 , n41709 );
not ( n70129 , n416760 );
buf ( n416762 , n70129 );
not ( n70131 , n416762 );
or ( n70132 , n70127 , n70131 );
buf ( n416765 , n69581 );
buf ( n416766 , n41664 );
nand ( n70135 , n416765 , n416766 );
buf ( n416768 , n70135 );
nand ( n70137 , n70132 , n416768 );
not ( n70138 , n70137 );
or ( n70139 , n70114 , n70138 );
not ( n70140 , n70113 );
not ( n70141 , n70140 );
not ( n70142 , n70137 );
not ( n70143 , n70142 );
or ( n70144 , n70141 , n70143 );
xor ( n70145 , n415019 , n415023 );
xor ( n70146 , n70145 , n415046 );
buf ( n416779 , n70146 );
xor ( n70148 , n413367 , n413383 );
xor ( n70149 , n70148 , n413386 );
xor ( n70150 , n68308 , n415038 );
xor ( n70151 , n70149 , n70150 );
buf ( n416784 , n62467 );
buf ( n416785 , n405215 );
and ( n70154 , n416784 , n416785 );
buf ( n416787 , n409468 );
buf ( n416788 , n58061 );
and ( n70157 , n416787 , n416788 );
nor ( n70158 , n70154 , n70157 );
buf ( n416791 , n70158 );
buf ( n416792 , n416791 );
buf ( n416793 , n403293 );
or ( n70162 , n416792 , n416793 );
buf ( n416795 , n414831 );
buf ( n416796 , n405476 );
or ( n70165 , n416795 , n416796 );
nand ( n70166 , n70162 , n70165 );
buf ( n416799 , n70166 );
buf ( n416800 , n416799 );
buf ( n416801 , n414714 );
buf ( n416802 , n401692 );
or ( n70171 , n416801 , n416802 );
buf ( n416804 , n67987 );
buf ( n416805 , n401689 );
or ( n70174 , n416804 , n416805 );
nand ( n70175 , n70171 , n70174 );
buf ( n416808 , n70175 );
buf ( n416809 , n416808 );
not ( n70178 , n416809 );
buf ( n416811 , n70178 );
buf ( n416812 , n416811 );
buf ( n416813 , n403158 );
or ( n70182 , n416812 , n416813 );
buf ( n416815 , n414751 );
buf ( n416816 , n403167 );
or ( n70185 , n416815 , n416816 );
nand ( n70186 , n70182 , n70185 );
buf ( n416819 , n70186 );
buf ( n416820 , n416819 );
nand ( n70189 , n54088 , n54224 );
not ( n70190 , n54110 );
not ( n70191 , n54219 );
or ( n70192 , n70190 , n70191 );
not ( n70193 , n54222 );
nand ( n70194 , n70192 , n70193 );
xnor ( n70195 , n70189 , n70194 );
buf ( n416828 , n70195 );
not ( n70197 , n416828 );
buf ( n416830 , n70197 );
buf ( n416831 , n416830 );
buf ( n416832 , n401623 );
or ( n70201 , n416831 , n416832 );
buf ( n416834 , n414729 );
buf ( n416835 , n403092 );
or ( n70204 , n416834 , n416835 );
nand ( n70205 , n70201 , n70204 );
buf ( n416838 , n70205 );
buf ( n416839 , n416838 );
xor ( n70208 , n416820 , n416839 );
and ( n70209 , n70193 , n54110 );
xor ( n70210 , n70209 , n54219 );
buf ( n416843 , n70210 );
not ( n70212 , n416843 );
buf ( n416845 , n70212 );
buf ( n416846 , n416845 );
buf ( n416847 , n403083 );
or ( n70216 , n416846 , n416847 );
buf ( n416849 , n416830 );
buf ( n416850 , n403092 );
or ( n70219 , n416849 , n416850 );
nand ( n70220 , n70216 , n70219 );
buf ( n416853 , n70220 );
buf ( n416854 , n416853 );
buf ( n416855 , n403164 );
not ( n70224 , n416855 );
buf ( n416857 , n416808 );
not ( n70226 , n416857 );
or ( n70227 , n70224 , n70226 );
buf ( n416860 , n401689 );
buf ( n416861 , n68002 );
and ( n70230 , n416860 , n416861 );
not ( n70231 , n416860 );
buf ( n416864 , n414729 );
and ( n70233 , n70231 , n416864 );
nor ( n70234 , n70230 , n70233 );
buf ( n416867 , n70234 );
buf ( n416868 , n416867 );
buf ( n416869 , n403158 );
or ( n70238 , n416868 , n416869 );
nand ( n70239 , n70227 , n70238 );
buf ( n416872 , n70239 );
buf ( n416873 , n416872 );
and ( n70242 , n416854 , n416873 );
buf ( n416875 , n70242 );
buf ( n416876 , n416875 );
and ( n70245 , n70208 , n416876 );
and ( n70246 , n416820 , n416839 );
or ( n70247 , n70245 , n70246 );
buf ( n416880 , n70247 );
buf ( n416881 , n416880 );
xor ( n70250 , n416800 , n416881 );
buf ( n416883 , n59435 );
buf ( n416884 , n59628 );
and ( n70253 , n416883 , n416884 );
buf ( n416886 , n406565 );
buf ( n416887 , n59457 );
and ( n70256 , n416886 , n416887 );
nor ( n70257 , n70253 , n70256 );
buf ( n416890 , n70257 );
or ( n70259 , n416890 , n59637 );
or ( n70260 , n68183 , n59467 );
nand ( n70261 , n70259 , n70260 );
buf ( n416894 , n70261 );
and ( n70263 , n70250 , n416894 );
and ( n70264 , n416800 , n416881 );
or ( n70265 , n70263 , n70264 );
buf ( n416898 , n70265 );
buf ( n416899 , n416898 );
xor ( n70268 , n414840 , n414857 );
xor ( n70269 , n70268 , n414883 );
buf ( n416902 , n70269 );
buf ( n416903 , n416902 );
xor ( n70272 , n416899 , n416903 );
xor ( n70273 , n68189 , n414916 );
xor ( n70274 , n70273 , n68209 );
buf ( n416907 , n70274 );
and ( n70276 , n70272 , n416907 );
and ( n70277 , n416899 , n416903 );
or ( n70278 , n70276 , n70277 );
buf ( n416911 , n70278 );
xor ( n70280 , n70151 , n416911 );
xor ( n70281 , n414937 , n415009 );
xor ( n70282 , n70281 , n415014 );
buf ( n416915 , n70282 );
and ( n70284 , n70280 , n416915 );
and ( n70285 , n70151 , n416911 );
or ( n70286 , n70284 , n70285 );
or ( n70287 , n416779 , n70286 );
not ( n70288 , n70287 );
xor ( n70289 , n414962 , n414979 );
xor ( n70290 , n70289 , n414999 );
buf ( n416923 , n70290 );
not ( n70292 , n409185 );
not ( n70293 , n68218 );
or ( n70294 , n70292 , n70293 );
buf ( n416927 , n58200 );
buf ( n416928 , n62177 );
and ( n70297 , n416927 , n416928 );
buf ( n416930 , n58201 );
buf ( n416931 , n62159 );
and ( n70300 , n416930 , n416931 );
nor ( n70301 , n70297 , n70300 );
buf ( n416934 , n70301 );
not ( n70303 , n416934 );
nand ( n70304 , n70303 , n409173 );
nand ( n70305 , n70294 , n70304 );
xor ( n70306 , n416923 , n70305 );
buf ( n416939 , n59596 );
buf ( n416940 , n59628 );
and ( n70309 , n416939 , n416940 );
buf ( n416942 , n409146 );
buf ( n416943 , n59457 );
and ( n70312 , n416942 , n416943 );
nor ( n70313 , n70309 , n70312 );
buf ( n416946 , n70313 );
buf ( n416947 , n416946 );
buf ( n416948 , n59637 );
or ( n70317 , n416947 , n416948 );
buf ( n416950 , n416890 );
buf ( n416951 , n59467 );
or ( n70320 , n416950 , n416951 );
nand ( n70321 , n70317 , n70320 );
buf ( n416954 , n70321 );
buf ( n416955 , n416954 );
buf ( n416956 , n62278 );
buf ( n416957 , n405391 );
and ( n70326 , n416956 , n416957 );
buf ( n416959 , n409474 );
buf ( n416960 , n414664 );
and ( n70329 , n416959 , n416960 );
nor ( n70330 , n70326 , n70329 );
buf ( n416963 , n70330 );
buf ( n416964 , n416963 );
buf ( n416965 , n405407 );
or ( n70334 , n416964 , n416965 );
buf ( n416967 , n414993 );
buf ( n416968 , n405384 );
or ( n70337 , n416967 , n416968 );
nand ( n70338 , n70334 , n70337 );
buf ( n416971 , n70338 );
buf ( n416972 , n416971 );
xor ( n70341 , n416955 , n416972 );
xor ( n70342 , n416854 , n416873 );
buf ( n416975 , n70342 );
buf ( n416976 , n416975 );
buf ( n416977 , n66359 );
buf ( n416978 , n55905 );
and ( n70347 , n416977 , n416978 );
buf ( n416980 , n413187 );
buf ( n416981 , n55895 );
and ( n70350 , n416980 , n416981 );
nor ( n70351 , n70347 , n70350 );
buf ( n416984 , n70351 );
buf ( n416985 , n416984 );
buf ( n416986 , n403120 );
or ( n70355 , n416985 , n416986 );
buf ( n416988 , n66270 );
buf ( n416989 , n55905 );
and ( n70358 , n416988 , n416989 );
buf ( n416991 , n413098 );
buf ( n416992 , n55895 );
and ( n70361 , n416991 , n416992 );
nor ( n70362 , n70358 , n70361 );
buf ( n416995 , n70362 );
buf ( n416996 , n416995 );
buf ( n416997 , n403133 );
or ( n70366 , n416996 , n416997 );
nand ( n70367 , n70355 , n70366 );
buf ( n417000 , n70367 );
buf ( n417001 , n417000 );
xor ( n70370 , n416976 , n417001 );
buf ( n417003 , n70195 );
buf ( n417004 , n401689 );
and ( n70373 , n417003 , n417004 );
buf ( n417006 , n416830 );
buf ( n417007 , n401692 );
and ( n70376 , n417006 , n417007 );
nor ( n70377 , n70373 , n70376 );
buf ( n417010 , n70377 );
buf ( n417011 , n417010 );
buf ( n417012 , n403158 );
or ( n70381 , n417011 , n417012 );
buf ( n417014 , n416867 );
buf ( n417015 , n403167 );
or ( n70384 , n417014 , n417015 );
nand ( n70385 , n70381 , n70384 );
buf ( n417018 , n70385 );
buf ( n417019 , n417018 );
and ( n70388 , n54218 , n54136 );
xor ( n70389 , n70388 , n54214 );
buf ( n417022 , n70389 );
not ( n70391 , n417022 );
buf ( n417024 , n70391 );
buf ( n417025 , n417024 );
buf ( n417026 , n403083 );
or ( n70395 , n417025 , n417026 );
buf ( n417028 , n416845 );
buf ( n417029 , n403092 );
or ( n70398 , n417028 , n417029 );
nand ( n70399 , n70395 , n70398 );
buf ( n417032 , n70399 );
buf ( n417033 , n417032 );
xor ( n70402 , n417019 , n417033 );
buf ( n417035 , n403123 );
not ( n70404 , n417035 );
buf ( n417037 , n67987 );
buf ( n417038 , n55905 );
and ( n70407 , n417037 , n417038 );
buf ( n417040 , n414714 );
buf ( n417041 , n55895 );
and ( n70410 , n417040 , n417041 );
nor ( n70411 , n70407 , n70410 );
buf ( n417044 , n70411 );
buf ( n417045 , n417044 );
not ( n70414 , n417045 );
buf ( n417047 , n70414 );
buf ( n417048 , n417047 );
not ( n70417 , n417048 );
or ( n70418 , n70404 , n70417 );
buf ( n417051 , n416984 );
buf ( n417052 , n403133 );
or ( n70421 , n417051 , n417052 );
nand ( n70422 , n70418 , n70421 );
buf ( n417055 , n70422 );
buf ( n417056 , n417055 );
and ( n70425 , n70402 , n417056 );
and ( n70426 , n417019 , n417033 );
or ( n70427 , n70425 , n70426 );
buf ( n417060 , n70427 );
buf ( n417061 , n417060 );
and ( n70430 , n70370 , n417061 );
and ( n70431 , n416976 , n417001 );
or ( n70432 , n70430 , n70431 );
buf ( n417065 , n70432 );
buf ( n417066 , n417065 );
and ( n70435 , n70341 , n417066 );
and ( n70436 , n416955 , n416972 );
or ( n70437 , n70435 , n70436 );
buf ( n417070 , n70437 );
and ( n70439 , n70306 , n417070 );
and ( n70440 , n416923 , n70305 );
or ( n70441 , n70439 , n70440 );
buf ( n417074 , n70441 );
buf ( n417075 , n55846 );
buf ( n417076 , n66411 );
and ( n70445 , n417075 , n417076 );
buf ( n417078 , n403079 );
buf ( n417079 , n62496 );
and ( n70448 , n417078 , n417079 );
nor ( n70449 , n70445 , n70448 );
buf ( n417082 , n70449 );
buf ( n417083 , n417082 );
buf ( n417084 , n410724 );
or ( n70453 , n417083 , n417084 );
buf ( n417086 , n414953 );
buf ( n417087 , n410721 );
or ( n70456 , n417086 , n417087 );
nand ( n70457 , n70453 , n70456 );
buf ( n417090 , n70457 );
buf ( n417091 , n417090 );
buf ( n417092 , n63564 );
buf ( n417093 , n405215 );
and ( n70462 , n417092 , n417093 );
buf ( n417095 , n413073 );
buf ( n417096 , n58061 );
and ( n70465 , n417095 , n417096 );
nor ( n70466 , n70462 , n70465 );
buf ( n417099 , n70466 );
buf ( n417100 , n417099 );
buf ( n417101 , n403293 );
or ( n70470 , n417100 , n417101 );
buf ( n417103 , n416791 );
buf ( n417104 , n405476 );
or ( n70473 , n417103 , n417104 );
nand ( n70474 , n70470 , n70473 );
buf ( n417107 , n70474 );
buf ( n417108 , n417107 );
buf ( n417109 , n416995 );
buf ( n417110 , n403120 );
or ( n70479 , n417109 , n417110 );
buf ( n417112 , n414970 );
buf ( n417113 , n403133 );
or ( n70482 , n417112 , n417113 );
nand ( n70483 , n70479 , n70482 );
buf ( n417116 , n70483 );
buf ( n417117 , n417116 );
xor ( n70486 , n417108 , n417117 );
xor ( n70487 , n416820 , n416839 );
xor ( n70488 , n70487 , n416876 );
buf ( n417121 , n70488 );
buf ( n417122 , n417121 );
and ( n70491 , n70486 , n417122 );
and ( n70492 , n417108 , n417117 );
or ( n70493 , n70491 , n70492 );
buf ( n417126 , n70493 );
buf ( n417127 , n417126 );
xor ( n70496 , n417091 , n417127 );
buf ( n417129 , n409507 );
not ( n70498 , n417129 );
buf ( n417131 , n58090 );
buf ( n417132 , n63625 );
and ( n70501 , n417131 , n417132 );
buf ( n417134 , n405335 );
buf ( n417135 , n63629 );
and ( n70504 , n417134 , n417135 );
nor ( n70505 , n70501 , n70504 );
buf ( n417138 , n70505 );
buf ( n417139 , n417138 );
not ( n70508 , n417139 );
buf ( n417141 , n70508 );
buf ( n417142 , n417141 );
not ( n70511 , n417142 );
or ( n70512 , n70498 , n70511 );
buf ( n417145 , n414926 );
buf ( n417146 , n409504 );
or ( n70515 , n417145 , n417146 );
nand ( n70516 , n70512 , n70515 );
buf ( n417149 , n70516 );
buf ( n417150 , n417149 );
and ( n70519 , n70496 , n417150 );
and ( n70520 , n417091 , n417127 );
or ( n70521 , n70519 , n70520 );
buf ( n417154 , n70521 );
buf ( n417155 , n417154 );
xor ( n70524 , n417074 , n417155 );
xor ( n70525 , n414945 , n414958 );
xor ( n70526 , n70525 , n415004 );
buf ( n417159 , n70526 );
buf ( n417160 , n417159 );
and ( n70529 , n70524 , n417160 );
and ( n70530 , n417074 , n417155 );
or ( n70531 , n70529 , n70530 );
buf ( n417164 , n70531 );
xor ( n70533 , n70151 , n416911 );
xor ( n70534 , n70533 , n416915 );
and ( n70535 , n417164 , n70534 );
or ( n70536 , n417082 , n410721 );
not ( n70537 , n410724 );
and ( n70538 , n58135 , n62495 );
and ( n70539 , n55984 , n62496 );
nor ( n70540 , n70538 , n70539 );
nand ( n70541 , n70537 , n70540 );
nand ( n70542 , n70536 , n70541 );
buf ( n417175 , n70542 );
buf ( n417176 , n58352 );
buf ( n417177 , n62177 );
and ( n70546 , n417176 , n417177 );
buf ( n417179 , n406571 );
buf ( n417180 , n62159 );
and ( n70549 , n417179 , n417180 );
nor ( n70550 , n70546 , n70549 );
buf ( n417183 , n70550 );
buf ( n417184 , n417183 );
buf ( n417185 , n409429 );
or ( n70554 , n417184 , n417185 );
buf ( n417187 , n416934 );
buf ( n417188 , n409170 );
or ( n70557 , n417187 , n417188 );
nand ( n70558 , n70554 , n70557 );
buf ( n417191 , n70558 );
buf ( n417192 , n417191 );
xor ( n70561 , n417175 , n417192 );
xor ( n70562 , n417108 , n417117 );
xor ( n70563 , n70562 , n417122 );
buf ( n417196 , n70563 );
buf ( n417197 , n417196 );
and ( n70566 , n70561 , n417197 );
and ( n70567 , n417175 , n417192 );
or ( n70568 , n70566 , n70567 );
buf ( n417201 , n70568 );
buf ( n417202 , n417201 );
xor ( n70571 , n416800 , n416881 );
xor ( n70572 , n70571 , n416894 );
buf ( n417205 , n70572 );
buf ( n417206 , n417205 );
xor ( n70575 , n417202 , n417206 );
xor ( n70576 , n417091 , n417127 );
xor ( n70577 , n70576 , n417150 );
buf ( n417210 , n70577 );
buf ( n417211 , n417210 );
and ( n70580 , n70575 , n417211 );
and ( n70581 , n417202 , n417206 );
or ( n70582 , n70580 , n70581 );
buf ( n417215 , n70582 );
xor ( n70584 , n416899 , n416903 );
xor ( n70585 , n70584 , n416907 );
buf ( n417218 , n70585 );
xor ( n70587 , n417215 , n417218 );
xor ( n70588 , n417074 , n417155 );
xor ( n70589 , n70588 , n417160 );
buf ( n417222 , n70589 );
and ( n70591 , n70587 , n417222 );
and ( n70592 , n417215 , n417218 );
or ( n70593 , n70591 , n70592 );
xor ( n70594 , n70151 , n416911 );
xor ( n70595 , n70594 , n416915 );
and ( n70596 , n70593 , n70595 );
and ( n70597 , n417164 , n70593 );
or ( n70598 , n70535 , n70596 , n70597 );
not ( n70599 , n70598 );
or ( n70600 , n70288 , n70599 );
nand ( n70601 , n416779 , n70286 );
nand ( n70602 , n70600 , n70601 );
nand ( n70603 , n70144 , n70602 );
nand ( n70604 , n70139 , n70603 );
buf ( n417237 , n70604 );
buf ( n417238 , n388803 );
not ( n70607 , n417238 );
buf ( n417240 , n416248 );
not ( n70609 , n417240 );
or ( n70610 , n70607 , n70609 );
and ( n70611 , n12480 , n388754 );
not ( n70612 , n12480 );
and ( n70613 , n70612 , n405736 );
or ( n70614 , n70611 , n70613 );
buf ( n417247 , n70614 );
buf ( n417248 , n388740 );
nand ( n70617 , n417247 , n417248 );
buf ( n417250 , n70617 );
buf ( n417251 , n417250 );
nand ( n70620 , n70610 , n417251 );
buf ( n417253 , n70620 );
buf ( n417254 , n417253 );
xor ( n70623 , n417237 , n417254 );
not ( n70624 , n391446 );
not ( n70625 , n40653 );
or ( n70626 , n70624 , n70625 );
buf ( n417259 , n407936 );
buf ( n417260 , n391443 );
nand ( n70629 , n417259 , n417260 );
buf ( n417262 , n70629 );
nand ( n70631 , n70626 , n417262 );
not ( n70632 , n70631 );
not ( n70633 , n60872 );
or ( n70634 , n70632 , n70633 );
buf ( n417267 , n415124 );
not ( n70636 , n417267 );
buf ( n417269 , n47726 );
nand ( n70638 , n70636 , n417269 );
buf ( n417271 , n70638 );
nand ( n70640 , n70634 , n417271 );
buf ( n417273 , n70640 );
and ( n70642 , n70623 , n417273 );
and ( n70643 , n417237 , n417254 );
or ( n70644 , n70642 , n70643 );
buf ( n417277 , n70644 );
buf ( n417278 , n417277 );
buf ( n417279 , n390362 );
not ( n70648 , n417279 );
buf ( n417281 , n415995 );
not ( n70650 , n417281 );
or ( n70651 , n70648 , n70650 );
and ( n70652 , n28644 , n40600 );
not ( n70653 , n28644 );
and ( n70654 , n70653 , n40601 );
or ( n70655 , n70652 , n70654 );
buf ( n417288 , n70655 );
buf ( n417289 , n40592 );
nand ( n70658 , n417288 , n417289 );
buf ( n417291 , n70658 );
buf ( n417292 , n417291 );
nand ( n70661 , n70651 , n417292 );
buf ( n417294 , n70661 );
buf ( n417295 , n417294 );
xor ( n70664 , n417278 , n417295 );
xor ( n70665 , n416269 , n416286 );
xor ( n70666 , n70665 , n416318 );
buf ( n417299 , n70666 );
buf ( n417300 , n417299 );
buf ( n417301 , n390362 );
not ( n70670 , n417301 );
buf ( n417303 , n70655 );
not ( n70672 , n417303 );
or ( n70673 , n70670 , n70672 );
buf ( n417306 , n40601 );
not ( n70675 , n417306 );
buf ( n417308 , n410400 );
not ( n70677 , n417308 );
or ( n70678 , n70675 , n70677 );
buf ( n417311 , n12471 );
buf ( n417312 , n40600 );
nand ( n70681 , n417311 , n417312 );
buf ( n417314 , n70681 );
buf ( n417315 , n417314 );
nand ( n70684 , n70678 , n417315 );
buf ( n417317 , n70684 );
buf ( n417318 , n417317 );
buf ( n417319 , n40592 );
nand ( n70688 , n417318 , n417319 );
buf ( n417321 , n70688 );
buf ( n417322 , n417321 );
nand ( n70691 , n70673 , n417322 );
buf ( n417324 , n70691 );
buf ( n417325 , n417324 );
xor ( n70694 , n417300 , n417325 );
not ( n70695 , n70140 );
not ( n70696 , n70602 );
or ( n70697 , n70695 , n70696 );
or ( n70698 , n70602 , n70140 );
nand ( n70699 , n70697 , n70698 );
and ( n70700 , n70137 , n70699 );
not ( n70701 , n70137 );
buf ( n417334 , n70699 );
not ( n70703 , n417334 );
buf ( n417336 , n70703 );
and ( n70705 , n70701 , n417336 );
nor ( n70706 , n70700 , n70705 );
buf ( n417339 , n70706 );
buf ( n417340 , n388803 );
not ( n70709 , n417340 );
buf ( n417342 , n70614 );
not ( n70711 , n417342 );
or ( n70712 , n70709 , n70711 );
buf ( n417345 , n405736 );
not ( n70714 , n417345 );
buf ( n417347 , n28353 );
not ( n70716 , n417347 );
buf ( n417349 , n70716 );
buf ( n417350 , n417349 );
not ( n70719 , n417350 );
or ( n70720 , n70714 , n70719 );
buf ( n417353 , n28353 );
buf ( n417354 , n388754 );
nand ( n70723 , n417353 , n417354 );
buf ( n417356 , n70723 );
buf ( n417357 , n417356 );
nand ( n70726 , n70720 , n417357 );
buf ( n417359 , n70726 );
buf ( n417360 , n417359 );
buf ( n417361 , n388740 );
nand ( n70730 , n417360 , n417361 );
buf ( n417363 , n70730 );
buf ( n417364 , n417363 );
nand ( n70733 , n70712 , n417364 );
buf ( n417366 , n70733 );
buf ( n417367 , n417366 );
xor ( n70736 , n417339 , n417367 );
buf ( n417369 , n389341 );
not ( n70738 , n417369 );
buf ( n417371 , n416292 );
not ( n70740 , n417371 );
or ( n70741 , n70738 , n70740 );
buf ( n417374 , n393185 );
buf ( n417375 , n416298 );
nand ( n70744 , n417374 , n417375 );
buf ( n417377 , n70744 );
buf ( n417378 , n417377 );
nand ( n70747 , n70741 , n417378 );
buf ( n417380 , n70747 );
buf ( n417381 , n417380 );
not ( n70750 , n417381 );
buf ( n417383 , n66128 );
not ( n70752 , n417383 );
or ( n70753 , n70750 , n70752 );
buf ( n417386 , n416305 );
buf ( n417387 , n412976 );
nand ( n70756 , n417386 , n417387 );
buf ( n417389 , n70756 );
buf ( n417390 , n417389 );
nand ( n70759 , n70753 , n417390 );
buf ( n417392 , n70759 );
buf ( n417393 , n417392 );
and ( n70762 , n70736 , n417393 );
and ( n70763 , n417339 , n417367 );
or ( n70764 , n70762 , n70763 );
buf ( n417397 , n70764 );
buf ( n417398 , n417397 );
and ( n70767 , n70694 , n417398 );
and ( n70768 , n417300 , n417325 );
or ( n70769 , n70767 , n70768 );
buf ( n417402 , n70769 );
buf ( n417403 , n417402 );
and ( n70772 , n70664 , n417403 );
and ( n70773 , n417278 , n417295 );
or ( n70774 , n70772 , n70773 );
buf ( n417407 , n70774 );
buf ( n417408 , n417407 );
buf ( n417409 , n45260 );
not ( n70778 , n417409 );
buf ( n417411 , n64136 );
not ( n70780 , n417411 );
buf ( n417413 , n388409 );
not ( n70782 , n417413 );
or ( n70783 , n70780 , n70782 );
buf ( n417416 , n388406 );
buf ( n417417 , n44776 );
nand ( n70786 , n417416 , n417417 );
buf ( n417419 , n70786 );
buf ( n417420 , n417419 );
nand ( n70789 , n70783 , n417420 );
buf ( n417422 , n70789 );
buf ( n417423 , n417422 );
not ( n70792 , n417423 );
or ( n70793 , n70778 , n70792 );
buf ( n417426 , n69262 );
buf ( n417427 , n413643 );
nand ( n70796 , n417426 , n417427 );
buf ( n417429 , n70796 );
buf ( n417430 , n417429 );
nand ( n70799 , n70793 , n417430 );
buf ( n417432 , n70799 );
buf ( n417433 , n417432 );
xor ( n70802 , n417408 , n417433 );
not ( n70803 , n37338 );
buf ( n417436 , n388905 );
not ( n70805 , n417436 );
buf ( n417438 , n399283 );
not ( n70807 , n417438 );
and ( n70808 , n70805 , n70807 );
buf ( n417441 , n395478 );
buf ( n417442 , n399283 );
and ( n70811 , n417441 , n417442 );
nor ( n70812 , n70808 , n70811 );
buf ( n417445 , n70812 );
buf ( n417446 , n417445 );
not ( n70815 , n417446 );
buf ( n417448 , n70815 );
not ( n70817 , n417448 );
or ( n70818 , n70803 , n70817 );
buf ( n417451 , n416348 );
buf ( n417452 , n37314 );
nand ( n70821 , n417451 , n417452 );
buf ( n417454 , n70821 );
nand ( n70823 , n70818 , n417454 );
buf ( n417456 , n70823 );
and ( n70825 , n70802 , n417456 );
and ( n70826 , n417408 , n417433 );
or ( n70827 , n70825 , n70826 );
buf ( n417460 , n70827 );
buf ( n417461 , n417460 );
nand ( n70830 , n70111 , n417461 );
buf ( n417463 , n70830 );
buf ( n417464 , n417463 );
nand ( n70833 , n70108 , n417464 );
buf ( n417466 , n70833 );
buf ( n417467 , n417466 );
and ( n70836 , n69997 , n417467 );
or ( n70838 , n70836 , C0 );
buf ( n417470 , n70838 );
buf ( n417471 , n417470 );
xor ( n70841 , n416622 , n417471 );
xor ( n70842 , n416075 , n416082 );
xor ( n70843 , n70842 , n416399 );
buf ( n417475 , n70843 );
buf ( n417476 , n417475 );
and ( n70846 , n70841 , n417476 );
and ( n70847 , n416622 , n417471 );
or ( n70848 , n70846 , n70847 );
buf ( n417480 , n70848 );
buf ( n417481 , n417480 );
and ( n70851 , n69963 , n417481 );
and ( n70852 , n416613 , n416617 );
or ( n70853 , n70851 , n70852 );
buf ( n417485 , n70853 );
buf ( n417486 , n417485 );
and ( n70856 , n69782 , n417486 );
and ( n70857 , n416469 , n416473 );
or ( n70858 , n70856 , n70857 );
buf ( n417490 , n70858 );
buf ( n417491 , n417490 );
or ( n70861 , n416462 , n417491 );
buf ( n417493 , n70861 );
buf ( n417494 , n417493 );
and ( n70864 , n415855 , n417494 );
buf ( n417496 , n69769 );
buf ( n417497 , n417490 );
and ( n70867 , n417496 , n417497 );
buf ( n417499 , n70867 );
buf ( n417500 , n417499 );
nor ( n70870 , n70864 , n417500 );
buf ( n417502 , n70870 );
buf ( n417503 , n417502 );
nand ( n70873 , n415849 , n417503 );
buf ( n417505 , n70873 );
buf ( n417506 , n417505 );
and ( n70876 , n415765 , n415845 , n417506 );
buf ( n417508 , n70876 );
not ( n70878 , n417508 );
buf ( n417510 , n413643 );
not ( n70880 , n417510 );
buf ( n417512 , n399986 );
not ( n70882 , n417512 );
buf ( n417514 , n388566 );
not ( n70884 , n417514 );
or ( n70885 , n70882 , n70884 );
buf ( n417517 , n27258 );
buf ( n417518 , n44776 );
nand ( n70888 , n417517 , n417518 );
buf ( n417520 , n70888 );
buf ( n417521 , n417520 );
nand ( n70891 , n70885 , n417521 );
buf ( n417523 , n70891 );
buf ( n417524 , n417523 );
not ( n70894 , n417524 );
or ( n70895 , n70880 , n70894 );
buf ( n417527 , n399986 );
not ( n70897 , n417527 );
buf ( n417529 , n403039 );
not ( n70899 , n417529 );
or ( n70900 , n70897 , n70899 );
buf ( n417532 , n388543 );
buf ( n417533 , n44776 );
nand ( n70903 , n417532 , n417533 );
buf ( n417535 , n70903 );
buf ( n417536 , n417535 );
nand ( n70906 , n70900 , n417536 );
buf ( n417538 , n70906 );
buf ( n417539 , n417538 );
buf ( n417540 , n44771 );
not ( n70910 , n417540 );
buf ( n417542 , n70910 );
buf ( n417543 , n417542 );
nand ( n70913 , n417539 , n417543 );
buf ( n417545 , n70913 );
buf ( n417546 , n417545 );
nand ( n70916 , n70895 , n417546 );
buf ( n417548 , n70916 );
buf ( n417549 , n417548 );
buf ( n417550 , n385473 );
buf ( n417551 , n49661 );
not ( n70921 , n417551 );
buf ( n417553 , n37919 );
not ( n70923 , n417553 );
or ( n70924 , n70921 , n70923 );
buf ( n417556 , n358975 );
nand ( n70926 , n70924 , n417556 );
buf ( n417558 , n70926 );
buf ( n417559 , n417558 );
buf ( n417560 , n37919 );
not ( n70930 , n417560 );
buf ( n417562 , n22982 );
nand ( n70932 , n70930 , n417562 );
buf ( n417564 , n70932 );
buf ( n417565 , n417564 );
and ( n70935 , n417550 , n417559 , n417565 );
buf ( n417567 , n70935 );
buf ( n417568 , n417567 );
xor ( n70938 , n417549 , n417568 );
buf ( n417570 , n394814 );
not ( n70940 , n417570 );
buf ( n417572 , n70940 );
buf ( n417573 , n417572 );
not ( n70943 , n417573 );
buf ( n417575 , n404601 );
not ( n70945 , n417575 );
or ( n70946 , n70943 , n70945 );
buf ( n417578 , n407936 );
buf ( n417579 , n394814 );
nand ( n70949 , n417578 , n417579 );
buf ( n417581 , n70949 );
buf ( n417582 , n417581 );
nand ( n70952 , n70946 , n417582 );
buf ( n417584 , n70952 );
buf ( n417585 , n417584 );
not ( n70955 , n417585 );
buf ( n417587 , n406422 );
not ( n70957 , n417587 );
or ( n70958 , n70955 , n70957 );
buf ( n417590 , n394210 );
not ( n70960 , n417590 );
buf ( n417592 , n409092 );
not ( n70962 , n417592 );
or ( n70963 , n70960 , n70962 );
buf ( n417595 , n407928 );
buf ( n417596 , n394219 );
nand ( n70966 , n417595 , n417596 );
buf ( n417598 , n70966 );
buf ( n417599 , n417598 );
nand ( n70969 , n70963 , n417599 );
buf ( n417601 , n70969 );
buf ( n417602 , n417601 );
buf ( n417603 , n409076 );
nand ( n70973 , n417602 , n417603 );
buf ( n417605 , n70973 );
buf ( n417606 , n417605 );
nand ( n70976 , n70958 , n417606 );
buf ( n417608 , n70976 );
buf ( n417609 , n417608 );
buf ( n417610 , n41861 );
not ( n70980 , n417610 );
buf ( n417612 , n388754 );
not ( n70982 , n417612 );
or ( n70983 , n70980 , n70982 );
buf ( n417615 , n371797 );
not ( n70985 , n417615 );
buf ( n417617 , n70985 );
buf ( n417618 , n417617 );
buf ( n417619 , n389353 );
nand ( n70989 , n417618 , n417619 );
buf ( n417621 , n70989 );
buf ( n417622 , n417621 );
nand ( n70992 , n70983 , n417622 );
buf ( n417624 , n70992 );
buf ( n417625 , n417624 );
buf ( n417626 , n388803 );
nand ( n70996 , n417625 , n417626 );
buf ( n417628 , n70996 );
not ( n70998 , n417628 );
buf ( n417630 , n389341 );
buf ( n417631 , n371800 );
and ( n71001 , n417630 , n417631 );
not ( n71002 , n417630 );
buf ( n417634 , n371797 );
and ( n71004 , n71002 , n417634 );
nor ( n71005 , n71001 , n71004 );
buf ( n417637 , n71005 );
not ( n71007 , n417637 );
nor ( n71008 , n71007 , n388737 );
nor ( n71009 , n70998 , n71008 );
buf ( n417641 , n58166 );
buf ( n417642 , n66411 );
and ( n71012 , n417641 , n417642 );
buf ( n417644 , n58205 );
buf ( n417645 , n62496 );
and ( n71015 , n417644 , n417645 );
nor ( n71016 , n71012 , n71015 );
buf ( n417648 , n71016 );
buf ( n417649 , n417648 );
buf ( n417650 , n410724 );
or ( n71020 , n417649 , n417650 );
buf ( n417652 , n58178 );
buf ( n417653 , n66411 );
and ( n71023 , n417652 , n417653 );
buf ( n417655 , n405335 );
buf ( n417656 , n62496 );
and ( n71026 , n417655 , n417656 );
nor ( n71027 , n71023 , n71026 );
buf ( n417659 , n71027 );
buf ( n417660 , n417659 );
buf ( n417661 , n410721 );
or ( n71031 , n417660 , n417661 );
nand ( n71032 , n71020 , n71031 );
buf ( n417664 , n71032 );
buf ( n417665 , n417664 );
buf ( n417666 , n63707 );
buf ( n417667 , n405391 );
and ( n71037 , n417666 , n417667 );
buf ( n417669 , n413104 );
buf ( n417670 , n405388 );
and ( n71040 , n417669 , n417670 );
nor ( n71041 , n71037 , n71040 );
buf ( n417673 , n71041 );
buf ( n417674 , n417673 );
buf ( n417675 , n405407 );
or ( n71045 , n417674 , n417675 );
buf ( n417677 , n63564 );
buf ( n417678 , n405391 );
and ( n71048 , n417677 , n417678 );
buf ( n417680 , n413073 );
buf ( n417681 , n414664 );
and ( n71051 , n417680 , n417681 );
nor ( n71052 , n71048 , n71051 );
buf ( n417684 , n71052 );
buf ( n417685 , n417684 );
buf ( n417686 , n405384 );
or ( n71056 , n417685 , n417686 );
nand ( n71057 , n71045 , n71056 );
buf ( n417689 , n71057 );
buf ( n417690 , n417689 );
buf ( n417691 , n70389 );
buf ( n417692 , n401689 );
and ( n71062 , n417691 , n417692 );
buf ( n417694 , n417024 );
buf ( n417695 , n401692 );
and ( n71065 , n417694 , n417695 );
nor ( n71066 , n71062 , n71065 );
buf ( n417698 , n71066 );
buf ( n417699 , n417698 );
buf ( n417700 , n403158 );
or ( n71070 , n417699 , n417700 );
buf ( n417702 , n70210 );
buf ( n417703 , n401689 );
and ( n71073 , n417702 , n417703 );
buf ( n417705 , n416845 );
buf ( n417706 , n401695 );
and ( n71076 , n417705 , n417706 );
nor ( n71077 , n71073 , n71076 );
buf ( n417709 , n71077 );
buf ( n417710 , n417709 );
buf ( n417711 , n403167 );
or ( n71081 , n417710 , n417711 );
nand ( n71082 , n71070 , n71081 );
buf ( n417714 , n71082 );
buf ( n417715 , n417714 );
buf ( n417716 , n401623 );
not ( n71086 , n54170 );
nor ( n71087 , n71086 , n54209 );
xor ( n71088 , n54206 , n71087 );
buf ( n417720 , n71088 );
not ( n71090 , n417720 );
buf ( n417722 , n71090 );
buf ( n417723 , n417722 );
or ( n71093 , n417716 , n417723 );
xor ( n71094 , n54150 , n54152 );
xor ( n71095 , n71094 , n54211 );
buf ( n417727 , n71095 );
not ( n71097 , n417727 );
buf ( n417729 , n71097 );
buf ( n417730 , n417729 );
buf ( n417731 , n403092 );
or ( n71101 , n417730 , n417731 );
nand ( n71102 , n71093 , n71101 );
buf ( n417734 , n71102 );
buf ( n417735 , n417734 );
xor ( n71105 , n417715 , n417735 );
buf ( n417737 , n55875 );
not ( n71107 , n417737 );
buf ( n417739 , n68002 );
buf ( n417740 , n55905 );
and ( n417741 , n417739 , n417740 );
buf ( n417742 , n414729 );
buf ( n417743 , n55895 );
and ( n71113 , n417742 , n417743 );
nor ( n71114 , n417741 , n71113 );
buf ( n417746 , n71114 );
buf ( n417747 , n417746 );
not ( n71117 , n417747 );
buf ( n417749 , n71117 );
buf ( n417750 , n417749 );
not ( n71120 , n417750 );
or ( n71121 , n71107 , n71120 );
buf ( n417753 , n70195 );
buf ( n417754 , n55905 );
and ( n71124 , n417753 , n417754 );
buf ( n417756 , n416830 );
buf ( n417757 , n55895 );
and ( n71127 , n417756 , n417757 );
nor ( n71128 , n71124 , n71127 );
buf ( n417760 , n71128 );
buf ( n417761 , n417760 );
buf ( n417762 , n403120 );
or ( n71132 , n417761 , n417762 );
nand ( n71133 , n71121 , n71132 );
buf ( n417765 , n71133 );
buf ( n417766 , n417765 );
and ( n71136 , n71105 , n417766 );
and ( n71137 , n417715 , n417735 );
or ( n71138 , n71136 , n71137 );
buf ( n417770 , n71138 );
buf ( n417771 , n417770 );
xor ( n71141 , n417690 , n417771 );
buf ( n417773 , n67987 );
buf ( n417774 , n405215 );
and ( n71144 , n417773 , n417774 );
buf ( n417776 , n414714 );
buf ( n417777 , n58061 );
and ( n71147 , n417776 , n417777 );
nor ( n71148 , n71144 , n71147 );
buf ( n417780 , n71148 );
buf ( n417781 , n417780 );
buf ( n417782 , n403293 );
or ( n71152 , n417781 , n417782 );
buf ( n417784 , n66359 );
buf ( n417785 , n405215 );
and ( n71155 , n417784 , n417785 );
buf ( n417787 , n413187 );
buf ( n417788 , n58061 );
and ( n71158 , n417787 , n417788 );
nor ( n71159 , n71155 , n71158 );
buf ( n417791 , n71159 );
buf ( n417792 , n417791 );
buf ( n417793 , n405476 );
or ( n71163 , n417792 , n417793 );
nand ( n71164 , n71152 , n71163 );
buf ( n417796 , n71164 );
buf ( n417797 , n417796 );
buf ( n417798 , n401623 );
not ( n71168 , n54203 );
nand ( n71169 , n71168 , n54205 );
xor ( n71170 , n71169 , n54199 );
buf ( n417802 , n71170 );
not ( n71172 , n417802 );
buf ( n417804 , n71172 );
buf ( n417805 , n417804 );
or ( n71175 , n417798 , n417805 );
buf ( n417807 , n403092 );
buf ( n417808 , n417722 );
or ( n71178 , n417807 , n417808 );
nand ( n71179 , n71175 , n71178 );
buf ( n417811 , n71179 );
buf ( n417812 , n417811 );
buf ( n417813 , n403164 );
not ( n71183 , n417813 );
buf ( n417815 , n417698 );
not ( n71185 , n417815 );
buf ( n417817 , n71185 );
buf ( n417818 , n417817 );
not ( n71188 , n417818 );
or ( n71189 , n71183 , n71188 );
buf ( n417821 , n401689 );
buf ( n417822 , n71095 );
and ( n71192 , n417821 , n417822 );
not ( n71193 , n417821 );
buf ( n417825 , n417729 );
and ( n71195 , n71193 , n417825 );
nor ( n71196 , n71192 , n71195 );
buf ( n417828 , n71196 );
buf ( n417829 , n417828 );
buf ( n417830 , n403158 );
or ( n71200 , n417829 , n417830 );
nand ( n71201 , n71189 , n71200 );
buf ( n417833 , n71201 );
buf ( n417834 , n417833 );
and ( n71204 , n417812 , n417834 );
buf ( n417836 , n71204 );
buf ( n417837 , n417836 );
xor ( n71207 , n417797 , n417837 );
xor ( n71208 , n417715 , n417735 );
xor ( n71209 , n71208 , n417766 );
buf ( n417841 , n71209 );
buf ( n417842 , n417841 );
and ( n71212 , n71207 , n417842 );
and ( n71213 , n417797 , n417837 );
or ( n71214 , n71212 , n71213 );
buf ( n417846 , n71214 );
buf ( n417847 , n417846 );
and ( n71217 , n71141 , n417847 );
and ( n71218 , n417690 , n417771 );
or ( n71219 , n71217 , n71218 );
buf ( n417851 , n71219 );
buf ( n417852 , n417851 );
xor ( n71222 , n417665 , n417852 );
buf ( n417854 , n62139 );
buf ( n417855 , n62177 );
and ( n71225 , n417854 , n417855 );
buf ( n417857 , n409140 );
buf ( n417858 , n62159 );
and ( n71228 , n417857 , n417858 );
nor ( n71229 , n71225 , n71228 );
buf ( n417861 , n71229 );
buf ( n417862 , n417861 );
buf ( n417863 , n409429 );
or ( n71233 , n417862 , n417863 );
buf ( n417865 , n59596 );
buf ( n417866 , n62177 );
and ( n71236 , n417865 , n417866 );
buf ( n417868 , n409146 );
buf ( n417869 , n62159 );
and ( n71239 , n417868 , n417869 );
nor ( n71240 , n71236 , n71239 );
buf ( n417872 , n71240 );
buf ( n417873 , n417872 );
buf ( n417874 , n409170 );
or ( n71244 , n417873 , n417874 );
nand ( n71245 , n71233 , n71244 );
buf ( n417877 , n71245 );
buf ( n417878 , n417877 );
buf ( n417879 , n62467 );
buf ( n417880 , n59628 );
and ( n71250 , n417879 , n417880 );
buf ( n417882 , n409468 );
buf ( n417883 , n59457 );
and ( n71253 , n417882 , n417883 );
nor ( n71254 , n71250 , n71253 );
buf ( n417886 , n71254 );
buf ( n417887 , n417886 );
buf ( n417888 , n59637 );
or ( n71258 , n417887 , n417888 );
buf ( n417890 , n62278 );
buf ( n417891 , n59628 );
and ( n71261 , n417890 , n417891 );
buf ( n417893 , n409474 );
buf ( n417894 , n59457 );
and ( n71264 , n417893 , n417894 );
nor ( n71265 , n71261 , n71264 );
buf ( n417897 , n71265 );
buf ( n417898 , n417897 );
buf ( n417899 , n59467 );
or ( n71269 , n417898 , n417899 );
nand ( n71270 , n71258 , n71269 );
buf ( n417902 , n71270 );
buf ( n417903 , n417902 );
xor ( n71273 , n417878 , n417903 );
buf ( n417905 , n401623 );
buf ( n417906 , n417729 );
or ( n71276 , n417905 , n417906 );
buf ( n417908 , n417024 );
buf ( n417909 , n403092 );
or ( n71279 , n417908 , n417909 );
nand ( n71280 , n71276 , n71279 );
buf ( n417912 , n71280 );
buf ( n417913 , n417912 );
buf ( n417914 , n417709 );
buf ( n417915 , n403158 );
or ( n71285 , n417914 , n417915 );
buf ( n417917 , n417010 );
buf ( n417918 , n403167 );
or ( n71288 , n417917 , n417918 );
nand ( n71289 , n71285 , n71288 );
buf ( n417921 , n71289 );
buf ( n417922 , n417921 );
xor ( n71292 , n417913 , n417922 );
buf ( n417924 , n71292 );
buf ( n417925 , n417924 );
buf ( n417926 , n417746 );
buf ( n417927 , n403120 );
or ( n71297 , n417926 , n417927 );
buf ( n417929 , n417044 );
buf ( n417930 , n403133 );
or ( n71300 , n417929 , n417930 );
nand ( n71301 , n71297 , n71300 );
buf ( n417933 , n71301 );
buf ( n417934 , n417933 );
xor ( n71304 , n417925 , n417934 );
buf ( n417936 , n417791 );
buf ( n417937 , n403293 );
or ( n71307 , n417936 , n417937 );
buf ( n417939 , n66270 );
buf ( n417940 , n405215 );
and ( n71310 , n417939 , n417940 );
buf ( n417942 , n413098 );
buf ( n417943 , n58061 );
and ( n71313 , n417942 , n417943 );
nor ( n71314 , n71310 , n71313 );
buf ( n417946 , n71314 );
buf ( n417947 , n417946 );
buf ( n417948 , n405476 );
or ( n71318 , n417947 , n417948 );
nand ( n71319 , n71307 , n71318 );
buf ( n417951 , n71319 );
buf ( n417952 , n417951 );
xor ( n71322 , n71304 , n417952 );
buf ( n417954 , n71322 );
buf ( n417955 , n417954 );
and ( n71325 , n71273 , n417955 );
and ( n71326 , n417878 , n417903 );
or ( n71327 , n71325 , n71326 );
buf ( n417959 , n71327 );
buf ( n417960 , n417959 );
and ( n71330 , n71222 , n417960 );
and ( n71331 , n417665 , n417852 );
or ( n71332 , n71330 , n71331 );
buf ( n417964 , n71332 );
buf ( n417965 , n58200 );
buf ( n417966 , n63625 );
and ( n71336 , n417965 , n417966 );
buf ( n417968 , n58201 );
buf ( n417969 , n63629 );
and ( n71339 , n417968 , n417969 );
nor ( n71340 , n71336 , n71339 );
buf ( n417972 , n71340 );
buf ( n417973 , n417972 );
buf ( n417974 , n410635 );
or ( n71344 , n417973 , n417974 );
buf ( n417976 , n58166 );
buf ( n417977 , n63625 );
and ( n71347 , n417976 , n417977 );
buf ( n417979 , n58205 );
buf ( n417980 , n63629 );
and ( n71350 , n417979 , n417980 );
nor ( n71351 , n71347 , n71350 );
buf ( n417983 , n71351 );
buf ( n417984 , n417983 );
buf ( n417985 , n409504 );
or ( n71355 , n417984 , n417985 );
nand ( n71356 , n71344 , n71355 );
buf ( n417988 , n71356 );
or ( n71358 , n417659 , n410724 );
not ( n71359 , n410721 );
nand ( n71360 , n71359 , n70540 );
nand ( n71361 , n71358 , n71360 );
xor ( n71362 , n417988 , n71361 );
xor ( n71363 , n417925 , n417934 );
and ( n71364 , n71363 , n417952 );
and ( n71365 , n417925 , n417934 );
or ( n71366 , n71364 , n71365 );
buf ( n417998 , n71366 );
buf ( n417999 , n417998 );
buf ( n418000 , n417684 );
buf ( n418001 , n405407 );
or ( n71371 , n418000 , n418001 );
buf ( n418003 , n62467 );
buf ( n418004 , n405391 );
and ( n71374 , n418003 , n418004 );
buf ( n418006 , n409468 );
buf ( n418007 , n414664 );
and ( n71377 , n418006 , n418007 );
nor ( n71378 , n71374 , n71377 );
buf ( n418010 , n71378 );
buf ( n418011 , n418010 );
buf ( n418012 , n405384 );
or ( n418013 , n418011 , n418012 );
nand ( n71383 , n71371 , n418013 );
buf ( n418015 , n71383 );
buf ( n418016 , n418015 );
xor ( n71386 , n417999 , n418016 );
buf ( n418018 , n417872 );
buf ( n418019 , n409429 );
or ( n71389 , n418018 , n418019 );
buf ( n418021 , n59435 );
buf ( n418022 , n62177 );
and ( n71392 , n418021 , n418022 );
buf ( n418024 , n406565 );
buf ( n418025 , n62159 );
and ( n71395 , n418024 , n418025 );
nor ( n71396 , n71392 , n71395 );
buf ( n418028 , n71396 );
buf ( n418029 , n418028 );
buf ( n418030 , n409170 );
or ( n71400 , n418029 , n418030 );
nand ( n71401 , n71389 , n71400 );
buf ( n418033 , n71401 );
buf ( n418034 , n418033 );
and ( n71404 , n71386 , n418034 );
and ( n71405 , n417999 , n418016 );
or ( n71406 , n71404 , n71405 );
buf ( n418038 , n71406 );
xor ( n71408 , n71362 , n418038 );
and ( n71409 , n417964 , n71408 );
buf ( n418041 , n417946 );
buf ( n418042 , n403293 );
or ( n71412 , n418041 , n418042 );
buf ( n418044 , n63707 );
buf ( n418045 , n405215 );
and ( n71415 , n418044 , n418045 );
buf ( n418047 , n413104 );
buf ( n418048 , n58061 );
and ( n71418 , n418047 , n418048 );
nor ( n71419 , n71415 , n71418 );
buf ( n418051 , n71419 );
buf ( n418052 , n418051 );
buf ( n418053 , n405476 );
or ( n71423 , n418052 , n418053 );
nand ( n71424 , n71412 , n71423 );
buf ( n418056 , n71424 );
buf ( n418057 , n418056 );
and ( n71427 , n417913 , n417922 );
buf ( n418059 , n71427 );
buf ( n418060 , n418059 );
xor ( n71430 , n418057 , n418060 );
xor ( n71431 , n417019 , n417033 );
xor ( n71432 , n71431 , n417056 );
buf ( n418064 , n71432 );
buf ( n418065 , n418064 );
xor ( n71435 , n71430 , n418065 );
buf ( n418067 , n71435 );
buf ( n418068 , n417897 );
buf ( n418069 , n59637 );
or ( n71439 , n418068 , n418069 );
buf ( n418071 , n62139 );
buf ( n418072 , n59628 );
and ( n71442 , n418071 , n418072 );
buf ( n418074 , n409140 );
buf ( n418075 , n59457 );
and ( n71445 , n418074 , n418075 );
nor ( n71446 , n71442 , n71445 );
buf ( n418078 , n71446 );
buf ( n418079 , n418078 );
buf ( n418080 , n59467 );
or ( n71450 , n418079 , n418080 );
nand ( n71451 , n71439 , n71450 );
buf ( n418083 , n71451 );
xor ( n71453 , n418067 , n418083 );
buf ( n418085 , n58352 );
buf ( n418086 , n63625 );
and ( n71456 , n418085 , n418086 );
buf ( n418088 , n406571 );
buf ( n418089 , n63629 );
and ( n71459 , n418088 , n418089 );
nor ( n71460 , n71456 , n71459 );
buf ( n418092 , n71460 );
buf ( n418093 , n418092 );
buf ( n418094 , n410635 );
or ( n71464 , n418093 , n418094 );
buf ( n418096 , n417972 );
buf ( n418097 , n409504 );
or ( n71467 , n418096 , n418097 );
nand ( n71468 , n71464 , n71467 );
buf ( n418100 , n71468 );
and ( n71470 , n71453 , n418100 );
and ( n71471 , n418067 , n418083 );
or ( n71472 , n71470 , n71471 );
buf ( n418104 , n71472 );
buf ( n418105 , n418010 );
buf ( n418106 , n405407 );
or ( n71476 , n418105 , n418106 );
buf ( n418108 , n416963 );
buf ( n418109 , n405384 );
or ( n71479 , n418108 , n418109 );
nand ( n71480 , n71476 , n71479 );
buf ( n418112 , n71480 );
buf ( n418113 , n418112 );
buf ( n418114 , n418051 );
buf ( n418115 , n403293 );
or ( n71485 , n418114 , n418115 );
buf ( n418117 , n417099 );
buf ( n418118 , n405476 );
or ( n71488 , n418117 , n418118 );
nand ( n71489 , n71485 , n71488 );
buf ( n418121 , n71489 );
buf ( n418122 , n418121 );
xor ( n71492 , n418113 , n418122 );
buf ( n418124 , n418078 );
buf ( n418125 , n59637 );
or ( n71495 , n418124 , n418125 );
buf ( n418127 , n416946 );
buf ( n418128 , n59467 );
or ( n71498 , n418127 , n418128 );
nand ( n71499 , n71495 , n71498 );
buf ( n418131 , n71499 );
buf ( n418132 , n418131 );
xor ( n71502 , n71492 , n418132 );
buf ( n418134 , n71502 );
buf ( n418135 , n418134 );
xor ( n71505 , n418104 , n418135 );
xor ( n71506 , n416976 , n417001 );
xor ( n71507 , n71506 , n417061 );
buf ( n418139 , n71507 );
buf ( n418140 , n418139 );
xor ( n71510 , n418057 , n418060 );
and ( n71511 , n71510 , n418065 );
and ( n71512 , n418057 , n418060 );
or ( n71513 , n71511 , n71512 );
buf ( n418145 , n71513 );
buf ( n418146 , n418145 );
xor ( n71516 , n418140 , n418146 );
buf ( n418148 , n418028 );
buf ( n418149 , n409429 );
or ( n71519 , n418148 , n418149 );
buf ( n418151 , n417183 );
buf ( n418152 , n409170 );
or ( n71522 , n418151 , n418152 );
nand ( n71523 , n71519 , n71522 );
buf ( n418155 , n71523 );
buf ( n418156 , n418155 );
xor ( n71526 , n71516 , n418156 );
buf ( n418158 , n71526 );
buf ( n418159 , n418158 );
xor ( n71529 , n71505 , n418159 );
buf ( n418161 , n71529 );
xor ( n71531 , n417988 , n71361 );
xor ( n71532 , n71531 , n418038 );
and ( n71533 , n418161 , n71532 );
and ( n71534 , n417964 , n418161 );
or ( n71535 , n71409 , n71533 , n71534 );
not ( n71536 , n71535 );
xor ( n71537 , n418104 , n418135 );
and ( n71538 , n71537 , n418159 );
and ( n71539 , n418104 , n418135 );
or ( n71540 , n71538 , n71539 );
buf ( n418172 , n71540 );
buf ( n418173 , n418172 );
xor ( n71543 , n418113 , n418122 );
and ( n71544 , n71543 , n418132 );
and ( n71545 , n418113 , n418122 );
or ( n71546 , n71544 , n71545 );
buf ( n418178 , n71546 );
buf ( n418179 , n418178 );
buf ( n418180 , n417983 );
buf ( n418181 , n410635 );
or ( n71551 , n418180 , n418181 );
buf ( n418183 , n417138 );
buf ( n418184 , n409504 );
or ( n71554 , n418183 , n418184 );
nand ( n71555 , n71551 , n71554 );
buf ( n418187 , n71555 );
buf ( n418188 , n418187 );
xor ( n71558 , n418179 , n418188 );
xor ( n71559 , n416955 , n416972 );
xor ( n71560 , n71559 , n417066 );
buf ( n418192 , n71560 );
buf ( n418193 , n418192 );
xor ( n71563 , n71558 , n418193 );
buf ( n418195 , n71563 );
buf ( n418196 , n418195 );
xor ( n71566 , n418173 , n418196 );
xor ( n71567 , n417988 , n71361 );
and ( n71568 , n71567 , n418038 );
and ( n71569 , n417988 , n71361 );
or ( n71570 , n71568 , n71569 );
buf ( n418202 , n71570 );
xor ( n71572 , n418140 , n418146 );
and ( n71573 , n71572 , n418156 );
and ( n71574 , n418140 , n418146 );
or ( n71575 , n71573 , n71574 );
buf ( n418207 , n71575 );
buf ( n418208 , n418207 );
xor ( n71578 , n418202 , n418208 );
xor ( n71579 , n417175 , n417192 );
xor ( n71580 , n71579 , n417197 );
buf ( n418212 , n71580 );
buf ( n418213 , n418212 );
xor ( n71583 , n71578 , n418213 );
buf ( n418215 , n71583 );
buf ( n418216 , n418215 );
xor ( n71586 , n71566 , n418216 );
buf ( n418218 , n71586 );
not ( n71588 , n418218 );
or ( n71589 , n71536 , n71588 );
not ( n71590 , n71535 );
not ( n71591 , n418218 );
and ( n71592 , n71590 , n71591 );
not ( n71593 , n71592 );
xor ( n71594 , n417988 , n71361 );
xor ( n71595 , n71594 , n418038 );
xor ( n71596 , n417964 , n418161 );
xor ( n71597 , n71595 , n71596 );
buf ( n418229 , n71597 );
xor ( n71599 , n417999 , n418016 );
xor ( n71600 , n71599 , n418034 );
buf ( n418232 , n71600 );
xor ( n71602 , n418067 , n418083 );
xor ( n71603 , n71602 , n418100 );
and ( n71604 , n418232 , n71603 );
buf ( n418236 , n59435 );
buf ( n418237 , n63625 );
and ( n71607 , n418236 , n418237 );
buf ( n418239 , n406565 );
buf ( n418240 , n63629 );
and ( n71610 , n418239 , n418240 );
nor ( n71611 , n71607 , n71610 );
buf ( n418243 , n71611 );
buf ( n418244 , n418243 );
buf ( n418245 , n410635 );
or ( n71615 , n418244 , n418245 );
buf ( n418247 , n418092 );
buf ( n418248 , n409504 );
or ( n71618 , n418247 , n418248 );
nand ( n71619 , n71615 , n71618 );
buf ( n418251 , n71619 );
buf ( n418252 , n418251 );
buf ( n418253 , n70210 );
buf ( n418254 , n55905 );
and ( n71624 , n418253 , n418254 );
buf ( n418256 , n416845 );
buf ( n418257 , n55895 );
and ( n71627 , n418256 , n418257 );
nor ( n71628 , n71624 , n71627 );
buf ( n418260 , n71628 );
buf ( n418261 , n418260 );
buf ( n418262 , n403120 );
or ( n71632 , n418261 , n418262 );
buf ( n418264 , n417760 );
buf ( n418265 , n403133 );
or ( n71635 , n418264 , n418265 );
nand ( n71636 , n71632 , n71635 );
buf ( n418268 , n71636 );
buf ( n418269 , n418268 );
buf ( n418270 , n403158 );
buf ( n418271 , n71088 );
buf ( n418272 , n401689 );
and ( n71642 , n418271 , n418272 );
buf ( n418274 , n417722 );
buf ( n418275 , n401678 );
and ( n71645 , n418274 , n418275 );
nor ( n71646 , n71642 , n71645 );
buf ( n418278 , n71646 );
buf ( n418279 , n418278 );
or ( n71649 , n418270 , n418279 );
buf ( n418281 , n417828 );
buf ( n418282 , n403167 );
or ( n71652 , n418281 , n418282 );
nand ( n71653 , n71649 , n71652 );
buf ( n418285 , n71653 );
buf ( n418286 , n401623 );
not ( n71656 , n54197 );
nor ( n71657 , n71656 , n54188 );
not ( n71658 , n71657 );
not ( n71659 , n54175 );
nor ( n71660 , n71659 , n54195 );
not ( n71661 , n71660 );
or ( n71662 , n71658 , n71661 );
or ( n71663 , n71660 , n71657 );
nand ( n71664 , n71662 , n71663 );
buf ( n418296 , n71664 );
not ( n71666 , n418296 );
buf ( n418298 , n71666 );
buf ( n418299 , n418298 );
or ( n71669 , n418286 , n418299 );
buf ( n418301 , n401619 );
buf ( n418302 , n417804 );
or ( n71672 , n418301 , n418302 );
nand ( n71673 , n71669 , n71672 );
buf ( n418305 , n71673 );
xor ( n71675 , n418285 , n418305 );
buf ( n418307 , n401623 );
not ( n71677 , n54195 );
or ( n71678 , n54192 , n621 );
nand ( n71679 , n71678 , n54193 , n54194 );
nand ( n71680 , n71677 , n71679 );
xnor ( n71681 , n71680 , n54174 );
buf ( n418313 , n71681 );
not ( n71683 , n418313 );
buf ( n418315 , n71683 );
buf ( n418316 , n418315 );
or ( n71686 , n418307 , n418316 );
buf ( n418318 , n401619 );
buf ( n418319 , n418298 );
or ( n71689 , n418318 , n418319 );
nand ( n71690 , n71686 , n71689 );
buf ( n418322 , n71690 );
buf ( n418323 , n418322 );
buf ( n418324 , n403158 );
buf ( n418325 , n401689 );
buf ( n418326 , n71170 );
and ( n71696 , n418325 , n418326 );
buf ( n418328 , n401678 );
buf ( n418329 , n417804 );
and ( n71699 , n418328 , n418329 );
nor ( n71700 , n71696 , n71699 );
buf ( n418332 , n71700 );
buf ( n418333 , n418332 );
or ( n71703 , n418324 , n418333 );
buf ( n418335 , n418278 );
buf ( n418336 , n401660 );
or ( n71706 , n418335 , n418336 );
nand ( n71707 , n71703 , n71706 );
buf ( n418339 , n71707 );
buf ( n418340 , n418339 );
and ( n71710 , n418323 , n418340 );
buf ( n418342 , n71710 );
and ( n71712 , n71675 , n418342 );
and ( n71713 , n418285 , n418305 );
or ( n71714 , n71712 , n71713 );
buf ( n418346 , n71714 );
xor ( n71716 , n418269 , n418346 );
xor ( n71717 , n417812 , n417834 );
buf ( n418349 , n71717 );
buf ( n418350 , n418349 );
and ( n71720 , n71716 , n418350 );
and ( n71721 , n418269 , n418346 );
or ( n71722 , n71720 , n71721 );
buf ( n418354 , n71722 );
buf ( n418355 , n66270 );
buf ( n418356 , n405391 );
and ( n71726 , n418355 , n418356 );
buf ( n418358 , n413098 );
buf ( n418359 , n414664 );
and ( n71729 , n418358 , n418359 );
nor ( n71730 , n71726 , n71729 );
buf ( n418362 , n71730 );
buf ( n418363 , n418362 );
buf ( n418364 , n405407 );
or ( n71734 , n418363 , n418364 );
buf ( n418366 , n417673 );
buf ( n418367 , n405384 );
or ( n71737 , n418366 , n418367 );
nand ( n71738 , n71734 , n71737 );
buf ( n418370 , n71738 );
xor ( n71740 , n418354 , n418370 );
buf ( n418372 , n63564 );
buf ( n418373 , n59628 );
and ( n71743 , n418372 , n418373 );
buf ( n418375 , n413073 );
buf ( n418376 , n59457 );
and ( n71746 , n418375 , n418376 );
nor ( n71747 , n71743 , n71746 );
buf ( n418379 , n71747 );
buf ( n418380 , n418379 );
buf ( n418381 , n59637 );
or ( n71751 , n418380 , n418381 );
buf ( n418383 , n417886 );
buf ( n418384 , n59467 );
or ( n71754 , n418383 , n418384 );
nand ( n71755 , n71751 , n71754 );
buf ( n418387 , n71755 );
and ( n71757 , n71740 , n418387 );
and ( n71758 , n418354 , n418370 );
or ( n71759 , n71757 , n71758 );
buf ( n418391 , n71759 );
xor ( n71761 , n418252 , n418391 );
xor ( n71762 , n417690 , n417771 );
xor ( n71763 , n71762 , n417847 );
buf ( n418395 , n71763 );
buf ( n418396 , n418395 );
and ( n71766 , n71761 , n418396 );
and ( n71767 , n418252 , n418391 );
or ( n71768 , n71766 , n71767 );
buf ( n418400 , n71768 );
xor ( n71770 , n418067 , n418083 );
xor ( n71771 , n71770 , n418100 );
and ( n71772 , n418400 , n71771 );
and ( n71773 , n418232 , n418400 );
or ( n71774 , n71604 , n71772 , n71773 );
buf ( n418406 , n71774 );
xor ( n71776 , n418229 , n418406 );
buf ( n418408 , n59596 );
buf ( n418409 , n63625 );
and ( n71779 , n418408 , n418409 );
buf ( n418411 , n409146 );
buf ( n418412 , n63629 );
and ( n71782 , n418411 , n418412 );
nor ( n71783 , n71779 , n71782 );
buf ( n418415 , n71783 );
buf ( n418416 , n418415 );
buf ( n418417 , n410635 );
or ( n71787 , n418416 , n418417 );
buf ( n418419 , n418243 );
buf ( n418420 , n409504 );
or ( n71790 , n418419 , n418420 );
nand ( n71791 , n71787 , n71790 );
buf ( n418423 , n71791 );
buf ( n418424 , n418423 );
xor ( n71794 , n417797 , n417837 );
xor ( n71795 , n71794 , n417842 );
buf ( n418427 , n71795 );
buf ( n418428 , n418427 );
xor ( n71798 , n418424 , n418428 );
buf ( n418430 , n66359 );
buf ( n418431 , n405391 );
and ( n71801 , n418430 , n418431 );
buf ( n418433 , n413187 );
buf ( n418434 , n414664 );
and ( n71804 , n418433 , n418434 );
nor ( n71805 , n71801 , n71804 );
buf ( n418437 , n71805 );
buf ( n418438 , n418437 );
buf ( n418439 , n405407 );
or ( n71809 , n418438 , n418439 );
buf ( n418441 , n418362 );
buf ( n418442 , n405384 );
or ( n71812 , n418441 , n418442 );
nand ( n71813 , n71809 , n71812 );
buf ( n418445 , n71813 );
buf ( n418446 , n418445 );
buf ( n418447 , n414729 );
buf ( n418448 , n58061 );
or ( n71818 , n418447 , n418448 );
buf ( n418450 , n68002 );
buf ( n418451 , n56041 );
or ( n71821 , n418450 , n418451 );
nand ( n71822 , n71818 , n71821 );
buf ( n418454 , n71822 );
buf ( n418455 , n418454 );
not ( n71825 , n418455 );
buf ( n418457 , n71825 );
buf ( n418458 , n418457 );
buf ( n418459 , n403293 );
or ( n71829 , n418458 , n418459 );
buf ( n418461 , n417780 );
buf ( n418462 , n405476 );
or ( n71832 , n418461 , n418462 );
nand ( n71833 , n71829 , n71832 );
buf ( n418465 , n71833 );
buf ( n418466 , n418465 );
xor ( n71836 , n418446 , n418466 );
buf ( n418468 , n70389 );
buf ( n418469 , n55905 );
and ( n71839 , n418468 , n418469 );
buf ( n418471 , n417024 );
buf ( n418472 , n55895 );
and ( n71842 , n418471 , n418472 );
nor ( n71843 , n71839 , n71842 );
buf ( n418475 , n71843 );
buf ( n418476 , n418475 );
buf ( n418477 , n403120 );
or ( n71847 , n418476 , n418477 );
buf ( n418479 , n418260 );
buf ( n418480 , n403133 );
or ( n71850 , n418479 , n418480 );
nand ( n71851 , n71847 , n71850 );
buf ( n418483 , n71851 );
xor ( n71853 , n418285 , n418305 );
xor ( n71854 , n71853 , n418342 );
and ( n71855 , n418483 , n71854 );
buf ( n418487 , n403305 );
not ( n71857 , n418487 );
buf ( n418489 , n418454 );
not ( n71859 , n418489 );
or ( n71860 , n71857 , n71859 );
buf ( n418492 , n70195 );
buf ( n418493 , n56041 );
and ( n71863 , n418492 , n418493 );
buf ( n418495 , n416830 );
buf ( n418496 , n58061 );
and ( n71866 , n418495 , n418496 );
nor ( n71867 , n71863 , n71866 );
buf ( n418499 , n71867 );
buf ( n418500 , n418499 );
buf ( n418501 , n403293 );
or ( n71871 , n418500 , n418501 );
nand ( n71872 , n71860 , n71871 );
buf ( n418504 , n71872 );
xor ( n71874 , n418285 , n418305 );
xor ( n71875 , n71874 , n418342 );
and ( n71876 , n418504 , n71875 );
and ( n71877 , n418483 , n418504 );
or ( n71878 , n71855 , n71876 , n71877 );
buf ( n418510 , n71878 );
and ( n71880 , n71836 , n418510 );
and ( n71881 , n418446 , n418466 );
or ( n71882 , n71880 , n71881 );
buf ( n418514 , n71882 );
buf ( n418515 , n418514 );
and ( n71885 , n71798 , n418515 );
and ( n71886 , n418424 , n418428 );
or ( n71887 , n71885 , n71886 );
buf ( n418519 , n71887 );
buf ( n418520 , n418519 );
buf ( n418521 , n58200 );
buf ( n418522 , n66411 );
and ( n71892 , n418521 , n418522 );
buf ( n418524 , n58201 );
buf ( n418525 , n62496 );
and ( n71895 , n418524 , n418525 );
nor ( n71896 , n71892 , n71895 );
buf ( n418528 , n71896 );
buf ( n418529 , n418528 );
buf ( n418530 , n410724 );
or ( n71900 , n418529 , n418530 );
buf ( n418532 , n417648 );
buf ( n418533 , n410721 );
or ( n71903 , n418532 , n418533 );
nand ( n71904 , n71900 , n71903 );
buf ( n418536 , n71904 );
buf ( n418537 , n418536 );
xor ( n71907 , n418520 , n418537 );
xor ( n418539 , n417878 , n417903 );
xor ( n71909 , n418539 , n417955 );
buf ( n418541 , n71909 );
buf ( n418542 , n418541 );
and ( n71912 , n71907 , n418542 );
and ( n71913 , n418520 , n418537 );
or ( n71914 , n71912 , n71913 );
buf ( n418546 , n71914 );
xor ( n71916 , n417665 , n417852 );
xor ( n71917 , n71916 , n417960 );
buf ( n418549 , n71917 );
xor ( n71919 , n418546 , n418549 );
xor ( n71920 , n418067 , n418083 );
xor ( n71921 , n71920 , n418100 );
xor ( n71922 , n418232 , n418400 );
xor ( n71923 , n71921 , n71922 );
and ( n71924 , n71919 , n71923 );
and ( n71925 , n418546 , n418549 );
or ( n71926 , n71924 , n71925 );
buf ( n418558 , n71926 );
and ( n71928 , n71776 , n418558 );
and ( n71929 , n418229 , n418406 );
or ( n71930 , n71928 , n71929 );
buf ( n418562 , n71930 );
nand ( n71932 , n71593 , n418562 );
nand ( n71933 , n71589 , n71932 );
xor ( n71934 , n418173 , n418196 );
and ( n71935 , n71934 , n418216 );
and ( n71936 , n418173 , n418196 );
or ( n71937 , n71935 , n71936 );
buf ( n418569 , n71937 );
xor ( n71939 , n416923 , n70305 );
xor ( n71940 , n71939 , n417070 );
xor ( n71941 , n418179 , n418188 );
and ( n71942 , n71941 , n418193 );
and ( n71943 , n418179 , n418188 );
or ( n71944 , n71942 , n71943 );
buf ( n418576 , n71944 );
xor ( n71946 , n417202 , n417206 );
xor ( n71947 , n71946 , n417211 );
buf ( n418579 , n71947 );
xor ( n71949 , n418576 , n418579 );
xor ( n71950 , n71940 , n71949 );
xor ( n71951 , n418202 , n418208 );
and ( n71952 , n71951 , n418213 );
and ( n71953 , n418202 , n418208 );
or ( n71954 , n71952 , n71953 );
buf ( n418586 , n71954 );
or ( n71956 , n71950 , n418586 );
not ( n71957 , n71956 );
and ( n71958 , n418569 , n71957 );
nand ( n71959 , n71950 , n418586 );
not ( n71960 , n71959 );
and ( n71961 , n71960 , n418569 );
nor ( n71962 , n71958 , n71961 );
not ( n71963 , n71950 );
not ( n71964 , n418569 );
nand ( n71965 , n71963 , n71964 , n418586 );
not ( n71966 , n418586 );
nand ( n71967 , n71966 , n71964 , n71950 );
and ( n71968 , n71962 , n71965 , n71967 );
and ( n71969 , n71933 , n71968 );
not ( n71970 , n71933 );
not ( n71971 , n71968 );
and ( n71972 , n71970 , n71971 );
nor ( n71973 , n71969 , n71972 );
and ( n71974 , n71009 , n71973 );
not ( n71975 , n71009 );
not ( n71976 , n71973 );
and ( n71977 , n71975 , n71976 );
nor ( n71978 , n71974 , n71977 );
buf ( n418610 , n71978 );
buf ( n418611 , n43515 );
not ( n71981 , n418611 );
buf ( n418613 , n391027 );
not ( n71983 , n418613 );
buf ( n418615 , n412920 );
not ( n71985 , n418615 );
or ( n71986 , n71983 , n71985 );
buf ( n418618 , n12480 );
buf ( n418619 , n391024 );
nand ( n71989 , n418618 , n418619 );
buf ( n418621 , n71989 );
buf ( n418622 , n418621 );
nand ( n71992 , n71986 , n418622 );
buf ( n418624 , n71992 );
buf ( n418625 , n418624 );
not ( n71995 , n418625 );
or ( n71996 , n71981 , n71995 );
buf ( n418628 , n391027 );
not ( n71998 , n418628 );
buf ( n418630 , n410127 );
not ( n72000 , n418630 );
or ( n72001 , n71998 , n72000 );
buf ( n418633 , n28353 );
buf ( n418634 , n391024 );
nand ( n72004 , n418633 , n418634 );
buf ( n418636 , n72004 );
buf ( n418637 , n418636 );
nand ( n72007 , n72001 , n418637 );
buf ( n418639 , n72007 );
buf ( n418640 , n418639 );
buf ( n418641 , n43536 );
nand ( n72011 , n418640 , n418641 );
buf ( n418643 , n72011 );
buf ( n418644 , n418643 );
nand ( n72014 , n71996 , n418644 );
buf ( n418646 , n72014 );
buf ( n418647 , n418646 );
xor ( n72017 , n418610 , n418647 );
and ( n72018 , n394210 , n41365 );
not ( n72019 , n394210 );
and ( n72020 , n72019 , n410407 );
nor ( n72021 , n72018 , n72020 );
not ( n72022 , n72021 );
not ( n72023 , n41373 );
or ( n72024 , n72022 , n72023 );
or ( n72025 , n41341 , n392887 );
or ( n72026 , n392884 , n23841 );
nand ( n72027 , n72025 , n72026 );
or ( n72028 , n41332 , n72027 );
nand ( n72029 , n72024 , n72028 );
buf ( n418661 , n72029 );
and ( n72031 , n72017 , n418661 );
and ( n72032 , n418610 , n418647 );
or ( n72033 , n72031 , n72032 );
buf ( n418665 , n72033 );
buf ( n418666 , n418665 );
xor ( n72036 , n417609 , n418666 );
buf ( n418668 , n413643 );
not ( n72038 , n418668 );
buf ( n418670 , n417538 );
not ( n72040 , n418670 );
or ( n72041 , n72038 , n72040 );
buf ( n418673 , n44775 );
not ( n72043 , n418673 );
buf ( n418675 , n410400 );
not ( n72045 , n418675 );
or ( n72046 , n72043 , n72045 );
buf ( n418678 , n12471 );
buf ( n418679 , n44776 );
nand ( n72049 , n418678 , n418679 );
buf ( n418681 , n72049 );
buf ( n418682 , n418681 );
nand ( n72052 , n72046 , n418682 );
buf ( n418684 , n72052 );
buf ( n418685 , n418684 );
buf ( n418686 , n417542 );
nand ( n72056 , n418685 , n418686 );
buf ( n418688 , n72056 );
buf ( n418689 , n418688 );
nand ( n72059 , n72041 , n418689 );
buf ( n418691 , n72059 );
buf ( n418692 , n418691 );
and ( n72062 , n72036 , n418692 );
and ( n72063 , n417609 , n418666 );
or ( n72064 , n72062 , n72063 );
buf ( n418696 , n72064 );
buf ( n418697 , n418696 );
xor ( n72067 , n70938 , n418697 );
buf ( n418699 , n72067 );
buf ( n418700 , n418699 );
xor ( n72070 , n71590 , n71591 );
xor ( n72071 , n72070 , n418562 );
buf ( n418703 , n388068 );
not ( n72073 , n418703 );
buf ( n418705 , n40601 );
not ( n72075 , n418705 );
not ( n72076 , n42066 );
buf ( n418708 , n72076 );
not ( n72078 , n418708 );
or ( n72079 , n72075 , n72078 );
buf ( n418711 , n42066 );
buf ( n418712 , n40600 );
nand ( n72082 , n418711 , n418712 );
buf ( n418714 , n72082 );
buf ( n418715 , n418714 );
nand ( n72085 , n72079 , n418715 );
buf ( n418717 , n72085 );
buf ( n418718 , n418717 );
not ( n72088 , n418718 );
or ( n72089 , n72073 , n72088 );
buf ( n418721 , n40592 );
buf ( n418722 , n388722 );
not ( n72092 , n418722 );
buf ( n418724 , n389353 );
not ( n72094 , n418724 );
or ( n72095 , n72092 , n72094 );
buf ( n418727 , n41861 );
not ( n72097 , n418727 );
buf ( n418729 , n72097 );
buf ( n418730 , n418729 );
not ( n72100 , n418730 );
buf ( n418732 , n388722 );
not ( n72102 , n418732 );
buf ( n418734 , n72102 );
buf ( n418735 , n418734 );
nand ( n72105 , n72100 , n418735 );
buf ( n418737 , n72105 );
buf ( n418738 , n418737 );
nand ( n72108 , n72095 , n418738 );
buf ( n418740 , n72108 );
buf ( n418741 , n418740 );
nand ( n72111 , n418721 , n418741 );
buf ( n418743 , n72111 );
buf ( n418744 , n418743 );
nand ( n72114 , n72089 , n418744 );
buf ( n418746 , n72114 );
xor ( n72116 , n72071 , n418746 );
buf ( n418748 , n391443 );
buf ( n418749 , n371797 );
and ( n72119 , n418748 , n418749 );
not ( n72120 , n418748 );
buf ( n418752 , n417617 );
and ( n72122 , n72120 , n418752 );
nor ( n72123 , n72119 , n72122 );
buf ( n418755 , n72123 );
buf ( n418756 , n418755 );
not ( n72126 , n418756 );
buf ( n418758 , n388740 );
not ( n72128 , n418758 );
or ( n72129 , n72126 , n72128 );
buf ( n418761 , n417637 );
buf ( n418762 , n388803 );
nand ( n72132 , n418761 , n418762 );
buf ( n418764 , n72132 );
buf ( n418765 , n418764 );
nand ( n72135 , n72129 , n418765 );
buf ( n418767 , n72135 );
xor ( n72137 , n72116 , n418767 );
not ( n72138 , n72137 );
not ( n72139 , n72138 );
not ( n72140 , n66128 );
buf ( n418772 , n417572 );
not ( n72142 , n418772 );
buf ( n418774 , n41341 );
not ( n72144 , n418774 );
or ( n72145 , n72142 , n72144 );
buf ( n418777 , n64780 );
buf ( n418778 , n394814 );
nand ( n72148 , n418777 , n418778 );
buf ( n418780 , n72148 );
buf ( n418781 , n418780 );
nand ( n72151 , n72145 , n418781 );
buf ( n418783 , n72151 );
not ( n72153 , n418783 );
or ( n72154 , n72140 , n72153 );
buf ( n418786 , n72021 );
buf ( n418787 , n412976 );
nand ( n72157 , n418786 , n418787 );
buf ( n418789 , n72157 );
nand ( n72159 , n72154 , n418789 );
not ( n72160 , n72159 );
not ( n72161 , n72160 );
and ( n418793 , n72139 , n72161 );
not ( n72163 , n72159 );
nand ( n72164 , n72163 , n72138 );
buf ( n418796 , n392608 );
not ( n72166 , n418796 );
buf ( n418798 , n371797 );
not ( n72168 , n418798 );
or ( n72169 , n72166 , n72168 );
buf ( n418801 , n371800 );
buf ( n418802 , n392608 );
not ( n72172 , n418802 );
buf ( n418804 , n72172 );
buf ( n418805 , n418804 );
nand ( n72175 , n418801 , n418805 );
buf ( n418807 , n72175 );
buf ( n418808 , n418807 );
nand ( n72178 , n72169 , n418808 );
buf ( n418810 , n72178 );
buf ( n418811 , n418810 );
not ( n72181 , n418811 );
buf ( n418813 , n388740 );
not ( n72183 , n418813 );
or ( n72184 , n72181 , n72183 );
buf ( n418816 , n418755 );
buf ( n418817 , n388803 );
nand ( n72187 , n418816 , n418817 );
buf ( n418819 , n72187 );
buf ( n418820 , n418819 );
nand ( n72190 , n72184 , n418820 );
buf ( n418822 , n72190 );
buf ( n418823 , n418822 );
xor ( n72193 , n418252 , n418391 );
xor ( n72194 , n72193 , n418396 );
buf ( n418826 , n72194 );
buf ( n418827 , n62278 );
buf ( n418828 , n62177 );
and ( n72198 , n418827 , n418828 );
buf ( n418830 , n409474 );
buf ( n418831 , n62159 );
and ( n72201 , n418830 , n418831 );
nor ( n72202 , n72198 , n72201 );
buf ( n418834 , n72202 );
buf ( n418835 , n418834 );
buf ( n418836 , n409429 );
or ( n72206 , n418835 , n418836 );
buf ( n418838 , n417861 );
buf ( n418839 , n409170 );
or ( n72209 , n418838 , n418839 );
nand ( n72210 , n72206 , n72209 );
buf ( n418842 , n72210 );
xor ( n72212 , n418354 , n418370 );
xor ( n72213 , n72212 , n418387 );
and ( n72214 , n418842 , n72213 );
buf ( n418846 , n58352 );
buf ( n418847 , n66411 );
and ( n72217 , n418846 , n418847 );
buf ( n418849 , n406571 );
buf ( n418850 , n62496 );
and ( n72220 , n418849 , n418850 );
nor ( n72221 , n72217 , n72220 );
buf ( n418853 , n72221 );
buf ( n418854 , n418853 );
buf ( n418855 , n410724 );
or ( n72225 , n418854 , n418855 );
buf ( n418857 , n418528 );
buf ( n418858 , n410721 );
or ( n72228 , n418857 , n418858 );
nand ( n72229 , n72225 , n72228 );
buf ( n418861 , n72229 );
xor ( n72231 , n418354 , n418370 );
xor ( n72232 , n72231 , n418387 );
and ( n72233 , n418861 , n72232 );
and ( n72234 , n418842 , n418861 );
or ( n72235 , n72214 , n72233 , n72234 );
xor ( n72236 , n418826 , n72235 );
xor ( n72237 , n418520 , n418537 );
xor ( n72238 , n72237 , n418542 );
buf ( n418870 , n72238 );
and ( n72240 , n72236 , n418870 );
and ( n72241 , n418826 , n72235 );
or ( n72242 , n72240 , n72241 );
xor ( n72243 , n418546 , n418549 );
xor ( n72244 , n72243 , n71923 );
and ( n72245 , n72242 , n72244 );
buf ( n418877 , n67987 );
buf ( n418878 , n405391 );
and ( n72248 , n418877 , n418878 );
buf ( n418880 , n414714 );
buf ( n418881 , n405388 );
and ( n72251 , n418880 , n418881 );
nor ( n72252 , n72248 , n72251 );
buf ( n418884 , n72252 );
buf ( n418885 , n418884 );
buf ( n418886 , n405407 );
or ( n72256 , n418885 , n418886 );
buf ( n418888 , n418437 );
buf ( n418889 , n405384 );
or ( n72259 , n418888 , n418889 );
nand ( n72260 , n72256 , n72259 );
buf ( n418892 , n72260 );
buf ( n418893 , n418892 );
buf ( n418894 , n417729 );
buf ( n418895 , n55895 );
or ( n72265 , n418894 , n418895 );
buf ( n418897 , n71095 );
buf ( n418898 , n15287 );
or ( n72268 , n418897 , n418898 );
nand ( n72269 , n72265 , n72268 );
buf ( n418901 , n72269 );
buf ( n418902 , n418901 );
not ( n72272 , n418902 );
buf ( n418904 , n72272 );
buf ( n418905 , n418904 );
buf ( n418906 , n403120 );
or ( n72276 , n418905 , n418906 );
buf ( n418908 , n418475 );
buf ( n418909 , n403133 );
or ( n72279 , n418908 , n418909 );
nand ( n72280 , n72276 , n72279 );
buf ( n418912 , n72280 );
buf ( n418913 , n418912 );
xor ( n72283 , n418323 , n418340 );
buf ( n418915 , n72283 );
buf ( n418916 , n418915 );
xor ( n72286 , n418913 , n418916 );
buf ( n418918 , n403158 );
buf ( n418919 , n401678 );
not ( n72289 , n418919 );
buf ( n418921 , n72289 );
buf ( n418922 , n418921 );
buf ( n418923 , n71664 );
and ( n72293 , n418922 , n418923 );
buf ( n418925 , n401678 );
buf ( n418926 , n418298 );
and ( n72296 , n418925 , n418926 );
nor ( n72297 , n72293 , n72296 );
buf ( n418929 , n72297 );
buf ( n418930 , n418929 );
or ( n72300 , n418918 , n418930 );
buf ( n418932 , n418332 );
buf ( n418933 , n401660 );
or ( n72303 , n418932 , n418933 );
nand ( n72304 , n72300 , n72303 );
buf ( n418936 , n72304 );
buf ( n418937 , n418936 );
buf ( n418938 , n401623 );
xor ( n72308 , n54173 , n54172 );
buf ( n418940 , n72308 );
not ( n72310 , n418940 );
buf ( n418942 , n72310 );
buf ( n418943 , n418942 );
or ( n72313 , n418938 , n418943 );
buf ( n418945 , n401619 );
buf ( n418946 , n418315 );
or ( n72316 , n418945 , n418946 );
nand ( n72317 , n72313 , n72316 );
buf ( n418949 , n72317 );
buf ( n418950 , n418949 );
xor ( n72320 , n418937 , n418950 );
buf ( n418952 , n55875 );
not ( n72322 , n418952 );
buf ( n418954 , n418901 );
not ( n72324 , n418954 );
or ( n72325 , n72322 , n72324 );
buf ( n418957 , n403120 );
buf ( n418958 , n71088 );
buf ( n418959 , n15287 );
and ( n72329 , n418958 , n418959 );
buf ( n418961 , n417722 );
buf ( n418962 , n15290 );
and ( n72332 , n418961 , n418962 );
nor ( n72333 , n72329 , n72332 );
buf ( n418965 , n72333 );
buf ( n418966 , n418965 );
or ( n72336 , n418957 , n418966 );
nand ( n72337 , n72325 , n72336 );
buf ( n418969 , n72337 );
buf ( n418970 , n418969 );
and ( n72340 , n72320 , n418970 );
and ( n72341 , n418937 , n418950 );
or ( n72342 , n72340 , n72341 );
buf ( n418974 , n72342 );
buf ( n418975 , n418974 );
and ( n72345 , n72286 , n418975 );
and ( n72346 , n418913 , n418916 );
or ( n72347 , n72345 , n72346 );
buf ( n418979 , n72347 );
buf ( n418980 , n418979 );
xor ( n72350 , n418893 , n418980 );
buf ( n418982 , n59471 );
not ( n72352 , n418982 );
buf ( n418984 , n63707 );
buf ( n418985 , n59628 );
and ( n72355 , n418984 , n418985 );
buf ( n418987 , n413104 );
buf ( n418988 , n59457 );
and ( n72358 , n418987 , n418988 );
nor ( n72359 , n72355 , n72358 );
buf ( n418991 , n72359 );
buf ( n418992 , n418991 );
not ( n72362 , n418992 );
buf ( n418994 , n72362 );
buf ( n418995 , n418994 );
not ( n72365 , n418995 );
or ( n72366 , n72352 , n72365 );
buf ( n418998 , n66270 );
buf ( n418999 , n59628 );
and ( n72369 , n418998 , n418999 );
buf ( n419001 , n413098 );
buf ( n419002 , n59457 );
and ( n72372 , n419001 , n419002 );
nor ( n72373 , n72369 , n72372 );
buf ( n419005 , n72373 );
buf ( n419006 , n419005 );
buf ( n419007 , n59637 );
or ( n72377 , n419006 , n419007 );
nand ( n72378 , n72366 , n72377 );
buf ( n419010 , n72378 );
buf ( n419011 , n419010 );
and ( n72381 , n72350 , n419011 );
and ( n72382 , n418893 , n418980 );
or ( n72383 , n72381 , n72382 );
buf ( n419015 , n72383 );
buf ( n419016 , n419015 );
buf ( n419017 , n62467 );
buf ( n419018 , n62177 );
and ( n72388 , n419017 , n419018 );
buf ( n419020 , n409468 );
buf ( n419021 , n62159 );
and ( n72391 , n419020 , n419021 );
nor ( n72392 , n72388 , n72391 );
buf ( n419024 , n72392 );
buf ( n419025 , n419024 );
buf ( n419026 , n409429 );
or ( n72396 , n419025 , n419026 );
buf ( n419028 , n418834 );
buf ( n419029 , n409170 );
or ( n72399 , n419028 , n419029 );
nand ( n72400 , n72396 , n72399 );
buf ( n419032 , n72400 );
buf ( n419033 , n419032 );
xor ( n72403 , n419016 , n419033 );
xor ( n72404 , n418446 , n418466 );
xor ( n72405 , n72404 , n418510 );
buf ( n419037 , n72405 );
buf ( n419038 , n419037 );
and ( n72408 , n72403 , n419038 );
and ( n72409 , n419016 , n419033 );
or ( n419041 , n72408 , n72409 );
buf ( n419042 , n419041 );
buf ( n419043 , n419042 );
buf ( n419044 , n418991 );
buf ( n419045 , n59637 );
or ( n72415 , n419044 , n419045 );
buf ( n419047 , n418379 );
buf ( n419048 , n59467 );
or ( n72418 , n419047 , n419048 );
nand ( n72419 , n72415 , n72418 );
buf ( n419051 , n72419 );
buf ( n419052 , n419051 );
xor ( n72422 , n418269 , n418346 );
xor ( n72423 , n72422 , n418350 );
buf ( n419055 , n72423 );
buf ( n419056 , n419055 );
xor ( n72426 , n419052 , n419056 );
buf ( n419058 , n409507 );
not ( n72428 , n419058 );
buf ( n419060 , n62139 );
buf ( n419061 , n63625 );
and ( n72431 , n419060 , n419061 );
buf ( n419063 , n409140 );
buf ( n419064 , n63629 );
and ( n72434 , n419063 , n419064 );
nor ( n72435 , n72431 , n72434 );
buf ( n419067 , n72435 );
buf ( n419068 , n419067 );
not ( n72438 , n419068 );
buf ( n419070 , n72438 );
buf ( n419071 , n419070 );
not ( n72441 , n419071 );
or ( n72442 , n72428 , n72441 );
buf ( n419074 , n418415 );
buf ( n419075 , n409504 );
or ( n72445 , n419074 , n419075 );
nand ( n72446 , n72442 , n72445 );
buf ( n419078 , n72446 );
buf ( n419079 , n419078 );
and ( n72449 , n72426 , n419079 );
and ( n72450 , n419052 , n419056 );
or ( n72451 , n72449 , n72450 );
buf ( n419083 , n72451 );
buf ( n419084 , n419083 );
xor ( n72454 , n419043 , n419084 );
xor ( n72455 , n418424 , n418428 );
xor ( n72456 , n72455 , n418515 );
buf ( n419088 , n72456 );
buf ( n419089 , n419088 );
and ( n72459 , n72454 , n419089 );
and ( n72460 , n419043 , n419084 );
or ( n72461 , n72459 , n72460 );
buf ( n419093 , n72461 );
xor ( n72463 , n418826 , n72235 );
xor ( n72464 , n72463 , n418870 );
and ( n72465 , n419093 , n72464 );
xor ( n72466 , n418354 , n418370 );
xor ( n72467 , n72466 , n418387 );
xor ( n72468 , n418842 , n418861 );
xor ( n72469 , n72467 , n72468 );
buf ( n419101 , n68002 );
buf ( n419102 , n405391 );
and ( n72472 , n419101 , n419102 );
buf ( n419104 , n414729 );
buf ( n419105 , n405388 );
and ( n72475 , n419104 , n419105 );
nor ( n72476 , n72472 , n72475 );
buf ( n419108 , n72476 );
buf ( n419109 , n419108 );
buf ( n419110 , n405407 );
or ( n72480 , n419109 , n419110 );
buf ( n419112 , n418884 );
buf ( n419113 , n405384 );
or ( n72483 , n419112 , n419113 );
nand ( n72484 , n72480 , n72483 );
buf ( n419116 , n72484 );
buf ( n419117 , n419116 );
buf ( n419118 , n70210 );
buf ( n419119 , n56041 );
and ( n72489 , n419118 , n419119 );
buf ( n419121 , n416845 );
buf ( n419122 , n403298 );
and ( n72492 , n419121 , n419122 );
nor ( n72493 , n72489 , n72492 );
buf ( n419125 , n72493 );
buf ( n419126 , n419125 );
buf ( n419127 , n403293 );
or ( n72497 , n419126 , n419127 );
buf ( n419129 , n418499 );
buf ( n419130 , n405476 );
or ( n72500 , n419129 , n419130 );
nand ( n72501 , n72497 , n72500 );
buf ( n419133 , n72501 );
buf ( n419134 , n419133 );
xor ( n72504 , n419117 , n419134 );
xor ( n72505 , n418913 , n418916 );
xor ( n72506 , n72505 , n418975 );
buf ( n419138 , n72506 );
buf ( n419139 , n419138 );
and ( n72509 , n72504 , n419139 );
and ( n72510 , n419117 , n419134 );
or ( n72511 , n72509 , n72510 );
buf ( n419143 , n72511 );
xor ( n72513 , n418285 , n418305 );
xor ( n72514 , n72513 , n418342 );
xor ( n72515 , n418483 , n418504 );
xor ( n72516 , n72514 , n72515 );
xor ( n72517 , n419143 , n72516 );
buf ( n419149 , n409173 );
not ( n72519 , n419149 );
buf ( n419151 , n63564 );
buf ( n419152 , n62177 );
and ( n72522 , n419151 , n419152 );
buf ( n419154 , n413073 );
buf ( n419155 , n62159 );
and ( n72525 , n419154 , n419155 );
nor ( n72526 , n72522 , n72525 );
buf ( n419158 , n72526 );
buf ( n419159 , n419158 );
not ( n72529 , n419159 );
buf ( n419161 , n72529 );
buf ( n419162 , n419161 );
not ( n72532 , n419162 );
or ( n72533 , n72519 , n72532 );
buf ( n419165 , n419024 );
buf ( n419166 , n409170 );
or ( n72536 , n419165 , n419166 );
nand ( n72537 , n72533 , n72536 );
buf ( n419169 , n72537 );
and ( n72539 , n72517 , n419169 );
and ( n72540 , n419143 , n72516 );
or ( n72541 , n72539 , n72540 );
buf ( n419173 , n72541 );
buf ( n419174 , n59435 );
buf ( n419175 , n66411 );
and ( n72545 , n419174 , n419175 );
buf ( n419177 , n406565 );
buf ( n419178 , n62496 );
and ( n72548 , n419177 , n419178 );
nor ( n72549 , n72545 , n72548 );
buf ( n419181 , n72549 );
buf ( n419182 , n419181 );
buf ( n419183 , n410724 );
or ( n72553 , n419182 , n419183 );
buf ( n419185 , n418853 );
buf ( n419186 , n410721 );
or ( n72556 , n419185 , n419186 );
nand ( n72557 , n72553 , n72556 );
buf ( n419189 , n72557 );
buf ( n419190 , n419189 );
xor ( n72560 , n419173 , n419190 );
xor ( n72561 , n419052 , n419056 );
xor ( n72562 , n72561 , n419079 );
buf ( n419194 , n72562 );
buf ( n419195 , n419194 );
and ( n72565 , n72560 , n419195 );
and ( n72566 , n419173 , n419190 );
or ( n72567 , n72565 , n72566 );
buf ( n419199 , n72567 );
xor ( n72569 , n72469 , n419199 );
xor ( n72570 , n419043 , n419084 );
xor ( n72571 , n72570 , n419089 );
buf ( n419203 , n72571 );
and ( n72573 , n72569 , n419203 );
and ( n72574 , n72469 , n419199 );
or ( n72575 , n72573 , n72574 );
xor ( n72576 , n418826 , n72235 );
xor ( n72577 , n72576 , n418870 );
and ( n72578 , n72575 , n72577 );
and ( n72579 , n419093 , n72575 );
or ( n72580 , n72465 , n72578 , n72579 );
xor ( n72581 , n418546 , n418549 );
xor ( n72582 , n72581 , n71923 );
and ( n72583 , n72580 , n72582 );
and ( n72584 , n72242 , n72580 );
or ( n72585 , n72245 , n72583 , n72584 );
buf ( n419217 , n72585 );
xor ( n72587 , n418229 , n418406 );
xor ( n72588 , n72587 , n418558 );
buf ( n419220 , n72588 );
buf ( n419221 , n419220 );
xor ( n72591 , n419217 , n419221 );
and ( n72592 , n389338 , n418734 );
not ( n72593 , n389338 );
and ( n72594 , n72593 , n388722 );
or ( n72595 , n72592 , n72594 );
buf ( n419227 , n72595 );
not ( n72597 , n419227 );
buf ( n419229 , n40592 );
not ( n72599 , n419229 );
or ( n72600 , n72597 , n72599 );
buf ( n419232 , n418740 );
buf ( n419233 , n388068 );
nand ( n72603 , n419232 , n419233 );
buf ( n419235 , n72603 );
buf ( n419236 , n419235 );
nand ( n72606 , n72600 , n419236 );
buf ( n419238 , n72606 );
buf ( n419239 , n419238 );
xor ( n72609 , n72591 , n419239 );
buf ( n419241 , n72609 );
buf ( n419242 , n419241 );
xor ( n72612 , n418823 , n419242 );
buf ( n419244 , n43515 );
not ( n72614 , n419244 );
buf ( n419246 , n391018 );
not ( n72616 , n419246 );
buf ( n419248 , n27320 );
not ( n72618 , n419248 );
buf ( n419250 , n72618 );
buf ( n419251 , n419250 );
not ( n72621 , n419251 );
or ( n72622 , n72616 , n72621 );
buf ( n419254 , n412892 );
not ( n72624 , n419254 );
buf ( n419256 , n391021 );
nand ( n72626 , n72624 , n419256 );
buf ( n419258 , n72626 );
buf ( n419259 , n419258 );
nand ( n72629 , n72622 , n419259 );
buf ( n419261 , n72629 );
buf ( n419262 , n419261 );
not ( n72632 , n419262 );
or ( n72633 , n72614 , n72632 );
buf ( n419265 , n391018 );
not ( n72635 , n419265 );
buf ( n419267 , n42065 );
not ( n72637 , n419267 );
or ( n72638 , n72635 , n72637 );
not ( n72639 , n42065 );
buf ( n419271 , n72639 );
buf ( n419272 , n391021 );
nand ( n72642 , n419271 , n419272 );
buf ( n419274 , n72642 );
buf ( n419275 , n419274 );
nand ( n72645 , n72638 , n419275 );
buf ( n419277 , n72645 );
buf ( n419278 , n419277 );
buf ( n419279 , n43536 );
nand ( n72649 , n419278 , n419279 );
buf ( n419281 , n72649 );
buf ( n419282 , n419281 );
nand ( n419283 , n72633 , n419282 );
buf ( n419284 , n419283 );
buf ( n419285 , n419284 );
and ( n72655 , n72612 , n419285 );
and ( n72656 , n418823 , n419242 );
or ( n72657 , n72655 , n72656 );
buf ( n419289 , n72657 );
buf ( n72659 , n419289 );
and ( n72660 , n72164 , n72659 );
nor ( n72661 , n418793 , n72660 );
buf ( n419293 , n72661 );
not ( n72663 , n419293 );
buf ( n419295 , n72663 );
buf ( n419296 , n419295 );
not ( n72666 , n419296 );
buf ( n419298 , n413643 );
not ( n72668 , n419298 );
buf ( n419300 , n418684 );
not ( n72670 , n419300 );
or ( n72671 , n72668 , n72670 );
buf ( n419303 , n44775 );
not ( n72673 , n419303 );
buf ( n419305 , n388227 );
not ( n72675 , n419305 );
or ( n72676 , n72673 , n72675 );
buf ( n419308 , n406821 );
buf ( n419309 , n44776 );
nand ( n72679 , n419308 , n419309 );
buf ( n419311 , n72679 );
buf ( n419312 , n419311 );
nand ( n72682 , n72676 , n419312 );
buf ( n419314 , n72682 );
buf ( n419315 , n419314 );
buf ( n419316 , n417542 );
nand ( n72686 , n419315 , n419316 );
buf ( n419318 , n72686 );
buf ( n419319 , n419318 );
nand ( n72689 , n72671 , n419319 );
buf ( n419321 , n72689 );
buf ( n419322 , n419321 );
not ( n72692 , n419322 );
or ( n72693 , n72666 , n72692 );
buf ( n419325 , n419321 );
buf ( n419326 , n419295 );
or ( n72696 , n419325 , n419326 );
xor ( n72697 , n418610 , n418647 );
xor ( n72698 , n72697 , n418661 );
buf ( n419330 , n72698 );
buf ( n419331 , n419330 );
nand ( n72701 , n72696 , n419331 );
buf ( n419333 , n72701 );
buf ( n419334 , n419333 );
nand ( n72704 , n72693 , n419334 );
buf ( n419336 , n72704 );
buf ( n419337 , n419336 );
buf ( n419338 , n399274 );
buf ( n419339 , n399167 );
and ( n72709 , n419338 , n419339 );
not ( n72710 , n419338 );
buf ( n419342 , n398298 );
and ( n72712 , n72710 , n419342 );
or ( n72713 , n72709 , n72712 );
buf ( n419345 , n72713 );
buf ( n419346 , n419345 );
not ( n72716 , n419346 );
buf ( n419348 , n72716 );
buf ( n419349 , n419348 );
not ( n72719 , n419349 );
buf ( n419351 , n389122 );
not ( n72721 , n419351 );
or ( n72722 , n72719 , n72721 );
buf ( n419354 , n55543 );
not ( n72724 , n419354 );
buf ( n419356 , n398298 );
not ( n72726 , n419356 );
or ( n72727 , n72724 , n72726 );
buf ( n419359 , n24049 );
buf ( n419360 , n51185 );
nand ( n72730 , n419359 , n419360 );
buf ( n419362 , n72730 );
buf ( n419363 , n419362 );
nand ( n72733 , n72727 , n419363 );
buf ( n419365 , n72733 );
buf ( n419366 , n419365 );
buf ( n419367 , n46921 );
nand ( n72737 , n419366 , n419367 );
buf ( n419369 , n72737 );
buf ( n419370 , n419369 );
nand ( n72740 , n72722 , n419370 );
buf ( n419372 , n72740 );
buf ( n419373 , n419372 );
xor ( n72743 , n419337 , n419373 );
buf ( n419375 , n395362 );
not ( n72745 , n419375 );
buf ( n419377 , n47863 );
not ( n72747 , n419377 );
buf ( n419379 , n388373 );
not ( n72749 , n419379 );
or ( n72750 , n72747 , n72749 );
buf ( n419382 , n397077 );
buf ( n419383 , n47863 );
not ( n72753 , n419383 );
buf ( n419385 , n72753 );
buf ( n419386 , n419385 );
nand ( n72756 , n419382 , n419386 );
buf ( n419388 , n72756 );
buf ( n419389 , n419388 );
nand ( n72759 , n72750 , n419389 );
buf ( n419391 , n72759 );
buf ( n419392 , n419391 );
not ( n72762 , n419392 );
or ( n72763 , n72745 , n72762 );
buf ( n419395 , n47863 );
not ( n72765 , n419395 );
buf ( n419397 , n394330 );
not ( n72767 , n419397 );
or ( n72768 , n72765 , n72767 );
buf ( n419400 , n388646 );
buf ( n419401 , n419385 );
nand ( n72771 , n419400 , n419401 );
buf ( n419403 , n72771 );
buf ( n419404 , n419403 );
nand ( n72774 , n72768 , n419404 );
buf ( n419406 , n72774 );
buf ( n419407 , n419406 );
buf ( n419408 , n395349 );
nand ( n72778 , n419407 , n419408 );
buf ( n419410 , n72778 );
buf ( n419411 , n419410 );
nand ( n72781 , n72763 , n419411 );
buf ( n419413 , n72781 );
buf ( n419414 , n419413 );
and ( n72784 , n72743 , n419414 );
and ( n72785 , n419337 , n419373 );
or ( n72786 , n72784 , n72785 );
buf ( n419418 , n72786 );
buf ( n419419 , n419418 );
xor ( n72789 , n418700 , n419419 );
buf ( n419421 , n61577 );
not ( n72791 , n419421 );
buf ( n419423 , n42825 );
not ( n72793 , n419423 );
not ( n72794 , n47891 );
buf ( n419426 , n72794 );
not ( n72796 , n419426 );
and ( n72797 , n72793 , n72796 );
buf ( n419429 , n42825 );
buf ( n419430 , n72794 );
and ( n72800 , n419429 , n419430 );
nor ( n72801 , n72797 , n72800 );
buf ( n419433 , n72801 );
buf ( n419434 , n419433 );
not ( n72804 , n419434 );
buf ( n419436 , n72804 );
buf ( n419437 , n419436 );
not ( n72807 , n419437 );
or ( n72808 , n72791 , n72807 );
and ( n72809 , n47891 , n388445 );
not ( n72810 , n47891 );
and ( n72811 , n72810 , n40819 );
or ( n72812 , n72809 , n72811 );
buf ( n419444 , n72812 );
buf ( n419445 , n50579 );
nand ( n72815 , n419444 , n419445 );
buf ( n419447 , n72815 );
buf ( n419448 , n419447 );
nand ( n72818 , n72808 , n419448 );
buf ( n419450 , n72818 );
buf ( n419451 , n419450 );
xor ( n72821 , n72789 , n419451 );
buf ( n419453 , n72821 );
buf ( n419454 , n419453 );
xor ( n72824 , n417609 , n418666 );
xor ( n72825 , n72824 , n418692 );
buf ( n419457 , n72825 );
buf ( n419458 , n419457 );
buf ( n419459 , n55055 );
not ( n72829 , n419459 );
buf ( n419461 , n46906 );
not ( n72831 , n419461 );
or ( n72832 , n72829 , n72831 );
buf ( n419464 , n49653 );
buf ( n419465 , n404855 );
nand ( n72835 , n419464 , n419465 );
buf ( n419467 , n72835 );
buf ( n419468 , n419467 );
nand ( n72838 , n72832 , n419468 );
buf ( n419470 , n72838 );
buf ( n419471 , n419470 );
not ( n72841 , n419471 );
buf ( n419473 , n399031 );
not ( n72843 , n419473 );
or ( n72844 , n72841 , n72843 );
buf ( n419476 , n400042 );
buf ( n419477 , n54957 );
and ( n72847 , n419476 , n419477 );
not ( n72848 , n419476 );
buf ( n419480 , n49660 );
and ( n72850 , n72848 , n419480 );
nor ( n72851 , n72847 , n72850 );
buf ( n419483 , n72851 );
buf ( n419484 , n419483 );
buf ( n419485 , n395199 );
nand ( n72855 , n419484 , n419485 );
buf ( n419487 , n72855 );
buf ( n419488 , n419487 );
nand ( n72858 , n72844 , n419488 );
buf ( n419490 , n72858 );
buf ( n419491 , n419490 );
xor ( n72861 , n419458 , n419491 );
buf ( n419493 , n388068 );
not ( n72863 , n419493 );
and ( n72864 , n40601 , n417349 );
not ( n72865 , n40601 );
and ( n72866 , n72865 , n28353 );
or ( n72867 , n72864 , n72866 );
buf ( n419499 , n72867 );
not ( n72869 , n419499 );
or ( n72870 , n72863 , n72869 );
buf ( n419502 , n40601 );
not ( n72872 , n419502 );
buf ( n419504 , n419250 );
not ( n72874 , n419504 );
or ( n72875 , n72872 , n72874 );
nand ( n72876 , n27320 , n40600 );
buf ( n419508 , n72876 );
nand ( n72878 , n72875 , n419508 );
buf ( n419510 , n72878 );
buf ( n419511 , n419510 );
buf ( n419512 , n40592 );
nand ( n72882 , n419511 , n419512 );
buf ( n419514 , n72882 );
buf ( n419515 , n419514 );
nand ( n72885 , n72870 , n419515 );
buf ( n419517 , n72885 );
buf ( n419518 , n419517 );
not ( n419519 , n71971 );
not ( n72889 , n71009 );
not ( n72890 , n72889 );
or ( n72891 , n419519 , n72890 );
not ( n72892 , n71008 );
nand ( n72893 , n72892 , n417628 , n71968 );
nand ( n72894 , n72893 , n71933 );
nand ( n72895 , n72891 , n72894 );
buf ( n419527 , n72895 );
xor ( n72897 , n419518 , n419527 );
buf ( n419529 , n66128 );
not ( n72899 , n419529 );
buf ( n419531 , n72899 );
buf ( n419532 , n419531 );
buf ( n419533 , n72027 );
or ( n72903 , n419532 , n419533 );
buf ( n419535 , n392611 );
buf ( n419536 , n410407 );
xnor ( n72906 , n419535 , n419536 );
buf ( n419538 , n72906 );
buf ( n419539 , n419538 );
not ( n72909 , n419539 );
buf ( n419541 , n72909 );
buf ( n419542 , n419541 );
buf ( n419543 , n41332 );
or ( n72913 , n419542 , n419543 );
nand ( n72914 , n72903 , n72913 );
buf ( n419546 , n72914 );
buf ( n419547 , n419546 );
xor ( n72917 , n72897 , n419547 );
buf ( n419549 , n72917 );
buf ( n419550 , n419549 );
buf ( n419551 , n397489 );
not ( n72921 , n419551 );
buf ( n419553 , n56919 );
not ( n72923 , n419553 );
or ( n72924 , n72921 , n72923 );
buf ( n419556 , n41559 );
buf ( n419557 , n397492 );
nand ( n72927 , n419556 , n419557 );
buf ( n419559 , n72927 );
buf ( n419560 , n419559 );
nand ( n72930 , n72924 , n419560 );
buf ( n419562 , n72930 );
buf ( n419563 , n419562 );
not ( n72933 , n419563 );
buf ( n419565 , n390432 );
not ( n72935 , n419565 );
or ( n72936 , n72933 , n72935 );
buf ( n419568 , n49117 );
not ( n72938 , n419568 );
buf ( n419570 , n51822 );
not ( n72940 , n419570 );
or ( n72941 , n72938 , n72940 );
buf ( n419573 , n57505 );
buf ( n419574 , n67126 );
nand ( n72944 , n419573 , n419574 );
buf ( n419576 , n72944 );
buf ( n419577 , n419576 );
nand ( n72947 , n72941 , n419577 );
buf ( n419579 , n72947 );
buf ( n419580 , n419579 );
buf ( n419581 , n42924 );
nand ( n72951 , n419580 , n419581 );
buf ( n419583 , n72951 );
buf ( n419584 , n419583 );
nand ( n72954 , n72936 , n419584 );
buf ( n419586 , n72954 );
buf ( n419587 , n419586 );
xor ( n72957 , n419550 , n419587 );
xor ( n72958 , n419217 , n419221 );
and ( n72959 , n72958 , n419239 );
and ( n72960 , n419217 , n419221 );
or ( n72961 , n72959 , n72960 );
buf ( n419593 , n72961 );
buf ( n419594 , n419593 );
buf ( n419595 , n392884 );
not ( n72965 , n419595 );
buf ( n419597 , n62006 );
not ( n72967 , n419597 );
or ( n72968 , n72965 , n72967 );
buf ( n419600 , n64268 );
buf ( n419601 , n392881 );
nand ( n72971 , n419600 , n419601 );
buf ( n419603 , n72971 );
buf ( n419604 , n419603 );
nand ( n72974 , n72968 , n419604 );
buf ( n419606 , n72974 );
buf ( n419607 , n419606 );
not ( n72977 , n419607 );
buf ( n419609 , n45076 );
not ( n72979 , n419609 );
or ( n72980 , n72977 , n72979 );
and ( n72981 , n392611 , n68376 );
not ( n72982 , n392611 );
and ( n72983 , n72982 , n64268 );
or ( n72984 , n72981 , n72983 );
buf ( n419616 , n72984 );
buf ( n419617 , n41664 );
nand ( n72987 , n419616 , n419617 );
buf ( n419619 , n72987 );
buf ( n419620 , n419619 );
nand ( n72990 , n72980 , n419620 );
buf ( n419622 , n72990 );
buf ( n419623 , n419622 );
xor ( n72993 , n419594 , n419623 );
buf ( n419625 , n43515 );
not ( n72995 , n419625 );
buf ( n419627 , n418639 );
not ( n72997 , n419627 );
or ( n72998 , n72995 , n72997 );
buf ( n419630 , n419261 );
buf ( n419631 , n43536 );
nand ( n73001 , n419630 , n419631 );
buf ( n419633 , n73001 );
buf ( n419634 , n419633 );
nand ( n73004 , n72998 , n419634 );
buf ( n419636 , n73004 );
buf ( n419637 , n419636 );
and ( n73007 , n72993 , n419637 );
and ( n73008 , n419594 , n419623 );
or ( n73009 , n73007 , n73008 );
buf ( n419641 , n73009 );
buf ( n419642 , n419641 );
buf ( n419643 , n388068 );
not ( n73013 , n419643 );
buf ( n419645 , n419510 );
not ( n73015 , n419645 );
or ( n73016 , n73013 , n73015 );
buf ( n419648 , n418717 );
buf ( n419649 , n40592 );
nand ( n73019 , n419648 , n419649 );
buf ( n419651 , n73019 );
buf ( n419652 , n419651 );
nand ( n73022 , n73016 , n419652 );
buf ( n419654 , n73022 );
buf ( n419655 , n72984 );
not ( n73025 , n419655 );
not ( n73026 , n41707 );
buf ( n419658 , n73026 );
not ( n73028 , n419658 );
or ( n73029 , n73025 , n73028 );
buf ( n419661 , n391446 );
not ( n73031 , n419661 );
buf ( n419663 , n62006 );
not ( n73033 , n419663 );
or ( n73034 , n73031 , n73033 );
buf ( n419666 , n24116 );
buf ( n419667 , n391443 );
nand ( n73037 , n419666 , n419667 );
buf ( n419669 , n73037 );
buf ( n419670 , n419669 );
nand ( n73040 , n73034 , n419670 );
buf ( n419672 , n73040 );
buf ( n419673 , n419672 );
buf ( n419674 , n41664 );
nand ( n73044 , n419673 , n419674 );
buf ( n419676 , n73044 );
buf ( n419677 , n419676 );
nand ( n73047 , n73029 , n419677 );
buf ( n419679 , n73047 );
xor ( n73049 , n419654 , n419679 );
xor ( n73050 , n72071 , n418746 );
and ( n73051 , n73050 , n418767 );
and ( n73052 , n72071 , n418746 );
or ( n73053 , n73051 , n73052 );
xor ( n73054 , n73049 , n73053 );
buf ( n419686 , n73054 );
xor ( n73056 , n419642 , n419686 );
buf ( n419688 , n49117 );
not ( n73058 , n419688 );
buf ( n419690 , n40653 );
not ( n73060 , n419690 );
or ( n73061 , n73058 , n73060 );
buf ( n419693 , n407936 );
buf ( n419694 , n67126 );
nand ( n73064 , n419693 , n419694 );
buf ( n419696 , n73064 );
buf ( n419697 , n419696 );
nand ( n73067 , n73061 , n419697 );
buf ( n419699 , n73067 );
buf ( n419700 , n419699 );
not ( n73070 , n419700 );
buf ( n419702 , n406422 );
not ( n73072 , n419702 );
or ( n73073 , n73070 , n73072 );
buf ( n419705 , n417584 );
buf ( n419706 , n409076 );
nand ( n73076 , n419705 , n419706 );
buf ( n419708 , n73076 );
buf ( n419709 , n419708 );
nand ( n73079 , n73073 , n419709 );
buf ( n419711 , n73079 );
buf ( n419712 , n419711 );
and ( n73082 , n73056 , n419712 );
and ( n73083 , n419642 , n419686 );
or ( n73084 , n73082 , n73083 );
buf ( n419716 , n73084 );
buf ( n419717 , n419716 );
xor ( n73087 , n72957 , n419717 );
buf ( n419719 , n73087 );
buf ( n419720 , n419719 );
and ( n73090 , n72861 , n419720 );
and ( n73091 , n419458 , n419491 );
or ( n73092 , n73090 , n73091 );
buf ( n419724 , n73092 );
buf ( n419725 , n419724 );
buf ( n419726 , n419365 );
not ( n73096 , n419726 );
buf ( n419728 , n389122 );
not ( n73098 , n419728 );
or ( n73099 , n73096 , n73098 );
buf ( n419731 , n397489 );
not ( n73101 , n419731 );
buf ( n419733 , n45391 );
not ( n73103 , n419733 );
or ( n73104 , n73101 , n73103 );
buf ( n419736 , n24049 );
buf ( n419737 , n397492 );
nand ( n73107 , n419736 , n419737 );
buf ( n419739 , n73107 );
buf ( n419740 , n419739 );
nand ( n73110 , n73104 , n419740 );
buf ( n419742 , n73110 );
buf ( n419743 , n419742 );
buf ( n419744 , n41563 );
nand ( n73114 , n419743 , n419744 );
buf ( n419746 , n73114 );
buf ( n419747 , n419746 );
nand ( n73117 , n73099 , n419747 );
buf ( n419749 , n73117 );
not ( n73119 , n419749 );
buf ( n419751 , n45954 );
not ( n73121 , n419751 );
buf ( n419753 , n393369 );
not ( n73123 , n419753 );
buf ( n419755 , n27301 );
not ( n73125 , n419755 );
buf ( n419757 , n73125 );
buf ( n419758 , n419757 );
not ( n73128 , n419758 );
or ( n73129 , n73123 , n73128 );
buf ( n419761 , n393154 );
buf ( n419762 , n393381 );
nand ( n73132 , n419761 , n419762 );
buf ( n419764 , n73132 );
buf ( n419765 , n419764 );
nand ( n73135 , n73129 , n419765 );
buf ( n419767 , n73135 );
buf ( n419768 , n419767 );
not ( n73138 , n419768 );
or ( n73139 , n73121 , n73138 );
buf ( n419771 , n393381 );
buf ( n419772 , n46478 );
and ( n73142 , n419771 , n419772 );
not ( n73143 , n419771 );
buf ( n419775 , n49686 );
and ( n73145 , n73143 , n419775 );
or ( n73146 , n73142 , n73145 );
buf ( n419778 , n73146 );
buf ( n419779 , n419778 );
not ( n73149 , n419779 );
buf ( n419781 , n45949 );
nand ( n73151 , n73149 , n419781 );
buf ( n419783 , n73151 );
buf ( n419784 , n419783 );
nand ( n73154 , n73139 , n419784 );
buf ( n419786 , n73154 );
not ( n73156 , n419786 );
xor ( n73157 , n73119 , n73156 );
not ( n73158 , n395469 );
and ( n73159 , n49661 , n399274 );
not ( n73160 , n49661 );
and ( n73161 , n73160 , n399283 );
or ( n73162 , n73159 , n73161 );
not ( n73163 , n73162 );
or ( n73164 , n73158 , n73163 );
nand ( n73165 , n419483 , n397102 );
nand ( n73166 , n73164 , n73165 );
xor ( n73167 , n73157 , n73166 );
buf ( n419799 , n73167 );
xor ( n73169 , n419725 , n419799 );
buf ( n419801 , C0 );
buf ( n419802 , n419801 );
xor ( n73196 , n73169 , n419802 );
buf ( n419804 , n73196 );
buf ( n419805 , n419804 );
xor ( n73199 , n419454 , n419805 );
buf ( n419807 , n393381 );
not ( n73201 , n419807 );
buf ( n419809 , n403042 );
not ( n73203 , n419809 );
or ( n73204 , n73201 , n73203 );
buf ( n419812 , n28644 );
not ( n73206 , n419812 );
buf ( n419814 , n393369 );
nand ( n73208 , n73206 , n419814 );
buf ( n419816 , n73208 );
buf ( n419817 , n419816 );
nand ( n73211 , n73204 , n419817 );
buf ( n419819 , n73211 );
and ( n73213 , n419819 , n45954 );
and ( n73214 , n410400 , n393369 );
not ( n73215 , n410400 );
and ( n73216 , n73215 , n393381 );
or ( n73217 , n73214 , n73216 );
and ( n73218 , n73217 , n45949 );
nor ( n73219 , n73213 , n73218 );
buf ( n419827 , n73219 );
not ( n73221 , n419827 );
buf ( n419829 , n395199 );
buf ( n419830 , n358975 );
nand ( n73224 , n419829 , n419830 );
buf ( n419832 , n73224 );
buf ( n419833 , n419832 );
not ( n73227 , n419833 );
or ( n73228 , n73221 , n73227 );
and ( n73229 , n399274 , n51822 );
not ( n73230 , n399274 );
and ( n73231 , n73230 , n53252 );
or ( n73232 , n73229 , n73231 );
buf ( n419840 , n73232 );
not ( n73234 , n419840 );
buf ( n419842 , n390429 );
not ( n73236 , n419842 );
or ( n73237 , n73234 , n73236 );
and ( n73238 , n55543 , n24071 );
not ( n73239 , n55543 );
and ( n73240 , n73239 , n41559 );
or ( n73241 , n73238 , n73240 );
buf ( n419849 , n73241 );
buf ( n419850 , n42924 );
nand ( n73244 , n419849 , n419850 );
buf ( n419852 , n73244 );
buf ( n419853 , n419852 );
nand ( n73247 , n73237 , n419853 );
buf ( n419855 , n73247 );
buf ( n419856 , n419855 );
nand ( n73250 , n73228 , n419856 );
buf ( n419858 , n73250 );
buf ( n419859 , n419858 );
buf ( n419860 , n73219 );
not ( n73254 , n419860 );
buf ( n419862 , n419832 );
not ( n73256 , n419862 );
buf ( n419864 , n73256 );
buf ( n419865 , n419864 );
nand ( n73259 , n73254 , n419865 );
buf ( n419867 , n73259 );
buf ( n419868 , n419867 );
nand ( n73262 , n419859 , n419868 );
buf ( n419870 , n73262 );
buf ( n419871 , n419870 );
and ( n73265 , n419321 , n72661 );
not ( n73266 , n419321 );
and ( n73267 , n73266 , n419295 );
or ( n73268 , n73265 , n73267 );
xor ( n73269 , n73268 , n419330 );
buf ( n419877 , n73269 );
xor ( n73271 , n419871 , n419877 );
and ( n73272 , n24116 , n394814 );
not ( n73273 , n24116 );
and ( n73274 , n73273 , n417572 );
or ( n73275 , n73272 , n73274 );
buf ( n419883 , n73275 );
not ( n73277 , n419883 );
buf ( n419885 , n416762 );
not ( n73279 , n419885 );
or ( n73280 , n73277 , n73279 );
buf ( n419888 , n394210 );
not ( n73282 , n419888 );
buf ( n419890 , n41323 );
not ( n73284 , n419890 );
or ( n73285 , n73282 , n73284 );
buf ( n419893 , n41324 );
buf ( n419894 , n394219 );
nand ( n73288 , n419893 , n419894 );
buf ( n419896 , n73288 );
buf ( n419897 , n419896 );
nand ( n73291 , n73285 , n419897 );
buf ( n419899 , n73291 );
buf ( n419900 , n419899 );
buf ( n419901 , n41664 );
nand ( n73295 , n419900 , n419901 );
buf ( n419903 , n73295 );
buf ( n419904 , n419903 );
nand ( n73298 , n73280 , n419904 );
buf ( n419906 , n73298 );
buf ( n419907 , n419906 );
xor ( n73301 , n418546 , n418549 );
xor ( n73302 , n73301 , n71923 );
xor ( n73303 , n72242 , n72580 );
xor ( n73304 , n73302 , n73303 );
buf ( n419912 , n73304 );
and ( n73306 , n391440 , n388722 );
not ( n73307 , n391440 );
and ( n73308 , n73307 , n388080 );
nor ( n73309 , n73306 , n73308 );
buf ( n419917 , n73309 );
not ( n73311 , n419917 );
buf ( n419919 , n73311 );
buf ( n419920 , n419919 );
not ( n73314 , n419920 );
buf ( n419922 , n40592 );
not ( n73316 , n419922 );
or ( n73317 , n73314 , n73316 );
buf ( n419925 , n72595 );
buf ( n419926 , n388068 );
nand ( n73320 , n419925 , n419926 );
buf ( n419928 , n73320 );
buf ( n419929 , n419928 );
nand ( n73323 , n73317 , n419929 );
buf ( n419931 , n73323 );
buf ( n419932 , n419931 );
xor ( n73326 , n419912 , n419932 );
buf ( n419934 , n43515 );
not ( n73328 , n419934 );
buf ( n419936 , n419277 );
not ( n73330 , n419936 );
or ( n73331 , n73328 , n73330 );
buf ( n419939 , n391018 );
not ( n73333 , n419939 );
buf ( n419941 , n418729 );
not ( n73335 , n419941 );
or ( n73336 , n73333 , n73335 );
buf ( n419944 , n41861 );
buf ( n419945 , n391021 );
nand ( n73339 , n419944 , n419945 );
buf ( n419947 , n73339 );
buf ( n419948 , n419947 );
nand ( n419949 , n73336 , n419948 );
buf ( n419950 , n419949 );
buf ( n419951 , n419950 );
buf ( n419952 , n43536 );
nand ( n73346 , n419951 , n419952 );
buf ( n419954 , n73346 );
buf ( n419955 , n419954 );
nand ( n73349 , n73331 , n419955 );
buf ( n419957 , n73349 );
buf ( n419958 , n419957 );
xor ( n73352 , n73326 , n419958 );
buf ( n419960 , n73352 );
buf ( n419961 , n419960 );
xor ( n73355 , n419907 , n419961 );
buf ( n419963 , n413643 );
not ( n73357 , n419963 );
and ( n73358 , n44775 , n417349 );
not ( n73359 , n44775 );
and ( n73360 , n73359 , n28353 );
or ( n73361 , n73358 , n73360 );
buf ( n419969 , n73361 );
not ( n73363 , n419969 );
or ( n73364 , n73357 , n73363 );
and ( n73365 , n44775 , n412892 );
not ( n73366 , n44775 );
and ( n73367 , n73366 , n27320 );
or ( n73368 , n73365 , n73367 );
buf ( n419976 , n73368 );
buf ( n419977 , n417542 );
nand ( n73371 , n419976 , n419977 );
buf ( n419979 , n73371 );
buf ( n419980 , n419979 );
nand ( n73374 , n73364 , n419980 );
buf ( n419982 , n73374 );
buf ( n419983 , n419982 );
and ( n73377 , n73355 , n419983 );
and ( n73378 , n419907 , n419961 );
or ( n73379 , n73377 , n73378 );
buf ( n419987 , n73379 );
buf ( n419988 , n419987 );
buf ( n419989 , n55543 );
not ( n73383 , n419989 );
buf ( n419991 , n404601 );
not ( n73385 , n419991 );
or ( n73386 , n73383 , n73385 );
buf ( n419994 , n407928 );
buf ( n419995 , n51185 );
nand ( n73389 , n419994 , n419995 );
buf ( n419997 , n73389 );
buf ( n419998 , n419997 );
nand ( n73392 , n73386 , n419998 );
buf ( n420000 , n73392 );
buf ( n420001 , n420000 );
not ( n73395 , n420001 );
buf ( n420003 , n409082 );
not ( n73397 , n420003 );
or ( n73398 , n73395 , n73397 );
buf ( n420006 , n397489 );
not ( n73400 , n420006 );
buf ( n420008 , n404601 );
not ( n73402 , n420008 );
or ( n73403 , n73400 , n73402 );
buf ( n420011 , n407928 );
buf ( n420012 , n397492 );
nand ( n73406 , n420011 , n420012 );
buf ( n420014 , n73406 );
buf ( n420015 , n420014 );
nand ( n73409 , n73403 , n420015 );
buf ( n420017 , n73409 );
buf ( n420018 , n420017 );
buf ( n420019 , n409076 );
nand ( n73413 , n420018 , n420019 );
buf ( n420021 , n73413 );
buf ( n420022 , n420021 );
nand ( n73416 , n73398 , n420022 );
buf ( n420024 , n73416 );
buf ( n420025 , n420024 );
xor ( n73419 , n419988 , n420025 );
xor ( n73420 , n419912 , n419932 );
and ( n73421 , n73420 , n419958 );
and ( n73422 , n419912 , n419932 );
or ( n73423 , n73421 , n73422 );
buf ( n420031 , n73423 );
buf ( n420032 , n420031 );
buf ( n420033 , n419899 );
not ( n73427 , n420033 );
buf ( n420035 , n73026 );
not ( n73429 , n420035 );
or ( n73430 , n73427 , n73429 );
buf ( n420038 , n419606 );
buf ( n420039 , n41664 );
nand ( n73433 , n420038 , n420039 );
buf ( n420041 , n73433 );
buf ( n420042 , n420041 );
nand ( n73436 , n73430 , n420042 );
buf ( n420044 , n73436 );
buf ( n420045 , n420044 );
xor ( n73439 , n420032 , n420045 );
xor ( n73440 , n418823 , n419242 );
xor ( n73441 , n73440 , n419285 );
buf ( n420049 , n73441 );
buf ( n420050 , n420049 );
xor ( n73444 , n73439 , n420050 );
buf ( n420052 , n73444 );
buf ( n420053 , n420052 );
and ( n73447 , n73419 , n420053 );
and ( n73448 , n419988 , n420025 );
or ( n73449 , n73447 , n73448 );
buf ( n420057 , n73449 );
buf ( n420058 , n420057 );
buf ( n420059 , n395359 );
not ( n73453 , n420059 );
buf ( n420061 , n47863 );
not ( n73455 , n420061 );
buf ( n420063 , n46478 );
not ( n73457 , n420063 );
or ( n73458 , n73455 , n73457 );
buf ( n420066 , n49686 );
buf ( n420067 , n419385 );
nand ( n73461 , n420066 , n420067 );
buf ( n420069 , n73461 );
buf ( n420070 , n420069 );
nand ( n73464 , n73458 , n420070 );
buf ( n420072 , n73464 );
buf ( n420073 , n420072 );
not ( n73467 , n420073 );
or ( n73468 , n73453 , n73467 );
buf ( n420076 , n47863 );
not ( n73470 , n420076 );
buf ( n420078 , n388566 );
not ( n73472 , n420078 );
or ( n73473 , n73470 , n73472 );
buf ( n420081 , n402836 );
not ( n73475 , n420081 );
buf ( n420083 , n419385 );
nand ( n73477 , n73475 , n420083 );
buf ( n420085 , n73477 );
buf ( n420086 , n420085 );
nand ( n73480 , n73473 , n420086 );
buf ( n420088 , n73480 );
buf ( n420089 , n420088 );
buf ( n420090 , n395346 );
nand ( n73484 , n420089 , n420090 );
buf ( n420092 , n73484 );
buf ( n420093 , n420092 );
nand ( n73487 , n73468 , n420093 );
buf ( n420095 , n73487 );
buf ( n420096 , n420095 );
xor ( n73490 , n420058 , n420096 );
xor ( n73491 , n419594 , n419623 );
xor ( n73492 , n73491 , n419637 );
buf ( n420100 , n73492 );
buf ( n420101 , n420100 );
buf ( n420102 , n420017 );
not ( n73496 , n420102 );
buf ( n420104 , n60872 );
not ( n73498 , n420104 );
or ( n73499 , n73496 , n73498 );
buf ( n420107 , n419699 );
buf ( n420108 , n47726 );
nand ( n73502 , n420107 , n420108 );
buf ( n420110 , n73502 );
buf ( n420111 , n420110 );
nand ( n73505 , n73499 , n420111 );
buf ( n420113 , n73505 );
buf ( n420114 , n420113 );
xor ( n73508 , n420101 , n420114 );
buf ( n420116 , n413643 );
not ( n73510 , n420116 );
buf ( n420118 , n419314 );
not ( n73512 , n420118 );
or ( n73513 , n73510 , n73512 );
buf ( n420121 , n412920 );
not ( n73515 , n420121 );
buf ( n420123 , n44776 );
nand ( n73517 , n73515 , n420123 );
buf ( n420125 , n73517 );
not ( n73519 , n420125 );
nand ( n73520 , n412920 , n44775 );
not ( n73521 , n73520 );
or ( n73522 , n73519 , n73521 );
nand ( n73523 , n73522 , n417542 );
buf ( n420131 , n73523 );
nand ( n73525 , n73513 , n420131 );
buf ( n420133 , n73525 );
buf ( n420134 , n420133 );
xor ( n73528 , n73508 , n420134 );
buf ( n420136 , n73528 );
buf ( n420137 , n420136 );
and ( n73531 , n73490 , n420137 );
and ( n73532 , n420058 , n420096 );
or ( n73533 , n73531 , n73532 );
buf ( n420141 , n73533 );
buf ( n420142 , n420141 );
and ( n73536 , n73271 , n420142 );
and ( n73537 , n419871 , n419877 );
or ( n73538 , n73536 , n73537 );
buf ( n420146 , n73538 );
buf ( n420147 , n420146 );
not ( n73541 , n420147 );
buf ( n420149 , n45954 );
not ( n73543 , n420149 );
not ( n73544 , n393369 );
not ( n73545 , n388566 );
or ( n73546 , n73544 , n73545 );
buf ( n420154 , n27258 );
buf ( n420155 , n393381 );
nand ( n73549 , n420154 , n420155 );
buf ( n420157 , n73549 );
nand ( n73551 , n73546 , n420157 );
buf ( n420159 , n73551 );
not ( n73553 , n420159 );
or ( n73554 , n73543 , n73553 );
buf ( n420162 , n419819 );
buf ( n420163 , n45949 );
nand ( n73557 , n420162 , n420163 );
buf ( n420165 , n73557 );
buf ( n420166 , n420165 );
nand ( n420167 , n73554 , n420166 );
buf ( n420168 , n420167 );
buf ( n420169 , n420168 );
not ( n73563 , n420169 );
buf ( n420171 , n38956 );
not ( n73565 , n420171 );
buf ( n420173 , n398298 );
not ( n73567 , n420173 );
or ( n73568 , n73565 , n73567 );
buf ( n420176 , n358975 );
nand ( n73570 , n73568 , n420176 );
buf ( n420178 , n73570 );
buf ( n420179 , n420178 );
buf ( n420180 , n22982 );
buf ( n420181 , n24049 );
buf ( n420182 , n23988 );
nand ( n73576 , n420181 , n420182 );
buf ( n420184 , n73576 );
buf ( n420185 , n420184 );
nand ( n73579 , n420179 , n420180 , n420185 );
buf ( n420187 , n73579 );
buf ( n420188 , n420187 );
nand ( n73582 , n73563 , n420188 );
buf ( n420190 , n73582 );
not ( n73584 , n420190 );
buf ( n420192 , n73241 );
not ( n73586 , n420192 );
buf ( n420194 , n390432 );
not ( n73588 , n420194 );
or ( n73589 , n73586 , n73588 );
buf ( n420197 , n419562 );
buf ( n420198 , n42924 );
nand ( n73592 , n420197 , n420198 );
buf ( n420200 , n73592 );
buf ( n420201 , n420200 );
nand ( n73595 , n73589 , n420201 );
buf ( n420203 , n73595 );
not ( n73597 , n420203 );
or ( n73598 , n73584 , n73597 );
buf ( n420206 , n420187 );
not ( n73600 , n420206 );
buf ( n420208 , n420168 );
nand ( n73602 , n73600 , n420208 );
buf ( n420210 , n73602 );
nand ( n73604 , n73598 , n420210 );
buf ( n420212 , n73604 );
xor ( n73606 , n417215 , n417218 );
xor ( n73607 , n73606 , n417222 );
xor ( n73608 , n416923 , n70305 );
xor ( n73609 , n73608 , n417070 );
and ( n73610 , n418576 , n73609 );
xor ( n73611 , n416923 , n70305 );
xor ( n73612 , n73611 , n417070 );
and ( n73613 , n418579 , n73612 );
and ( n73614 , n418576 , n418579 );
or ( n73615 , n73610 , n73613 , n73614 );
not ( n73616 , n418569 );
not ( n73617 , n71956 );
or ( n73618 , n73616 , n73617 );
nand ( n73619 , n73618 , n71959 );
xor ( n73620 , n73615 , n73619 );
xor ( n73621 , n73607 , n73620 );
buf ( n420229 , n73621 );
buf ( n420230 , n417624 );
not ( n73624 , n420230 );
buf ( n420232 , n388740 );
not ( n73626 , n420232 );
or ( n73627 , n73624 , n73626 );
buf ( n420235 , n371784 );
buf ( n420236 , n72639 );
and ( n73630 , n420235 , n420236 );
not ( n73631 , n420235 );
buf ( n420239 , n42065 );
and ( n73633 , n73631 , n420239 );
nor ( n73634 , n73630 , n73633 );
buf ( n420242 , n73634 );
buf ( n420243 , n420242 );
buf ( n420244 , n388803 );
nand ( n73638 , n420243 , n420244 );
buf ( n420246 , n73638 );
buf ( n420247 , n420246 );
nand ( n73641 , n73627 , n420247 );
buf ( n420249 , n73641 );
buf ( n420250 , n420249 );
xor ( n73644 , n420229 , n420250 );
buf ( n420252 , n419672 );
not ( n73646 , n420252 );
buf ( n420254 , n416762 );
not ( n73648 , n420254 );
or ( n73649 , n73646 , n73648 );
buf ( n420257 , n389341 );
not ( n73651 , n420257 );
buf ( n420259 , n68376 );
not ( n73653 , n420259 );
or ( n73654 , n73651 , n73653 );
buf ( n420262 , n24116 );
buf ( n420263 , n393185 );
nand ( n73657 , n420262 , n420263 );
buf ( n420265 , n73657 );
buf ( n420266 , n420265 );
nand ( n73660 , n73654 , n420266 );
buf ( n420268 , n73660 );
buf ( n420269 , n420268 );
buf ( n420270 , n41664 );
nand ( n73664 , n420269 , n420270 );
buf ( n420272 , n73664 );
buf ( n420273 , n420272 );
nand ( n73667 , n73649 , n420273 );
buf ( n420275 , n73667 );
buf ( n420276 , n420275 );
xor ( n73670 , n73644 , n420276 );
buf ( n420278 , n73670 );
buf ( n420279 , n420278 );
not ( n73673 , n419679 );
not ( n73674 , n419654 );
nand ( n73675 , n73673 , n73674 );
not ( n73676 , n73675 );
not ( n73677 , n73053 );
or ( n73678 , n73676 , n73677 );
not ( n73679 , n73674 );
nand ( n73680 , n73679 , n419679 );
nand ( n73681 , n73678 , n73680 );
buf ( n420289 , n73681 );
xor ( n73683 , n420279 , n420289 );
buf ( n420291 , n43515 );
not ( n73685 , n420291 );
buf ( n420293 , n411504 );
not ( n73687 , n420293 );
buf ( n420295 , n406824 );
not ( n73689 , n420295 );
or ( n73690 , n73687 , n73689 );
buf ( n420298 , n388230 );
buf ( n420299 , n391024 );
nand ( n73693 , n420298 , n420299 );
buf ( n420301 , n73693 );
buf ( n420302 , n420301 );
nand ( n73696 , n73690 , n420302 );
buf ( n420304 , n73696 );
buf ( n420305 , n420304 );
not ( n73699 , n420305 );
or ( n73700 , n73685 , n73699 );
buf ( n420308 , n418624 );
buf ( n420309 , n43536 );
nand ( n73703 , n420308 , n420309 );
buf ( n420311 , n73703 );
buf ( n420312 , n420311 );
nand ( n73706 , n73700 , n420312 );
buf ( n420314 , n73706 );
buf ( n420315 , n420314 );
xor ( n73709 , n73683 , n420315 );
buf ( n420317 , n73709 );
buf ( n420318 , n420317 );
buf ( n420319 , n37923 );
buf ( n420320 , n402819 );
nor ( n73714 , n420319 , n420320 );
buf ( n420322 , n73714 );
buf ( n420323 , n420322 );
xor ( n73717 , n420318 , n420323 );
buf ( n420325 , n45949 );
not ( n73719 , n420325 );
buf ( n420327 , n73551 );
not ( n73721 , n420327 );
or ( n73722 , n73719 , n73721 );
buf ( n420330 , n419778 );
buf ( n420331 , n393409 );
or ( n73725 , n420330 , n420331 );
nand ( n73726 , n73722 , n73725 );
buf ( n420334 , n73726 );
buf ( n420335 , n420334 );
xor ( n73729 , n73717 , n420335 );
buf ( n420337 , n73729 );
buf ( n420338 , n420337 );
xor ( n73732 , n420212 , n420338 );
buf ( n420340 , n50579 );
not ( n73734 , n420340 );
buf ( n420342 , n47891 );
buf ( n420343 , n390673 );
and ( n73737 , n420342 , n420343 );
not ( n73738 , n420342 );
buf ( n420346 , n388409 );
and ( n73740 , n73738 , n420346 );
nor ( n73741 , n73737 , n73740 );
buf ( n420349 , n73741 );
buf ( n420350 , n420349 );
not ( n73744 , n420350 );
or ( n73745 , n73734 , n73744 );
buf ( n420353 , n72812 );
buf ( n420354 , n61577 );
nand ( n73748 , n420353 , n420354 );
buf ( n420356 , n73748 );
buf ( n420357 , n420356 );
nand ( n73751 , n73745 , n420357 );
buf ( n420359 , n73751 );
buf ( n420360 , n420359 );
xor ( n73754 , n73732 , n420360 );
buf ( n420362 , n73754 );
buf ( n420363 , n420362 );
not ( n73757 , n420363 );
or ( n73758 , n73541 , n73757 );
buf ( n420366 , n420146 );
buf ( n420367 , n420362 );
or ( n73761 , n420366 , n420367 );
nand ( n73762 , n420190 , n420210 );
xor ( n73763 , n73762 , n420203 );
buf ( n420371 , n73763 );
not ( n73765 , n420371 );
buf ( n420373 , n61577 );
not ( n73767 , n420373 );
buf ( n420375 , n420349 );
not ( n73769 , n420375 );
or ( n73770 , n73767 , n73769 );
buf ( n420378 , n72794 );
buf ( n420379 , n397072 );
and ( n73773 , n420378 , n420379 );
not ( n73774 , n420378 );
buf ( n420382 , n388370 );
and ( n73776 , n73774 , n420382 );
nor ( n73777 , n73773 , n73776 );
buf ( n420385 , n73777 );
buf ( n420386 , n420385 );
buf ( n420387 , n50579 );
nand ( n73781 , n420386 , n420387 );
buf ( n420389 , n73781 );
buf ( n420390 , n420389 );
nand ( n73784 , n73770 , n420390 );
buf ( n420392 , n73784 );
buf ( n420393 , n420392 );
not ( n73787 , n420393 );
buf ( n420395 , n73787 );
buf ( n420396 , n420395 );
not ( n73790 , n420396 );
or ( n73791 , n73765 , n73790 );
xor ( n73792 , n420101 , n420114 );
and ( n73793 , n73792 , n420134 );
and ( n73794 , n420101 , n420114 );
or ( n73795 , n73793 , n73794 );
buf ( n420403 , n73795 );
buf ( n420404 , n420403 );
xor ( n73798 , n419642 , n419686 );
xor ( n73799 , n73798 , n419712 );
buf ( n420407 , n73799 );
buf ( n420408 , n420407 );
xor ( n73802 , n420404 , n420408 );
xor ( n73803 , n420032 , n420045 );
and ( n73804 , n73803 , n420050 );
and ( n73805 , n420032 , n420045 );
or ( n73806 , n73804 , n73805 );
buf ( n420414 , n73806 );
and ( n73808 , n72138 , n419289 );
not ( n73809 , n72138 );
not ( n73810 , n419289 );
and ( n73811 , n73809 , n73810 );
nor ( n73812 , n73808 , n73811 );
and ( n73813 , n73812 , n72160 );
not ( n73814 , n73812 );
and ( n73815 , n73814 , n72159 );
nor ( n73816 , n73813 , n73815 );
xor ( n73817 , n420414 , n73816 );
buf ( n420425 , n392884 );
not ( n73819 , n420425 );
buf ( n420427 , n371787 );
not ( n73821 , n420427 );
or ( n73822 , n73819 , n73821 );
buf ( n420430 , n371784 );
buf ( n420431 , n392881 );
nand ( n73825 , n420430 , n420431 );
buf ( n420433 , n73825 );
buf ( n420434 , n420433 );
nand ( n73828 , n73822 , n420434 );
buf ( n420436 , n73828 );
not ( n73830 , n420436 );
not ( n73831 , n388740 );
or ( n73832 , n73830 , n73831 );
buf ( n420440 , n418810 );
buf ( n420441 , n388803 );
nand ( n73835 , n420440 , n420441 );
buf ( n420443 , n73835 );
nand ( n73837 , n73832 , n420443 );
not ( n73838 , n73837 );
xor ( n73839 , n418826 , n72235 );
xor ( n73840 , n73839 , n418870 );
xor ( n73841 , n419093 , n72575 );
xor ( n73842 , n73840 , n73841 );
buf ( n420450 , n73842 );
xor ( n73844 , n419016 , n419033 );
xor ( n73845 , n73844 , n419038 );
buf ( n420453 , n73845 );
buf ( n420454 , n420453 );
buf ( n420455 , n62278 );
buf ( n420456 , n63625 );
and ( n73850 , n420455 , n420456 );
buf ( n420458 , n409474 );
buf ( n420459 , n63629 );
and ( n73853 , n420458 , n420459 );
nor ( n73854 , n73850 , n73853 );
buf ( n420462 , n73854 );
buf ( n420463 , n420462 );
buf ( n420464 , n410635 );
or ( n73858 , n420463 , n420464 );
buf ( n420466 , n419067 );
buf ( n420467 , n409504 );
or ( n73861 , n420466 , n420467 );
nand ( n73862 , n73858 , n73861 );
buf ( n420470 , n73862 );
buf ( n420471 , n420470 );
xor ( n73865 , n418893 , n418980 );
xor ( n73866 , n73865 , n419011 );
buf ( n420474 , n73866 );
buf ( n420475 , n420474 );
xor ( n73869 , n420471 , n420475 );
buf ( n420477 , n348158 );
not ( n73871 , n420477 );
buf ( n420479 , n419181 );
not ( n73873 , n420479 );
buf ( n420481 , n73873 );
buf ( n420482 , n420481 );
not ( n73876 , n420482 );
or ( n73877 , n73871 , n73876 );
buf ( n420485 , n59596 );
buf ( n420486 , n66411 );
and ( n73880 , n420485 , n420486 );
buf ( n420488 , n409146 );
buf ( n420489 , n62496 );
and ( n73883 , n420488 , n420489 );
nor ( n73884 , n73880 , n73883 );
buf ( n420492 , n73884 );
buf ( n420493 , n420492 );
buf ( n420494 , n410724 );
or ( n73888 , n420493 , n420494 );
nand ( n73889 , n73877 , n73888 );
buf ( n420497 , n73889 );
buf ( n420498 , n420497 );
and ( n73892 , n73869 , n420498 );
and ( n73893 , n420471 , n420475 );
or ( n73894 , n73892 , n73893 );
buf ( n420502 , n73894 );
buf ( n420503 , n420502 );
xor ( n73897 , n420454 , n420503 );
buf ( n420505 , n66359 );
buf ( n420506 , n59628 );
and ( n73900 , n420505 , n420506 );
buf ( n420508 , n413187 );
buf ( n420509 , n59457 );
and ( n73903 , n420508 , n420509 );
nor ( n73904 , n73900 , n73903 );
buf ( n420512 , n73904 );
buf ( n420513 , n420512 );
buf ( n420514 , n59637 );
or ( n73908 , n420513 , n420514 );
buf ( n420516 , n419005 );
buf ( n420517 , n59467 );
or ( n73911 , n420516 , n420517 );
nand ( n73912 , n73908 , n73911 );
buf ( n420520 , n73912 );
buf ( n420521 , n420520 );
buf ( n420522 , n70389 );
buf ( n420523 , n56041 );
and ( n73917 , n420522 , n420523 );
buf ( n420525 , n417024 );
buf ( n420526 , n403298 );
and ( n73920 , n420525 , n420526 );
nor ( n73921 , n73917 , n73920 );
buf ( n420529 , n73921 );
buf ( n420530 , n420529 );
buf ( n420531 , n403293 );
or ( n73925 , n420530 , n420531 );
buf ( n420533 , n419125 );
buf ( n420534 , n405476 );
or ( n73928 , n420533 , n420534 );
nand ( n73929 , n73925 , n73928 );
buf ( n420537 , n73929 );
buf ( n420538 , n420537 );
buf ( n420539 , n403158 );
buf ( n420540 , n401689 );
buf ( n420541 , n71681 );
and ( n73935 , n420540 , n420541 );
buf ( n420543 , n401678 );
buf ( n420544 , n418315 );
and ( n73938 , n420543 , n420544 );
nor ( n73939 , n73935 , n73938 );
buf ( n420547 , n73939 );
buf ( n420548 , n420547 );
or ( n73942 , n420539 , n420548 );
buf ( n420550 , n418929 );
buf ( n420551 , n403167 );
or ( n73945 , n420550 , n420551 );
nand ( n73946 , n73942 , n73945 );
buf ( n420554 , n73946 );
buf ( n420555 , n420554 );
buf ( n420556 , n15287 );
buf ( n420557 , n71170 );
and ( n73951 , n420556 , n420557 );
buf ( n420559 , n55895 );
buf ( n420560 , n417804 );
and ( n73954 , n420559 , n420560 );
nor ( n73955 , n73951 , n73954 );
buf ( n420563 , n73955 );
buf ( n420564 , n420563 );
not ( n73958 , n420564 );
buf ( n420566 , n73958 );
buf ( n420567 , n420566 );
not ( n73961 , n420567 );
buf ( n420569 , n403123 );
not ( n73963 , n420569 );
or ( n73964 , n73961 , n73963 );
buf ( n420572 , n418965 );
buf ( n420573 , n403133 );
or ( n73967 , n420572 , n420573 );
nand ( n73968 , n73964 , n73967 );
buf ( n420576 , n73968 );
buf ( n420577 , n420576 );
and ( n73971 , n420555 , n420577 );
buf ( n420579 , n73971 );
buf ( n420580 , n420579 );
xor ( n73974 , n420538 , n420580 );
xor ( n73975 , n418937 , n418950 );
xor ( n73976 , n73975 , n418970 );
buf ( n420584 , n73976 );
buf ( n420585 , n420584 );
and ( n73979 , n73974 , n420585 );
and ( n73980 , n420538 , n420580 );
or ( n73981 , n73979 , n73980 );
buf ( n420589 , n73981 );
buf ( n420590 , n420589 );
xor ( n73984 , n420521 , n420590 );
buf ( n420592 , n71095 );
buf ( n420593 , n56041 );
and ( n73987 , n420592 , n420593 );
buf ( n420595 , n417729 );
buf ( n420596 , n403298 );
and ( n73990 , n420595 , n420596 );
nor ( n73991 , n73987 , n73990 );
buf ( n420599 , n73991 );
buf ( n420600 , n420599 );
buf ( n420601 , n403293 );
or ( n73995 , n420600 , n420601 );
buf ( n420603 , n420529 );
buf ( n420604 , n405476 );
or ( n73998 , n420603 , n420604 );
nand ( n73999 , n73995 , n73998 );
buf ( n420607 , n73999 );
buf ( n420608 , n401623 );
and ( n74002 , n54173 , n622 );
buf ( n420610 , n74002 );
not ( n74004 , n420610 );
buf ( n420612 , n74004 );
buf ( n420613 , n420612 );
or ( n74007 , n420608 , n420613 );
buf ( n420615 , n403092 );
buf ( n420616 , n418942 );
or ( n74010 , n420615 , n420616 );
nand ( n74011 , n74007 , n74010 );
buf ( n420619 , n74011 );
xor ( n74013 , n420607 , n420619 );
xor ( n74014 , n420555 , n420577 );
buf ( n420622 , n74014 );
and ( n74016 , n74013 , n420622 );
and ( n74017 , n420607 , n420619 );
or ( n74018 , n74016 , n74017 );
buf ( n420626 , n70195 );
buf ( n420627 , n405391 );
and ( n74021 , n420626 , n420627 );
buf ( n420629 , n416830 );
buf ( n420630 , n405388 );
and ( n74024 , n420629 , n420630 );
nor ( n74025 , n74021 , n74024 );
buf ( n420633 , n74025 );
buf ( n420634 , n420633 );
buf ( n420635 , n405407 );
or ( n74029 , n420634 , n420635 );
buf ( n420637 , n419108 );
buf ( n420638 , n405384 );
or ( n74032 , n420637 , n420638 );
nand ( n74033 , n74029 , n74032 );
buf ( n420641 , n74033 );
xor ( n74035 , n74018 , n420641 );
buf ( n420643 , n59468 );
not ( n74037 , n420643 );
buf ( n420645 , n414714 );
buf ( n420646 , n58223 );
or ( n74040 , n420645 , n420646 );
buf ( n420648 , n67987 );
buf ( n420649 , n14083 );
or ( n74043 , n420648 , n420649 );
nand ( n74044 , n74040 , n74043 );
buf ( n420652 , n74044 );
buf ( n420653 , n420652 );
not ( n74047 , n420653 );
or ( n74048 , n74037 , n74047 );
buf ( n420656 , n420512 );
buf ( n420657 , n59467 );
or ( n74051 , n420656 , n420657 );
nand ( n74052 , n74048 , n74051 );
buf ( n420660 , n74052 );
and ( n74054 , n74035 , n420660 );
and ( n74055 , n74018 , n420641 );
or ( n74056 , n74054 , n74055 );
buf ( n420664 , n74056 );
and ( n74058 , n73984 , n420664 );
and ( n74059 , n420521 , n420590 );
or ( n74060 , n74058 , n74059 );
buf ( n420668 , n74060 );
xor ( n74062 , n419143 , n72516 );
xor ( n74063 , n74062 , n419169 );
and ( n74064 , n420668 , n74063 );
xor ( n74065 , n419117 , n419134 );
xor ( n74066 , n74065 , n419139 );
buf ( n420674 , n74066 );
buf ( n420675 , n420674 );
buf ( n420676 , n63707 );
buf ( n420677 , n62177 );
and ( n74071 , n420676 , n420677 );
buf ( n420679 , n413104 );
buf ( n420680 , n62159 );
and ( n74074 , n420679 , n420680 );
nor ( n74075 , n74071 , n74074 );
buf ( n420683 , n74075 );
buf ( n420684 , n420683 );
buf ( n420685 , n409429 );
or ( n74079 , n420684 , n420685 );
buf ( n420687 , n419158 );
buf ( n420688 , n409170 );
or ( n74082 , n420687 , n420688 );
nand ( n74083 , n74079 , n74082 );
buf ( n420691 , n74083 );
buf ( n420692 , n420691 );
xor ( n74086 , n420675 , n420692 );
buf ( n420694 , n348158 );
not ( n74088 , n420694 );
buf ( n420696 , n420492 );
not ( n74090 , n420696 );
buf ( n420698 , n74090 );
buf ( n420699 , n420698 );
not ( n74093 , n420699 );
or ( n74094 , n74088 , n74093 );
buf ( n420702 , n62139 );
buf ( n420703 , n66411 );
and ( n74097 , n420702 , n420703 );
buf ( n420705 , n409140 );
buf ( n420706 , n62496 );
and ( n74100 , n420705 , n420706 );
nor ( n74101 , n74097 , n74100 );
buf ( n420709 , n74101 );
buf ( n420710 , n420709 );
buf ( n420711 , n410724 );
or ( n74105 , n420710 , n420711 );
nand ( n74106 , n74094 , n74105 );
buf ( n420714 , n74106 );
buf ( n420715 , n420714 );
and ( n74109 , n74086 , n420715 );
and ( n74110 , n420675 , n420692 );
or ( n74111 , n74109 , n74110 );
buf ( n420719 , n74111 );
xor ( n74113 , n419143 , n72516 );
xor ( n74114 , n74113 , n419169 );
and ( n74115 , n420719 , n74114 );
and ( n74116 , n420668 , n420719 );
or ( n74117 , n74064 , n74115 , n74116 );
buf ( n420725 , n74117 );
and ( n74119 , n73897 , n420725 );
and ( n74120 , n420454 , n420503 );
or ( n74121 , n74119 , n74120 );
buf ( n420729 , n74121 );
xor ( n74123 , n72469 , n419199 );
xor ( n74124 , n74123 , n419203 );
and ( n74125 , n420729 , n74124 );
xor ( n74126 , n420471 , n420475 );
xor ( n74127 , n74126 , n420498 );
buf ( n420735 , n74127 );
buf ( n420736 , n62467 );
buf ( n420737 , n63625 );
and ( n74131 , n420736 , n420737 );
buf ( n420739 , n409468 );
buf ( n420740 , n63629 );
and ( n74134 , n420739 , n420740 );
nor ( n74135 , n74131 , n74134 );
buf ( n420743 , n74135 );
buf ( n420744 , n420743 );
buf ( n420745 , n410635 );
or ( n74139 , n420744 , n420745 );
buf ( n420747 , n420462 );
buf ( n420748 , n409504 );
or ( n74142 , n420747 , n420748 );
nand ( n74143 , n74139 , n74142 );
buf ( n420751 , n74143 );
buf ( n420752 , n420751 );
buf ( n420753 , n66270 );
buf ( n420754 , n62177 );
and ( n74148 , n420753 , n420754 );
buf ( n420756 , n413098 );
buf ( n420757 , n62159 );
and ( n74151 , n420756 , n420757 );
nor ( n74152 , n74148 , n74151 );
buf ( n420760 , n74152 );
buf ( n420761 , n420760 );
buf ( n420762 , n409429 );
or ( n74156 , n420761 , n420762 );
buf ( n420764 , n420683 );
buf ( n420765 , n409170 );
or ( n74159 , n420764 , n420765 );
nand ( n74160 , n74156 , n74159 );
buf ( n420768 , n74160 );
buf ( n420769 , n420768 );
xor ( n74163 , n420538 , n420580 );
xor ( n74164 , n74163 , n420585 );
buf ( n420772 , n74164 );
buf ( n420773 , n420772 );
xor ( n74167 , n420769 , n420773 );
buf ( n420775 , n70210 );
buf ( n420776 , n405391 );
and ( n74170 , n420775 , n420776 );
buf ( n420778 , n416845 );
buf ( n420779 , n405388 );
and ( n74173 , n420778 , n420779 );
nor ( n74174 , n74170 , n74173 );
buf ( n420782 , n74174 );
buf ( n420783 , n420782 );
buf ( n420784 , n405407 );
or ( n420785 , n420783 , n420784 );
buf ( n420786 , n420633 );
buf ( n420787 , n405384 );
or ( n74181 , n420786 , n420787 );
nand ( n74182 , n420785 , n74181 );
buf ( n420790 , n74182 );
buf ( n420791 , n420790 );
buf ( n420792 , n403158 );
buf ( n420793 , n401689 );
buf ( n420794 , n72308 );
and ( n74188 , n420793 , n420794 );
buf ( n420796 , n401678 );
buf ( n420797 , n418942 );
and ( n74191 , n420796 , n420797 );
nor ( n74192 , n74188 , n74191 );
buf ( n420800 , n74192 );
buf ( n420801 , n420800 );
or ( n74195 , n420792 , n420801 );
buf ( n420803 , n420547 );
buf ( n420804 , n401660 );
or ( n74198 , n420803 , n420804 );
nand ( n74199 , n74195 , n74198 );
buf ( n420807 , n74199 );
buf ( n420808 , n420807 );
buf ( n420809 , n401619 );
buf ( n420810 , n420612 );
nor ( n74204 , n420809 , n420810 );
buf ( n420812 , n74204 );
buf ( n420813 , n420812 );
xor ( n74207 , n420808 , n420813 );
buf ( n420815 , n403120 );
buf ( n420816 , n55905 );
buf ( n420817 , n71664 );
and ( n74211 , n420816 , n420817 );
buf ( n420819 , n15290 );
buf ( n420820 , n418298 );
and ( n74214 , n420819 , n420820 );
nor ( n74215 , n74211 , n74214 );
buf ( n420823 , n74215 );
buf ( n420824 , n420823 );
or ( n74218 , n420815 , n420824 );
buf ( n420826 , n420563 );
buf ( n420827 , n403133 );
or ( n74221 , n420826 , n420827 );
nand ( n74222 , n74218 , n74221 );
buf ( n420830 , n74222 );
buf ( n420831 , n420830 );
and ( n74225 , n74207 , n420831 );
and ( n74226 , n420808 , n420813 );
or ( n74227 , n74225 , n74226 );
buf ( n420835 , n74227 );
buf ( n420836 , n420835 );
xor ( n74230 , n420791 , n420836 );
buf ( n420838 , n59471 );
not ( n74232 , n420838 );
buf ( n420840 , n420652 );
not ( n74234 , n420840 );
or ( n74235 , n74232 , n74234 );
buf ( n420843 , n68002 );
buf ( n420844 , n59628 );
and ( n74238 , n420843 , n420844 );
buf ( n420846 , n414729 );
buf ( n420847 , n58223 );
and ( n74241 , n420846 , n420847 );
nor ( n74242 , n74238 , n74241 );
buf ( n420850 , n74242 );
buf ( n420851 , n420850 );
buf ( n420852 , n59637 );
or ( n74246 , n420851 , n420852 );
nand ( n74247 , n74235 , n74246 );
buf ( n420855 , n74247 );
buf ( n420856 , n420855 );
and ( n74250 , n74230 , n420856 );
and ( n74251 , n420791 , n420836 );
or ( n74252 , n74250 , n74251 );
buf ( n420860 , n74252 );
buf ( n420861 , n420860 );
and ( n74255 , n74167 , n420861 );
and ( n74256 , n420769 , n420773 );
or ( n74257 , n74255 , n74256 );
buf ( n420865 , n74257 );
buf ( n420866 , n420865 );
xor ( n74260 , n420752 , n420866 );
xor ( n74261 , n420521 , n420590 );
xor ( n74262 , n74261 , n420664 );
buf ( n420870 , n74262 );
buf ( n420871 , n420870 );
and ( n74265 , n74260 , n420871 );
and ( n74266 , n420752 , n420866 );
or ( n74267 , n74265 , n74266 );
buf ( n420875 , n74267 );
xor ( n74269 , n420735 , n420875 );
xor ( n74270 , n419143 , n72516 );
xor ( n74271 , n74270 , n419169 );
xor ( n74272 , n420668 , n420719 );
xor ( n74273 , n74271 , n74272 );
and ( n74274 , n74269 , n74273 );
and ( n74275 , n420735 , n420875 );
or ( n74276 , n74274 , n74275 );
buf ( n420884 , n74276 );
xor ( n74278 , n419173 , n419190 );
xor ( n74279 , n74278 , n419195 );
buf ( n420887 , n74279 );
buf ( n420888 , n420887 );
xor ( n74282 , n420884 , n420888 );
xor ( n74283 , n420454 , n420503 );
xor ( n74284 , n74283 , n420725 );
buf ( n420892 , n74284 );
buf ( n420893 , n420892 );
and ( n74287 , n74282 , n420893 );
and ( n74288 , n420884 , n420888 );
or ( n74289 , n74287 , n74288 );
buf ( n420897 , n74289 );
xor ( n74291 , n72469 , n419199 );
xor ( n74292 , n74291 , n419203 );
and ( n74293 , n420897 , n74292 );
and ( n74294 , n420729 , n420897 );
or ( n74295 , n74125 , n74293 , n74294 );
buf ( n420903 , n74295 );
xor ( n74297 , n420450 , n420903 );
buf ( n420905 , n40591 );
buf ( n420906 , n372471 );
not ( n74300 , n420906 );
buf ( n420908 , n74300 );
buf ( n420909 , n420908 );
not ( n74303 , n420909 );
buf ( n420911 , n74303 );
buf ( n420912 , n420911 );
not ( n74306 , n420912 );
buf ( n420914 , n388080 );
not ( n74308 , n420914 );
or ( n74309 , n74306 , n74308 );
buf ( n420917 , n388080 );
not ( n74311 , n420917 );
buf ( n420919 , n74311 );
buf ( n420920 , n420919 );
buf ( n420921 , n418804 );
nand ( n74315 , n420920 , n420921 );
buf ( n420923 , n74315 );
buf ( n420924 , n420923 );
nand ( n74318 , n74309 , n420924 );
buf ( n420926 , n74318 );
buf ( n420927 , n420926 );
not ( n74321 , n420927 );
buf ( n420929 , n74321 );
buf ( n420930 , n420929 );
or ( n74324 , n420905 , n420930 );
buf ( n420932 , n73309 );
buf ( n420933 , n388071 );
or ( n74327 , n420932 , n420933 );
nand ( n74328 , n74324 , n74327 );
buf ( n420936 , n74328 );
buf ( n420937 , n420936 );
and ( n74331 , n74297 , n420937 );
and ( n74332 , n420450 , n420903 );
or ( n74333 , n74331 , n74332 );
buf ( n420941 , n74333 );
not ( n74335 , n420941 );
nand ( n74336 , n73838 , n74335 );
not ( n74337 , n74336 );
buf ( n420945 , n43515 );
not ( n74339 , n420945 );
buf ( n420947 , n419950 );
not ( n74341 , n420947 );
or ( n74342 , n74339 , n74341 );
buf ( n420950 , n388064 );
not ( n74344 , n420950 );
buf ( n420952 , n372527 );
not ( n74346 , n420952 );
buf ( n420954 , n74346 );
buf ( n420955 , n420954 );
not ( n74349 , n420955 );
or ( n74350 , n74344 , n74349 );
buf ( n420958 , n389338 );
buf ( n420959 , n371876 );
nand ( n74353 , n420958 , n420959 );
buf ( n420961 , n74353 );
buf ( n420962 , n420961 );
nand ( n74356 , n74350 , n420962 );
buf ( n420964 , n74356 );
buf ( n420965 , n420964 );
buf ( n420966 , n43536 );
nand ( n74360 , n420965 , n420966 );
buf ( n420968 , n74360 );
buf ( n420969 , n420968 );
nand ( n74363 , n74342 , n420969 );
buf ( n420971 , n74363 );
buf ( n420972 , n420971 );
not ( n74366 , n420972 );
buf ( n420974 , n43515 );
not ( n74368 , n420974 );
buf ( n420976 , n420964 );
not ( n74370 , n420976 );
or ( n74371 , n74368 , n74370 );
nand ( n420979 , n390997 , n23725 );
not ( n74373 , n420979 );
nor ( n74374 , n74373 , n43533 );
buf ( n74375 , n74374 );
buf ( n420983 , n74375 );
buf ( n420984 , n388064 );
not ( n74378 , n420984 );
buf ( n420986 , n74378 );
buf ( n420987 , n420986 );
not ( n74381 , n420987 );
buf ( n420989 , n24887 );
not ( n74383 , n420989 );
or ( n74384 , n74381 , n74383 );
buf ( n420992 , n24887 );
buf ( n74386 , n420992 );
buf ( n420994 , n74386 );
buf ( n420995 , n420994 );
not ( n74389 , n420995 );
buf ( n420997 , n74389 );
buf ( n420998 , n420997 );
buf ( n420999 , n371879 );
nand ( n74393 , n420998 , n420999 );
buf ( n421001 , n74393 );
buf ( n421002 , n421001 );
nand ( n74396 , n74384 , n421002 );
buf ( n421004 , n74396 );
buf ( n421005 , n421004 );
nand ( n74399 , n420983 , n421005 );
buf ( n421007 , n74399 );
buf ( n421008 , n421007 );
nand ( n74402 , n74371 , n421008 );
buf ( n421010 , n74402 );
not ( n74404 , n421010 );
not ( n74405 , n74404 );
xor ( n74406 , n72469 , n419199 );
xor ( n74407 , n74406 , n419203 );
xor ( n74408 , n420729 , n420897 );
xor ( n74409 , n74407 , n74408 );
not ( n74410 , n74409 );
not ( n74411 , n74410 );
or ( n74412 , n74405 , n74411 );
buf ( n421020 , n392884 );
not ( n74414 , n421020 );
buf ( n421022 , n24226 );
not ( n74416 , n421022 );
buf ( n421024 , n74416 );
buf ( n421025 , n421024 );
not ( n74419 , n421025 );
or ( n74420 , n74414 , n74419 );
buf ( n421028 , n420919 );
buf ( n421029 , n392881 );
nand ( n74423 , n421028 , n421029 );
buf ( n421031 , n74423 );
buf ( n421032 , n421031 );
nand ( n74426 , n74420 , n421032 );
buf ( n421034 , n74426 );
not ( n74428 , n421034 );
not ( n74429 , n67042 );
or ( n74430 , n74428 , n74429 );
buf ( n421038 , n420926 );
buf ( n421039 , n388068 );
nand ( n74433 , n421038 , n421039 );
buf ( n421041 , n74433 );
nand ( n74435 , n74430 , n421041 );
nand ( n74436 , n74412 , n74435 );
not ( n74437 , n74410 );
nand ( n74438 , n74437 , n421010 );
nand ( n74439 , n74436 , n74438 );
buf ( n421047 , n74439 );
not ( n74441 , n421047 );
or ( n74442 , n74366 , n74441 );
buf ( n421050 , n74439 );
buf ( n421051 , n420971 );
or ( n74445 , n421050 , n421051 );
xor ( n74446 , n420450 , n420903 );
xor ( n74447 , n74446 , n420937 );
buf ( n421055 , n74447 );
buf ( n421056 , n421055 );
nand ( n74450 , n74445 , n421056 );
buf ( n421058 , n74450 );
buf ( n421059 , n421058 );
nand ( n74453 , n74442 , n421059 );
buf ( n421061 , n74453 );
not ( n74455 , n421061 );
or ( n74456 , n74337 , n74455 );
nand ( n74457 , n73837 , n420941 );
nand ( n74458 , n74456 , n74457 );
buf ( n421066 , n74458 );
not ( n74460 , n413643 );
nand ( n74461 , n420125 , n73520 );
not ( n74462 , n74461 );
or ( n74463 , n74460 , n74462 );
buf ( n421071 , n73361 );
buf ( n421072 , n417542 );
nand ( n74466 , n421071 , n421072 );
buf ( n421074 , n74466 );
nand ( n74468 , n74463 , n421074 );
buf ( n421076 , n74468 );
xor ( n74470 , n421066 , n421076 );
buf ( n421078 , n49117 );
not ( n74472 , n421078 );
buf ( n421080 , n41341 );
not ( n74474 , n421080 );
or ( n74475 , n74472 , n74474 );
buf ( n421083 , n41365 );
buf ( n421084 , n67126 );
nand ( n74478 , n421083 , n421084 );
buf ( n421086 , n74478 );
buf ( n421087 , n421086 );
nand ( n74481 , n74475 , n421087 );
buf ( n421089 , n74481 );
buf ( n421090 , n421089 );
not ( n74484 , n421090 );
buf ( n421092 , n66128 );
not ( n74486 , n421092 );
or ( n74487 , n74484 , n74486 );
buf ( n421095 , n418783 );
buf ( n421096 , n412976 );
nand ( n74490 , n421095 , n421096 );
buf ( n421098 , n74490 );
buf ( n421099 , n421098 );
nand ( n74493 , n74487 , n421099 );
buf ( n421101 , n74493 );
buf ( n421102 , n421101 );
and ( n74496 , n74470 , n421102 );
and ( n74497 , n421066 , n421076 );
or ( n74498 , n74496 , n74497 );
buf ( n421106 , n74498 );
and ( n74500 , n73817 , n421106 );
and ( n74501 , n420414 , n73816 );
or ( n74502 , n74500 , n74501 );
buf ( n421110 , n74502 );
xor ( n74504 , n73802 , n421110 );
buf ( n421112 , n74504 );
buf ( n421113 , n421112 );
nand ( n74507 , n73791 , n421113 );
buf ( n421115 , n74507 );
buf ( n421116 , n421115 );
buf ( n421117 , n73763 );
not ( n74511 , n421117 );
buf ( n421119 , n420392 );
nand ( n74513 , n74511 , n421119 );
buf ( n421121 , n74513 );
buf ( n421122 , n421121 );
nand ( n74516 , n421116 , n421122 );
buf ( n421124 , n74516 );
buf ( n421125 , n421124 );
nand ( n74519 , n73761 , n421125 );
buf ( n421127 , n74519 );
buf ( n421128 , n421127 );
nand ( n74522 , n73758 , n421128 );
buf ( n421130 , n74522 );
buf ( n421131 , n421130 );
xor ( n74525 , n73199 , n421131 );
buf ( n421133 , n74525 );
buf ( n421134 , n421133 );
not ( n74528 , n421134 );
buf ( n421136 , n74528 );
buf ( n421137 , n421136 );
not ( n74531 , n421137 );
xor ( n74532 , n419518 , n419527 );
and ( n74533 , n74532 , n419547 );
and ( n74534 , n419518 , n419527 );
or ( n74535 , n74533 , n74534 );
buf ( n421143 , n74535 );
buf ( n421144 , n421143 );
buf ( n74538 , n41709 );
buf ( n421146 , n74538 );
buf ( n421147 , n420268 );
not ( n74541 , n421147 );
buf ( n421149 , n74541 );
buf ( n421150 , n421149 );
or ( n74544 , n421146 , n421150 );
buf ( n421152 , n41861 );
not ( n74546 , n421152 );
buf ( n421154 , n24117 );
not ( n74548 , n421154 );
or ( n74549 , n74546 , n74548 );
buf ( n421157 , n24116 );
buf ( n421158 , n389353 );
nand ( n74552 , n421157 , n421158 );
buf ( n421160 , n74552 );
buf ( n421161 , n421160 );
nand ( n74555 , n74549 , n421161 );
buf ( n421163 , n74555 );
buf ( n421164 , n421163 );
not ( n74558 , n421164 );
buf ( n421166 , n74558 );
buf ( n421167 , n421166 );
buf ( n74561 , n41663 );
buf ( n421169 , n74561 );
or ( n74563 , n421167 , n421169 );
nand ( n74564 , n74544 , n74563 );
buf ( n421172 , n74564 );
buf ( n421173 , n421172 );
xor ( n74567 , n70151 , n416911 );
xor ( n74568 , n74567 , n416915 );
xor ( n74569 , n417164 , n70593 );
xor ( n74570 , n74568 , n74569 );
buf ( n421178 , n74570 );
xor ( n74572 , n417215 , n417218 );
xor ( n74573 , n74572 , n417222 );
and ( n74574 , n73615 , n74573 );
xor ( n74575 , n417215 , n417218 );
xor ( n74576 , n74575 , n417222 );
and ( n74577 , n73619 , n74576 );
and ( n74578 , n73615 , n73619 );
or ( n74579 , n74574 , n74577 , n74578 );
buf ( n421187 , n74579 );
xor ( n74581 , n421178 , n421187 );
buf ( n421189 , n388803 );
not ( n74583 , n421189 );
buf ( n421191 , n371800 );
not ( n74585 , n421191 );
buf ( n421193 , n412892 );
not ( n74587 , n421193 );
or ( n74588 , n74585 , n74587 );
buf ( n421196 , n417617 );
not ( n74590 , n421196 );
buf ( n421198 , n27320 );
nand ( n74592 , n74590 , n421198 );
buf ( n421200 , n74592 );
buf ( n421201 , n421200 );
nand ( n74595 , n74588 , n421201 );
buf ( n421203 , n74595 );
buf ( n421204 , n421203 );
not ( n74598 , n421204 );
or ( n74599 , n74583 , n74598 );
buf ( n421207 , n388740 );
buf ( n421208 , n420242 );
nand ( n74602 , n421207 , n421208 );
buf ( n421210 , n74602 );
buf ( n421211 , n421210 );
nand ( n74605 , n74599 , n421211 );
buf ( n421213 , n74605 );
buf ( n421214 , n421213 );
xor ( n74608 , n74581 , n421214 );
buf ( n421216 , n74608 );
buf ( n421217 , n421216 );
xor ( n74611 , n421173 , n421217 );
buf ( n421219 , n419538 );
not ( n74613 , n421219 );
buf ( n421221 , n66128 );
not ( n74615 , n421221 );
or ( n74616 , n74613 , n74615 );
buf ( n421224 , n391446 );
not ( n74618 , n421224 );
buf ( n421226 , n66132 );
not ( n74620 , n421226 );
or ( n74621 , n74618 , n74620 );
buf ( n421229 , n416298 );
buf ( n421230 , n391443 );
nand ( n74624 , n421229 , n421230 );
buf ( n421232 , n74624 );
buf ( n421233 , n421232 );
nand ( n74627 , n74621 , n421233 );
buf ( n421235 , n74627 );
buf ( n421236 , n421235 );
buf ( n421237 , n412976 );
nand ( n74631 , n421236 , n421237 );
buf ( n421239 , n74631 );
buf ( n421240 , n421239 );
nand ( n74634 , n74616 , n421240 );
buf ( n421242 , n74634 );
buf ( n421243 , n421242 );
xor ( n74637 , n74611 , n421243 );
buf ( n421245 , n74637 );
buf ( n421246 , n421245 );
xor ( n74640 , n421144 , n421246 );
not ( n74641 , n420304 );
not ( n74642 , n43536 );
or ( n74643 , n74641 , n74642 );
buf ( n421251 , n411504 );
not ( n74645 , n421251 );
buf ( n421253 , n410400 );
not ( n74647 , n421253 );
or ( n74648 , n74645 , n74647 );
buf ( n421256 , n12471 );
buf ( n421257 , n391024 );
nand ( n74651 , n421256 , n421257 );
buf ( n421259 , n74651 );
buf ( n421260 , n421259 );
nand ( n74654 , n74648 , n421260 );
buf ( n421262 , n74654 );
buf ( n421263 , n421262 );
not ( n74657 , n421263 );
buf ( n421265 , n74657 );
or ( n74659 , n421265 , n43516 );
nand ( n74660 , n74643 , n74659 );
buf ( n421268 , n74660 );
xor ( n74662 , n74640 , n421268 );
buf ( n421270 , n74662 );
buf ( n421271 , n421270 );
xor ( n74665 , n419550 , n419587 );
and ( n74666 , n74665 , n419717 );
and ( n74667 , n419550 , n419587 );
or ( n74668 , n74666 , n74667 );
buf ( n421276 , n74668 );
buf ( n421277 , n421276 );
xor ( n74671 , n421271 , n421277 );
buf ( n421279 , n419579 );
not ( n74673 , n421279 );
buf ( n421281 , n52812 );
not ( n74675 , n421281 );
or ( n74676 , n74673 , n74675 );
buf ( n421284 , n394817 );
not ( n74678 , n421284 );
buf ( n421286 , n41555 );
not ( n74680 , n421286 );
or ( n74681 , n74678 , n74680 );
buf ( n421289 , n60880 );
buf ( n421290 , n394814 );
nand ( n74684 , n421289 , n421290 );
buf ( n421292 , n74684 );
buf ( n421293 , n421292 );
nand ( n74687 , n74681 , n421293 );
buf ( n421295 , n74687 );
buf ( n421296 , n421295 );
buf ( n421297 , n42924 );
nand ( n74691 , n421296 , n421297 );
buf ( n421299 , n74691 );
buf ( n421300 , n421299 );
nand ( n74694 , n74676 , n421300 );
buf ( n421302 , n74694 );
buf ( n421303 , n421302 );
not ( n74697 , n421303 );
buf ( n421305 , n74697 );
xor ( n74699 , n420279 , n420289 );
and ( n74700 , n74699 , n420315 );
and ( n74701 , n420279 , n420289 );
or ( n74702 , n74700 , n74701 );
buf ( n421310 , n74702 );
xor ( n74704 , n421305 , n421310 );
buf ( n421312 , n417601 );
not ( n74706 , n421312 );
buf ( n421314 , n409082 );
not ( n74708 , n421314 );
or ( n74709 , n74706 , n74708 );
buf ( n421317 , n392884 );
not ( n74711 , n421317 );
buf ( n421319 , n409092 );
not ( n74713 , n421319 );
or ( n74714 , n74711 , n74713 );
buf ( n421322 , n407928 );
buf ( n421323 , n392887 );
nand ( n74717 , n421322 , n421323 );
buf ( n421325 , n74717 );
buf ( n421326 , n421325 );
nand ( n74720 , n74714 , n421326 );
buf ( n421328 , n74720 );
buf ( n421329 , n421328 );
buf ( n421330 , n409076 );
nand ( n74724 , n421329 , n421330 );
buf ( n421332 , n74724 );
buf ( n421333 , n421332 );
nand ( n74727 , n74709 , n421333 );
buf ( n421335 , n74727 );
not ( n74729 , n72867 );
not ( n74730 , n40592 );
or ( n74731 , n74729 , n74730 );
buf ( n421339 , n12480 );
buf ( n421340 , n40601 );
xnor ( n74734 , n421339 , n421340 );
buf ( n421342 , n74734 );
or ( n74736 , n421342 , n388071 );
nand ( n74737 , n74731 , n74736 );
buf ( n421345 , n74737 );
not ( n74739 , n421345 );
xor ( n74740 , n420229 , n420250 );
and ( n74741 , n74740 , n420276 );
and ( n421349 , n420229 , n420250 );
or ( n74743 , n74741 , n421349 );
buf ( n421351 , n74743 );
buf ( n421352 , n421351 );
not ( n74746 , n421352 );
buf ( n421354 , n74746 );
buf ( n421355 , n421354 );
not ( n74749 , n421355 );
and ( n74750 , n74739 , n74749 );
buf ( n421358 , n74737 );
buf ( n421359 , n421354 );
and ( n74753 , n421358 , n421359 );
nor ( n74754 , n74750 , n74753 );
buf ( n421362 , n74754 );
xor ( n74756 , n421335 , n421362 );
xor ( n74757 , n74704 , n74756 );
buf ( n421365 , n74757 );
xor ( n74759 , n74671 , n421365 );
buf ( n421367 , n74759 );
xor ( n74761 , n420212 , n420338 );
and ( n74762 , n74761 , n420360 );
and ( n74763 , n420212 , n420338 );
or ( n74764 , n74762 , n74763 );
buf ( n421372 , n74764 );
xor ( n74766 , n421367 , n421372 );
buf ( n421374 , n74766 );
xor ( n74768 , n420318 , n420323 );
and ( n74769 , n74768 , n420335 );
and ( n74770 , n420318 , n420323 );
or ( n74771 , n74769 , n74770 );
buf ( n421379 , n74771 );
buf ( n421380 , n395362 );
not ( n74774 , n421380 );
buf ( n421382 , n47863 );
not ( n74776 , n421382 );
buf ( n421384 , n41194 );
not ( n74778 , n421384 );
or ( n74779 , n74776 , n74778 );
buf ( n421387 , n28250 );
buf ( n421388 , n419385 );
nand ( n74782 , n421387 , n421388 );
buf ( n421390 , n74782 );
buf ( n421391 , n421390 );
nand ( n74785 , n74779 , n421391 );
buf ( n421393 , n74785 );
buf ( n421394 , n421393 );
not ( n74788 , n421394 );
or ( n74789 , n74774 , n74788 );
buf ( n421397 , n419391 );
buf ( n421398 , n395349 );
nand ( n74792 , n421397 , n421398 );
buf ( n421400 , n74792 );
buf ( n421401 , n421400 );
nand ( n74795 , n74789 , n421401 );
buf ( n421403 , n74795 );
buf ( n421404 , n421403 );
not ( n74798 , n421404 );
buf ( n421406 , n74798 );
and ( n74800 , n421379 , n421406 );
not ( n74801 , n421379 );
and ( n74802 , n74801 , n421403 );
or ( n74803 , n74800 , n74802 );
buf ( n421411 , n74803 );
buf ( n421412 , n358975 );
buf ( n421413 , n388962 );
and ( n74807 , n421412 , n421413 );
not ( n74808 , n421412 );
buf ( n421416 , n385488 );
and ( n74810 , n74808 , n421416 );
nor ( n74811 , n74807 , n74810 );
buf ( n421419 , n74811 );
buf ( n421420 , n421419 );
not ( n74814 , n421420 );
buf ( n421422 , n391553 );
not ( n74816 , n421422 );
or ( n74817 , n74814 , n74816 );
buf ( n421425 , n55055 );
not ( n74819 , n421425 );
buf ( n421427 , n388965 );
not ( n74821 , n421427 );
or ( n74822 , n74819 , n74821 );
buf ( n421430 , n385473 );
buf ( n421431 , n55054 );
nand ( n74825 , n421430 , n421431 );
buf ( n421433 , n74825 );
buf ( n421434 , n421433 );
nand ( n74828 , n74822 , n421434 );
buf ( n421436 , n74828 );
buf ( n421437 , n421436 );
buf ( n421438 , n49166 );
nand ( n74832 , n421437 , n421438 );
buf ( n421440 , n74832 );
buf ( n421441 , n421440 );
nand ( n74835 , n74817 , n421441 );
buf ( n421443 , n74835 );
buf ( n421444 , n421443 );
not ( n74838 , n421444 );
buf ( n421446 , n74838 );
buf ( n421447 , n421446 );
and ( n74841 , n421411 , n421447 );
not ( n74842 , n421411 );
buf ( n421450 , n421443 );
and ( n74844 , n74842 , n421450 );
nor ( n74845 , n74841 , n74844 );
buf ( n421453 , n74845 );
buf ( n421454 , n421453 );
not ( n74848 , n421454 );
buf ( n421456 , n74848 );
buf ( n421457 , n421456 );
and ( n74851 , n421374 , n421457 );
not ( n74852 , n421374 );
buf ( n421460 , n421453 );
and ( n74854 , n74852 , n421460 );
nor ( n74855 , n74851 , n74854 );
buf ( n421463 , n74855 );
buf ( n421464 , n421463 );
not ( n74858 , n421464 );
buf ( n421466 , n74858 );
buf ( n421467 , n421466 );
not ( n74861 , n421467 );
buf ( n421469 , n38630 );
not ( n74869 , n421469 );
buf ( n421471 , n74869 );
xor ( n74886 , n420404 , n420408 );
and ( n74887 , n74886 , n421110 );
and ( n74888 , n420404 , n420408 );
or ( n74889 , n74887 , n74888 );
buf ( n421476 , n74889 );
buf ( n421477 , n421476 );
buf ( n421478 , n389122 );
not ( n74893 , n421478 );
buf ( n421480 , n74893 );
buf ( n421481 , n421480 );
buf ( n421482 , n400042 );
buf ( n421483 , n24049 );
and ( n74898 , n421482 , n421483 );
not ( n74899 , n421482 );
buf ( n421486 , n45391 );
and ( n74901 , n74899 , n421486 );
nor ( n74902 , n74898 , n74901 );
buf ( n421489 , n74902 );
buf ( n421490 , n421489 );
or ( n74905 , n421481 , n421490 );
buf ( n421492 , n419345 );
buf ( n421493 , n41562 );
or ( n74908 , n421492 , n421493 );
nand ( n74909 , n74905 , n74908 );
buf ( n421496 , n74909 );
buf ( n421497 , n421496 );
buf ( n421498 , n45102 );
buf ( n421499 , n358975 );
or ( n74914 , n421498 , n421499 );
buf ( n421501 , n22982 );
buf ( n421502 , n402819 );
or ( n74917 , n421501 , n421502 );
nand ( n421504 , n74914 , n74917 );
buf ( n421505 , n421504 );
buf ( n421506 , n421505 );
not ( n74921 , n421506 );
buf ( n421508 , n38961 );
not ( n74923 , n421508 );
or ( n74924 , n74921 , n74923 );
buf ( n421511 , n419470 );
buf ( n421512 , n393127 );
nand ( n74927 , n421511 , n421512 );
buf ( n421514 , n74927 );
buf ( n421515 , n421514 );
nand ( n74930 , n74924 , n421515 );
buf ( n421517 , n74930 );
buf ( n421518 , n421517 );
xor ( n74933 , n421497 , n421518 );
buf ( n421520 , n419406 );
not ( n74935 , n421520 );
buf ( n421522 , n74935 );
buf ( n421523 , n421522 );
buf ( n421524 , n395365 );
or ( n74939 , n421523 , n421524 );
buf ( n421526 , n420072 );
buf ( n421527 , n395346 );
nand ( n74942 , n421526 , n421527 );
buf ( n421529 , n74942 );
buf ( n421530 , n421529 );
nand ( n74945 , n74939 , n421530 );
buf ( n421532 , n74945 );
buf ( n421533 , n421532 );
and ( n74948 , n74933 , n421533 );
and ( n74949 , n421497 , n421518 );
or ( n74950 , n74948 , n74949 );
buf ( n421537 , n74950 );
buf ( n421538 , n421537 );
not ( n74955 , n42825 );
buf ( n421540 , C0 );
buf ( n421541 , n421540 );
and ( n74973 , n421477 , n421538 );
or ( n74974 , C0 , n74973 );
buf ( n421544 , n74974 );
buf ( n421545 , n421544 );
buf ( n421546 , C1 );
buf ( n421547 , n421546 );
nand ( n74987 , n421545 , n421547 );
buf ( n421549 , n74987 );
buf ( n421550 , n421549 );
nand ( n74990 , C1 , n421550 );
buf ( n421552 , n74990 );
buf ( n421553 , n421552 );
buf ( n421554 , C0 );
buf ( n421555 , n421554 );
xor ( n75013 , n419337 , n419373 );
xor ( n75014 , n75013 , n419414 );
buf ( n421558 , n75014 );
buf ( n421559 , n421558 );
or ( n75017 , n421555 , n421559 );
xor ( n75018 , n419458 , n419491 );
xor ( n75019 , n75018 , n419720 );
buf ( n421563 , n75019 );
buf ( n421564 , n421563 );
nand ( n75022 , n75017 , n421564 );
buf ( n421566 , n75022 );
buf ( n421567 , n421566 );
buf ( n421568 , C1 );
buf ( n421569 , n421568 );
and ( n75030 , n421567 , n421569 );
buf ( n421571 , n75030 );
buf ( n421572 , n421571 );
and ( n75033 , n421553 , n421572 );
not ( n75034 , n421553 );
buf ( n421575 , n421571 );
not ( n75036 , n421575 );
buf ( n421577 , n75036 );
buf ( n421578 , n421577 );
and ( n75039 , n75034 , n421578 );
nor ( n75040 , n75033 , n75039 );
buf ( n421581 , n75040 );
buf ( n421582 , n421581 );
not ( n75043 , n421582 );
buf ( n421584 , n75043 );
buf ( n421585 , n421584 );
not ( n75046 , n421585 );
or ( n75047 , n74861 , n75046 );
buf ( n421588 , n421581 );
buf ( n421589 , n421463 );
nand ( n75050 , n421588 , n421589 );
buf ( n421591 , n75050 );
buf ( n421592 , n421591 );
nand ( n75053 , n75047 , n421592 );
buf ( n421594 , n75053 );
buf ( n421595 , n421594 );
xor ( n75056 , n421477 , n421538 );
xor ( n75057 , n75056 , n421541 );
buf ( n421598 , n75057 );
buf ( n421599 , n421598 );
xor ( n75060 , n421497 , n421518 );
xor ( n75061 , n75060 , n421533 );
buf ( n421602 , n75061 );
buf ( n421603 , n421602 );
buf ( n421604 , C0 );
buf ( n421605 , n421604 );
xor ( n75084 , n421603 , n421605 );
xor ( n75085 , n419871 , n419877 );
xor ( n75086 , n75085 , n420142 );
buf ( n421609 , n75086 );
buf ( n421610 , n421609 );
and ( n75089 , n75084 , n421610 );
or ( n75091 , n75089 , C0 );
buf ( n421613 , n75091 );
buf ( n421614 , n421613 );
xor ( n75094 , n421599 , n421614 );
xor ( n75095 , n420414 , n73816 );
xor ( n75096 , n75095 , n421106 );
buf ( n421618 , n75096 );
not ( n75098 , n45954 );
not ( n75099 , n73217 );
or ( n75100 , n75098 , n75099 );
buf ( n421622 , n393369 );
not ( n75102 , n421622 );
buf ( n421624 , n388227 );
not ( n75104 , n421624 );
or ( n75105 , n75102 , n75104 );
buf ( n421627 , n406821 );
buf ( n421628 , n393381 );
nand ( n75108 , n421627 , n421628 );
buf ( n421630 , n75108 );
buf ( n421631 , n421630 );
nand ( n75111 , n75105 , n421631 );
buf ( n421633 , n75111 );
buf ( n421634 , n421633 );
buf ( n421635 , n45949 );
nand ( n75115 , n421634 , n421635 );
buf ( n421637 , n75115 );
nand ( n75117 , n75100 , n421637 );
buf ( n421639 , n394219 );
not ( n75119 , n421639 );
buf ( n421641 , n371784 );
not ( n75121 , n421641 );
or ( n75122 , n75119 , n75121 );
buf ( n421644 , n388751 );
not ( n75124 , n421644 );
buf ( n421646 , n75124 );
buf ( n421647 , n421646 );
not ( n75127 , n421647 );
buf ( n421649 , n394210 );
nand ( n75129 , n75127 , n421649 );
buf ( n421651 , n75129 );
buf ( n421652 , n421651 );
nand ( n75132 , n75122 , n421652 );
buf ( n421654 , n75132 );
buf ( n421655 , n421654 );
not ( n75135 , n421655 );
buf ( n421657 , n388740 );
not ( n75137 , n421657 );
or ( n75138 , n75135 , n75137 );
buf ( n421660 , n420436 );
buf ( n421661 , n388803 );
nand ( n75141 , n421660 , n421661 );
buf ( n421663 , n75141 );
buf ( n421664 , n421663 );
nand ( n75144 , n75138 , n421664 );
buf ( n421666 , n75144 );
buf ( n421667 , n421666 );
buf ( n421668 , n413643 );
not ( n75148 , n421668 );
buf ( n421670 , n73368 );
not ( n75150 , n421670 );
or ( n75151 , n75148 , n75150 );
buf ( n421673 , n44775 );
buf ( n421674 , n42066 );
and ( n75154 , n421673 , n421674 );
not ( n75155 , n421673 );
buf ( n421677 , n42065 );
and ( n75157 , n75155 , n421677 );
or ( n75158 , n75154 , n75157 );
buf ( n421680 , n75158 );
buf ( n421681 , n421680 );
not ( n75161 , n421681 );
buf ( n421683 , n417542 );
nand ( n75163 , n75161 , n421683 );
buf ( n421685 , n75163 );
buf ( n421686 , n421685 );
nand ( n75166 , n75151 , n421686 );
buf ( n421688 , n75166 );
buf ( n421689 , n421688 );
xor ( n75169 , n421667 , n421689 );
buf ( n421691 , n49117 );
not ( n75171 , n421691 );
buf ( n421693 , n41323 );
not ( n75173 , n421693 );
or ( n75174 , n75171 , n75173 );
buf ( n421696 , n24116 );
buf ( n421697 , n67126 );
nand ( n75177 , n421696 , n421697 );
buf ( n421699 , n75177 );
buf ( n421700 , n421699 );
nand ( n75180 , n75174 , n421700 );
buf ( n421702 , n75180 );
buf ( n421703 , n421702 );
not ( n75183 , n421703 );
buf ( n421705 , n73026 );
not ( n75185 , n421705 );
or ( n75186 , n75183 , n75185 );
buf ( n421708 , n73275 );
buf ( n421709 , n41664 );
nand ( n75189 , n421708 , n421709 );
buf ( n421711 , n75189 );
buf ( n421712 , n421711 );
nand ( n75192 , n75186 , n421712 );
buf ( n421714 , n75192 );
buf ( n421715 , n421714 );
and ( n75195 , n75169 , n421715 );
and ( n75196 , n421667 , n421689 );
or ( n75197 , n75195 , n75196 );
buf ( n421719 , n75197 );
not ( n75199 , n421719 );
and ( n75200 , n73838 , n74335 );
not ( n75201 , n73838 );
and ( n75202 , n75201 , n420941 );
nor ( n75203 , n75200 , n75202 );
xor ( n75204 , n421061 , n75203 );
not ( n75205 , n75204 );
or ( n75206 , n75199 , n75205 );
or ( n75207 , n421719 , n75204 );
buf ( n421729 , n397489 );
not ( n75209 , n421729 );
buf ( n421731 , n416292 );
not ( n75211 , n421731 );
or ( n75212 , n75209 , n75211 );
buf ( n421734 , n67832 );
buf ( n421735 , n397492 );
nand ( n75215 , n421734 , n421735 );
buf ( n421737 , n75215 );
buf ( n421738 , n421737 );
nand ( n75218 , n75212 , n421738 );
buf ( n421740 , n75218 );
buf ( n421741 , n421740 );
not ( n75221 , n421741 );
buf ( n421743 , n66128 );
not ( n75223 , n421743 );
or ( n75224 , n75221 , n75223 );
buf ( n421746 , n421089 );
buf ( n421747 , n412976 );
nand ( n75227 , n421746 , n421747 );
buf ( n421749 , n75227 );
buf ( n421750 , n421749 );
nand ( n75230 , n75224 , n421750 );
buf ( n421752 , n75230 );
nand ( n75232 , n75207 , n421752 );
nand ( n75233 , n75206 , n75232 );
xor ( n75234 , n75117 , n75233 );
buf ( n75235 , n53252 );
buf ( n421757 , n75235 );
buf ( n421758 , n389107 );
not ( n75238 , n421758 );
buf ( n421760 , n75238 );
buf ( n421761 , n421760 );
nand ( n75241 , n421757 , n421761 );
buf ( n421763 , n75241 );
buf ( n421764 , n421760 );
buf ( n421765 , n51821 );
or ( n75245 , n421764 , n421765 );
buf ( n421767 , n358975 );
nand ( n75247 , n75245 , n421767 );
buf ( n421769 , n75247 );
and ( n75249 , n421763 , n421769 , n24049 );
and ( n75250 , n75234 , n75249 );
and ( n75251 , n75117 , n75233 );
or ( n421773 , n75250 , n75251 );
buf ( n421774 , n421773 );
xor ( n75254 , n421618 , n421774 );
buf ( n421776 , n50579 );
not ( n75256 , n421776 );
buf ( n421778 , n47891 );
not ( n75258 , n421778 );
buf ( n421780 , n396585 );
not ( n75260 , n421780 );
or ( n75261 , n75258 , n75260 );
buf ( n421783 , n388643 );
buf ( n421784 , n72794 );
nand ( n75264 , n421783 , n421784 );
buf ( n421786 , n75264 );
buf ( n421787 , n421786 );
nand ( n75267 , n75261 , n421787 );
buf ( n421789 , n75267 );
buf ( n421790 , n421789 );
not ( n75270 , n421790 );
or ( n75271 , n75256 , n75270 );
buf ( n421793 , n420385 );
buf ( n421794 , n61577 );
nand ( n75274 , n421793 , n421794 );
buf ( n421796 , n75274 );
buf ( n421797 , n421796 );
nand ( n75277 , n75271 , n421797 );
buf ( n421799 , n75277 );
buf ( n421800 , n421799 );
and ( n75280 , n75254 , n421800 );
and ( n75281 , n421618 , n421774 );
or ( n75282 , n75280 , n75281 );
buf ( n421804 , n75282 );
buf ( n421805 , n421804 );
buf ( n421806 , n55055 );
buf ( n421807 , n41577 );
and ( n75287 , n421806 , n421807 );
not ( n75288 , n421806 );
buf ( n421810 , n45391 );
and ( n75290 , n75288 , n421810 );
nor ( n75291 , n75287 , n75290 );
buf ( n421813 , n75291 );
buf ( n421814 , n421813 );
not ( n75294 , n421814 );
buf ( n421816 , n396622 );
not ( n75296 , n421816 );
or ( n75297 , n75294 , n75296 );
buf ( n421819 , n421489 );
not ( n75299 , n421819 );
buf ( n421821 , n41565 );
nand ( n75301 , n75299 , n421821 );
buf ( n421823 , n75301 );
buf ( n421824 , n421823 );
nand ( n75304 , n75297 , n421824 );
buf ( n421826 , n75304 );
buf ( n421827 , n421826 );
buf ( n421828 , n400033 );
not ( n75308 , n421828 );
buf ( n421830 , n24071 );
not ( n75310 , n421830 );
or ( n75311 , n75308 , n75310 );
buf ( n421833 , n53252 );
buf ( n421834 , n400042 );
nand ( n75314 , n421833 , n421834 );
buf ( n421836 , n75314 );
buf ( n421837 , n421836 );
nand ( n75317 , n75311 , n421837 );
buf ( n421839 , n75317 );
buf ( n421840 , n421839 );
not ( n75320 , n421840 );
buf ( n421842 , n390432 );
not ( n75322 , n421842 );
or ( n75323 , n75320 , n75322 );
buf ( n421845 , n73232 );
buf ( n421846 , n42924 );
nand ( n75326 , n421845 , n421846 );
buf ( n421848 , n75326 );
buf ( n421849 , n421848 );
nand ( n75329 , n75323 , n421849 );
buf ( n421851 , n75329 );
buf ( n421852 , n421851 );
xor ( n75332 , n421066 , n421076 );
xor ( n75333 , n75332 , n421102 );
buf ( n421855 , n75333 );
buf ( n421856 , n421855 );
xor ( n75336 , n421852 , n421856 );
buf ( n421858 , n395362 );
not ( n75338 , n421858 );
buf ( n421860 , n420088 );
not ( n75340 , n421860 );
or ( n75341 , n75338 , n75340 );
buf ( n421863 , n47863 );
not ( n75343 , n421863 );
buf ( n421865 , n403039 );
not ( n75345 , n421865 );
or ( n75346 , n75343 , n75345 );
buf ( n421868 , n28644 );
buf ( n421869 , n47863 );
not ( n75349 , n421869 );
buf ( n421871 , n75349 );
buf ( n421872 , n421871 );
nand ( n75352 , n421868 , n421872 );
buf ( n421874 , n75352 );
buf ( n421875 , n421874 );
nand ( n75355 , n75346 , n421875 );
buf ( n421877 , n75355 );
buf ( n421878 , n421877 );
buf ( n421879 , n395346 );
nand ( n75359 , n421878 , n421879 );
buf ( n421881 , n75359 );
buf ( n421882 , n421881 );
nand ( n75362 , n75341 , n421882 );
buf ( n421884 , n75362 );
buf ( n421885 , n421884 );
and ( n75365 , n75336 , n421885 );
and ( n75366 , n421852 , n421856 );
or ( n75367 , n75365 , n75366 );
buf ( n421889 , n75367 );
buf ( n421890 , n421889 );
xor ( n75370 , n421827 , n421890 );
buf ( n421892 , n73219 );
not ( n75372 , n421892 );
buf ( n421894 , n419855 );
not ( n75374 , n421894 );
or ( n75375 , n75372 , n75374 );
buf ( n421897 , n419855 );
buf ( n421898 , n73219 );
or ( n75378 , n421897 , n421898 );
nand ( n75379 , n75375 , n75378 );
buf ( n421901 , n75379 );
buf ( n421902 , n421901 );
buf ( n421903 , n419864 );
and ( n75383 , n421902 , n421903 );
not ( n75384 , n421902 );
buf ( n421906 , n419832 );
and ( n75386 , n75384 , n421906 );
nor ( n75387 , n75383 , n75386 );
buf ( n421909 , n75387 );
buf ( n421910 , n421909 );
and ( n75390 , n75370 , n421910 );
and ( n75391 , n421827 , n421890 );
or ( n75392 , n75390 , n75391 );
buf ( n421914 , n75392 );
buf ( n421915 , n421914 );
buf ( n421916 , C0 );
buf ( n421917 , n421916 );
and ( n75417 , n421805 , n421915 );
or ( n75418 , C0 , n75417 );
buf ( n421920 , n75418 );
buf ( n421921 , n421920 );
and ( n75421 , n75094 , n421921 );
and ( n75422 , n421599 , n421614 );
or ( n75423 , n75421 , n75422 );
buf ( n421925 , n75423 );
buf ( n421926 , n421925 );
not ( n75426 , n421926 );
buf ( n421928 , n75426 );
buf ( n421929 , n421928 );
and ( n75429 , n421595 , n421929 );
not ( n75430 , n421595 );
buf ( n421932 , n421925 );
and ( n75432 , n75430 , n421932 );
nor ( n75433 , n75429 , n75432 );
buf ( n421935 , n75433 );
buf ( n421936 , n421935 );
not ( n75436 , n421936 );
or ( n75437 , n74531 , n75436 );
xor ( n75438 , n421563 , n421554 );
xnor ( n75439 , n75438 , n421558 );
buf ( n421941 , n75439 );
not ( n75441 , n421941 );
buf ( n421943 , n420146 );
buf ( n421944 , n421124 );
xor ( n75444 , n421943 , n421944 );
buf ( n421946 , n420362 );
xnor ( n75446 , n75444 , n421946 );
buf ( n421948 , n75446 );
buf ( n421949 , n421948 );
not ( n75449 , n421949 );
or ( n75450 , n75441 , n75449 );
buf ( n421952 , n45954 );
not ( n75452 , n421952 );
buf ( n421954 , n421633 );
not ( n75454 , n421954 );
or ( n75455 , n75452 , n75454 );
buf ( n421957 , n393369 );
not ( n75457 , n421957 );
buf ( n421959 , n412920 );
not ( n75459 , n421959 );
or ( n75460 , n75457 , n75459 );
buf ( n421962 , n12480 );
buf ( n421963 , n393381 );
nand ( n75463 , n421962 , n421963 );
buf ( n421965 , n75463 );
buf ( n421966 , n421965 );
nand ( n75466 , n75460 , n421966 );
buf ( n421968 , n75466 );
buf ( n421969 , n421968 );
buf ( n421970 , n45949 );
nand ( n75470 , n421969 , n421970 );
buf ( n421972 , n75470 );
buf ( n421973 , n421972 );
nand ( n75473 , n75455 , n421973 );
buf ( n421975 , n75473 );
buf ( n421976 , n421975 );
not ( n75476 , n421976 );
buf ( n421978 , n399274 );
buf ( n421979 , n40653 );
and ( n75479 , n421978 , n421979 );
not ( n75480 , n421978 );
buf ( n421982 , n407936 );
and ( n75482 , n75480 , n421982 );
nor ( n75483 , n75479 , n75482 );
buf ( n421985 , n75483 );
buf ( n421986 , n421985 );
not ( n75486 , n421986 );
buf ( n421988 , n75486 );
buf ( n421989 , n421988 );
not ( n75489 , n421989 );
buf ( n421991 , n60872 );
not ( n75491 , n421991 );
or ( n75492 , n75489 , n75491 );
buf ( n421994 , n420000 );
buf ( n421995 , n409076 );
nand ( n75495 , n421994 , n421995 );
buf ( n421997 , n75495 );
buf ( n421998 , n421997 );
nand ( n75498 , n75492 , n421998 );
buf ( n422000 , n75498 );
buf ( n422001 , n422000 );
not ( n75501 , n422001 );
or ( n75502 , n75476 , n75501 );
buf ( n422004 , n422000 );
buf ( n422005 , n421975 );
or ( n75505 , n422004 , n422005 );
xor ( n75506 , n419907 , n419961 );
xor ( n75507 , n75506 , n419983 );
buf ( n422009 , n75507 );
buf ( n422010 , n422009 );
nand ( n75510 , n75505 , n422010 );
buf ( n422012 , n75510 );
buf ( n422013 , n422012 );
nand ( n75513 , n75502 , n422013 );
buf ( n422015 , n75513 );
buf ( n422016 , n422015 );
xor ( n75516 , n419988 , n420025 );
xor ( n75517 , n75516 , n420053 );
buf ( n422019 , n75517 );
buf ( n422020 , n422019 );
xor ( n75520 , n422016 , n422020 );
buf ( n422022 , n55543 );
not ( n75522 , n422022 );
buf ( n422024 , n66132 );
not ( n75524 , n422024 );
or ( n75525 , n75522 , n75524 );
buf ( n422027 , n41365 );
buf ( n422028 , n51185 );
nand ( n75528 , n422027 , n422028 );
buf ( n422030 , n75528 );
buf ( n422031 , n422030 );
nand ( n75531 , n75525 , n422031 );
buf ( n422033 , n75531 );
buf ( n422034 , n422033 );
not ( n75534 , n422034 );
buf ( n422036 , n66128 );
not ( n75536 , n422036 );
or ( n75537 , n75534 , n75536 );
buf ( n422039 , n421740 );
buf ( n422040 , n412976 );
nand ( n75540 , n422039 , n422040 );
buf ( n422042 , n75540 );
buf ( n422043 , n422042 );
nand ( n75543 , n75537 , n422043 );
buf ( n422045 , n75543 );
buf ( n422046 , n422045 );
buf ( n422047 , n45954 );
not ( n75547 , n422047 );
buf ( n422049 , n421968 );
not ( n75549 , n422049 );
or ( n75550 , n75547 , n75549 );
buf ( n422052 , n393369 );
not ( n75552 , n422052 );
buf ( n422054 , n412964 );
not ( n75554 , n422054 );
or ( n75555 , n75552 , n75554 );
buf ( n422057 , n28353 );
buf ( n422058 , n393381 );
nand ( n75558 , n422057 , n422058 );
buf ( n422060 , n75558 );
buf ( n422061 , n422060 );
nand ( n75561 , n75555 , n422061 );
buf ( n422063 , n75561 );
buf ( n422064 , n422063 );
buf ( n422065 , n45949 );
nand ( n75565 , n422064 , n422065 );
buf ( n422067 , n75565 );
buf ( n422068 , n422067 );
nand ( n75568 , n75550 , n422068 );
buf ( n422070 , n75568 );
buf ( n422071 , n422070 );
xor ( n75571 , n422046 , n422071 );
xor ( n75572 , n421667 , n421689 );
xor ( n75573 , n75572 , n421715 );
buf ( n422075 , n75573 );
buf ( n422076 , n422075 );
and ( n75576 , n75571 , n422076 );
and ( n75577 , n422046 , n422071 );
or ( n75578 , n75576 , n75577 );
buf ( n422080 , n75578 );
buf ( n422081 , n422080 );
not ( n75581 , n422081 );
buf ( n422083 , n75581 );
not ( n75583 , n422083 );
buf ( n422085 , n395359 );
not ( n75585 , n422085 );
buf ( n422087 , n421877 );
not ( n75587 , n422087 );
or ( n75588 , n75585 , n75587 );
buf ( n422090 , n47863 );
not ( n75590 , n422090 );
buf ( n422092 , n410400 );
not ( n75592 , n422092 );
or ( n75593 , n75590 , n75592 );
buf ( n422095 , n12471 );
buf ( n422096 , n421871 );
nand ( n75596 , n422095 , n422096 );
buf ( n422098 , n75596 );
buf ( n422099 , n422098 );
nand ( n75599 , n75593 , n422099 );
buf ( n422101 , n75599 );
buf ( n422102 , n422101 );
buf ( n422103 , n395346 );
nand ( n75603 , n422102 , n422103 );
buf ( n422105 , n75603 );
buf ( n422106 , n422105 );
nand ( n75606 , n75588 , n422106 );
buf ( n422108 , n75606 );
nor ( n75608 , n75583 , n422108 );
buf ( n422110 , n394814 );
not ( n75610 , n422110 );
buf ( n422112 , n417617 );
not ( n75612 , n422112 );
or ( n75613 , n75610 , n75612 );
buf ( n422115 , n371784 );
not ( n75615 , n422115 );
buf ( n422117 , n417572 );
nand ( n75617 , n75615 , n422117 );
buf ( n422119 , n75617 );
buf ( n422120 , n422119 );
nand ( n75620 , n75613 , n422120 );
buf ( n422122 , n75620 );
buf ( n422123 , n422122 );
not ( n75623 , n422123 );
buf ( n422125 , n388740 );
not ( n75625 , n422125 );
or ( n75626 , n75623 , n75625 );
buf ( n422128 , n421654 );
buf ( n422129 , n388803 );
nand ( n75629 , n422128 , n422129 );
buf ( n422131 , n75629 );
buf ( n422132 , n422131 );
nand ( n75632 , n75626 , n422132 );
buf ( n422134 , n75632 );
buf ( n422135 , n422134 );
not ( n75635 , n422135 );
buf ( n422137 , n75635 );
buf ( n422138 , n422137 );
not ( n75638 , n422138 );
and ( n75639 , n397489 , n68376 );
not ( n75640 , n397489 );
and ( n75641 , n75640 , n41324 );
or ( n75642 , n75639 , n75641 );
buf ( n422144 , n75642 );
not ( n75644 , n422144 );
buf ( n422146 , n73026 );
not ( n75646 , n422146 );
or ( n75647 , n75644 , n75646 );
buf ( n422149 , n421702 );
buf ( n422150 , n41664 );
nand ( n75650 , n422149 , n422150 );
buf ( n422152 , n75650 );
buf ( n422153 , n422152 );
nand ( n75653 , n75647 , n422153 );
buf ( n422155 , n75653 );
buf ( n422156 , n422155 );
not ( n75656 , n422156 );
buf ( n422158 , n75656 );
buf ( n422159 , n422158 );
not ( n75659 , n422159 );
or ( n75660 , n75638 , n75659 );
xor ( n75661 , n74409 , n74435 );
xnor ( n75662 , n75661 , n421010 );
buf ( n422164 , n75662 );
not ( n75664 , n422164 );
buf ( n422166 , n75664 );
buf ( n422167 , n422166 );
nand ( n75667 , n75660 , n422167 );
buf ( n422169 , n75667 );
buf ( n422170 , n422169 );
buf ( n422171 , n422155 );
buf ( n422172 , n422134 );
nand ( n75672 , n422171 , n422172 );
buf ( n422174 , n75672 );
buf ( n422175 , n422174 );
nand ( n75675 , n422170 , n422175 );
buf ( n422177 , n75675 );
buf ( n422178 , n422177 );
not ( n75678 , n422178 );
buf ( n422180 , n75678 );
not ( n75680 , n422180 );
buf ( n422182 , n420971 );
buf ( n422183 , n74439 );
xor ( n75683 , n422182 , n422183 );
buf ( n422185 , n421055 );
xnor ( n75685 , n75683 , n422185 );
buf ( n422187 , n75685 );
not ( n75687 , n422187 );
and ( n75688 , n75680 , n75687 );
buf ( n422190 , n422180 );
buf ( n422191 , n422187 );
nand ( n75691 , n422190 , n422191 );
buf ( n422193 , n75691 );
xor ( n75693 , n420884 , n420888 );
xor ( n75694 , n75693 , n420893 );
buf ( n422196 , n75694 );
buf ( n422197 , n392608 );
not ( n75697 , n422197 );
buf ( n422199 , n420986 );
not ( n75699 , n422199 );
or ( n75700 , n75697 , n75699 );
buf ( n422202 , n371879 );
buf ( n422203 , n420908 );
nand ( n75703 , n422202 , n422203 );
buf ( n422205 , n75703 );
buf ( n422206 , n422205 );
nand ( n75706 , n75700 , n422206 );
buf ( n422208 , n75706 );
not ( n422209 , n422208 );
not ( n75709 , n74375 );
or ( n75710 , n422209 , n75709 );
buf ( n422212 , n421004 );
buf ( n422213 , n43515 );
nand ( n75713 , n422212 , n422213 );
buf ( n422215 , n75713 );
nand ( n75715 , n75710 , n422215 );
or ( n75716 , n422196 , n75715 );
xor ( n75717 , n420675 , n420692 );
xor ( n75718 , n75717 , n420715 );
buf ( n422220 , n75718 );
buf ( n422221 , n63564 );
buf ( n422222 , n63625 );
and ( n75722 , n422221 , n422222 );
buf ( n422224 , n413073 );
buf ( n422225 , n63629 );
and ( n75725 , n422224 , n422225 );
nor ( n75726 , n75722 , n75725 );
buf ( n422228 , n75726 );
buf ( n422229 , n422228 );
buf ( n422230 , n410635 );
or ( n75730 , n422229 , n422230 );
buf ( n422232 , n420743 );
buf ( n422233 , n409504 );
or ( n75733 , n422232 , n422233 );
nand ( n75734 , n75730 , n75733 );
buf ( n422236 , n75734 );
xor ( n75736 , n74018 , n420641 );
xor ( n75737 , n75736 , n420660 );
and ( n75738 , n422236 , n75737 );
buf ( n422240 , n348158 );
not ( n75740 , n422240 );
buf ( n422242 , n420709 );
not ( n75742 , n422242 );
buf ( n422244 , n75742 );
buf ( n422245 , n422244 );
not ( n75745 , n422245 );
or ( n75746 , n75740 , n75745 );
buf ( n422248 , n62278 );
buf ( n422249 , n66411 );
and ( n75749 , n422248 , n422249 );
buf ( n422251 , n409474 );
buf ( n422252 , n62496 );
and ( n75752 , n422251 , n422252 );
nor ( n75753 , n75749 , n75752 );
buf ( n422255 , n75753 );
buf ( n422256 , n422255 );
buf ( n422257 , n410724 );
or ( n75757 , n422256 , n422257 );
nand ( n75758 , n75746 , n75757 );
buf ( n422260 , n75758 );
xor ( n75760 , n74018 , n420641 );
xor ( n75761 , n75760 , n420660 );
and ( n75762 , n422260 , n75761 );
and ( n75763 , n422236 , n422260 );
or ( n75764 , n75738 , n75762 , n75763 );
xor ( n75765 , n422220 , n75764 );
xor ( n75766 , n420791 , n420836 );
xor ( n75767 , n75766 , n420856 );
buf ( n422269 , n75767 );
buf ( n422270 , n66359 );
buf ( n422271 , n62177 );
and ( n75771 , n422270 , n422271 );
buf ( n422273 , n413187 );
buf ( n422274 , n62159 );
and ( n75774 , n422273 , n422274 );
nor ( n75775 , n75771 , n75774 );
buf ( n422277 , n75775 );
buf ( n422278 , n422277 );
buf ( n422279 , n409429 );
or ( n75779 , n422278 , n422279 );
buf ( n422281 , n420760 );
buf ( n422282 , n409170 );
or ( n75782 , n422281 , n422282 );
nand ( n75783 , n75779 , n75782 );
buf ( n422285 , n75783 );
xor ( n75785 , n422269 , n422285 );
buf ( n422287 , n409507 );
not ( n75787 , n422287 );
buf ( n422289 , n63707 );
buf ( n422290 , n63625 );
and ( n75790 , n422289 , n422290 );
buf ( n422292 , n413104 );
buf ( n422293 , n63629 );
and ( n75793 , n422292 , n422293 );
nor ( n75794 , n75790 , n75793 );
buf ( n422296 , n75794 );
buf ( n422297 , n422296 );
not ( n75797 , n422297 );
buf ( n422299 , n75797 );
buf ( n422300 , n422299 );
not ( n75800 , n422300 );
or ( n75801 , n75787 , n75800 );
buf ( n422303 , n422228 );
buf ( n422304 , n409504 );
or ( n75804 , n422303 , n422304 );
nand ( n75805 , n75801 , n75804 );
buf ( n422307 , n75805 );
and ( n75807 , n75785 , n422307 );
and ( n75808 , n422269 , n422285 );
or ( n75809 , n75807 , n75808 );
buf ( n422311 , n75809 );
buf ( n422312 , n401623 );
buf ( n422313 , n623 );
not ( n75813 , n422313 );
buf ( n422315 , n75813 );
buf ( n422316 , n422315 );
nor ( n75816 , n422312 , n422316 );
buf ( n422318 , n75816 );
buf ( n422319 , n422318 );
buf ( n422320 , n56041 );
buf ( n422321 , n71170 );
and ( n75821 , n422320 , n422321 );
buf ( n422323 , n403298 );
buf ( n422324 , n417804 );
and ( n75824 , n422323 , n422324 );
nor ( n75825 , n75821 , n75824 );
buf ( n422327 , n75825 );
buf ( n422328 , n422327 );
buf ( n422329 , n403293 );
or ( n75829 , n422328 , n422329 );
buf ( n422331 , n71088 );
buf ( n422332 , n56041 );
and ( n75832 , n422331 , n422332 );
buf ( n422334 , n417722 );
buf ( n422335 , n403298 );
and ( n75835 , n422334 , n422335 );
nor ( n75836 , n75832 , n75835 );
buf ( n422338 , n75836 );
buf ( n422339 , n422338 );
buf ( n422340 , n405476 );
or ( n75840 , n422339 , n422340 );
nand ( n75841 , n75829 , n75840 );
buf ( n422343 , n75841 );
buf ( n422344 , n422343 );
and ( n75844 , n422319 , n422344 );
buf ( n422346 , n75844 );
buf ( n422347 , n422346 );
buf ( n422348 , n403293 );
buf ( n422349 , n422338 );
or ( n75849 , n422348 , n422349 );
buf ( n422351 , n420599 );
buf ( n422352 , n405476 );
or ( n75852 , n422351 , n422352 );
nand ( n75853 , n75849 , n75852 );
buf ( n422355 , n75853 );
buf ( n422356 , n422355 );
xor ( n75856 , n422347 , n422356 );
buf ( n422358 , n405381 );
not ( n75858 , n422358 );
buf ( n422360 , n420782 );
not ( n75860 , n422360 );
buf ( n422362 , n75860 );
buf ( n422363 , n422362 );
not ( n75863 , n422363 );
or ( n75864 , n75858 , n75863 );
buf ( n422366 , n70389 );
buf ( n422367 , n405391 );
and ( n75867 , n422366 , n422367 );
buf ( n422369 , n417024 );
buf ( n422370 , n405388 );
and ( n75870 , n422369 , n422370 );
nor ( n75871 , n75867 , n75870 );
buf ( n422373 , n75871 );
buf ( n422374 , n422373 );
buf ( n422375 , n405407 );
or ( n75875 , n422374 , n422375 );
nand ( n75876 , n75864 , n75875 );
buf ( n422378 , n75876 );
buf ( n422379 , n422378 );
and ( n75879 , n75856 , n422379 );
and ( n75880 , n422347 , n422356 );
or ( n75881 , n75879 , n75880 );
buf ( n422383 , n75881 );
xor ( n75883 , n420607 , n420619 );
xor ( n75884 , n75883 , n420622 );
and ( n75885 , n422383 , n75884 );
buf ( n422387 , n403120 );
buf ( n422388 , n15287 );
buf ( n422389 , n71681 );
and ( n75889 , n422388 , n422389 );
buf ( n422391 , n55895 );
buf ( n422392 , n418315 );
and ( n75892 , n422391 , n422392 );
nor ( n75893 , n75889 , n75892 );
buf ( n422395 , n75893 );
buf ( n422396 , n422395 );
or ( n75896 , n422387 , n422396 );
buf ( n422398 , n420823 );
buf ( n422399 , n403108 );
or ( n75899 , n422398 , n422399 );
nand ( n75900 , n75896 , n75899 );
buf ( n422402 , n75900 );
buf ( n422403 , n422402 );
buf ( n422404 , n403158 );
buf ( n422405 , n418921 );
buf ( n422406 , n74002 );
and ( n75906 , n422405 , n422406 );
buf ( n422408 , n401678 );
buf ( n422409 , n420612 );
and ( n75909 , n422408 , n422409 );
nor ( n75910 , n75906 , n75909 );
buf ( n422412 , n75910 );
buf ( n422413 , n422412 );
or ( n75913 , n422404 , n422413 );
buf ( n422415 , n420800 );
buf ( n422416 , n403167 );
or ( n75916 , n422415 , n422416 );
nand ( n75917 , n75913 , n75916 );
buf ( n422419 , n75917 );
buf ( n422420 , n422419 );
xor ( n75920 , n422403 , n422420 );
buf ( n422422 , n401650 );
buf ( n422423 , n623 );
and ( n75923 , n422422 , n422423 );
buf ( n422425 , n75923 );
buf ( n422426 , n422425 );
buf ( n422427 , n403293 );
buf ( n422428 , n56041 );
buf ( n422429 , n71664 );
and ( n75929 , n422428 , n422429 );
buf ( n422431 , n403298 );
buf ( n422432 , n418298 );
and ( n75932 , n422431 , n422432 );
nor ( n75933 , n75929 , n75932 );
buf ( n422435 , n75933 );
buf ( n422436 , n422435 );
or ( n75936 , n422427 , n422436 );
buf ( n422438 , n422327 );
buf ( n422439 , n403290 );
or ( n75939 , n422438 , n422439 );
nand ( n75940 , n75936 , n75939 );
buf ( n422442 , n75940 );
buf ( n422443 , n422442 );
and ( n75943 , n422426 , n422443 );
buf ( n422445 , n75943 );
buf ( n422446 , n422445 );
and ( n75946 , n75920 , n422446 );
and ( n75947 , n422403 , n422420 );
or ( n75948 , n75946 , n75947 );
buf ( n422450 , n75948 );
xor ( n75950 , n420808 , n420813 );
xor ( n75951 , n75950 , n420831 );
buf ( n422453 , n75951 );
xor ( n75953 , n422450 , n422453 );
buf ( n422455 , n59471 );
not ( n75955 , n422455 );
buf ( n422457 , n420850 );
not ( n75957 , n422457 );
buf ( n422459 , n75957 );
buf ( n422460 , n422459 );
not ( n75960 , n422460 );
or ( n75961 , n75955 , n75960 );
buf ( n422463 , n70195 );
buf ( n422464 , n59628 );
and ( n75964 , n422463 , n422464 );
buf ( n422466 , n416830 );
buf ( n422467 , n58223 );
and ( n75967 , n422466 , n422467 );
nor ( n75968 , n75964 , n75967 );
buf ( n422470 , n75968 );
buf ( n422471 , n422470 );
buf ( n422472 , n59637 );
or ( n75972 , n422471 , n422472 );
nand ( n75973 , n75961 , n75972 );
buf ( n422475 , n75973 );
and ( n75975 , n75953 , n422475 );
and ( n75976 , n422450 , n422453 );
or ( n75977 , n75975 , n75976 );
xor ( n75978 , n420607 , n420619 );
xor ( n75979 , n75978 , n420622 );
and ( n75980 , n75977 , n75979 );
and ( n75981 , n422383 , n75977 );
or ( n422483 , n75885 , n75980 , n75981 );
buf ( n422484 , n422483 );
xor ( n75984 , n422311 , n422484 );
xor ( n75985 , n420769 , n420773 );
xor ( n75986 , n75985 , n420861 );
buf ( n422488 , n75986 );
buf ( n422489 , n422488 );
and ( n75989 , n75984 , n422489 );
and ( n75990 , n422311 , n422484 );
or ( n75991 , n75989 , n75990 );
buf ( n422493 , n75991 );
and ( n75993 , n75765 , n422493 );
and ( n75994 , n422220 , n75764 );
or ( n75995 , n75993 , n75994 );
xor ( n75996 , n420735 , n420875 );
xor ( n75997 , n75996 , n74273 );
and ( n75998 , n75995 , n75997 );
xor ( n75999 , n420752 , n420866 );
xor ( n76000 , n75999 , n420871 );
buf ( n422502 , n76000 );
xor ( n76002 , n422220 , n75764 );
xor ( n76003 , n76002 , n422493 );
and ( n76004 , n422502 , n76003 );
xor ( n76005 , n74018 , n420641 );
xor ( n76006 , n76005 , n420660 );
xor ( n76007 , n422236 , n422260 );
xor ( n76008 , n76006 , n76007 );
buf ( n422510 , n62467 );
buf ( n422511 , n66411 );
and ( n76011 , n422510 , n422511 );
buf ( n422513 , n409468 );
buf ( n422514 , n62496 );
and ( n76014 , n422513 , n422514 );
nor ( n76015 , n76011 , n76014 );
buf ( n422517 , n76015 );
buf ( n422518 , n422517 );
buf ( n422519 , n410724 );
or ( n76019 , n422518 , n422519 );
buf ( n422521 , n422255 );
buf ( n422522 , n410721 );
or ( n76022 , n422521 , n422522 );
nand ( n76023 , n76019 , n76022 );
buf ( n422525 , n76023 );
buf ( n422526 , n422525 );
xor ( n76026 , n422347 , n422356 );
xor ( n76027 , n76026 , n422379 );
buf ( n422529 , n76027 );
buf ( n422530 , n422529 );
buf ( n422531 , n56050 );
buf ( n422532 , n71095 );
and ( n76032 , n422531 , n422532 );
not ( n76033 , n422531 );
buf ( n422535 , n417729 );
and ( n76035 , n76033 , n422535 );
nor ( n76036 , n76032 , n76035 );
buf ( n422538 , n76036 );
buf ( n422539 , n422538 );
not ( n76039 , n422539 );
buf ( n422541 , n76039 );
buf ( n422542 , n422541 );
buf ( n422543 , n405407 );
or ( n76043 , n422542 , n422543 );
buf ( n422545 , n422373 );
buf ( n422546 , n405378 );
or ( n76046 , n422545 , n422546 );
nand ( n76047 , n76043 , n76046 );
buf ( n422549 , n76047 );
buf ( n422550 , n422549 );
xor ( n76050 , n422319 , n422344 );
buf ( n422552 , n76050 );
buf ( n422553 , n422552 );
xor ( n76053 , n422550 , n422553 );
buf ( n422555 , n422412 );
buf ( n422556 , n401660 );
or ( n76056 , n422555 , n422556 );
buf ( n422558 , n401681 );
nand ( n76058 , n76056 , n422558 );
buf ( n422560 , n76058 );
buf ( n422561 , n422560 );
buf ( n422562 , n403120 );
buf ( n422563 , n55905 );
buf ( n422564 , n72308 );
and ( n76064 , n422563 , n422564 );
buf ( n422566 , n55895 );
buf ( n422567 , n418942 );
and ( n76067 , n422566 , n422567 );
nor ( n76068 , n76064 , n76067 );
buf ( n422570 , n76068 );
buf ( n422571 , n422570 );
or ( n76071 , n422562 , n422571 );
buf ( n422573 , n422395 );
buf ( n422574 , n403108 );
or ( n76074 , n422573 , n422574 );
nand ( n76075 , n76071 , n76074 );
buf ( n422577 , n76075 );
buf ( n422578 , n422577 );
xor ( n76078 , n422561 , n422578 );
buf ( n422580 , n405381 );
not ( n76080 , n422580 );
buf ( n422582 , n422538 );
not ( n76082 , n422582 );
or ( n76083 , n76080 , n76082 );
buf ( n422585 , n405407 );
buf ( n422586 , n403283 );
buf ( n422587 , n71088 );
and ( n76087 , n422586 , n422587 );
buf ( n422589 , n417722 );
buf ( n422590 , n56050 );
and ( n76090 , n422589 , n422590 );
nor ( n76091 , n76087 , n76090 );
buf ( n422593 , n76091 );
buf ( n422594 , n422593 );
or ( n76094 , n422585 , n422594 );
nand ( n76095 , n76083 , n76094 );
buf ( n422597 , n76095 );
buf ( n422598 , n422597 );
and ( n76098 , n76078 , n422598 );
and ( n76099 , n422561 , n422578 );
or ( n76100 , n76098 , n76099 );
buf ( n422602 , n76100 );
buf ( n422603 , n422602 );
and ( n76103 , n76053 , n422603 );
and ( n76104 , n422550 , n422553 );
or ( n76105 , n76103 , n76104 );
buf ( n422607 , n76105 );
buf ( n422608 , n422607 );
xor ( n76108 , n422530 , n422608 );
buf ( n422610 , n409173 );
not ( n422611 , n422610 );
buf ( n422612 , n414714 );
buf ( n422613 , n62159 );
or ( n76113 , n422612 , n422613 );
buf ( n422615 , n67987 );
buf ( n422616 , n62177 );
or ( n76116 , n422615 , n422616 );
nand ( n76117 , n76113 , n76116 );
buf ( n422619 , n76117 );
buf ( n422620 , n422619 );
not ( n76120 , n422620 );
or ( n76121 , n422611 , n76120 );
buf ( n422623 , n422277 );
buf ( n422624 , n409170 );
or ( n76124 , n422623 , n422624 );
nand ( n76125 , n76121 , n76124 );
buf ( n422627 , n76125 );
buf ( n422628 , n422627 );
and ( n76128 , n76108 , n422628 );
and ( n76129 , n422530 , n422608 );
or ( n76130 , n76128 , n76129 );
buf ( n422632 , n76130 );
buf ( n422633 , n422632 );
xor ( n76133 , n422526 , n422633 );
xor ( n76134 , n420607 , n420619 );
xor ( n76135 , n76134 , n420622 );
xor ( n76136 , n422383 , n75977 );
xor ( n76137 , n76135 , n76136 );
buf ( n422639 , n76137 );
and ( n76139 , n76133 , n422639 );
and ( n76140 , n422526 , n422633 );
or ( n76141 , n76139 , n76140 );
buf ( n422643 , n76141 );
xor ( n76143 , n76008 , n422643 );
xor ( n76144 , n422311 , n422484 );
xor ( n76145 , n76144 , n422489 );
buf ( n422647 , n76145 );
and ( n76147 , n76143 , n422647 );
and ( n76148 , n76008 , n422643 );
or ( n76149 , n76147 , n76148 );
xor ( n76150 , n422220 , n75764 );
xor ( n76151 , n76150 , n422493 );
and ( n76152 , n76149 , n76151 );
and ( n76153 , n422502 , n76149 );
or ( n76154 , n76004 , n76152 , n76153 );
xor ( n76155 , n420735 , n420875 );
xor ( n76156 , n76155 , n74273 );
and ( n76157 , n76154 , n76156 );
and ( n76158 , n75995 , n76154 );
or ( n76159 , n75998 , n76157 , n76158 );
nand ( n76160 , n75716 , n76159 );
nand ( n76161 , n75715 , n422196 );
nand ( n76162 , n76160 , n76161 );
buf ( n422664 , n76162 );
buf ( n422665 , n44775 );
not ( n76165 , n422665 );
buf ( n422667 , n418729 );
not ( n76167 , n422667 );
or ( n76168 , n76165 , n76167 );
buf ( n422670 , n41861 );
buf ( n422671 , n44775 );
not ( n76171 , n422671 );
buf ( n422673 , n76171 );
buf ( n422674 , n422673 );
nand ( n76174 , n422670 , n422674 );
buf ( n422676 , n76174 );
buf ( n422677 , n422676 );
nand ( n76177 , n76168 , n422677 );
buf ( n422679 , n76177 );
not ( n76179 , n422679 );
not ( n76180 , n417542 );
or ( n76181 , n76179 , n76180 );
or ( n76182 , n421680 , n392224 );
nand ( n76183 , n76181 , n76182 );
buf ( n422685 , n76183 );
xor ( n76185 , n422664 , n422685 );
buf ( n422687 , n394210 );
not ( n76187 , n422687 );
buf ( n422689 , n418734 );
not ( n76189 , n422689 );
or ( n76190 , n76187 , n76189 );
buf ( n422692 , n388722 );
buf ( n422693 , n394219 );
nand ( n76193 , n422692 , n422693 );
buf ( n422695 , n76193 );
buf ( n422696 , n422695 );
nand ( n76196 , n76190 , n422696 );
buf ( n422698 , n76196 );
buf ( n422699 , n422698 );
not ( n76199 , n422699 );
buf ( n422701 , n67042 );
not ( n76201 , n422701 );
or ( n76202 , n76199 , n76201 );
buf ( n422704 , n421034 );
buf ( n422705 , n388068 );
nand ( n76205 , n422704 , n422705 );
buf ( n422707 , n76205 );
buf ( n422708 , n422707 );
nand ( n76208 , n76202 , n422708 );
buf ( n422710 , n76208 );
buf ( n422711 , n422710 );
not ( n76211 , n75715 );
buf ( n422713 , n76159 );
buf ( n422714 , n422196 );
xnor ( n76214 , n422713 , n422714 );
buf ( n422716 , n76214 );
not ( n76216 , n422716 );
or ( n76217 , n76211 , n76216 );
or ( n76218 , n75715 , n422716 );
nand ( n76219 , n76217 , n76218 );
buf ( n422721 , n76219 );
xor ( n76221 , n422711 , n422721 );
buf ( n422723 , n413643 );
not ( n76223 , n422723 );
buf ( n422725 , n422679 );
not ( n76225 , n422725 );
or ( n76226 , n76223 , n76225 );
buf ( n422728 , n44775 );
not ( n76228 , n422728 );
buf ( n422730 , n420954 );
not ( n76230 , n422730 );
or ( n76231 , n76228 , n76230 );
buf ( n422733 , n389338 );
buf ( n422734 , n422673 );
nand ( n76234 , n422733 , n422734 );
buf ( n422736 , n76234 );
buf ( n422737 , n422736 );
nand ( n76237 , n76231 , n422737 );
buf ( n422739 , n76237 );
buf ( n422740 , n422739 );
buf ( n422741 , n417542 );
nand ( n76241 , n422740 , n422741 );
buf ( n422743 , n76241 );
buf ( n422744 , n422743 );
nand ( n76244 , n76226 , n422744 );
buf ( n422746 , n76244 );
buf ( n422747 , n422746 );
and ( n76247 , n76221 , n422747 );
and ( n76248 , n422711 , n422721 );
or ( n76249 , n76247 , n76248 );
buf ( n422751 , n76249 );
buf ( n422752 , n422751 );
and ( n76252 , n76185 , n422752 );
and ( n76253 , n422664 , n422685 );
or ( n76254 , n76252 , n76253 );
buf ( n422756 , n76254 );
and ( n76256 , n422193 , n422756 );
nor ( n76257 , n75688 , n76256 );
or ( n76258 , n75608 , n76257 );
nand ( n76259 , n422108 , n422080 );
nand ( n76260 , n76258 , n76259 );
buf ( n422762 , n76260 );
and ( n76262 , n75520 , n422762 );
and ( n76263 , n422016 , n422020 );
or ( n76264 , n76262 , n76263 );
buf ( n422766 , n76264 );
xor ( n76279 , n422766 , C0 );
xor ( n76280 , n420058 , n420096 );
xor ( n76281 , n76280 , n420137 );
buf ( n422770 , n76281 );
and ( n76283 , n76279 , n422770 );
or ( n76285 , n76283 , C0 );
buf ( n422773 , n76285 );
buf ( n422774 , C0 );
buf ( n422775 , n422774 );
buf ( n422776 , n61577 );
not ( n76310 , n422776 );
buf ( n422778 , n421789 );
not ( n76312 , n422778 );
or ( n76313 , n76310 , n76312 );
buf ( n422781 , n47891 );
buf ( n422782 , n46481 );
and ( n76316 , n422781 , n422782 );
not ( n76317 , n422781 );
buf ( n422785 , n46478 );
and ( n76319 , n76317 , n422785 );
nor ( n76320 , n76316 , n76319 );
buf ( n422788 , n76320 );
buf ( n422789 , n422788 );
buf ( n422790 , n50579 );
nand ( n76324 , n422789 , n422790 );
buf ( n422792 , n76324 );
buf ( n422793 , n422792 );
nand ( n76327 , n76313 , n422793 );
buf ( n422795 , n76327 );
buf ( n422796 , n422795 );
xor ( n76330 , n75117 , n75233 );
xor ( n76331 , n76330 , n75249 );
buf ( n422799 , n76331 );
xor ( n76333 , n422796 , n422799 );
buf ( n422801 , n41563 );
buf ( n422802 , n358975 );
nand ( n76336 , n422801 , n422802 );
buf ( n422804 , n76336 );
buf ( n422805 , n422804 );
not ( n76339 , n422805 );
buf ( n422807 , n55055 );
not ( n76341 , n422807 );
buf ( n422809 , n56919 );
not ( n76343 , n422809 );
or ( n76344 , n76341 , n76343 );
buf ( n422812 , n41559 );
buf ( n422813 , n404855 );
nand ( n76347 , n422812 , n422813 );
buf ( n422815 , n76347 );
buf ( n422816 , n422815 );
nand ( n76350 , n76344 , n422816 );
buf ( n422818 , n76350 );
buf ( n422819 , n422818 );
not ( n76353 , n422819 );
buf ( n422821 , n52812 );
not ( n76355 , n422821 );
or ( n76356 , n76353 , n76355 );
buf ( n422824 , n421839 );
buf ( n422825 , n400143 );
nand ( n76359 , n422824 , n422825 );
buf ( n422827 , n76359 );
buf ( n422828 , n422827 );
nand ( n76362 , n76356 , n422828 );
buf ( n422830 , n76362 );
buf ( n422831 , n422830 );
not ( n76365 , n422831 );
buf ( n422833 , n76365 );
buf ( n422834 , n422833 );
not ( n76368 , n422834 );
or ( n76369 , n76339 , n76368 );
xor ( n76370 , n421719 , n75204 );
xor ( n76371 , n76370 , n421752 );
buf ( n422839 , n76371 );
nand ( n76373 , n76369 , n422839 );
buf ( n422841 , n76373 );
buf ( n422842 , n422841 );
buf ( n422843 , n422804 );
not ( n76377 , n422843 );
buf ( n422845 , n422830 );
nand ( n76379 , n76377 , n422845 );
buf ( n422847 , n76379 );
buf ( n422848 , n422847 );
nand ( n76382 , n422842 , n422848 );
buf ( n422850 , n76382 );
buf ( n422851 , n422850 );
and ( n76385 , n76333 , n422851 );
and ( n76386 , n422796 , n422799 );
or ( n76387 , n76385 , n76386 );
buf ( n422855 , n76387 );
buf ( n422856 , n422855 );
xor ( n76390 , n422775 , n422856 );
xor ( n76391 , n421618 , n421774 );
xor ( n76392 , n76391 , n421800 );
buf ( n422860 , n76392 );
buf ( n422861 , n422860 );
and ( n76395 , n76390 , n422861 );
or ( n76397 , n76395 , C0 );
buf ( n422864 , n76397 );
buf ( n422865 , n422864 );
xor ( n76400 , n422773 , n422865 );
xor ( n76401 , n73763 , n421112 );
xor ( n76402 , n76401 , n420395 );
buf ( n422869 , n76402 );
and ( n76404 , n76400 , n422869 );
and ( n76405 , n422773 , n422865 );
or ( n76406 , n76404 , n76405 );
buf ( n422873 , n76406 );
buf ( n422874 , n422873 );
nand ( n76409 , n75450 , n422874 );
buf ( n422876 , n76409 );
buf ( n422877 , n422876 );
not ( n76412 , n422877 );
buf ( n422879 , n75439 );
not ( n76414 , n422879 );
buf ( n422881 , n76414 );
buf ( n422882 , n422881 );
buf ( n422883 , n421948 );
not ( n76418 , n422883 );
buf ( n422885 , n76418 );
buf ( n422886 , n422885 );
and ( n76421 , n422882 , n422886 );
buf ( n422888 , n76421 );
buf ( n422889 , n422888 );
nor ( n76424 , n76412 , n422889 );
buf ( n422891 , n76424 );
buf ( n422892 , n422891 );
not ( n76427 , n422892 );
buf ( n422894 , n76427 );
buf ( n422895 , n422894 );
nand ( n76430 , n75437 , n422895 );
buf ( n422897 , n76430 );
buf ( n422898 , n422897 );
buf ( n422899 , n421935 );
not ( n76434 , n422899 );
buf ( n422901 , n421133 );
nand ( n76436 , n76434 , n422901 );
buf ( n422903 , n76436 );
buf ( n422904 , n422903 );
nand ( n76439 , n422898 , n422904 );
buf ( n422906 , n76439 );
buf ( n422907 , n422906 );
buf ( n422908 , n413643 );
not ( n76443 , n422908 );
buf ( n422910 , n399986 );
not ( n76445 , n422910 );
buf ( n422912 , n46478 );
not ( n76447 , n422912 );
or ( n76448 , n76445 , n76447 );
buf ( n422915 , n49686 );
buf ( n422916 , n44776 );
nand ( n76451 , n422915 , n422916 );
buf ( n422918 , n76451 );
buf ( n422919 , n422918 );
nand ( n76454 , n76448 , n422919 );
buf ( n422921 , n76454 );
buf ( n422922 , n422921 );
not ( n76457 , n422922 );
or ( n422924 , n76443 , n76457 );
buf ( n422925 , n417523 );
buf ( n422926 , n417542 );
nand ( n76461 , n422925 , n422926 );
buf ( n422928 , n76461 );
buf ( n422929 , n422928 );
nand ( n76464 , n422924 , n422929 );
buf ( n422931 , n76464 );
buf ( n422932 , n422931 );
buf ( n422933 , n419742 );
not ( n76468 , n422933 );
buf ( n422935 , n389122 );
not ( n76470 , n422935 );
or ( n76471 , n76468 , n76470 );
buf ( n422938 , n49117 );
not ( n76473 , n422938 );
buf ( n422940 , n398298 );
not ( n76475 , n422940 );
or ( n76476 , n76473 , n76475 );
buf ( n422943 , n24049 );
buf ( n422944 , n67126 );
nand ( n76479 , n422943 , n422944 );
buf ( n422946 , n76479 );
buf ( n422947 , n422946 );
nand ( n76482 , n76476 , n422947 );
buf ( n422949 , n76482 );
buf ( n422950 , n422949 );
buf ( n422951 , n46921 );
nand ( n76486 , n422950 , n422951 );
buf ( n422953 , n76486 );
buf ( n422954 , n422953 );
nand ( n76489 , n76471 , n422954 );
buf ( n422956 , n76489 );
buf ( n422957 , n422956 );
xor ( n76492 , n422932 , n422957 );
buf ( n422959 , n73162 );
not ( n76494 , n422959 );
buf ( n422961 , n38961 );
not ( n76496 , n422961 );
or ( n76497 , n76494 , n76496 );
and ( n76498 , n51183 , n22982 );
not ( n76499 , n51183 );
and ( n76500 , n76499 , n49661 );
nor ( n76501 , n76498 , n76500 );
nand ( n76502 , n76501 , n395199 );
buf ( n422969 , n76502 );
nand ( n76504 , n76497 , n422969 );
buf ( n422971 , n76504 );
buf ( n422972 , n422971 );
xor ( n76507 , n76492 , n422972 );
buf ( n422974 , n76507 );
buf ( n422975 , n422974 );
buf ( n422976 , C0 );
buf ( n422977 , n422976 );
xor ( n76538 , n422975 , n422977 );
buf ( n422979 , n421443 );
not ( n76540 , n422979 );
buf ( n422981 , n421403 );
not ( n76542 , n422981 );
or ( n76543 , n76540 , n76542 );
buf ( n422984 , n421446 );
not ( n76545 , n422984 );
buf ( n422986 , n421406 );
not ( n76547 , n422986 );
or ( n76548 , n76545 , n76547 );
buf ( n422989 , n421379 );
nand ( n76550 , n76548 , n422989 );
buf ( n422991 , n76550 );
buf ( n422992 , n422991 );
nand ( n76553 , n76543 , n422992 );
buf ( n422994 , n76553 );
buf ( n422995 , n422994 );
xor ( n76556 , n76538 , n422995 );
buf ( n422997 , n76556 );
buf ( n422998 , n422997 );
buf ( n422999 , n421367 );
not ( n76560 , n422999 );
buf ( n423001 , n421453 );
nand ( n423002 , n76560 , n423001 );
buf ( n423003 , n423002 );
buf ( n423004 , n423003 );
buf ( n423005 , n421372 );
and ( n76566 , n423004 , n423005 );
buf ( n423007 , n421367 );
not ( n76568 , n423007 );
buf ( n423009 , n421453 );
nor ( n76570 , n76568 , n423009 );
buf ( n423011 , n76570 );
buf ( n423012 , n423011 );
nor ( n76573 , n76566 , n423012 );
buf ( n423014 , n76573 );
buf ( n423015 , n423014 );
not ( n76576 , n423015 );
buf ( n423017 , n76576 );
buf ( n423018 , n423017 );
xor ( n76579 , n422998 , n423018 );
buf ( n423020 , n421295 );
not ( n76581 , n423020 );
buf ( n423022 , n52812 );
not ( n76583 , n423022 );
or ( n76584 , n76581 , n76583 );
buf ( n423025 , n394210 );
not ( n76586 , n423025 );
buf ( n423027 , n51822 );
not ( n76588 , n423027 );
or ( n76589 , n76586 , n76588 );
buf ( n423030 , n60880 );
buf ( n423031 , n394207 );
nand ( n76592 , n423030 , n423031 );
buf ( n423033 , n76592 );
buf ( n423034 , n423033 );
nand ( n76595 , n76589 , n423034 );
buf ( n423036 , n76595 );
buf ( n423037 , n423036 );
buf ( n423038 , n42924 );
nand ( n76599 , n423037 , n423038 );
buf ( n423040 , n76599 );
buf ( n423041 , n423040 );
nand ( n76602 , n76584 , n423041 );
buf ( n423043 , n76602 );
buf ( n423044 , n43515 );
not ( n76605 , n423044 );
and ( n76606 , n28644 , n391024 );
not ( n76607 , n28644 );
and ( n76608 , n76607 , n411504 );
or ( n76609 , n76606 , n76608 );
buf ( n423050 , n76609 );
not ( n76611 , n423050 );
or ( n76612 , n76605 , n76611 );
buf ( n423053 , n421262 );
buf ( n423054 , n43536 );
nand ( n76615 , n423053 , n423054 );
buf ( n423056 , n76615 );
buf ( n423057 , n423056 );
nand ( n76618 , n76612 , n423057 );
buf ( n423059 , n76618 );
xor ( n76620 , n423043 , n423059 );
xor ( n76621 , n421178 , n421187 );
and ( n76622 , n76621 , n421214 );
and ( n76623 , n421178 , n421187 );
or ( n76624 , n76622 , n76623 );
buf ( n423065 , n76624 );
buf ( n423066 , n423065 );
buf ( n423067 , n421235 );
not ( n76628 , n423067 );
buf ( n423069 , n66128 );
not ( n76630 , n423069 );
or ( n76631 , n76628 , n76630 );
buf ( n423072 , n417380 );
buf ( n423073 , n412976 );
nand ( n76634 , n423072 , n423073 );
buf ( n423075 , n76634 );
buf ( n423076 , n423075 );
nand ( n76637 , n76631 , n423076 );
buf ( n423078 , n76637 );
buf ( n423079 , n423078 );
xor ( n76640 , n423066 , n423079 );
not ( n76641 , n70287 );
and ( n76642 , n70598 , n76641 );
not ( n76643 , n70601 );
and ( n76644 , n70598 , n76643 );
nor ( n76645 , n76642 , n76644 );
not ( n76646 , n416779 );
not ( n76647 , n70598 );
nand ( n76648 , n76646 , n76647 , n70286 );
not ( n76649 , n70286 );
nand ( n76650 , n76649 , n76647 , n416779 );
nand ( n76651 , n76645 , n76648 , n76650 );
buf ( n423092 , n421163 );
not ( n76653 , n423092 );
buf ( n423094 , n416762 );
not ( n76655 , n423094 );
or ( n76656 , n76653 , n76655 );
buf ( n423097 , n416758 );
buf ( n423098 , n41664 );
nand ( n76659 , n423097 , n423098 );
buf ( n423100 , n76659 );
buf ( n423101 , n423100 );
nand ( n76662 , n76656 , n423101 );
buf ( n423103 , n76662 );
xor ( n76664 , n76651 , n423103 );
buf ( n423105 , n388803 );
not ( n76666 , n423105 );
buf ( n423107 , n417359 );
not ( n76668 , n423107 );
or ( n76669 , n76666 , n76668 );
buf ( n423110 , n421203 );
buf ( n423111 , n388740 );
nand ( n76672 , n423110 , n423111 );
buf ( n423113 , n76672 );
buf ( n423114 , n423113 );
nand ( n76675 , n76669 , n423114 );
buf ( n423116 , n76675 );
xor ( n76677 , n76664 , n423116 );
buf ( n423118 , n76677 );
xnor ( n76679 , n76640 , n423118 );
buf ( n423120 , n76679 );
xnor ( n76681 , n76620 , n423120 );
buf ( n423122 , n76681 );
buf ( n423123 , n395349 );
not ( n76684 , n423123 );
buf ( n423125 , n421393 );
not ( n76686 , n423125 );
or ( n76687 , n76684 , n76686 );
buf ( n423128 , n47863 );
not ( n76689 , n423128 );
buf ( n423130 , n50317 );
not ( n76691 , n423130 );
or ( n76692 , n76689 , n76691 );
buf ( n423133 , n40818 );
buf ( n423134 , n419385 );
nand ( n76695 , n423133 , n423134 );
buf ( n423136 , n76695 );
buf ( n423137 , n423136 );
nand ( n76698 , n76692 , n423137 );
buf ( n423139 , n76698 );
buf ( n423140 , n423139 );
buf ( n423141 , n395362 );
nand ( n76702 , n423140 , n423141 );
buf ( n423143 , n76702 );
buf ( n423144 , n423143 );
nand ( n76705 , n76687 , n423144 );
buf ( n423146 , n76705 );
buf ( n423147 , n423146 );
xor ( n76708 , n423122 , n423147 );
xor ( n76709 , n417549 , n417568 );
and ( n76710 , n76709 , n418697 );
and ( n76711 , n417549 , n417568 );
or ( n76712 , n76710 , n76711 );
buf ( n423153 , n76712 );
buf ( n423154 , n423153 );
xor ( n76715 , n76708 , n423154 );
buf ( n423156 , n76715 );
buf ( n423157 , n423156 );
buf ( n423158 , C0 );
xor ( n76735 , n423157 , n423158 );
xor ( n76736 , n418700 , n419419 );
and ( n76737 , n76736 , n419451 );
and ( n76738 , n418700 , n419419 );
or ( n76739 , n76737 , n76738 );
buf ( n423164 , n76739 );
buf ( n423165 , n423164 );
xor ( n76742 , n76735 , n423165 );
buf ( n423167 , n76742 );
buf ( n423168 , n423167 );
xor ( n76745 , n76579 , n423168 );
buf ( n423170 , n76745 );
buf ( n423171 , n423170 );
buf ( n423172 , n421463 );
not ( n76749 , n423172 );
buf ( n423174 , n421584 );
not ( n76751 , n423174 );
or ( n423176 , n76749 , n76751 );
buf ( n423177 , n421466 );
not ( n76754 , n423177 );
buf ( n423179 , n421581 );
not ( n76756 , n423179 );
or ( n76757 , n76754 , n76756 );
buf ( n423182 , n421925 );
nand ( n76759 , n76757 , n423182 );
buf ( n423184 , n76759 );
buf ( n423185 , n423184 );
nand ( n76762 , n423176 , n423185 );
buf ( n423187 , n76762 );
buf ( n423188 , n423187 );
xor ( n76765 , n423171 , n423188 );
buf ( n423190 , n421571 );
not ( n76774 , n423190 );
or ( n76775 , C0 , n76774 );
buf ( n423193 , n421544 );
nand ( n76777 , n76775 , n423193 );
buf ( n423195 , n76777 );
buf ( n423196 , n423195 );
nand ( n76780 , C1 , n423196 );
buf ( n423198 , n76780 );
buf ( n423199 , n423198 );
xor ( n76783 , n419454 , n419805 );
and ( n76784 , n76783 , n421131 );
and ( n76785 , n419454 , n419805 );
or ( n76786 , n76784 , n76785 );
buf ( n423204 , n76786 );
buf ( n423205 , n423204 );
xor ( n76789 , n423199 , n423205 );
buf ( n423207 , n421436 );
not ( n76791 , n423207 );
buf ( n423209 , n393544 );
not ( n76793 , n423209 );
or ( n76794 , n76791 , n76793 );
buf ( n423212 , n400033 );
not ( n76796 , n423212 );
buf ( n423214 , n388965 );
not ( n76798 , n423214 );
or ( n76799 , n76796 , n76798 );
buf ( n423217 , n385473 );
buf ( n423218 , n400042 );
nand ( n76802 , n423217 , n423218 );
buf ( n423220 , n76802 );
buf ( n423221 , n423220 );
nand ( n76805 , n76799 , n423221 );
buf ( n423223 , n76805 );
buf ( n423224 , n423223 );
buf ( n423225 , n41447 );
nand ( n76809 , n423224 , n423225 );
buf ( n423227 , n76809 );
buf ( n423228 , n423227 );
nand ( n76812 , n76794 , n423228 );
buf ( n423230 , n76812 );
buf ( n423231 , n423230 );
buf ( n423232 , n421335 );
buf ( n423233 , n74737 );
or ( n76817 , n423232 , n423233 );
buf ( n423235 , n421351 );
nand ( n76819 , n76817 , n423235 );
buf ( n423237 , n76819 );
buf ( n423238 , n423237 );
buf ( n423239 , n421335 );
buf ( n423240 , n74737 );
nand ( n76824 , n423239 , n423240 );
buf ( n423242 , n76824 );
buf ( n423243 , n423242 );
nand ( n76827 , n423238 , n423243 );
buf ( n423245 , n76827 );
buf ( n423246 , n423245 );
buf ( n423247 , n390362 );
not ( n76831 , n423247 );
buf ( n423249 , n40601 );
not ( n76833 , n423249 );
buf ( n423251 , n406824 );
not ( n76835 , n423251 );
or ( n76836 , n76833 , n76835 );
buf ( n423254 , n406821 );
buf ( n423255 , n40600 );
nand ( n76839 , n423254 , n423255 );
buf ( n423257 , n76839 );
buf ( n423258 , n423257 );
nand ( n76842 , n76836 , n423258 );
buf ( n423260 , n76842 );
buf ( n423261 , n423260 );
not ( n76845 , n423261 );
or ( n76846 , n76831 , n76845 );
buf ( n423264 , n421342 );
not ( n76848 , n423264 );
buf ( n423266 , n40592 );
nand ( n76850 , n76848 , n423266 );
buf ( n423268 , n76850 );
buf ( n423269 , n423268 );
nand ( n76853 , n76846 , n423269 );
buf ( n423271 , n76853 );
buf ( n423272 , n423271 );
buf ( n423273 , n421328 );
not ( n76857 , n423273 );
buf ( n423275 , n60872 );
not ( n76859 , n423275 );
or ( n76860 , n76857 , n76859 );
buf ( n423278 , n392611 );
buf ( n423279 , n407936 );
and ( n76863 , n423278 , n423279 );
not ( n76864 , n423278 );
buf ( n423282 , n40653 );
and ( n76866 , n76864 , n423282 );
nor ( n76867 , n76863 , n76866 );
buf ( n423285 , n76867 );
buf ( n423286 , n423285 );
buf ( n423287 , n409076 );
nand ( n76871 , n423286 , n423287 );
buf ( n423289 , n76871 );
buf ( n423290 , n423289 );
nand ( n76874 , n76860 , n423290 );
buf ( n423292 , n76874 );
buf ( n423293 , n423292 );
xor ( n76877 , n423272 , n423293 );
xor ( n76878 , n421173 , n421217 );
and ( n76879 , n76878 , n421243 );
and ( n76880 , n421173 , n421217 );
or ( n76881 , n76879 , n76880 );
buf ( n423299 , n76881 );
buf ( n423300 , n423299 );
xor ( n76884 , n76877 , n423300 );
buf ( n423302 , n76884 );
buf ( n423303 , n423302 );
xor ( n76887 , n423246 , n423303 );
xor ( n76888 , n421144 , n421246 );
and ( n76889 , n76888 , n421268 );
and ( n76890 , n421144 , n421246 );
or ( n76891 , n76889 , n76890 );
buf ( n423309 , n76891 );
buf ( n423310 , n423309 );
xor ( n76894 , n76887 , n423310 );
buf ( n423312 , n76894 );
buf ( n423313 , n423312 );
xor ( n76897 , n423231 , n423313 );
buf ( n423315 , n419433 );
buf ( n423316 , n50580 );
or ( n76900 , n423315 , n423316 );
buf ( n423318 , n72794 );
buf ( n423319 , n40778 );
and ( n76903 , n423318 , n423319 );
not ( n76904 , n423318 );
buf ( n423322 , n40759 );
and ( n76906 , n76904 , n423322 );
nor ( n76907 , n76903 , n76906 );
buf ( n423325 , n76907 );
buf ( n423326 , n423325 );
buf ( n423327 , n50564 );
or ( n76911 , n423326 , n423327 );
nand ( n76912 , n76900 , n76911 );
buf ( n423330 , n76912 );
buf ( n423331 , n423330 );
xor ( n76915 , n76897 , n423331 );
buf ( n423333 , n76915 );
buf ( n423334 , n423333 );
and ( n76920 , n419725 , n419799 );
or ( n76921 , C0 , n76920 );
buf ( n423337 , n76921 );
buf ( n423338 , n423337 );
xor ( n76924 , n423334 , n423338 );
not ( n76925 , n73119 );
not ( n76926 , n73156 );
or ( n76927 , n76925 , n76926 );
nand ( n76928 , n76927 , n73166 );
not ( n76929 , n73156 );
nand ( n76930 , n76929 , n419749 );
nand ( n76931 , n76928 , n76930 );
buf ( n423347 , n76931 );
not ( n76933 , n423347 );
buf ( n423349 , n76933 );
and ( n76935 , n358975 , n393100 );
not ( n76936 , n421305 );
not ( n76937 , n74756 );
and ( n76938 , n76936 , n76937 );
buf ( n423354 , n421305 );
buf ( n423355 , n74756 );
nand ( n76941 , n423354 , n423355 );
buf ( n423357 , n76941 );
and ( n76943 , n423357 , n421310 );
nor ( n76944 , n76938 , n76943 );
xor ( n76945 , n76935 , n76944 );
buf ( n423361 , n419767 );
buf ( n423362 , n45949 );
and ( n76948 , n423361 , n423362 );
buf ( n423364 , n393369 );
not ( n76950 , n423364 );
buf ( n423366 , n388367 );
not ( n76952 , n423366 );
or ( n76953 , n76950 , n76952 );
buf ( n423369 , n397069 );
buf ( n423370 , n393381 );
nand ( n76956 , n423369 , n423370 );
buf ( n423372 , n76956 );
buf ( n423373 , n423372 );
nand ( n76959 , n76953 , n423373 );
buf ( n423375 , n76959 );
buf ( n423376 , n423375 );
buf ( n423377 , n45954 );
and ( n76963 , n423376 , n423377 );
nor ( n76964 , n76948 , n76963 );
buf ( n423380 , n76964 );
buf ( n76966 , n423380 );
xnor ( n76967 , n76945 , n76966 );
xor ( n76968 , n423349 , n76967 );
xor ( n76969 , n421271 , n421277 );
and ( n76970 , n76969 , n421365 );
and ( n76971 , n421271 , n421277 );
or ( n76972 , n76970 , n76971 );
buf ( n423388 , n76972 );
xor ( n76974 , n76968 , n423388 );
buf ( n423390 , n76974 );
xor ( n76976 , n76924 , n423390 );
buf ( n423392 , n76976 );
buf ( n423393 , n423392 );
xor ( n76979 , n76789 , n423393 );
buf ( n423395 , n76979 );
buf ( n423396 , n423395 );
xor ( n76982 , n76765 , n423396 );
buf ( n423398 , n76982 );
buf ( n423399 , n423398 );
xor ( n76985 , n422907 , n423399 );
buf ( n423401 , n402819 );
buf ( n423402 , n45391 );
and ( n76988 , n423401 , n423402 );
not ( n76989 , n423401 );
buf ( n423405 , n24050 );
and ( n76991 , n76989 , n423405 );
nor ( n423407 , n76988 , n76991 );
buf ( n423408 , n423407 );
buf ( n423409 , n423408 );
not ( n76995 , n423409 );
buf ( n423411 , n389122 );
not ( n76997 , n423411 );
or ( n76998 , n76995 , n76997 );
buf ( n423414 , n421813 );
buf ( n423415 , n41565 );
nand ( n77001 , n423414 , n423415 );
buf ( n423417 , n77001 );
buf ( n423418 , n423417 );
nand ( n77004 , n76998 , n423418 );
buf ( n423420 , n77004 );
buf ( n423421 , n423420 );
buf ( n423422 , C0 );
buf ( n423423 , n423422 );
xor ( n77035 , n423421 , n423423 );
xor ( n77036 , n421852 , n421856 );
xor ( n77037 , n77036 , n421885 );
buf ( n423427 , n77037 );
buf ( n423428 , n423427 );
and ( n77040 , n77035 , n423428 );
or ( n77042 , n77040 , C0 );
buf ( n423431 , n77042 );
buf ( n423432 , n423431 );
xor ( n77045 , n421827 , n421890 );
xor ( n77046 , n77045 , n421910 );
buf ( n423435 , n77046 );
buf ( n423436 , n423435 );
and ( n77049 , n423432 , n423436 );
not ( n77050 , n423432 );
buf ( n423439 , n423435 );
not ( n77052 , n423439 );
buf ( n423441 , n77052 );
buf ( n423442 , n423441 );
and ( n77055 , n77050 , n423442 );
nor ( n77056 , n77049 , n77055 );
buf ( n423445 , n77056 );
buf ( n423446 , n423445 );
buf ( n423447 , n59916 );
not ( n423448 , n423447 );
buf ( n423449 , n422788 );
not ( n77062 , n423449 );
or ( n77063 , n423448 , n77062 );
and ( n77064 , n47891 , n394663 );
not ( n77065 , n47891 );
and ( n77066 , n77065 , n27258 );
or ( n77067 , n77064 , n77066 );
buf ( n423456 , n77067 );
buf ( n423457 , n50579 );
nand ( n77070 , n423456 , n423457 );
buf ( n423459 , n77070 );
buf ( n423460 , n423459 );
nand ( n77073 , n77063 , n423460 );
buf ( n423462 , n77073 );
not ( n77075 , n423462 );
xor ( n77076 , n421975 , n422009 );
xor ( n77077 , n77076 , n422000 );
not ( n77078 , n77077 );
or ( n77079 , n77075 , n77078 );
buf ( n423468 , n77077 );
buf ( n423469 , n423462 );
or ( n77082 , n423468 , n423469 );
buf ( n423471 , n47411 );
buf ( n423472 , n388192 );
not ( n77085 , n423472 );
buf ( n423474 , n390389 );
nand ( n77087 , n77085 , n423474 );
buf ( n423476 , n77087 );
buf ( n423477 , n423476 );
buf ( n423478 , n358975 );
and ( n77091 , n423477 , n423478 );
buf ( n423480 , n407936 );
buf ( n423481 , n371522 );
and ( n77094 , n423480 , n423481 );
nor ( n77095 , n77091 , n77094 );
buf ( n423484 , n77095 );
buf ( n423485 , n423484 );
nand ( n77098 , n423471 , n423485 );
buf ( n423487 , n77098 );
buf ( n423488 , n423487 );
not ( n77101 , n423488 );
buf ( n77102 , n63906 );
buf ( n423491 , n77102 );
not ( n77104 , n423491 );
buf ( n423493 , n400042 );
buf ( n423494 , n407928 );
and ( n77107 , n423493 , n423494 );
not ( n77108 , n423493 );
buf ( n423497 , n404601 );
and ( n77110 , n77108 , n423497 );
nor ( n77111 , n77107 , n77110 );
buf ( n423500 , n77111 );
buf ( n423501 , n423500 );
not ( n77114 , n423501 );
and ( n77115 , n77104 , n77114 );
buf ( n423504 , n421985 );
buf ( n423505 , n40640 );
nor ( n77118 , n423504 , n423505 );
buf ( n423507 , n77118 );
buf ( n423508 , n423507 );
nor ( n77121 , n77115 , n423508 );
buf ( n423510 , n77121 );
buf ( n423511 , n423510 );
not ( n77124 , n423511 );
or ( n77125 , n77101 , n77124 );
buf ( n423514 , n45954 );
not ( n77127 , n423514 );
buf ( n423516 , n422063 );
not ( n77129 , n423516 );
or ( n77130 , n77127 , n77129 );
and ( n77131 , n27320 , n393381 );
not ( n77132 , n27320 );
and ( n77133 , n77132 , n393369 );
or ( n77134 , n77131 , n77133 );
buf ( n423523 , n77134 );
buf ( n423524 , n45949 );
nand ( n77137 , n423523 , n423524 );
buf ( n423526 , n77137 );
buf ( n423527 , n423526 );
nand ( n77140 , n77130 , n423527 );
buf ( n423529 , n77140 );
buf ( n423530 , n423529 );
xor ( n77143 , n422664 , n422685 );
xor ( n77144 , n77143 , n422752 );
buf ( n423533 , n77144 );
buf ( n423534 , n423533 );
xor ( n77147 , n423530 , n423534 );
xor ( n77148 , n420735 , n420875 );
xor ( n77149 , n77148 , n74273 );
xor ( n77150 , n75995 , n76154 );
xor ( n77151 , n77149 , n77150 );
buf ( n423540 , n77151 );
buf ( n423541 , n392884 );
not ( n77154 , n423541 );
buf ( n423543 , n391021 );
not ( n77156 , n423543 );
or ( n77157 , n77154 , n77156 );
buf ( n423546 , n388064 );
buf ( n423547 , n392881 );
nand ( n77160 , n423546 , n423547 );
buf ( n423549 , n77160 );
buf ( n423550 , n423549 );
nand ( n77163 , n77157 , n423550 );
buf ( n423552 , n77163 );
buf ( n423553 , n423552 );
not ( n77166 , n423553 );
buf ( n423555 , n74375 );
not ( n77168 , n423555 );
or ( n77169 , n77166 , n77168 );
buf ( n423558 , n422208 );
buf ( n423559 , n43515 );
nand ( n77172 , n423558 , n423559 );
buf ( n423561 , n77172 );
buf ( n423562 , n423561 );
nand ( n77175 , n77169 , n423562 );
buf ( n423564 , n77175 );
buf ( n423565 , n423564 );
xor ( n423566 , n423540 , n423565 );
buf ( n423567 , n417572 );
not ( n77180 , n423567 );
buf ( n423569 , n388722 );
not ( n77182 , n423569 );
buf ( n423571 , n77182 );
buf ( n423572 , n423571 );
not ( n77185 , n423572 );
or ( n77186 , n77180 , n77185 );
buf ( n423575 , n421024 );
not ( n77188 , n423575 );
buf ( n423577 , n394814 );
nand ( n77190 , n77188 , n423577 );
buf ( n423579 , n77190 );
buf ( n423580 , n423579 );
nand ( n77193 , n77186 , n423580 );
buf ( n423582 , n77193 );
buf ( n423583 , n423582 );
not ( n77196 , n423583 );
buf ( n423585 , n67042 );
not ( n77198 , n423585 );
or ( n77199 , n77196 , n77198 );
buf ( n423588 , n422698 );
buf ( n423589 , n388068 );
nand ( n77202 , n423588 , n423589 );
buf ( n423591 , n77202 );
buf ( n423592 , n423591 );
nand ( n77205 , n77199 , n423592 );
buf ( n423594 , n77205 );
buf ( n423595 , n423594 );
and ( n77208 , n423566 , n423595 );
and ( n77209 , n423540 , n423565 );
or ( n77210 , n77208 , n77209 );
buf ( n423599 , n77210 );
buf ( n423600 , n423599 );
and ( n77213 , n49117 , n388751 );
not ( n77214 , n49117 );
and ( n77215 , n77214 , n371784 );
or ( n77216 , n77213 , n77215 );
buf ( n423605 , n77216 );
not ( n77218 , n423605 );
buf ( n423607 , n388740 );
not ( n77220 , n423607 );
or ( n77221 , n77218 , n77220 );
buf ( n423610 , n422122 );
buf ( n423611 , n388803 );
nand ( n77224 , n423610 , n423611 );
buf ( n423613 , n77224 );
buf ( n423614 , n423613 );
nand ( n77227 , n77221 , n423614 );
buf ( n423616 , n77227 );
buf ( n423617 , n423616 );
xor ( n77230 , n423600 , n423617 );
buf ( n423619 , n45954 );
not ( n77232 , n423619 );
buf ( n423621 , n77134 );
not ( n77234 , n423621 );
or ( n77235 , n77232 , n77234 );
buf ( n423624 , n393369 );
not ( n77237 , n423624 );
buf ( n423626 , n72076 );
not ( n77239 , n423626 );
or ( n77240 , n77237 , n77239 );
buf ( n423629 , n72639 );
buf ( n423630 , n393381 );
nand ( n77243 , n423629 , n423630 );
buf ( n423632 , n77243 );
buf ( n423633 , n423632 );
nand ( n77246 , n77240 , n423633 );
buf ( n423635 , n77246 );
buf ( n423636 , n423635 );
buf ( n423637 , n45949 );
nand ( n77250 , n423636 , n423637 );
buf ( n423639 , n77250 );
buf ( n423640 , n423639 );
nand ( n77253 , n77235 , n423640 );
buf ( n423642 , n77253 );
buf ( n423643 , n423642 );
and ( n77256 , n77230 , n423643 );
and ( n77257 , n423600 , n423617 );
or ( n77258 , n77256 , n77257 );
buf ( n423647 , n77258 );
buf ( n423648 , n423647 );
and ( n77261 , n77147 , n423648 );
and ( n77262 , n423530 , n423534 );
or ( n77263 , n77261 , n77262 );
buf ( n423652 , n77263 );
buf ( n423653 , n423652 );
nand ( n77266 , n77125 , n423653 );
buf ( n423655 , n77266 );
buf ( n423656 , n423655 );
buf ( n423657 , n423487 );
not ( n77270 , n423657 );
buf ( n423659 , n77270 );
buf ( n423660 , n423659 );
buf ( n423661 , n423510 );
not ( n77274 , n423661 );
buf ( n423663 , n77274 );
buf ( n423664 , n423663 );
nand ( n77277 , n423660 , n423664 );
buf ( n423666 , n77277 );
buf ( n423667 , n423666 );
nand ( n77280 , n423656 , n423667 );
buf ( n423669 , n77280 );
buf ( n423670 , n423669 );
nand ( n77283 , n77082 , n423670 );
buf ( n423672 , n77283 );
nand ( n77285 , n77079 , n423672 );
not ( n77286 , n77285 );
not ( n77287 , n77286 );
or ( n77297 , n77287 , C0 );
buf ( n423677 , n76257 );
not ( n77299 , n423677 );
buf ( n423679 , n422108 );
not ( n77301 , n423679 );
or ( n77302 , n77299 , n77301 );
buf ( n423682 , n422108 );
buf ( n423683 , n76257 );
or ( n77305 , n423682 , n423683 );
nand ( n77306 , n77302 , n77305 );
buf ( n423686 , n77306 );
buf ( n423687 , n423686 );
not ( n77309 , n423687 );
buf ( n423689 , n422083 );
not ( n77311 , n423689 );
and ( n77312 , n77309 , n77311 );
buf ( n423692 , n423686 );
buf ( n423693 , n422083 );
and ( n77315 , n423692 , n423693 );
nor ( n77316 , n77312 , n77315 );
buf ( n423696 , n77316 );
buf ( n423697 , n423696 );
not ( n77319 , n423697 );
buf ( n423699 , n77319 );
buf ( n423700 , C0 );
buf ( n423701 , n423700 );
buf ( n423702 , n423699 );
or ( n77352 , n423701 , n423702 );
buf ( n423704 , n422177 );
not ( n77354 , n423704 );
buf ( n423706 , n422756 );
not ( n77356 , n423706 );
buf ( n423708 , n422187 );
not ( n77358 , n423708 );
and ( n77359 , n77356 , n77358 );
buf ( n423711 , n422187 );
buf ( n423712 , n422756 );
and ( n77362 , n423711 , n423712 );
nor ( n77363 , n77359 , n77362 );
buf ( n423715 , n77363 );
buf ( n423716 , n423715 );
not ( n77366 , n423716 );
or ( n77367 , n77354 , n77366 );
buf ( n423719 , n422177 );
buf ( n423720 , n423715 );
or ( n77370 , n423719 , n423720 );
nand ( n77371 , n77367 , n77370 );
buf ( n423723 , n77371 );
buf ( n423724 , n423723 );
buf ( n423725 , n395359 );
not ( n77375 , n423725 );
buf ( n423727 , n422101 );
not ( n77377 , n423727 );
or ( n77378 , n77375 , n77377 );
buf ( n423730 , n47863 );
not ( n77380 , n423730 );
buf ( n423732 , n406824 );
not ( n77382 , n423732 );
or ( n77383 , n77380 , n77382 );
buf ( n423735 , n406821 );
buf ( n423736 , n421871 );
nand ( n77386 , n423735 , n423736 );
buf ( n423738 , n77386 );
buf ( n423739 , n423738 );
nand ( n77389 , n77383 , n423739 );
buf ( n423741 , n77389 );
buf ( n423742 , n423741 );
buf ( n423743 , n395346 );
nand ( n77393 , n423742 , n423743 );
buf ( n423745 , n77393 );
buf ( n423746 , n423745 );
nand ( n77396 , n77378 , n423746 );
buf ( n423748 , n77396 );
buf ( n423749 , n423748 );
xor ( n77399 , n423724 , n423749 );
buf ( n423751 , n422155 );
not ( n77401 , n423751 );
buf ( n423753 , n75662 );
not ( n77403 , n423753 );
buf ( n423755 , n422134 );
not ( n77405 , n423755 );
and ( n77406 , n77403 , n77405 );
buf ( n423758 , n75662 );
buf ( n423759 , n422134 );
and ( n77409 , n423758 , n423759 );
nor ( n423761 , n77406 , n77409 );
buf ( n423762 , n423761 );
buf ( n423763 , n423762 );
not ( n77413 , n423763 );
and ( n77414 , n77401 , n77413 );
buf ( n423766 , n422155 );
buf ( n423767 , n423762 );
and ( n77417 , n423766 , n423767 );
nor ( n77418 , n77414 , n77417 );
buf ( n423770 , n77418 );
buf ( n423771 , n423770 );
not ( n423772 , n423771 );
buf ( n423773 , n423772 );
buf ( n423774 , n423773 );
not ( n77424 , n423774 );
buf ( n423776 , n399274 );
not ( n423777 , n423776 );
buf ( n423778 , n66132 );
not ( n77428 , n423778 );
or ( n77429 , n423777 , n77428 );
buf ( n423781 , n67832 );
buf ( n423782 , n399283 );
nand ( n77432 , n423781 , n423782 );
buf ( n423784 , n77432 );
buf ( n423785 , n423784 );
nand ( n423786 , n77429 , n423785 );
buf ( n423787 , n423786 );
buf ( n423788 , n423787 );
not ( n77438 , n423788 );
buf ( n423790 , n66128 );
not ( n423791 , n423790 );
or ( n423792 , n77438 , n423791 );
buf ( n423793 , n41332 );
not ( n77443 , n423793 );
buf ( n423795 , n422033 );
nand ( n423796 , n77443 , n423795 );
buf ( n423797 , n423796 );
buf ( n423798 , n423797 );
nand ( n77448 , n423792 , n423798 );
buf ( n423800 , n77448 );
buf ( n423801 , n423800 );
not ( n423802 , n423801 );
or ( n77452 , n77424 , n423802 );
buf ( n423804 , n423800 );
buf ( n423805 , n423773 );
or ( n423806 , n423804 , n423805 );
xor ( n423807 , n422711 , n422721 );
xor ( n77457 , n423807 , n422747 );
buf ( n423809 , n77457 );
buf ( n423810 , n423809 );
buf ( n423811 , n413643 );
not ( n423812 , n423811 );
buf ( n423813 , n422739 );
not ( n77463 , n423813 );
or ( n77464 , n423812 , n77463 );
buf ( n423816 , n44775 );
not ( n423817 , n423816 );
buf ( n423818 , n391440 );
not ( n77468 , n423818 );
or ( n77469 , n423817 , n77468 );
buf ( n423821 , n420994 );
buf ( n423822 , n44776 );
nand ( n77472 , n423821 , n423822 );
buf ( n423824 , n77472 );
buf ( n423825 , n423824 );
nand ( n423826 , n77469 , n423825 );
buf ( n423827 , n423826 );
buf ( n423828 , n423827 );
buf ( n423829 , n417542 );
nand ( n77479 , n423828 , n423829 );
buf ( n423831 , n77479 );
buf ( n423832 , n423831 );
nand ( n77482 , n77464 , n423832 );
buf ( n423834 , n77482 );
buf ( n423835 , n423834 );
not ( n423836 , n423835 );
buf ( n423837 , n413643 );
not ( n77487 , n423837 );
buf ( n423839 , n423827 );
not ( n77489 , n423839 );
or ( n423841 , n77487 , n77489 );
buf ( n423842 , n44775 );
not ( n77492 , n423842 );
buf ( n423844 , n420908 );
not ( n77494 , n423844 );
or ( n423846 , n77492 , n77494 );
buf ( n423847 , n420911 );
buf ( n423848 , n44776 );
nand ( n77498 , n423847 , n423848 );
buf ( n423850 , n77498 );
buf ( n423851 , n423850 );
nand ( n423852 , n423846 , n423851 );
buf ( n423853 , n423852 );
buf ( n423854 , n423853 );
buf ( n423855 , n417542 );
nand ( n423856 , n423854 , n423855 );
buf ( n423857 , n423856 );
buf ( n423858 , n423857 );
nand ( n77508 , n423841 , n423858 );
buf ( n423860 , n77508 );
buf ( n423861 , n423860 );
xor ( n423862 , n422220 , n75764 );
xor ( n77512 , n423862 , n422493 );
xor ( n77513 , n422502 , n76149 );
xor ( n77514 , n77512 , n77513 );
buf ( n423866 , n77514 );
or ( n423867 , n423861 , n423866 );
buf ( n423868 , n66270 );
buf ( n423869 , n63625 );
and ( n77519 , n423868 , n423869 );
buf ( n423871 , n413098 );
buf ( n423872 , n63629 );
and ( n77522 , n423871 , n423872 );
nor ( n77523 , n77519 , n77522 );
buf ( n423875 , n77523 );
buf ( n423876 , n423875 );
buf ( n423877 , n410635 );
or ( n77527 , n423876 , n423877 );
buf ( n423879 , n422296 );
buf ( n423880 , n409504 );
or ( n423881 , n423879 , n423880 );
nand ( n423882 , n77527 , n423881 );
buf ( n423883 , n423882 );
xor ( n77533 , n422450 , n422453 );
xor ( n77534 , n77533 , n422475 );
and ( n423886 , n423883 , n77534 );
xor ( n423887 , n422403 , n422420 );
xor ( n77537 , n423887 , n422446 );
buf ( n423889 , n77537 );
buf ( n423890 , n70210 );
buf ( n423891 , n59628 );
and ( n423892 , n423890 , n423891 );
buf ( n423893 , n416845 );
buf ( n423894 , n59457 );
and ( n77544 , n423893 , n423894 );
nor ( n423896 , n423892 , n77544 );
buf ( n423897 , n423896 );
buf ( n423898 , n423897 );
buf ( n423899 , n59637 );
or ( n77549 , n423898 , n423899 );
buf ( n423901 , n422470 );
buf ( n423902 , n59467 );
or ( n77552 , n423901 , n423902 );
nand ( n77553 , n77549 , n77552 );
buf ( n423905 , n77553 );
xor ( n423906 , n423889 , n423905 );
buf ( n423907 , n409185 );
not ( n77557 , n423907 );
buf ( n423909 , n422619 );
not ( n77559 , n423909 );
or ( n423911 , n77557 , n77559 );
buf ( n423912 , n414729 );
buf ( n423913 , n409178 );
or ( n77563 , n423912 , n423913 );
buf ( n423915 , n68002 );
buf ( n423916 , n59463 );
or ( n423917 , n423915 , n423916 );
nand ( n77567 , n77563 , n423917 );
buf ( n423919 , n77567 );
buf ( n423920 , n423919 );
not ( n423921 , n423920 );
buf ( n423922 , n423921 );
buf ( n423923 , n423922 );
buf ( n423924 , n409429 );
or ( n77574 , n423923 , n423924 );
nand ( n423926 , n423911 , n77574 );
buf ( n423927 , n423926 );
and ( n77577 , n423906 , n423927 );
and ( n77578 , n423889 , n423905 );
or ( n77579 , n77577 , n77578 );
xor ( n423931 , n422450 , n422453 );
xor ( n423932 , n423931 , n422475 );
and ( n77582 , n77579 , n423932 );
and ( n77583 , n423883 , n77579 );
or ( n77584 , n423886 , n77582 , n77583 );
xor ( n423936 , n422269 , n422285 );
xor ( n423937 , n423936 , n422307 );
and ( n77587 , n77584 , n423937 );
xor ( n77588 , n422550 , n422553 );
xor ( n77589 , n77588 , n422603 );
buf ( n423941 , n77589 );
buf ( n423942 , n405407 );
buf ( n423943 , n403283 );
buf ( n423944 , n71170 );
and ( n77594 , n423943 , n423944 );
buf ( n423946 , n56050 );
buf ( n423947 , n417804 );
and ( n77597 , n423946 , n423947 );
nor ( n77598 , n77594 , n77597 );
buf ( n423950 , n77598 );
buf ( n423951 , n423950 );
or ( n423952 , n423942 , n423951 );
buf ( n423953 , n422593 );
buf ( n423954 , n405378 );
or ( n77604 , n423953 , n423954 );
nand ( n423956 , n423952 , n77604 );
buf ( n423957 , n423956 );
buf ( n423958 , n54346 );
buf ( n423959 , n623 );
and ( n77609 , n423958 , n423959 );
buf ( n423961 , n54346 );
not ( n423962 , n423961 );
buf ( n423963 , n423962 );
buf ( n423964 , n423963 );
buf ( n423965 , n422315 );
and ( n423966 , n423964 , n423965 );
buf ( n423967 , n15287 );
nor ( n77617 , n423966 , n423967 );
buf ( n423969 , n77617 );
buf ( n423970 , n423969 );
buf ( n423971 , n401612 );
nor ( n423972 , n77609 , n423970 , n423971 );
buf ( n423973 , n423972 );
xor ( n77623 , n423957 , n423973 );
buf ( n423975 , n403293 );
buf ( n423976 , n56041 );
buf ( n423977 , n71681 );
and ( n77627 , n423976 , n423977 );
buf ( n423979 , n403298 );
buf ( n423980 , n418315 );
and ( n423981 , n423979 , n423980 );
nor ( n423982 , n77627 , n423981 );
buf ( n423983 , n423982 );
buf ( n423984 , n423983 );
or ( n77634 , n423975 , n423984 );
buf ( n423986 , n422435 );
buf ( n423987 , n405476 );
or ( n77637 , n423986 , n423987 );
nand ( n77638 , n77634 , n77637 );
buf ( n423990 , n77638 );
and ( n423991 , n77623 , n423990 );
and ( n423992 , n423957 , n423973 );
or ( n77642 , n423991 , n423992 );
buf ( n423994 , n77642 );
xor ( n77644 , n422426 , n422443 );
buf ( n423996 , n77644 );
buf ( n423997 , n423996 );
xor ( n77647 , n423994 , n423997 );
buf ( n423999 , n59468 );
not ( n77649 , n423999 );
buf ( n424001 , n70389 );
buf ( n424002 , n14083 );
and ( n77652 , n424001 , n424002 );
buf ( n424004 , n417024 );
buf ( n424005 , n59457 );
and ( n424006 , n424004 , n424005 );
nor ( n424007 , n77652 , n424006 );
buf ( n424008 , n424007 );
buf ( n424009 , n424008 );
not ( n77659 , n424009 );
buf ( n424011 , n77659 );
buf ( n424012 , n424011 );
not ( n77662 , n424012 );
or ( n77663 , n77649 , n77662 );
buf ( n424015 , n423897 );
buf ( n424016 , n59467 );
or ( n424017 , n424015 , n424016 );
nand ( n77667 , n77663 , n424017 );
buf ( n424019 , n77667 );
buf ( n424020 , n424019 );
and ( n424021 , n77647 , n424020 );
and ( n424022 , n423994 , n423997 );
or ( n77672 , n424021 , n424022 );
buf ( n424024 , n77672 );
xor ( n77674 , n423941 , n424024 );
buf ( n424026 , n409516 );
not ( n424027 , n424026 );
buf ( n424028 , n423875 );
not ( n77678 , n424028 );
buf ( n424030 , n77678 );
buf ( n424031 , n424030 );
not ( n424032 , n424031 );
or ( n77682 , n424027 , n424032 );
buf ( n424034 , n66359 );
buf ( n424035 , n63625 );
and ( n424036 , n424034 , n424035 );
buf ( n424037 , n413187 );
buf ( n424038 , n63629 );
and ( n77688 , n424037 , n424038 );
nor ( n77689 , n424036 , n77688 );
buf ( n424041 , n77689 );
buf ( n424042 , n424041 );
buf ( n424043 , n410635 );
or ( n77693 , n424042 , n424043 );
nand ( n77694 , n77682 , n77693 );
buf ( n424046 , n77694 );
and ( n424047 , n77674 , n424046 );
and ( n77697 , n423941 , n424024 );
or ( n77698 , n424047 , n77697 );
buf ( n424050 , n77698 );
buf ( n424051 , n63564 );
buf ( n424052 , n66411 );
and ( n77702 , n424051 , n424052 );
buf ( n424054 , n413073 );
buf ( n424055 , n62496 );
and ( n424056 , n424054 , n424055 );
nor ( n424057 , n77702 , n424056 );
buf ( n424058 , n424057 );
buf ( n424059 , n424058 );
buf ( n424060 , n410724 );
or ( n424061 , n424059 , n424060 );
buf ( n424062 , n422517 );
buf ( n424063 , n410721 );
or ( n77713 , n424062 , n424063 );
nand ( n77714 , n424061 , n77713 );
buf ( n424066 , n77714 );
buf ( n424067 , n424066 );
xor ( n77717 , n424050 , n424067 );
xor ( n77718 , n422530 , n422608 );
xor ( n77719 , n77718 , n422628 );
buf ( n424071 , n77719 );
buf ( n424072 , n424071 );
and ( n77722 , n77717 , n424072 );
and ( n77723 , n424050 , n424067 );
or ( n77724 , n77722 , n77723 );
buf ( n424076 , n77724 );
xor ( n424077 , n422269 , n422285 );
xor ( n77727 , n424077 , n422307 );
and ( n77728 , n424076 , n77727 );
and ( n77729 , n77584 , n424076 );
or ( n424081 , n77587 , n77728 , n77729 );
xor ( n424082 , n76008 , n422643 );
xor ( n77732 , n424082 , n422647 );
and ( n77733 , n424081 , n77732 );
xor ( n77734 , n422450 , n422453 );
xor ( n424086 , n77734 , n422475 );
xor ( n424087 , n423883 , n77579 );
xor ( n77737 , n424086 , n424087 );
buf ( n424089 , n401681 );
buf ( n424090 , n623 );
or ( n424091 , n424089 , n424090 );
buf ( n424092 , n401674 );
buf ( n424093 , n418921 );
buf ( n424094 , n623 );
and ( n77744 , n424092 , n424093 , n424094 );
buf ( n424096 , n401664 );
nor ( n424097 , n77744 , n424096 );
buf ( n424098 , n424097 );
buf ( n424099 , n424098 );
nand ( n77749 , n424091 , n424099 );
buf ( n424101 , n77749 );
buf ( n424102 , n403120 );
buf ( n424103 , n15287 );
buf ( n424104 , n74002 );
and ( n77754 , n424103 , n424104 );
buf ( n424106 , n15290 );
buf ( n424107 , n420612 );
and ( n77757 , n424106 , n424107 );
nor ( n77758 , n77754 , n77757 );
buf ( n424110 , n77758 );
buf ( n424111 , n424110 );
or ( n424112 , n424102 , n424111 );
buf ( n424113 , n422570 );
buf ( n424114 , n403108 );
or ( n77764 , n424113 , n424114 );
nand ( n424116 , n424112 , n77764 );
buf ( n424117 , n424116 );
xor ( n77767 , n424101 , n424117 );
buf ( n424119 , n401660 );
buf ( n424120 , n422315 );
nor ( n424121 , n424119 , n424120 );
buf ( n424122 , n424121 );
buf ( n424123 , n424122 );
buf ( n424124 , n405388 );
buf ( n424125 , n418298 );
or ( n424126 , n424124 , n424125 );
buf ( n424127 , n403283 );
buf ( n424128 , n71664 );
or ( n77778 , n424127 , n424128 );
nand ( n77779 , n424126 , n77778 );
buf ( n424131 , n77779 );
buf ( n424132 , n424131 );
not ( n77782 , n424132 );
buf ( n424134 , n405410 );
not ( n77784 , n424134 );
or ( n424136 , n77782 , n77784 );
buf ( n424137 , n423950 );
buf ( n424138 , n405378 );
or ( n77788 , n424137 , n424138 );
nand ( n77789 , n424136 , n77788 );
buf ( n424141 , n77789 );
buf ( n424142 , n424141 );
and ( n77792 , n424123 , n424142 );
buf ( n424144 , n77792 );
and ( n77794 , n77767 , n424144 );
and ( n424146 , n424101 , n424117 );
or ( n424147 , n77794 , n424146 );
xor ( n77797 , n422561 , n422578 );
xor ( n77798 , n77797 , n422598 );
buf ( n424150 , n77798 );
xor ( n424151 , n424147 , n424150 );
buf ( n424152 , n409185 );
not ( n77802 , n424152 );
buf ( n424154 , n423919 );
not ( n77804 , n424154 );
or ( n424156 , n77802 , n77804 );
buf ( n424157 , n70195 );
buf ( n424158 , n59463 );
and ( n77808 , n424157 , n424158 );
buf ( n424160 , n416830 );
buf ( n424161 , n62159 );
and ( n424162 , n424160 , n424161 );
nor ( n77812 , n77808 , n424162 );
buf ( n424164 , n77812 );
buf ( n424165 , n424164 );
buf ( n424166 , n409429 );
or ( n424167 , n424165 , n424166 );
nand ( n77817 , n424156 , n424167 );
buf ( n424169 , n77817 );
and ( n77819 , n424151 , n424169 );
and ( n424171 , n424147 , n424150 );
or ( n424172 , n77819 , n424171 );
xor ( n77822 , n423889 , n423905 );
xor ( n77823 , n77822 , n423927 );
and ( n77824 , n424172 , n77823 );
buf ( n424176 , n348158 );
not ( n424177 , n424176 );
buf ( n424178 , n424058 );
not ( n77828 , n424178 );
buf ( n424180 , n77828 );
buf ( n424181 , n424180 );
not ( n424182 , n424181 );
or ( n77832 , n424177 , n424182 );
buf ( n424184 , n63707 );
buf ( n424185 , n62499 );
and ( n424186 , n424184 , n424185 );
buf ( n424187 , n413104 );
buf ( n424188 , n410717 );
and ( n77838 , n424187 , n424188 );
nor ( n77839 , n424186 , n77838 );
buf ( n424191 , n77839 );
buf ( n424192 , n424191 );
buf ( n424193 , n410724 );
or ( n77843 , n424192 , n424193 );
nand ( n77844 , n77832 , n77843 );
buf ( n424196 , n77844 );
xor ( n424197 , n423889 , n423905 );
xor ( n77847 , n424197 , n423927 );
and ( n77848 , n424196 , n77847 );
and ( n77849 , n424172 , n424196 );
or ( n424201 , n77824 , n77848 , n77849 );
xor ( n424202 , n77737 , n424201 );
xor ( n77852 , n424050 , n424067 );
xor ( n77853 , n77852 , n424072 );
buf ( n424205 , n77853 );
and ( n424206 , n424202 , n424205 );
and ( n424207 , n77737 , n424201 );
or ( n77857 , n424206 , n424207 );
buf ( n424209 , n77857 );
xor ( n77859 , n422526 , n422633 );
xor ( n424211 , n77859 , n422639 );
buf ( n424212 , n424211 );
buf ( n424213 , n424212 );
xor ( n77863 , n424209 , n424213 );
xor ( n77864 , n422269 , n422285 );
xor ( n424216 , n77864 , n422307 );
xor ( n424217 , n77584 , n424076 );
xor ( n77867 , n424216 , n424217 );
buf ( n424219 , n77867 );
and ( n77869 , n77863 , n424219 );
and ( n424221 , n424209 , n424213 );
or ( n424222 , n77869 , n424221 );
buf ( n424223 , n424222 );
xor ( n77873 , n76008 , n422643 );
xor ( n77874 , n77873 , n422647 );
and ( n424226 , n424223 , n77874 );
and ( n424227 , n424081 , n424223 );
or ( n77877 , n77733 , n424226 , n424227 );
buf ( n424229 , n77877 );
nand ( n77879 , n423867 , n424229 );
buf ( n424231 , n77879 );
buf ( n424232 , n424231 );
buf ( n424233 , n423860 );
buf ( n424234 , n77514 );
nand ( n77884 , n424233 , n424234 );
buf ( n424236 , n77884 );
buf ( n424237 , n424236 );
and ( n77887 , n424232 , n424237 );
buf ( n424239 , n77887 );
buf ( n424240 , n424239 );
nand ( n424241 , n423836 , n424240 );
buf ( n424242 , n424241 );
buf ( n424243 , n424242 );
not ( n77893 , n424243 );
xor ( n77894 , n423540 , n423565 );
xor ( n424246 , n77894 , n423595 );
buf ( n424247 , n424246 );
buf ( n424248 , n424247 );
not ( n77898 , n424248 );
or ( n77899 , n77893 , n77898 );
buf ( n424251 , n424239 );
not ( n424252 , n424251 );
buf ( n424253 , n423834 );
nand ( n77903 , n424252 , n424253 );
buf ( n424255 , n77903 );
buf ( n424256 , n424255 );
nand ( n424257 , n77899 , n424256 );
buf ( n424258 , n424257 );
buf ( n424259 , n424258 );
xor ( n77909 , n423810 , n424259 );
buf ( n424261 , n55543 );
not ( n424262 , n424261 );
buf ( n424263 , n68376 );
not ( n77913 , n424263 );
or ( n77914 , n424262 , n77913 );
buf ( n424266 , n24116 );
buf ( n424267 , n51185 );
nand ( n77917 , n424266 , n424267 );
buf ( n424269 , n77917 );
buf ( n424270 , n424269 );
nand ( n424271 , n77914 , n424270 );
buf ( n424272 , n424271 );
buf ( n424273 , n424272 );
not ( n77923 , n424273 );
buf ( n424275 , n416762 );
not ( n424276 , n424275 );
or ( n424277 , n77923 , n424276 );
buf ( n424278 , n75642 );
buf ( n424279 , n41664 );
nand ( n77929 , n424278 , n424279 );
buf ( n424281 , n77929 );
buf ( n424282 , n424281 );
nand ( n77932 , n424277 , n424282 );
buf ( n424284 , n77932 );
buf ( n424285 , n424284 );
and ( n424286 , n77909 , n424285 );
and ( n424287 , n423810 , n424259 );
or ( n77937 , n424286 , n424287 );
buf ( n424289 , n77937 );
buf ( n424290 , n424289 );
nand ( n424291 , n423806 , n424290 );
buf ( n424292 , n424291 );
buf ( n424293 , n424292 );
nand ( n77943 , n77452 , n424293 );
buf ( n424295 , n77943 );
buf ( n424296 , n424295 );
and ( n424297 , n77399 , n424296 );
and ( n77947 , n423724 , n423749 );
or ( n77948 , n424297 , n77947 );
buf ( n424300 , n77948 );
buf ( n424301 , n424300 );
nand ( n424302 , n77352 , n424301 );
buf ( n424303 , n424302 );
buf ( n424304 , n424303 );
nand ( n77954 , C1 , n424304 );
buf ( n424306 , n77954 );
nand ( n424307 , n77297 , n424306 );
buf ( n424308 , n424307 );
buf ( n424309 , C1 );
nand ( n424310 , n424308 , n424309 );
buf ( n424311 , n424310 );
buf ( n424312 , n424311 );
not ( n77963 , n424312 );
buf ( n424314 , n77963 );
buf ( n424315 , n424314 );
and ( n424316 , n423446 , n424315 );
not ( n77967 , n423446 );
buf ( n424318 , n424311 );
and ( n77969 , n77967 , n424318 );
nor ( n424320 , n424316 , n77969 );
buf ( n424321 , n424320 );
buf ( n424322 , n424321 );
buf ( n424323 , n53251 );
not ( n77974 , n424323 );
buf ( n424325 , n358975 );
not ( n424326 , n424325 );
or ( n77977 , n77974 , n424326 );
buf ( n424328 , n47411 );
buf ( n424329 , n402819 );
nand ( n424330 , n424328 , n424329 );
buf ( n424331 , n424330 );
buf ( n424332 , n424331 );
nand ( n77983 , n77977 , n424332 );
buf ( n424334 , n77983 );
buf ( n424335 , n424334 );
not ( n424336 , n424335 );
buf ( n424337 , n52812 );
not ( n77988 , n424337 );
or ( n77989 , n424336 , n77988 );
buf ( n424340 , n422818 );
buf ( n424341 , n42924 );
nand ( n77992 , n424340 , n424341 );
buf ( n424343 , n77992 );
buf ( n424344 , n424343 );
nand ( n424345 , n77989 , n424344 );
buf ( n424346 , n424345 );
buf ( n424347 , n424346 );
not ( n77998 , n424347 );
buf ( n424349 , n59916 );
not ( n424350 , n424349 );
buf ( n424351 , n77067 );
not ( n78002 , n424351 );
or ( n78003 , n424350 , n78002 );
buf ( n424354 , n47891 );
not ( n424355 , n424354 );
buf ( n424356 , n403039 );
not ( n78007 , n424356 );
or ( n78008 , n424355 , n78007 );
buf ( n424359 , n28644 );
buf ( n424360 , n72794 );
nand ( n424361 , n424359 , n424360 );
buf ( n424362 , n424361 );
buf ( n424363 , n424362 );
nand ( n78014 , n78008 , n424363 );
buf ( n424365 , n78014 );
buf ( n424366 , n424365 );
buf ( n424367 , n50579 );
nand ( n78018 , n424366 , n424367 );
buf ( n424369 , n78018 );
buf ( n424370 , n424369 );
nand ( n424371 , n78003 , n424370 );
buf ( n424372 , n424371 );
buf ( n424373 , n424372 );
not ( n78024 , n424373 );
buf ( n424375 , n78024 );
buf ( n424376 , n424375 );
nand ( n78027 , n77998 , n424376 );
buf ( n424378 , n78027 );
xor ( n78029 , n422046 , n422071 );
xor ( n424380 , n78029 , n422076 );
buf ( n424381 , n424380 );
and ( n78032 , n424378 , n424381 );
and ( n78033 , n424372 , n424346 );
nor ( n78034 , n78032 , n78033 );
buf ( n424385 , n78034 );
buf ( n424386 , n422804 );
buf ( n424387 , n76371 );
xor ( n78038 , n424386 , n424387 );
buf ( n424389 , n422830 );
xor ( n424390 , n78038 , n424389 );
buf ( n424391 , n424390 );
buf ( n424392 , n424391 );
xor ( n78043 , n424385 , n424392 );
buf ( n424394 , C1 );
and ( n78059 , n78043 , n424394 );
and ( n78060 , n424385 , n424392 );
or ( n424397 , n78059 , n78060 );
buf ( n424398 , n424397 );
buf ( n424399 , n424398 );
not ( n78064 , n424399 );
not ( n78066 , n77286 );
and ( n78067 , n78066 , C1 );
nor ( n78068 , C0 , n78067 );
and ( n424404 , n78068 , n424306 );
not ( n78070 , n78068 );
not ( n78071 , n424306 );
and ( n78072 , n78070 , n78071 );
nor ( n78073 , n424404 , n78072 );
buf ( n424409 , n78073 );
not ( n78075 , n424409 );
or ( n78076 , n78064 , n78075 );
buf ( n424412 , n423669 );
buf ( n424413 , n423462 );
xor ( n78079 , n424412 , n424413 );
buf ( n424415 , n77077 );
xnor ( n78081 , n78079 , n424415 );
buf ( n424417 , n78081 );
not ( n78083 , n424417 );
buf ( n424419 , n397489 );
not ( n78085 , n424419 );
buf ( n424421 , n371787 );
not ( n78087 , n424421 );
or ( n78088 , n78085 , n78087 );
buf ( n424424 , n371784 );
buf ( n424425 , n397486 );
nand ( n78091 , n424424 , n424425 );
buf ( n424427 , n78091 );
buf ( n424428 , n424427 );
nand ( n78094 , n78088 , n424428 );
buf ( n424430 , n78094 );
buf ( n424431 , n424430 );
not ( n424432 , n424431 );
buf ( n424433 , n388740 );
not ( n78099 , n424433 );
or ( n78100 , n424432 , n78099 );
buf ( n424436 , n77216 );
buf ( n424437 , n388803 );
nand ( n78103 , n424436 , n424437 );
buf ( n424439 , n78103 );
buf ( n424440 , n424439 );
nand ( n78106 , n78100 , n424440 );
buf ( n424442 , n78106 );
buf ( n424443 , n424442 );
buf ( n424444 , n394210 );
buf ( n424445 , n391018 );
and ( n78111 , n424444 , n424445 );
not ( n78112 , n424444 );
buf ( n424448 , n420986 );
and ( n78114 , n78112 , n424448 );
nor ( n424450 , n78111 , n78114 );
buf ( n424451 , n424450 );
buf ( n424452 , n424451 );
not ( n78118 , n424452 );
buf ( n424454 , n43536 );
not ( n424455 , n424454 );
or ( n78121 , n78118 , n424455 );
buf ( n424457 , n423552 );
buf ( n424458 , n43515 );
nand ( n78124 , n424457 , n424458 );
buf ( n424460 , n78124 );
buf ( n424461 , n424460 );
nand ( n78127 , n78121 , n424461 );
buf ( n424463 , n78127 );
buf ( n424464 , n424463 );
buf ( n424465 , n71095 );
buf ( n424466 , n14083 );
and ( n78132 , n424465 , n424466 );
buf ( n424468 , n417729 );
buf ( n424469 , n59457 );
and ( n78135 , n424468 , n424469 );
nor ( n78136 , n78132 , n78135 );
buf ( n424472 , n78136 );
buf ( n424473 , n424472 );
buf ( n424474 , n59637 );
or ( n78140 , n424473 , n424474 );
buf ( n424476 , n424008 );
buf ( n424477 , n59467 );
or ( n78143 , n424476 , n424477 );
nand ( n78144 , n78140 , n78143 );
buf ( n424480 , n78144 );
xor ( n78146 , n423957 , n423973 );
xor ( n78147 , n78146 , n423990 );
and ( n78148 , n424480 , n78147 );
buf ( n424484 , n424110 );
buf ( n424485 , n403108 );
or ( n78151 , n424484 , n424485 );
buf ( n424487 , n403128 );
nand ( n78153 , n78151 , n424487 );
buf ( n424489 , n78153 );
buf ( n424490 , n424489 );
buf ( n424491 , n403293 );
buf ( n424492 , n56041 );
buf ( n424493 , n72308 );
and ( n78159 , n424492 , n424493 );
buf ( n424495 , n403298 );
buf ( n424496 , n418942 );
and ( n78162 , n424495 , n424496 );
nor ( n78163 , n78159 , n78162 );
buf ( n424499 , n78163 );
buf ( n424500 , n424499 );
or ( n424501 , n424491 , n424500 );
buf ( n424502 , n423983 );
buf ( n424503 , n403290 );
or ( n78169 , n424502 , n424503 );
nand ( n78170 , n424501 , n78169 );
buf ( n424506 , n78170 );
buf ( n424507 , n424506 );
xor ( n78173 , n424490 , n424507 );
buf ( n424509 , n71088 );
buf ( n424510 , n14083 );
and ( n78176 , n424509 , n424510 );
buf ( n424512 , n417722 );
buf ( n424513 , n59457 );
and ( n78179 , n424512 , n424513 );
nor ( n78180 , n78176 , n78179 );
buf ( n424516 , n78180 );
buf ( n424517 , n424516 );
not ( n78183 , n424517 );
buf ( n424519 , n78183 );
buf ( n424520 , n424519 );
not ( n78186 , n424520 );
buf ( n424522 , n59468 );
not ( n78188 , n424522 );
or ( n78189 , n78186 , n78188 );
buf ( n424525 , n424472 );
buf ( n424526 , n59467 );
or ( n78192 , n424525 , n424526 );
nand ( n78193 , n78189 , n78192 );
buf ( n424529 , n78193 );
buf ( n424530 , n424529 );
and ( n78196 , n78173 , n424530 );
and ( n78197 , n424490 , n424507 );
or ( n78198 , n78196 , n78197 );
buf ( n424534 , n78198 );
xor ( n78200 , n423957 , n423973 );
xor ( n78201 , n78200 , n423990 );
and ( n78202 , n424534 , n78201 );
and ( n78203 , n424480 , n424534 );
or ( n78204 , n78148 , n78202 , n78203 );
buf ( n424540 , n78204 );
buf ( n424541 , n67987 );
buf ( n424542 , n63625 );
and ( n78208 , n424541 , n424542 );
buf ( n424544 , n414714 );
buf ( n424545 , n63629 );
and ( n78211 , n424544 , n424545 );
nor ( n78212 , n78208 , n78211 );
buf ( n424548 , n78212 );
buf ( n424549 , n424548 );
buf ( n424550 , n410635 );
or ( n78216 , n424549 , n424550 );
buf ( n424552 , n424041 );
buf ( n424553 , n409504 );
or ( n78219 , n424552 , n424553 );
nand ( n78220 , n78216 , n78219 );
buf ( n424556 , n78220 );
buf ( n424557 , n424556 );
xor ( n78223 , n424540 , n424557 );
xor ( n78224 , n423994 , n423997 );
xor ( n78225 , n78224 , n424020 );
buf ( n424561 , n78225 );
buf ( n424562 , n424561 );
and ( n78228 , n78223 , n424562 );
and ( n78229 , n424540 , n424557 );
or ( n78230 , n78228 , n78229 );
buf ( n424566 , n78230 );
xor ( n78232 , n423941 , n424024 );
xor ( n78233 , n78232 , n424046 );
and ( n424569 , n424566 , n78233 );
buf ( n424570 , n66270 );
buf ( n424571 , n62499 );
and ( n78237 , n424570 , n424571 );
buf ( n424573 , n413098 );
buf ( n424574 , n62496 );
and ( n78240 , n424573 , n424574 );
nor ( n78241 , n78237 , n78240 );
buf ( n424577 , n78241 );
buf ( n424578 , n424577 );
buf ( n424579 , n410724 );
or ( n78245 , n424578 , n424579 );
buf ( n424581 , n424191 );
buf ( n424582 , n410721 );
or ( n78248 , n424581 , n424582 );
nand ( n78249 , n78245 , n78248 );
buf ( n424585 , n78249 );
xor ( n424586 , n424147 , n424150 );
xor ( n78252 , n424586 , n424169 );
and ( n78253 , n424585 , n78252 );
buf ( n424589 , n70210 );
buf ( n424590 , n62177 );
and ( n78256 , n424589 , n424590 );
buf ( n424592 , n416845 );
buf ( n424593 , n62159 );
and ( n78259 , n424592 , n424593 );
nor ( n424595 , n78256 , n78259 );
buf ( n424596 , n424595 );
buf ( n424597 , n424596 );
buf ( n424598 , n409429 );
or ( n78264 , n424597 , n424598 );
buf ( n424600 , n424164 );
buf ( n424601 , n409170 );
or ( n78267 , n424600 , n424601 );
nand ( n78268 , n78264 , n78267 );
buf ( n424604 , n78268 );
xor ( n78270 , n424101 , n424117 );
xor ( n78271 , n78270 , n424144 );
and ( n78272 , n424604 , n78271 );
buf ( n424608 , n409507 );
not ( n78274 , n424608 );
buf ( n424610 , n68002 );
buf ( n424611 , n63625 );
and ( n78277 , n424610 , n424611 );
buf ( n424613 , n414729 );
buf ( n424614 , n63629 );
and ( n78280 , n424613 , n424614 );
nor ( n78281 , n78277 , n78280 );
buf ( n424617 , n78281 );
not ( n78283 , n424617 );
buf ( n424619 , n78283 );
not ( n78285 , n424619 );
or ( n78286 , n78274 , n78285 );
buf ( n424622 , n424548 );
buf ( n424623 , n409504 );
or ( n78289 , n424622 , n424623 );
nand ( n78290 , n78286 , n78289 );
buf ( n424626 , n78290 );
xor ( n78292 , n424101 , n424117 );
xor ( n78293 , n78292 , n424144 );
and ( n78294 , n424626 , n78293 );
and ( n78295 , n424604 , n424626 );
or ( n78296 , n78272 , n78294 , n78295 );
xor ( n78297 , n424147 , n424150 );
xor ( n78298 , n78297 , n424169 );
and ( n78299 , n78296 , n78298 );
and ( n78300 , n424585 , n78296 );
or ( n78301 , n78253 , n78299 , n78300 );
xor ( n78302 , n423941 , n424024 );
xor ( n78303 , n78302 , n424046 );
and ( n78304 , n78301 , n78303 );
and ( n78305 , n424566 , n78301 );
or ( n78306 , n424569 , n78304 , n78305 );
xor ( n78307 , n77737 , n424201 );
xor ( n78308 , n78307 , n424205 );
and ( n78309 , n78306 , n78308 );
xor ( n78310 , n424540 , n424557 );
xor ( n78311 , n78310 , n424562 );
buf ( n424647 , n78311 );
buf ( n424648 , n66359 );
buf ( n424649 , n62499 );
and ( n78315 , n424648 , n424649 );
buf ( n424651 , n413187 );
buf ( n424652 , n62496 );
and ( n78318 , n424651 , n424652 );
nor ( n78319 , n78315 , n78318 );
buf ( n424655 , n78319 );
buf ( n424656 , n424655 );
buf ( n424657 , n410724 );
or ( n78323 , n424656 , n424657 );
buf ( n424659 , n424577 );
buf ( n424660 , n410721 );
or ( n78326 , n424659 , n424660 );
nand ( n78327 , n78323 , n78326 );
buf ( n424663 , n78327 );
buf ( n424664 , n424663 );
buf ( n424665 , n59637 );
buf ( n424666 , n14083 );
buf ( n424667 , n71170 );
and ( n78333 , n424666 , n424667 );
buf ( n424669 , n417804 );
buf ( n424670 , n59457 );
and ( n78336 , n424669 , n424670 );
nor ( n78337 , n78333 , n78336 );
buf ( n424673 , n78337 );
buf ( n424674 , n424673 );
or ( n78340 , n424665 , n424674 );
buf ( n424676 , n424516 );
buf ( n424677 , n59467 );
or ( n78343 , n424676 , n424677 );
nand ( n424679 , n78340 , n78343 );
buf ( n424680 , n424679 );
buf ( n424681 , n15626 );
buf ( n424682 , n623 );
and ( n78348 , n424681 , n424682 );
buf ( n424684 , n353695 );
buf ( n424685 , n422315 );
and ( n78351 , n424684 , n424685 );
buf ( n424687 , n56041 );
nor ( n78353 , n78351 , n424687 );
buf ( n424689 , n78353 );
buf ( n424690 , n424689 );
buf ( n424691 , n15287 );
nor ( n78357 , n78348 , n424690 , n424691 );
buf ( n424693 , n78357 );
xor ( n78359 , n424680 , n424693 );
buf ( n424695 , n403293 );
buf ( n424696 , n56041 );
buf ( n424697 , n74002 );
and ( n78363 , n424696 , n424697 );
buf ( n424699 , n403298 );
buf ( n424700 , n420612 );
and ( n78366 , n424699 , n424700 );
nor ( n78367 , n78363 , n78366 );
buf ( n424703 , n78367 );
buf ( n424704 , n424703 );
or ( n78370 , n424695 , n424704 );
buf ( n424706 , n424499 );
buf ( n424707 , n405476 );
or ( n78373 , n424706 , n424707 );
nand ( n78374 , n78370 , n78373 );
buf ( n424710 , n78374 );
and ( n78376 , n78359 , n424710 );
and ( n78377 , n424680 , n424693 );
or ( n78378 , n78376 , n78377 );
buf ( n424714 , n78378 );
xor ( n78380 , n424123 , n424142 );
buf ( n424716 , n78380 );
buf ( n424717 , n424716 );
xor ( n78383 , n424714 , n424717 );
buf ( n424719 , n409173 );
not ( n78385 , n424719 );
buf ( n424721 , n417024 );
buf ( n424722 , n409178 );
or ( n78388 , n424721 , n424722 );
buf ( n424724 , n70389 );
buf ( n424725 , n62177 );
or ( n78391 , n424724 , n424725 );
nand ( n78392 , n78388 , n78391 );
buf ( n424728 , n78392 );
buf ( n424729 , n424728 );
not ( n78395 , n424729 );
or ( n78396 , n78385 , n78395 );
buf ( n424732 , n424596 );
buf ( n424733 , n409170 );
or ( n78399 , n424732 , n424733 );
nand ( n78400 , n78396 , n78399 );
buf ( n424736 , n78400 );
buf ( n424737 , n424736 );
and ( n78403 , n78383 , n424737 );
and ( n78404 , n424714 , n424717 );
or ( n78405 , n78403 , n78404 );
buf ( n424741 , n78405 );
buf ( n424742 , n424741 );
xor ( n78408 , n424664 , n424742 );
xor ( n78409 , n423957 , n423973 );
xor ( n78410 , n78409 , n423990 );
xor ( n78411 , n424480 , n424534 );
xor ( n78412 , n78410 , n78411 );
buf ( n424748 , n78412 );
and ( n78414 , n78408 , n424748 );
and ( n78415 , n424664 , n424742 );
or ( n78416 , n78414 , n78415 );
buf ( n424752 , n78416 );
xor ( n78418 , n424647 , n424752 );
xor ( n78419 , n424147 , n424150 );
xor ( n78420 , n78419 , n424169 );
xor ( n78421 , n424585 , n78296 );
xor ( n78422 , n78420 , n78421 );
and ( n78423 , n78418 , n78422 );
and ( n78424 , n424647 , n424752 );
or ( n78425 , n78423 , n78424 );
buf ( n424761 , n78425 );
xor ( n78427 , n423889 , n423905 );
xor ( n78428 , n78427 , n423927 );
xor ( n78429 , n424172 , n424196 );
xor ( n78430 , n78428 , n78429 );
buf ( n424766 , n78430 );
xor ( n78432 , n424761 , n424766 );
xor ( n78433 , n423941 , n424024 );
xor ( n78434 , n78433 , n424046 );
xor ( n78435 , n424566 , n78301 );
xor ( n78436 , n78434 , n78435 );
buf ( n424772 , n78436 );
and ( n78438 , n78432 , n424772 );
and ( n424774 , n424761 , n424766 );
or ( n78440 , n78438 , n424774 );
buf ( n424776 , n78440 );
xor ( n78442 , n77737 , n424201 );
xor ( n78443 , n78442 , n424205 );
and ( n78444 , n424776 , n78443 );
and ( n78445 , n78306 , n424776 );
or ( n78446 , n78309 , n78444 , n78445 );
not ( n78447 , n78446 );
buf ( n424783 , n394210 );
not ( n78449 , n424783 );
buf ( n424785 , n390985 );
not ( n78451 , n424785 );
or ( n78452 , n78449 , n78451 );
buf ( n424788 , n390988 );
buf ( n424789 , n394207 );
nand ( n78455 , n424788 , n424789 );
buf ( n424791 , n78455 );
buf ( n424792 , n424791 );
nand ( n78458 , n78452 , n424792 );
buf ( n424794 , n78458 );
buf ( n424795 , n424794 );
not ( n78461 , n424795 );
buf ( n424797 , n44770 );
not ( n78463 , n424797 );
or ( n78464 , n78461 , n78463 );
buf ( n424800 , n44775 );
not ( n78466 , n424800 );
buf ( n424802 , n392878 );
not ( n78468 , n424802 );
or ( n78469 , n78466 , n78468 );
buf ( n424805 , n390985 );
buf ( n424806 , n392878 );
not ( n78472 , n424806 );
buf ( n424808 , n78472 );
buf ( n424809 , n424808 );
nand ( n78475 , n424805 , n424809 );
buf ( n424811 , n78475 );
buf ( n424812 , n424811 );
nand ( n78478 , n78469 , n424812 );
buf ( n424814 , n78478 );
buf ( n424815 , n424814 );
buf ( n424816 , n392740 );
nand ( n78482 , n424815 , n424816 );
buf ( n424818 , n78482 );
buf ( n424819 , n424818 );
nand ( n78485 , n78464 , n424819 );
buf ( n424821 , n78485 );
not ( n78487 , n424821 );
or ( n78488 , n78447 , n78487 );
buf ( n424824 , n424821 );
buf ( n424825 , n78446 );
or ( n78491 , n424824 , n424825 );
xor ( n78492 , n424209 , n424213 );
xor ( n78493 , n78492 , n424219 );
buf ( n424829 , n78493 );
buf ( n424830 , n424829 );
nand ( n78496 , n78491 , n424830 );
buf ( n424832 , n78496 );
nand ( n78498 , n78488 , n424832 );
not ( n78499 , n78498 );
xor ( n78500 , n76008 , n422643 );
xor ( n78501 , n78500 , n422647 );
xor ( n78502 , n424081 , n424223 );
xor ( n78503 , n78501 , n78502 );
buf ( n424839 , n78503 );
not ( n78505 , n424839 );
buf ( n424841 , n78505 );
buf ( n424842 , n423853 );
buf ( n424843 , n413643 );
and ( n78509 , n424842 , n424843 );
buf ( n424845 , n424814 );
not ( n78511 , n424845 );
buf ( n424847 , n44771 );
nor ( n78513 , n78511 , n424847 );
buf ( n424849 , n78513 );
buf ( n424850 , n424849 );
nor ( n78516 , n78509 , n424850 );
buf ( n424852 , n78516 );
nand ( n424853 , n424841 , n424852 );
not ( n78519 , n424853 );
or ( n78520 , n78499 , n78519 );
buf ( n424856 , n424852 );
not ( n78522 , n424856 );
buf ( n424858 , n78503 );
nand ( n78524 , n78522 , n424858 );
buf ( n424860 , n78524 );
nand ( n78526 , n78520 , n424860 );
buf ( n424862 , n78526 );
xor ( n78528 , n424464 , n424862 );
buf ( n424864 , n49117 );
not ( n78530 , n424864 );
buf ( n424866 , n423571 );
not ( n78532 , n424866 );
or ( n78533 , n78530 , n78532 );
buf ( n424869 , n388722 );
buf ( n424870 , n67126 );
nand ( n78536 , n424869 , n424870 );
buf ( n424872 , n78536 );
buf ( n424873 , n424872 );
nand ( n78539 , n78533 , n424873 );
buf ( n424875 , n78539 );
buf ( n424876 , n424875 );
not ( n78542 , n424876 );
buf ( n424878 , n40592 );
not ( n78544 , n424878 );
or ( n78545 , n78542 , n78544 );
buf ( n424881 , n423582 );
buf ( n424882 , n388068 );
nand ( n78548 , n424881 , n424882 );
buf ( n424884 , n78548 );
buf ( n424885 , n424884 );
nand ( n78551 , n78545 , n424885 );
buf ( n424887 , n78551 );
buf ( n424888 , n424887 );
and ( n78554 , n78528 , n424888 );
and ( n78555 , n424464 , n424862 );
or ( n78556 , n78554 , n78555 );
buf ( n424892 , n78556 );
buf ( n424893 , n424892 );
xor ( n78559 , n424443 , n424893 );
buf ( n424895 , n45954 );
not ( n78561 , n424895 );
buf ( n424897 , n423635 );
not ( n78563 , n424897 );
or ( n78564 , n78561 , n78563 );
buf ( n424900 , n393369 );
buf ( n424901 , n41861 );
and ( n78567 , n424900 , n424901 );
not ( n78568 , n424900 );
buf ( n424904 , n418729 );
and ( n78570 , n78568 , n424904 );
nor ( n78571 , n78567 , n78570 );
buf ( n424907 , n78571 );
buf ( n424908 , n424907 );
buf ( n424909 , n45949 );
nand ( n78575 , n424908 , n424909 );
buf ( n424911 , n78575 );
buf ( n424912 , n424911 );
nand ( n78578 , n78564 , n424912 );
buf ( n424914 , n78578 );
buf ( n424915 , n424914 );
and ( n78581 , n78559 , n424915 );
and ( n78582 , n424443 , n424893 );
or ( n78583 , n78581 , n78582 );
buf ( n424919 , n78583 );
buf ( n424920 , n424919 );
buf ( n424921 , n66132 );
not ( n78587 , n424921 );
buf ( n424923 , n388128 );
not ( n78589 , n424923 );
or ( n78590 , n78587 , n78589 );
buf ( n424926 , n358975 );
nand ( n78592 , n78590 , n424926 );
buf ( n424928 , n78592 );
buf ( n424929 , n424928 );
buf ( n424930 , n407928 );
buf ( n424931 , n41365 );
buf ( n424932 , n23900 );
nand ( n78598 , n424931 , n424932 );
buf ( n424934 , n78598 );
buf ( n424935 , n424934 );
and ( n78601 , n424929 , n424930 , n424935 );
buf ( n424937 , n78601 );
buf ( n424938 , n424937 );
xor ( n78604 , n424920 , n424938 );
xor ( n78605 , n423600 , n423617 );
xor ( n78606 , n78605 , n423643 );
buf ( n424942 , n78606 );
buf ( n424943 , n424942 );
and ( n78609 , n78604 , n424943 );
and ( n78610 , n424920 , n424938 );
or ( n78611 , n78609 , n78610 );
buf ( n424947 , n78611 );
buf ( n424948 , n424947 );
xor ( n78614 , n423530 , n423534 );
xor ( n78615 , n78614 , n423648 );
buf ( n424951 , n78615 );
buf ( n424952 , n424951 );
xor ( n78618 , n424948 , n424952 );
buf ( n424954 , n59916 );
not ( n78620 , n424954 );
buf ( n424956 , n424365 );
not ( n78622 , n424956 );
or ( n78623 , n78620 , n78622 );
buf ( n424959 , n47891 );
not ( n78625 , n424959 );
buf ( n424961 , n405126 );
not ( n78627 , n424961 );
or ( n424963 , n78625 , n78627 );
buf ( n424964 , n12471 );
buf ( n424965 , n72794 );
nand ( n78631 , n424964 , n424965 );
buf ( n424967 , n78631 );
buf ( n424968 , n424967 );
nand ( n78634 , n424963 , n424968 );
buf ( n424970 , n78634 );
buf ( n424971 , n424970 );
buf ( n424972 , n50579 );
nand ( n78638 , n424971 , n424972 );
buf ( n424974 , n78638 );
buf ( n424975 , n424974 );
nand ( n78641 , n78623 , n424975 );
buf ( n424977 , n78641 );
buf ( n424978 , n424977 );
and ( n78644 , n78618 , n424978 );
and ( n78645 , n424948 , n424952 );
or ( n78646 , n78644 , n78645 );
buf ( n424982 , n78646 );
buf ( n424983 , n424982 );
buf ( n424984 , n423659 );
buf ( n424985 , n423663 );
and ( n78651 , n424984 , n424985 );
not ( n78652 , n424984 );
buf ( n424988 , n423510 );
and ( n78654 , n78652 , n424988 );
nor ( n78655 , n78651 , n78654 );
buf ( n424991 , n78655 );
xor ( n78657 , n424991 , n423652 );
buf ( n424993 , n78657 );
not ( n78659 , n424993 );
buf ( n424995 , n78659 );
buf ( n424996 , n424995 );
nor ( n78662 , n42923 , n402819 );
buf ( n424998 , n78662 );
buf ( n424999 , n395359 );
not ( n78665 , n424999 );
buf ( n425001 , n423741 );
not ( n78667 , n425001 );
or ( n78668 , n78665 , n78667 );
and ( n78669 , n12480 , n421871 );
not ( n78670 , n12480 );
and ( n78671 , n78670 , n47863 );
or ( n78672 , n78669 , n78671 );
buf ( n425008 , n78672 );
buf ( n425009 , n395346 );
nand ( n78675 , n425008 , n425009 );
buf ( n425011 , n78675 );
buf ( n425012 , n425011 );
nand ( n78678 , n78668 , n425012 );
buf ( n425014 , n78678 );
buf ( n425015 , n425014 );
xor ( n78681 , n424998 , n425015 );
buf ( n425017 , n50041 );
buf ( n425018 , n404855 );
buf ( n425019 , n407928 );
and ( n78685 , n425018 , n425019 );
not ( n78686 , n425018 );
buf ( n425022 , n409092 );
and ( n78688 , n78686 , n425022 );
nor ( n78689 , n78685 , n78688 );
buf ( n425025 , n78689 );
buf ( n425026 , n425025 );
or ( n78692 , n425017 , n425026 );
buf ( n425028 , n423500 );
buf ( n425029 , n62075 );
or ( n78695 , n425028 , n425029 );
nand ( n78696 , n78692 , n78695 );
buf ( n425032 , n78696 );
buf ( n425033 , n425032 );
and ( n78699 , n78681 , n425033 );
and ( n78700 , n424998 , n425015 );
or ( n78701 , n78699 , n78700 );
buf ( n425037 , n78701 );
buf ( n425038 , n425037 );
not ( n78704 , n425038 );
buf ( n425040 , n78704 );
buf ( n425041 , n425040 );
nand ( n78707 , n424996 , n425041 );
buf ( n425043 , n78707 );
buf ( n425044 , n425043 );
and ( n78710 , n424983 , n425044 );
buf ( n425046 , n425040 );
buf ( n425047 , n424995 );
nor ( n78713 , n425046 , n425047 );
buf ( n425049 , n78713 );
buf ( n425050 , n425049 );
nor ( n78716 , n78710 , n425050 );
buf ( n425052 , n78716 );
not ( n78718 , n425052 );
or ( n78719 , n78083 , n78718 );
xor ( n78720 , n423770 , n423800 );
xor ( n78721 , n78720 , n424289 );
not ( n78722 , n78721 );
xor ( n78723 , n423834 , n424239 );
xnor ( n78724 , n78723 , n424247 );
buf ( n425060 , n78724 );
buf ( n425061 , n77514 );
buf ( n425062 , n77877 );
xnor ( n78728 , n425061 , n425062 );
buf ( n425064 , n78728 );
buf ( n425065 , n425064 );
not ( n78731 , n425065 );
buf ( n425067 , n423860 );
not ( n78733 , n425067 );
or ( n78734 , n78731 , n78733 );
buf ( n425070 , n423860 );
buf ( n425071 , n425064 );
or ( n78737 , n425070 , n425071 );
nand ( n78738 , n78734 , n78737 );
buf ( n425074 , n78738 );
buf ( n425075 , n425074 );
buf ( n425076 , n45954 );
not ( n78742 , n425076 );
buf ( n425078 , n424907 );
not ( n78744 , n425078 );
or ( n78745 , n78742 , n78744 );
buf ( n425081 , n393369 );
not ( n78747 , n425081 );
buf ( n425083 , n420954 );
not ( n78749 , n425083 );
or ( n78750 , n78747 , n78749 );
buf ( n425086 , n389338 );
buf ( n425087 , n393381 );
nand ( n78753 , n425086 , n425087 );
buf ( n425089 , n78753 );
buf ( n425090 , n425089 );
nand ( n78756 , n78750 , n425090 );
buf ( n425092 , n78756 );
buf ( n425093 , n425092 );
buf ( n425094 , n45949 );
nand ( n78760 , n425093 , n425094 );
buf ( n425096 , n78760 );
buf ( n425097 , n425096 );
nand ( n78763 , n78745 , n425097 );
buf ( n425099 , n78763 );
buf ( n425100 , n425099 );
xor ( n78766 , n425075 , n425100 );
buf ( n425102 , n417572 );
not ( n78768 , n425102 );
buf ( n425104 , n420986 );
not ( n78770 , n425104 );
or ( n78771 , n78768 , n78770 );
buf ( n425107 , n391018 );
buf ( n425108 , n394814 );
nand ( n78774 , n425107 , n425108 );
buf ( n425110 , n78774 );
buf ( n425111 , n425110 );
nand ( n78777 , n78771 , n425111 );
buf ( n425113 , n78777 );
buf ( n425114 , n425113 );
not ( n78780 , n425114 );
buf ( n425116 , n74375 );
not ( n78782 , n425116 );
or ( n78783 , n78780 , n78782 );
buf ( n425119 , n424451 );
buf ( n425120 , n43515 );
nand ( n78786 , n425119 , n425120 );
buf ( n425122 , n78786 );
buf ( n425123 , n425122 );
nand ( n78789 , n78783 , n425123 );
buf ( n425125 , n78789 );
buf ( n425126 , n425125 );
buf ( n425127 , n45954 );
not ( n78793 , n425127 );
buf ( n425129 , n425092 );
not ( n78795 , n425129 );
or ( n78796 , n78793 , n78795 );
buf ( n425132 , n393369 );
not ( n78798 , n425132 );
buf ( n425134 , n391440 );
not ( n78800 , n425134 );
or ( n78801 , n78798 , n78800 );
buf ( n425137 , n420994 );
buf ( n425138 , n393381 );
nand ( n78804 , n425137 , n425138 );
buf ( n425140 , n78804 );
buf ( n425141 , n425140 );
nand ( n78807 , n78801 , n425141 );
buf ( n425143 , n78807 );
buf ( n425144 , n425143 );
buf ( n425145 , n45949 );
nand ( n78811 , n425144 , n425145 );
buf ( n425147 , n78811 );
buf ( n425148 , n425147 );
nand ( n78814 , n78796 , n425148 );
buf ( n425150 , n78814 );
buf ( n425151 , n425150 );
xor ( n78817 , n425126 , n425151 );
buf ( n425153 , n397489 );
not ( n78819 , n425153 );
buf ( n425155 , n423571 );
not ( n78821 , n425155 );
or ( n78822 , n78819 , n78821 );
buf ( n425158 , n388722 );
buf ( n425159 , n397486 );
nand ( n78825 , n425158 , n425159 );
buf ( n425161 , n78825 );
buf ( n425162 , n425161 );
nand ( n78828 , n78822 , n425162 );
buf ( n425164 , n78828 );
buf ( n425165 , n425164 );
not ( n78831 , n425165 );
buf ( n425167 , n67042 );
not ( n78833 , n425167 );
or ( n78834 , n78831 , n78833 );
buf ( n425170 , n424875 );
buf ( n425171 , n388068 );
nand ( n78837 , n425170 , n425171 );
buf ( n425173 , n78837 );
buf ( n425174 , n425173 );
nand ( n78840 , n78834 , n425174 );
buf ( n425176 , n78840 );
buf ( n425177 , n425176 );
and ( n78843 , n78817 , n425177 );
and ( n78844 , n425126 , n425151 );
or ( n78845 , n78843 , n78844 );
buf ( n425181 , n78845 );
buf ( n425182 , n425181 );
and ( n78848 , n78766 , n425182 );
and ( n78849 , n425075 , n425100 );
or ( n78850 , n78848 , n78849 );
buf ( n425186 , n78850 );
buf ( n425187 , n425186 );
xor ( n78853 , n425060 , n425187 );
buf ( n425189 , n74538 );
buf ( n425190 , n399283 );
buf ( n425191 , n24116 );
and ( n78857 , n425190 , n425191 );
not ( n78858 , n425190 );
buf ( n425194 , n62006 );
and ( n78860 , n78858 , n425194 );
nor ( n78861 , n78857 , n78860 );
buf ( n425197 , n78861 );
buf ( n425198 , n425197 );
or ( n78864 , n425189 , n425198 );
buf ( n425200 , n424272 );
not ( n78866 , n425200 );
buf ( n425202 , n78866 );
buf ( n425203 , n425202 );
buf ( n425204 , n74561 );
or ( n78870 , n425203 , n425204 );
nand ( n78871 , n78864 , n78870 );
buf ( n425207 , n78871 );
buf ( n425208 , n425207 );
and ( n78874 , n78853 , n425208 );
and ( n78875 , n425060 , n425187 );
or ( n78876 , n78874 , n78875 );
buf ( n425212 , n78876 );
not ( n78878 , n425212 );
buf ( n425214 , n78672 );
buf ( n425215 , n395359 );
and ( n78881 , n425214 , n425215 );
buf ( n425217 , n47863 );
not ( n78883 , n425217 );
buf ( n425219 , n417349 );
not ( n78885 , n425219 );
or ( n78886 , n78883 , n78885 );
buf ( n425222 , n28353 );
buf ( n425223 , n421871 );
nand ( n78889 , n425222 , n425223 );
buf ( n425225 , n78889 );
buf ( n425226 , n425225 );
nand ( n78892 , n78886 , n425226 );
buf ( n425228 , n78892 );
buf ( n425229 , n425228 );
not ( n78895 , n425229 );
buf ( n425231 , n47904 );
nor ( n78897 , n78895 , n425231 );
buf ( n425233 , n78897 );
buf ( n425234 , n425233 );
nor ( n78900 , n78881 , n425234 );
buf ( n425236 , n78900 );
buf ( n425237 , n425236 );
buf ( n425238 , n400033 );
not ( n78904 , n425238 );
buf ( n425240 , n416292 );
not ( n78906 , n425240 );
or ( n78907 , n78904 , n78906 );
buf ( n425243 , n416298 );
buf ( n425244 , n400042 );
nand ( n425245 , n425243 , n425244 );
buf ( n425246 , n425245 );
buf ( n425247 , n425246 );
nand ( n78913 , n78907 , n425247 );
buf ( n425249 , n78913 );
not ( n78915 , n425249 );
not ( n78916 , n66128 );
or ( n78917 , n78915 , n78916 );
buf ( n425253 , n423787 );
buf ( n425254 , n412976 );
nand ( n78920 , n425253 , n425254 );
buf ( n425256 , n78920 );
nand ( n78922 , n78917 , n425256 );
not ( n78923 , n78922 );
buf ( n425259 , n78923 );
nand ( n78925 , n425237 , n425259 );
buf ( n425261 , n78925 );
not ( n78927 , n425261 );
or ( n78928 , n78878 , n78927 );
not ( n78929 , n425236 );
nand ( n78930 , n78929 , n78922 );
nand ( n78931 , n78928 , n78930 );
nand ( n78932 , n78722 , n78931 );
not ( n78933 , n78721 );
not ( n78934 , n78931 );
not ( n78935 , n78934 );
or ( n78936 , n78933 , n78935 );
xor ( n78937 , n423810 , n424259 );
xor ( n78938 , n78937 , n424285 );
buf ( n425274 , n78938 );
buf ( n425275 , n425274 );
buf ( n425276 , n395359 );
not ( n78942 , n425276 );
buf ( n425278 , n425228 );
not ( n78944 , n425278 );
or ( n78945 , n78942 , n78944 );
buf ( n425281 , n47863 );
not ( n78947 , n425281 );
buf ( n425283 , n27320 );
not ( n78949 , n425283 );
buf ( n425285 , n78949 );
buf ( n425286 , n425285 );
not ( n78952 , n425286 );
or ( n78953 , n78947 , n78952 );
buf ( n425289 , n27320 );
buf ( n425290 , n421871 );
nand ( n78956 , n425289 , n425290 );
buf ( n425292 , n78956 );
buf ( n425293 , n425292 );
nand ( n78959 , n78953 , n425293 );
buf ( n425295 , n78959 );
buf ( n425296 , n425295 );
buf ( n425297 , n395346 );
nand ( n78963 , n425296 , n425297 );
buf ( n425299 , n78963 );
buf ( n425300 , n425299 );
nand ( n78966 , n78945 , n425300 );
buf ( n425302 , n78966 );
buf ( n425303 , n425302 );
not ( n78969 , n425303 );
buf ( n425305 , n78969 );
buf ( n425306 , n425305 );
not ( n78972 , n425306 );
buf ( n425308 , n62075 );
not ( n78974 , n425308 );
buf ( n425310 , n358975 );
nand ( n78976 , n78974 , n425310 );
buf ( n425312 , n78976 );
buf ( n425313 , n425312 );
not ( n78979 , n425313 );
or ( n78980 , n78972 , n78979 );
xor ( n78981 , n424443 , n424893 );
xor ( n78982 , n78981 , n424915 );
buf ( n425318 , n78982 );
buf ( n425319 , n425318 );
nand ( n78985 , n78980 , n425319 );
buf ( n425321 , n78985 );
buf ( n425322 , n425321 );
buf ( n425323 , n425312 );
not ( n78989 , n425323 );
buf ( n425325 , n78989 );
buf ( n425326 , n425325 );
buf ( n425327 , n425302 );
nand ( n78993 , n425326 , n425327 );
buf ( n425329 , n78993 );
buf ( n425330 , n425329 );
nand ( n78996 , n425322 , n425330 );
buf ( n425332 , n78996 );
buf ( n425333 , n425332 );
xor ( n78999 , n425275 , n425333 );
xor ( n79000 , n424920 , n424938 );
xor ( n79001 , n79000 , n424943 );
buf ( n425337 , n79001 );
buf ( n425338 , n425337 );
and ( n79004 , n78999 , n425338 );
and ( n79005 , n425275 , n425333 );
or ( n79006 , n79004 , n79005 );
buf ( n425342 , n79006 );
nand ( n79008 , n78936 , n425342 );
nand ( n79009 , n78932 , n79008 );
buf ( n425345 , n79009 );
xor ( n79011 , n423724 , n423749 );
xor ( n79012 , n79011 , n424296 );
buf ( n425348 , n79012 );
buf ( n425349 , n425348 );
buf ( n425350 , C0 );
buf ( n425351 , n425350 );
and ( n79040 , n425345 , n425349 );
or ( n79041 , C0 , n79040 );
buf ( n425354 , n79041 );
nand ( n79043 , n78719 , n425354 );
buf ( n425356 , n424417 );
not ( n79045 , n425356 );
buf ( n425358 , n79045 );
buf ( n425359 , n425358 );
buf ( n425360 , n425052 );
not ( n79049 , n425360 );
buf ( n425362 , n79049 );
buf ( n425363 , n425362 );
nand ( n79052 , n425359 , n425363 );
buf ( n425365 , n79052 );
nand ( n79054 , n79043 , n425365 );
buf ( n425367 , n79054 );
nand ( n79056 , n78076 , n425367 );
buf ( n425369 , n79056 );
buf ( n425370 , n78073 );
buf ( n425371 , n424398 );
or ( n79060 , n425370 , n425371 );
buf ( n425373 , n79060 );
and ( n79062 , n425369 , n425373 );
buf ( n425375 , n79062 );
xor ( n79064 , n424322 , n425375 );
xor ( n79065 , n422766 , C0 );
xor ( n79066 , n79065 , n422770 );
buf ( n425379 , n79066 );
xor ( n79068 , n422775 , n422856 );
xor ( n79069 , n79068 , n422861 );
buf ( n425382 , n79069 );
buf ( n425383 , n425382 );
xor ( n79072 , n425379 , n425383 );
xor ( n79073 , n422016 , n422020 );
xor ( n79074 , n79073 , n422762 );
buf ( n425387 , n79074 );
buf ( n425388 , n425387 );
not ( n79077 , n425388 );
xor ( n79078 , n422796 , n422799 );
xor ( n79079 , n79078 , n422851 );
buf ( n425392 , n79079 );
buf ( n425393 , n425392 );
not ( n79082 , n425393 );
or ( n79083 , n79077 , n79082 );
xor ( n79084 , n423421 , n423423 );
xor ( n79085 , n79084 , n423428 );
buf ( n425398 , n79085 );
buf ( n425399 , n425398 );
buf ( n425400 , n425387 );
not ( n79089 , n425400 );
buf ( n425402 , n425392 );
not ( n79091 , n425402 );
buf ( n425404 , n79091 );
buf ( n425405 , n425404 );
nand ( n79094 , n79089 , n425405 );
buf ( n425407 , n79094 );
buf ( n425408 , n425407 );
nand ( n79097 , n425399 , n425408 );
buf ( n425410 , n79097 );
buf ( n425411 , n425410 );
nand ( n79100 , n79083 , n425411 );
buf ( n425413 , n79100 );
buf ( n425414 , n425413 );
xnor ( n79103 , n79072 , n425414 );
buf ( n425416 , n79103 );
buf ( n425417 , n425416 );
xor ( n79106 , n79064 , n425417 );
buf ( n425419 , n79106 );
buf ( n425420 , n425419 );
buf ( n425421 , C1 );
buf ( n425422 , n425421 );
buf ( n425423 , n424381 );
buf ( n425424 , n424346 );
xor ( n79130 , n425423 , n425424 );
buf ( n425426 , n424375 );
xor ( n79132 , n79130 , n425426 );
buf ( n425428 , n79132 );
buf ( n425429 , n425428 );
nand ( n79135 , n425422 , n425429 );
buf ( n425431 , n79135 );
buf ( n425432 , n425431 );
xor ( n79138 , n424998 , n425015 );
xor ( n79139 , n79138 , n425033 );
buf ( n425435 , n79139 );
buf ( n425436 , n425435 );
buf ( n425437 , C0 );
buf ( n425438 , n425437 );
xor ( n79166 , n425436 , n425438 );
buf ( n425440 , n50041 );
buf ( n425441 , n358975 );
buf ( n425442 , n388154 );
and ( n79170 , n425441 , n425442 );
not ( n79171 , n425441 );
buf ( n425445 , n405897 );
and ( n79173 , n79171 , n425445 );
nor ( n79174 , n79170 , n79173 );
buf ( n425448 , n79174 );
buf ( n425449 , n425448 );
or ( n79177 , n425440 , n425449 );
buf ( n425451 , n425025 );
buf ( n425452 , n62075 );
or ( n79180 , n425451 , n425452 );
nand ( n79181 , n79177 , n79180 );
buf ( n425455 , n79181 );
buf ( n425456 , n425455 );
buf ( n425457 , n395359 );
not ( n79185 , n425457 );
buf ( n425459 , n425295 );
not ( n79187 , n425459 );
or ( n79188 , n79185 , n79187 );
buf ( n425462 , n47863 );
not ( n79190 , n425462 );
buf ( n425464 , n72076 );
not ( n79192 , n425464 );
or ( n79193 , n79190 , n79192 );
buf ( n425467 , n42066 );
buf ( n425468 , n421871 );
nand ( n79196 , n425467 , n425468 );
buf ( n425470 , n79196 );
buf ( n425471 , n425470 );
nand ( n79199 , n79193 , n425471 );
buf ( n425473 , n79199 );
buf ( n425474 , n425473 );
buf ( n425475 , n395346 );
nand ( n79203 , n425474 , n425475 );
buf ( n425477 , n79203 );
buf ( n425478 , n425477 );
nand ( n79206 , n79188 , n425478 );
buf ( n425480 , n79206 );
buf ( n425481 , n425480 );
xor ( n79209 , n425075 , n425100 );
xor ( n79210 , n79209 , n425182 );
buf ( n425484 , n79210 );
buf ( n425485 , n425484 );
xor ( n79213 , n425481 , n425485 );
and ( n79214 , n424852 , n78503 );
not ( n79215 , n424852 );
and ( n79216 , n79215 , n424841 );
or ( n79217 , n79214 , n79216 );
xor ( n79218 , n79217 , n78498 );
xor ( n79219 , n424829 , n78446 );
xor ( n79220 , n79219 , n424821 );
buf ( n425494 , n79220 );
buf ( n425495 , n45954 );
not ( n79223 , n425495 );
buf ( n425497 , n425143 );
not ( n79225 , n425497 );
or ( n79226 , n79223 , n79225 );
buf ( n425500 , n393369 );
not ( n79228 , n425500 );
buf ( n425502 , n420908 );
not ( n79230 , n425502 );
or ( n79231 , n79228 , n79230 );
buf ( n425505 , n392608 );
buf ( n425506 , n393381 );
nand ( n79234 , n425505 , n425506 );
buf ( n425508 , n79234 );
buf ( n425509 , n425508 );
nand ( n79237 , n79231 , n425509 );
buf ( n425511 , n79237 );
buf ( n425512 , n425511 );
buf ( n425513 , n45949 );
nand ( n79241 , n425512 , n425513 );
buf ( n425515 , n79241 );
buf ( n425516 , n425515 );
nand ( n79244 , n79226 , n425516 );
buf ( n425518 , n79244 );
buf ( n425519 , n425518 );
xor ( n79247 , n425494 , n425519 );
buf ( n425521 , n49117 );
not ( n79249 , n425521 );
buf ( n425523 , n371879 );
not ( n79251 , n425523 );
buf ( n425525 , n79251 );
buf ( n425526 , n425525 );
not ( n79254 , n425526 );
or ( n79255 , n79249 , n79254 );
buf ( n425529 , n390997 );
buf ( n425530 , n67126 );
nand ( n79258 , n425529 , n425530 );
buf ( n425532 , n79258 );
buf ( n425533 , n425532 );
nand ( n79261 , n79255 , n425533 );
buf ( n425535 , n79261 );
buf ( n425536 , n425535 );
not ( n79264 , n425536 );
buf ( n425538 , n74375 );
not ( n79266 , n425538 );
or ( n79267 , n79264 , n79266 );
buf ( n425541 , n425113 );
buf ( n425542 , n43515 );
nand ( n79270 , n425541 , n425542 );
buf ( n425544 , n79270 );
buf ( n425545 , n425544 );
nand ( n79273 , n79267 , n425545 );
buf ( n425547 , n79273 );
buf ( n425548 , n425547 );
and ( n79276 , n79247 , n425548 );
and ( n79277 , n425494 , n425519 );
or ( n79278 , n79276 , n79277 );
buf ( n425552 , n79278 );
xor ( n79280 , n79218 , n425552 );
buf ( n425554 , n395359 );
not ( n79282 , n425554 );
buf ( n425556 , n425473 );
not ( n79284 , n425556 );
or ( n79285 , n79282 , n79284 );
buf ( n425559 , n47863 );
buf ( n425560 , n41861 );
and ( n79288 , n425559 , n425560 );
not ( n79289 , n425559 );
buf ( n425563 , n418729 );
and ( n79291 , n79289 , n425563 );
nor ( n79292 , n79288 , n79291 );
buf ( n425566 , n79292 );
buf ( n425567 , n425566 );
buf ( n425568 , n395346 );
nand ( n79296 , n425567 , n425568 );
buf ( n425570 , n79296 );
buf ( n425571 , n425570 );
nand ( n79299 , n79285 , n425571 );
buf ( n425573 , n79299 );
and ( n79301 , n79280 , n425573 );
and ( n79302 , n79218 , n425552 );
or ( n79303 , n79301 , n79302 );
buf ( n425577 , n79303 );
and ( n79305 , n79213 , n425577 );
and ( n79306 , n425481 , n425485 );
or ( n79307 , n79305 , n79306 );
buf ( n425581 , n79307 );
buf ( n425582 , n425581 );
xor ( n79310 , n424464 , n424862 );
xor ( n79311 , n79310 , n424888 );
buf ( n425585 , n79311 );
buf ( n425586 , n425585 );
buf ( n425587 , n55543 );
buf ( n425588 , n371800 );
and ( n79316 , n425587 , n425588 );
not ( n79317 , n425587 );
buf ( n425591 , n371787 );
and ( n79319 , n79317 , n425591 );
nor ( n79320 , n79316 , n79319 );
buf ( n425594 , n79320 );
buf ( n425595 , n425594 );
not ( n79323 , n425595 );
buf ( n425597 , n388740 );
not ( n79325 , n425597 );
or ( n79326 , n79323 , n79325 );
buf ( n425600 , n424430 );
buf ( n425601 , n388803 );
nand ( n79329 , n425600 , n425601 );
buf ( n425603 , n79329 );
buf ( n425604 , n425603 );
nand ( n79332 , n79326 , n425604 );
buf ( n425606 , n79332 );
buf ( n425607 , n425606 );
xor ( n79335 , n425586 , n425607 );
buf ( n425609 , n410407 );
not ( n79337 , n371420 );
not ( n79338 , n24116 );
or ( n79339 , n79337 , n79338 );
buf ( n425613 , n371420 );
buf ( n425614 , n24116 );
nor ( n79342 , n425613 , n425614 );
buf ( n425616 , n79342 );
or ( n79344 , n425616 , n402819 );
nand ( n79345 , n79339 , n79344 );
buf ( n425619 , n79345 );
nor ( n79347 , n425609 , n425619 );
buf ( n425621 , n79347 );
buf ( n425622 , n425621 );
and ( n79350 , n79335 , n425622 );
and ( n79351 , n425586 , n425607 );
or ( n79352 , n79350 , n79351 );
buf ( n425626 , n79352 );
buf ( n425627 , n425626 );
xor ( n79355 , n425582 , n425627 );
buf ( n425629 , n41374 );
buf ( n425630 , n55055 );
not ( n79358 , n425630 );
buf ( n425632 , n41341 );
not ( n79360 , n425632 );
or ( n79361 , n79358 , n79360 );
buf ( n425635 , n23841 );
buf ( n425636 , n55054 );
nand ( n79364 , n425635 , n425636 );
buf ( n425638 , n79364 );
buf ( n425639 , n425638 );
nand ( n79367 , n79361 , n425639 );
buf ( n425641 , n79367 );
buf ( n425642 , n425641 );
not ( n79370 , n425642 );
buf ( n425644 , n79370 );
buf ( n425645 , n425644 );
or ( n79373 , n425629 , n425645 );
buf ( n425647 , n425249 );
not ( n79375 , n425647 );
buf ( n425649 , n79375 );
buf ( n425650 , n425649 );
buf ( n425651 , n41332 );
or ( n79379 , n425650 , n425651 );
nand ( n79380 , n79373 , n79379 );
buf ( n425654 , n79380 );
buf ( n425655 , n425654 );
and ( n79383 , n79355 , n425655 );
and ( n79384 , n425582 , n425627 );
or ( n79385 , n79383 , n79384 );
buf ( n425659 , n79385 );
buf ( n425660 , n425659 );
xor ( n79388 , n425456 , n425660 );
buf ( n425662 , n61577 );
not ( n79390 , n425662 );
buf ( n425664 , n424970 );
not ( n79392 , n425664 );
or ( n79393 , n79390 , n79392 );
buf ( n425667 , n47891 );
not ( n79395 , n425667 );
buf ( n425669 , n388227 );
not ( n79397 , n425669 );
or ( n79398 , n79395 , n79397 );
buf ( n425672 , n406821 );
buf ( n425673 , n72794 );
nand ( n79401 , n425672 , n425673 );
buf ( n425675 , n79401 );
buf ( n425676 , n425675 );
nand ( n79404 , n79398 , n425676 );
buf ( n425678 , n79404 );
buf ( n425679 , n425678 );
buf ( n425680 , n50579 );
nand ( n79408 , n425679 , n425680 );
buf ( n425682 , n79408 );
buf ( n425683 , n425682 );
nand ( n79411 , n79393 , n425683 );
buf ( n425685 , n79411 );
buf ( n425686 , n425685 );
and ( n79414 , n79388 , n425686 );
and ( n79415 , n425456 , n425660 );
or ( n79416 , n79414 , n79415 );
buf ( n425690 , n79416 );
buf ( n425691 , n425690 );
and ( n79419 , n79166 , n425691 );
or ( n79421 , n79419 , C0 );
buf ( n425694 , n79421 );
buf ( n425695 , n425694 );
and ( n79424 , n425432 , n425695 );
buf ( n425697 , C0 );
buf ( n425698 , n425697 );
nor ( n79430 , n79424 , n425698 );
buf ( n425700 , n79430 );
not ( n79432 , n425700 );
xor ( n79433 , n424385 , n424392 );
xor ( n79434 , n79433 , n424394 );
buf ( n425704 , n79434 );
not ( n79436 , n425704 );
or ( n79437 , n79432 , n79436 );
or ( n79438 , n425704 , n425700 );
xor ( n79439 , n423700 , n424300 );
xnor ( n79440 , n79439 , n423696 );
not ( n79441 , n79440 );
nand ( n79442 , n79438 , n79441 );
nand ( n79443 , n79437 , n79442 );
buf ( n425713 , n425387 );
buf ( n425714 , n425404 );
and ( n79446 , n425713 , n425714 );
not ( n79447 , n425713 );
buf ( n425717 , n425392 );
and ( n79449 , n79447 , n425717 );
nor ( n79450 , n79446 , n79449 );
buf ( n425720 , n79450 );
xor ( n79452 , n425720 , n425398 );
xor ( n79453 , n79443 , n79452 );
xor ( n79454 , n424398 , n79054 );
xnor ( n79455 , n79454 , n78073 );
and ( n79456 , n79453 , n79455 );
and ( n79457 , n79443 , n79452 );
or ( n79458 , n79456 , n79457 );
buf ( n425728 , n79458 );
nand ( n79460 , n425420 , n425728 );
buf ( n425730 , n79460 );
not ( n79462 , n425730 );
xor ( n79463 , n79443 , n79452 );
xor ( n79464 , n79463 , n79455 );
buf ( n425734 , n79464 );
not ( n79466 , n425734 );
buf ( n425736 , n79466 );
buf ( n425737 , n425736 );
buf ( n425738 , n425358 );
not ( n79470 , n425738 );
buf ( n425740 , n425052 );
not ( n79472 , n425740 );
or ( n79473 , n79470 , n79472 );
buf ( n425743 , n424417 );
buf ( n425744 , n425362 );
nand ( n79476 , n425743 , n425744 );
buf ( n425746 , n79476 );
buf ( n425747 , n425746 );
nand ( n79479 , n79473 , n425747 );
buf ( n425749 , n79479 );
buf ( n425750 , n425749 );
buf ( n425751 , n425354 );
buf ( n79483 , n425751 );
buf ( n425753 , n79483 );
buf ( n425754 , n425753 );
xnor ( n79486 , n425750 , n425754 );
buf ( n425756 , n79486 );
not ( n79488 , n425756 );
not ( n79489 , n425704 );
xor ( n79490 , n79440 , n79489 );
xnor ( n79491 , n79490 , n425700 );
not ( n79492 , n79491 );
not ( n79493 , n79492 );
or ( n79494 , n79488 , n79493 );
buf ( n425764 , n425037 );
buf ( n425765 , n78657 );
xor ( n79497 , n425764 , n425765 );
buf ( n425767 , n424982 );
xor ( n79499 , n79497 , n425767 );
buf ( n425769 , n79499 );
not ( n79501 , n425769 );
xor ( n79502 , n424948 , n424952 );
xor ( n79503 , n79502 , n424978 );
buf ( n425773 , n79503 );
buf ( n425774 , n425773 );
not ( n79506 , n425342 );
not ( n79507 , n78721 );
not ( n79508 , n78931 );
and ( n79509 , n79507 , n79508 );
and ( n79510 , n78721 , n78931 );
nor ( n79511 , n79509 , n79510 );
not ( n79512 , n79511 );
or ( n79513 , n79506 , n79512 );
or ( n79514 , n79511 , n425342 );
nand ( n79515 , n79513 , n79514 );
buf ( n425785 , n79515 );
buf ( n425786 , C0 );
buf ( n425787 , n425786 );
and ( n79533 , n425774 , n425785 );
or ( n79534 , C0 , n79533 );
buf ( n425790 , n79534 );
not ( n79536 , n425790 );
or ( n79537 , n79501 , n79536 );
not ( n79538 , n425769 );
not ( n79539 , n79538 );
not ( n79540 , n425790 );
not ( n79541 , n79540 );
or ( n79542 , n79539 , n79541 );
xor ( n79543 , n425345 , n425349 );
xor ( n79544 , n79543 , n425351 );
buf ( n425800 , n79544 );
nand ( n79546 , n79542 , n425800 );
nand ( n79547 , n79537 , n79546 );
nand ( n79548 , n79494 , n79547 );
buf ( n425804 , n79548 );
buf ( n425805 , n425756 );
not ( n79551 , n425805 );
buf ( n425807 , n79491 );
nand ( n79553 , n79551 , n425807 );
buf ( n425809 , n79553 );
buf ( n425810 , n425809 );
and ( n79556 , n425804 , n425810 );
buf ( n425812 , n79556 );
buf ( n425813 , n425812 );
not ( n79559 , n425813 );
buf ( n425815 , n79559 );
buf ( n425816 , n425815 );
nand ( n79562 , n425737 , n425816 );
buf ( n425818 , n79562 );
buf ( n425819 , n425818 );
not ( n79565 , n79491 );
not ( n79566 , n425769 );
not ( n79567 , n425790 );
or ( n79568 , n79566 , n79567 );
nand ( n79569 , n79568 , n79546 );
not ( n79570 , n79569 );
not ( n79571 , n425756 );
or ( n79572 , n79570 , n79571 );
or ( n79573 , n425756 , n79547 );
nand ( n79574 , n79572 , n79573 );
or ( n79575 , n79565 , n79574 );
not ( n79576 , n79491 );
nand ( n79577 , n79576 , n79574 );
nand ( n79578 , n79575 , n79577 );
xnor ( n79579 , n425421 , n425428 );
xor ( n79580 , n425694 , n79579 );
not ( n79581 , n79580 );
xnor ( n79582 , n425236 , n425212 );
buf ( n425838 , n79582 );
buf ( n425839 , n78922 );
and ( n79585 , n425838 , n425839 );
not ( n79586 , n425838 );
buf ( n425842 , n78923 );
and ( n79588 , n79586 , n425842 );
nor ( n79589 , n79585 , n79588 );
buf ( n425845 , n79589 );
buf ( n425846 , n425845 );
xor ( n79592 , n425060 , n425187 );
xor ( n79593 , n79592 , n425208 );
buf ( n425849 , n79593 );
buf ( n425850 , n425849 );
buf ( n425851 , n59916 );
not ( n79597 , n425851 );
buf ( n425853 , n425678 );
not ( n79599 , n425853 );
or ( n79600 , n79597 , n79599 );
buf ( n425856 , n47891 );
not ( n79602 , n425856 );
buf ( n425858 , n388215 );
not ( n79604 , n425858 );
or ( n79605 , n79602 , n79604 );
buf ( n425861 , n12480 );
buf ( n425862 , n72794 );
nand ( n79608 , n425861 , n425862 );
buf ( n425864 , n79608 );
buf ( n425865 , n425864 );
nand ( n79611 , n79605 , n425865 );
buf ( n425867 , n79611 );
buf ( n425868 , n425867 );
buf ( n425869 , n50579 );
nand ( n79615 , n425868 , n425869 );
buf ( n425871 , n79615 );
buf ( n425872 , n425871 );
nand ( n79618 , n79600 , n425872 );
buf ( n425874 , n79618 );
buf ( n425875 , n425874 );
xor ( n79621 , n425850 , n425875 );
xor ( n79622 , n425126 , n425151 );
xor ( n79623 , n79622 , n425177 );
buf ( n425879 , n79623 );
buf ( n425880 , n425879 );
buf ( n425881 , n399274 );
not ( n79627 , n425881 );
buf ( n425883 , n371797 );
not ( n79629 , n425883 );
or ( n79630 , n79627 , n79629 );
buf ( n425886 , n399283 );
buf ( n425887 , n371784 );
nand ( n79633 , n425886 , n425887 );
buf ( n425889 , n79633 );
buf ( n425890 , n425889 );
nand ( n79636 , n79630 , n425890 );
buf ( n425892 , n79636 );
buf ( n425893 , n425892 );
not ( n79639 , n425893 );
buf ( n425895 , n388740 );
not ( n79641 , n425895 );
or ( n79642 , n79639 , n79641 );
buf ( n425898 , n425594 );
buf ( n425899 , n388803 );
nand ( n79645 , n425898 , n425899 );
buf ( n425901 , n79645 );
buf ( n425902 , n425901 );
nand ( n79648 , n79642 , n425902 );
buf ( n425904 , n79648 );
buf ( n425905 , n425904 );
xor ( n79651 , n425880 , n425905 );
xor ( n79652 , n77737 , n424201 );
xor ( n79653 , n79652 , n424205 );
xor ( n79654 , n78306 , n424776 );
xor ( n79655 , n79653 , n79654 );
buf ( n425911 , n79655 );
buf ( n425912 , n417572 );
not ( n79658 , n425912 );
buf ( n425914 , n422673 );
not ( n79660 , n425914 );
or ( n79661 , n79658 , n79660 );
buf ( n425917 , n394814 );
buf ( n425918 , n44775 );
nand ( n79664 , n425917 , n425918 );
buf ( n425920 , n79664 );
buf ( n425921 , n425920 );
nand ( n79667 , n79661 , n425921 );
buf ( n425923 , n79667 );
buf ( n425924 , n425923 );
not ( n79670 , n425924 );
buf ( n425926 , n44770 );
not ( n79672 , n425926 );
or ( n79673 , n79670 , n79672 );
buf ( n425929 , n424794 );
buf ( n425930 , n413643 );
nand ( n79676 , n425929 , n425930 );
buf ( n425932 , n79676 );
buf ( n425933 , n425932 );
nand ( n79679 , n79673 , n425933 );
buf ( n425935 , n79679 );
buf ( n425936 , n425935 );
xor ( n79682 , n425911 , n425936 );
buf ( n425938 , n45954 );
not ( n79684 , n425938 );
buf ( n425940 , n425511 );
not ( n79686 , n425940 );
or ( n79687 , n79684 , n79686 );
buf ( n425943 , n393369 );
not ( n79689 , n425943 );
buf ( n425945 , n392881 );
not ( n79691 , n425945 );
or ( n79692 , n79689 , n79691 );
buf ( n425948 , n424808 );
buf ( n425949 , n393381 );
nand ( n79695 , n425948 , n425949 );
buf ( n425951 , n79695 );
buf ( n425952 , n425951 );
nand ( n79698 , n79692 , n425952 );
buf ( n425954 , n79698 );
buf ( n425955 , n425954 );
buf ( n425956 , n45949 );
nand ( n79702 , n425955 , n425956 );
buf ( n425958 , n79702 );
buf ( n425959 , n425958 );
nand ( n79705 , n79687 , n425959 );
buf ( n425961 , n79705 );
buf ( n425962 , n425961 );
and ( n79708 , n79682 , n425962 );
and ( n79709 , n425911 , n425936 );
or ( n79710 , n79708 , n79709 );
buf ( n425966 , n79710 );
buf ( n425967 , n425966 );
buf ( n425968 , n55543 );
not ( n79714 , n425968 );
buf ( n425970 , n423571 );
not ( n79716 , n425970 );
or ( n79717 , n79714 , n79716 );
buf ( n425973 , n388722 );
buf ( n425974 , n51185 );
nand ( n79720 , n425973 , n425974 );
buf ( n425976 , n79720 );
buf ( n425977 , n425976 );
nand ( n79723 , n79717 , n425977 );
buf ( n425979 , n79723 );
buf ( n425980 , n425979 );
not ( n79726 , n425980 );
buf ( n425982 , n40592 );
not ( n79728 , n425982 );
or ( n79729 , n79726 , n79728 );
buf ( n425985 , n425164 );
buf ( n425986 , n388068 );
nand ( n79732 , n425985 , n425986 );
buf ( n425988 , n79732 );
buf ( n425989 , n425988 );
nand ( n79735 , n79729 , n425989 );
buf ( n425991 , n79735 );
buf ( n425992 , n425991 );
xor ( n79738 , n425967 , n425992 );
xor ( n79739 , n425494 , n425519 );
xor ( n79740 , n79739 , n425548 );
buf ( n425996 , n79740 );
buf ( n425997 , n425996 );
and ( n79743 , n79738 , n425997 );
and ( n79744 , n425967 , n425992 );
or ( n79745 , n79743 , n79744 );
buf ( n426001 , n79745 );
buf ( n426002 , n426001 );
and ( n79748 , n79651 , n426002 );
and ( n79749 , n425880 , n425905 );
or ( n79750 , n79748 , n79749 );
buf ( n426006 , n79750 );
buf ( n426007 , n426006 );
buf ( n426008 , n400033 );
not ( n79754 , n426008 );
buf ( n426010 , n62006 );
not ( n79756 , n426010 );
or ( n79757 , n79754 , n79756 );
buf ( n426013 , n24116 );
buf ( n426014 , n400042 );
nand ( n79760 , n426013 , n426014 );
buf ( n426016 , n79760 );
buf ( n426017 , n426016 );
nand ( n79763 , n79757 , n426017 );
buf ( n426019 , n79763 );
buf ( n426020 , n426019 );
not ( n79766 , n426020 );
buf ( n426022 , n73026 );
not ( n79768 , n426022 );
or ( n79769 , n79766 , n79768 );
buf ( n426025 , n425197 );
not ( n79771 , n426025 );
buf ( n426027 , n41664 );
nand ( n79773 , n79771 , n426027 );
buf ( n426029 , n79773 );
buf ( n426030 , n426029 );
nand ( n79776 , n79769 , n426030 );
buf ( n426032 , n79776 );
buf ( n426033 , n426032 );
xor ( n79779 , n426007 , n426033 );
xor ( n79780 , n425586 , n425607 );
xor ( n79781 , n79780 , n425622 );
buf ( n426037 , n79781 );
buf ( n426038 , n426037 );
and ( n79784 , n79779 , n426038 );
and ( n79785 , n426007 , n426033 );
or ( n79786 , n79784 , n79785 );
buf ( n426042 , n79786 );
buf ( n426043 , n426042 );
and ( n79789 , n79621 , n426043 );
and ( n79790 , n425850 , n425875 );
or ( n79791 , n79789 , n79790 );
buf ( n426047 , n79791 );
buf ( n426048 , n426047 );
buf ( n426049 , C0 );
buf ( n426050 , n426049 );
and ( n79821 , n425846 , n426048 );
or ( n79822 , C0 , n79821 );
buf ( n426053 , n79822 );
not ( n79824 , n426053 );
not ( n79825 , n79824 );
not ( n79826 , n79825 );
xor ( n79827 , n425275 , n425333 );
xor ( n79828 , n79827 , n425338 );
buf ( n426059 , n79828 );
buf ( n426060 , n426059 );
xnor ( n79831 , n425305 , n425318 );
buf ( n426062 , n79831 );
buf ( n426063 , n425325 );
and ( n79834 , n426062 , n426063 );
not ( n79835 , n426062 );
buf ( n426066 , n425312 );
and ( n79837 , n79835 , n426066 );
nor ( n79838 , n79834 , n79837 );
buf ( n426069 , n79838 );
buf ( n426070 , n426069 );
buf ( n426071 , C0 );
buf ( n426072 , n426071 );
xor ( n79862 , n426070 , n426072 );
buf ( n426074 , n358975 );
not ( n79864 , n426074 );
buf ( n426076 , n41330 );
nor ( n79866 , n79864 , n426076 );
buf ( n426078 , n79866 );
buf ( n426079 , n426078 );
buf ( n426080 , n397489 );
not ( n79870 , n426080 );
buf ( n426082 , n371876 );
not ( n79872 , n426082 );
or ( n79873 , n79870 , n79872 );
buf ( n426085 , n388064 );
buf ( n426086 , n397486 );
nand ( n79876 , n426085 , n426086 );
buf ( n426088 , n79876 );
buf ( n426089 , n426088 );
nand ( n79879 , n79873 , n426089 );
buf ( n426091 , n79879 );
buf ( n426092 , n426091 );
not ( n79882 , n426092 );
buf ( n426094 , n74375 );
not ( n79884 , n426094 );
or ( n79885 , n79882 , n79884 );
buf ( n426097 , n43515 );
buf ( n426098 , n425535 );
nand ( n79888 , n426097 , n426098 );
buf ( n426100 , n79888 );
buf ( n426101 , n426100 );
nand ( n79891 , n79885 , n426101 );
buf ( n426103 , n79891 );
buf ( n426104 , n426103 );
xor ( n79894 , n424101 , n424117 );
xor ( n79895 , n79894 , n424144 );
xor ( n79896 , n424604 , n424626 );
xor ( n79897 , n79895 , n79896 );
buf ( n426109 , n79897 );
not ( n79899 , n68043 );
not ( n79900 , n78283 );
or ( n79901 , n79899 , n79900 );
not ( n79902 , n410635 );
not ( n79903 , n63629 );
not ( n79904 , n416830 );
or ( n79905 , n79903 , n79904 );
nand ( n79906 , n63625 , n70195 );
nand ( n79907 , n79905 , n79906 );
nand ( n79908 , n79902 , n79907 );
nand ( n79909 , n79901 , n79908 );
buf ( n426121 , n403133 );
buf ( n426122 , n422315 );
nor ( n79912 , n426121 , n426122 );
buf ( n426124 , n79912 );
buf ( n426125 , n426124 );
buf ( n426126 , n59637 );
buf ( n426127 , n14083 );
buf ( n426128 , n71664 );
and ( n79918 , n426127 , n426128 );
buf ( n426130 , n59457 );
buf ( n426131 , n418298 );
and ( n79921 , n426130 , n426131 );
nor ( n79922 , n79918 , n79921 );
buf ( n426134 , n79922 );
buf ( n426135 , n426134 );
or ( n79925 , n426126 , n426135 );
buf ( n426137 , n424673 );
buf ( n426138 , n59467 );
or ( n79928 , n426137 , n426138 );
nand ( n79929 , n79925 , n79928 );
buf ( n426141 , n79929 );
buf ( n426142 , n426141 );
and ( n79932 , n426125 , n426142 );
buf ( n426144 , n79932 );
buf ( n426145 , n405407 );
buf ( n426146 , n405391 );
buf ( n426147 , n71681 );
and ( n79937 , n426146 , n426147 );
buf ( n426149 , n405388 );
buf ( n426150 , n418315 );
and ( n79940 , n426149 , n426150 );
nor ( n79941 , n79937 , n79940 );
buf ( n426153 , n79941 );
buf ( n426154 , n426153 );
or ( n79944 , n426145 , n426154 );
buf ( n426156 , n424131 );
not ( n79946 , n426156 );
buf ( n426158 , n79946 );
buf ( n426159 , n426158 );
buf ( n426160 , n405378 );
or ( n79950 , n426159 , n426160 );
nand ( n79951 , n79944 , n79950 );
buf ( n426163 , n79951 );
xor ( n79953 , n426144 , n426163 );
buf ( n426165 , n403128 );
buf ( n426166 , n623 );
or ( n79956 , n426165 , n426166 );
buf ( n426168 , n403123 );
buf ( n426169 , n55905 );
buf ( n426170 , n623 );
and ( n79960 , n426168 , n426169 , n426170 );
buf ( n426172 , n403138 );
nor ( n79962 , n79960 , n426172 );
buf ( n426174 , n79962 );
buf ( n426175 , n426174 );
nand ( n79965 , n79956 , n426175 );
buf ( n426177 , n79965 );
and ( n79967 , n79953 , n426177 );
and ( n79968 , n426144 , n426163 );
or ( n79969 , n79967 , n79968 );
xor ( n79970 , n79909 , n79969 );
xor ( n79971 , n424490 , n424507 );
xor ( n79972 , n79971 , n424530 );
buf ( n426184 , n79972 );
and ( n79974 , n79970 , n426184 );
and ( n79975 , n79909 , n79969 );
or ( n79976 , n79974 , n79975 );
buf ( n426188 , n79976 );
xor ( n79978 , n426109 , n426188 );
buf ( n426190 , n71095 );
buf ( n426191 , n59463 );
and ( n79981 , n426190 , n426191 );
buf ( n426193 , n417729 );
buf ( n426194 , n62159 );
and ( n79984 , n426193 , n426194 );
nor ( n79985 , n79981 , n79984 );
buf ( n426197 , n79985 );
buf ( n426198 , n426197 );
buf ( n426199 , n409429 );
or ( n79989 , n426198 , n426199 );
buf ( n426201 , n424728 );
not ( n79991 , n426201 );
buf ( n426203 , n79991 );
buf ( n426204 , n426203 );
buf ( n426205 , n409170 );
or ( n79995 , n426204 , n426205 );
nand ( n79996 , n79989 , n79995 );
buf ( n426208 , n79996 );
xor ( n79998 , n424680 , n424693 );
xor ( n79999 , n79998 , n424710 );
and ( n80000 , n426208 , n79999 );
buf ( n426212 , n71088 );
buf ( n426213 , n62177 );
and ( n80003 , n426212 , n426213 );
buf ( n426215 , n417722 );
buf ( n426216 , n409178 );
and ( n80006 , n426215 , n426216 );
nor ( n80007 , n80003 , n80006 );
buf ( n426219 , n80007 );
buf ( n426220 , n426219 );
buf ( n426221 , n409429 );
or ( n80011 , n426220 , n426221 );
buf ( n426223 , n426197 );
buf ( n426224 , n409170 );
or ( n80014 , n426223 , n426224 );
nand ( n80015 , n80011 , n80014 );
buf ( n426227 , n80015 );
buf ( n426228 , n426227 );
buf ( n426229 , n405391 );
buf ( n426230 , n72308 );
and ( n80020 , n426229 , n426230 );
buf ( n426232 , n405388 );
buf ( n426233 , n418942 );
and ( n80023 , n426232 , n426233 );
nor ( n80024 , n80020 , n80023 );
buf ( n426236 , n80024 );
buf ( n426237 , n426236 );
buf ( n426238 , n405407 );
or ( n80028 , n426237 , n426238 );
buf ( n426240 , n426153 );
buf ( n426241 , n405378 );
or ( n80031 , n426240 , n426241 );
nand ( n80032 , n80028 , n80031 );
buf ( n426244 , n80032 );
buf ( n426245 , n426244 );
xor ( n80035 , n426228 , n426245 );
buf ( n426247 , n424703 );
buf ( n426248 , n405476 );
or ( n80038 , n426247 , n426248 );
buf ( n426250 , n403301 );
nand ( n80040 , n80038 , n426250 );
buf ( n426252 , n80040 );
buf ( n426253 , n426252 );
and ( n80043 , n80035 , n426253 );
and ( n80044 , n426228 , n426245 );
or ( n80045 , n80043 , n80044 );
buf ( n426257 , n80045 );
xor ( n80047 , n424680 , n424693 );
xor ( n80048 , n80047 , n424710 );
and ( n426260 , n426257 , n80048 );
and ( n426261 , n426208 , n426257 );
or ( n80051 , n80000 , n426260 , n426261 );
buf ( n426263 , n80051 );
buf ( n426264 , n67987 );
buf ( n426265 , n66411 );
and ( n426266 , n426264 , n426265 );
buf ( n426267 , n414714 );
buf ( n426268 , n62496 );
and ( n426269 , n426267 , n426268 );
nor ( n426270 , n426266 , n426269 );
buf ( n426271 , n426270 );
buf ( n426272 , n426271 );
buf ( n426273 , n410724 );
or ( n80063 , n426272 , n426273 );
buf ( n426275 , n424655 );
buf ( n426276 , n410721 );
or ( n80066 , n426275 , n426276 );
nand ( n426278 , n80063 , n80066 );
buf ( n426279 , n426278 );
buf ( n426280 , n426279 );
xor ( n426281 , n426263 , n426280 );
xor ( n426282 , n424714 , n424717 );
xor ( n80072 , n426282 , n424737 );
buf ( n426284 , n80072 );
buf ( n426285 , n426284 );
and ( n80075 , n426281 , n426285 );
and ( n426287 , n426263 , n426280 );
or ( n426288 , n80075 , n426287 );
buf ( n426289 , n426288 );
buf ( n426290 , n426289 );
and ( n426291 , n79978 , n426290 );
and ( n80081 , n426109 , n426188 );
or ( n426293 , n426291 , n80081 );
buf ( n426294 , n426293 );
xor ( n80084 , n424647 , n424752 );
xor ( n426296 , n80084 , n78422 );
and ( n426297 , n426294 , n426296 );
buf ( n426298 , n70210 );
buf ( n426299 , n63625 );
and ( n426300 , n426298 , n426299 );
buf ( n426301 , n416845 );
buf ( n426302 , n63629 );
and ( n426303 , n426301 , n426302 );
nor ( n80093 , n426300 , n426303 );
buf ( n426305 , n80093 );
or ( n426306 , n426305 , n410635 );
nand ( n80096 , n79907 , n68043 );
nand ( n426308 , n426306 , n80096 );
xor ( n426309 , n426144 , n426163 );
xor ( n80099 , n426309 , n426177 );
and ( n80100 , n426308 , n80099 );
buf ( n426312 , n68002 );
buf ( n426313 , n66411 );
and ( n80103 , n426312 , n426313 );
buf ( n426315 , n414729 );
buf ( n426316 , n62496 );
and ( n80106 , n426315 , n426316 );
nor ( n80107 , n80103 , n80106 );
buf ( n426319 , n80107 );
buf ( n426320 , n426319 );
buf ( n426321 , n410724 );
or ( n80111 , n426320 , n426321 );
buf ( n426323 , n426271 );
buf ( n426324 , n410721 );
or ( n80114 , n426323 , n426324 );
nand ( n80115 , n80111 , n80114 );
buf ( n426327 , n80115 );
xor ( n80117 , n426144 , n426163 );
xor ( n80118 , n80117 , n426177 );
and ( n80119 , n426327 , n80118 );
and ( n80120 , n426308 , n426327 );
or ( n80121 , n80100 , n80119 , n80120 );
xor ( n80122 , n79909 , n79969 );
xor ( n80123 , n80122 , n426184 );
and ( n80124 , n80121 , n80123 );
xor ( n80125 , n426263 , n426280 );
xor ( n80126 , n80125 , n426285 );
buf ( n426338 , n80126 );
xor ( n80128 , n79909 , n79969 );
xor ( n80129 , n80128 , n426184 );
and ( n80130 , n426338 , n80129 );
and ( n80131 , n80121 , n426338 );
or ( n80132 , n80124 , n80130 , n80131 );
buf ( n426344 , n80132 );
xor ( n80134 , n424664 , n424742 );
xor ( n80135 , n80134 , n424748 );
buf ( n426347 , n80135 );
buf ( n426348 , n426347 );
xor ( n80138 , n426344 , n426348 );
xor ( n80139 , n426109 , n426188 );
xor ( n80140 , n80139 , n426290 );
buf ( n426352 , n80140 );
buf ( n426353 , n426352 );
and ( n80143 , n80138 , n426353 );
and ( n80144 , n426344 , n426348 );
or ( n426356 , n80143 , n80144 );
buf ( n426357 , n426356 );
xor ( n80147 , n424647 , n424752 );
xor ( n80148 , n80147 , n78422 );
and ( n80149 , n426357 , n80148 );
and ( n426361 , n426294 , n426357 );
or ( n426362 , n426297 , n80149 , n426361 );
buf ( n426363 , n426362 );
xor ( n80153 , n424761 , n424766 );
xor ( n80154 , n80153 , n424772 );
buf ( n426366 , n80154 );
buf ( n426367 , n426366 );
xor ( n80157 , n426363 , n426367 );
not ( n80158 , n49116 );
not ( n426370 , n80158 );
not ( n426371 , n422673 );
or ( n80161 , n426370 , n426371 );
buf ( n426373 , n390988 );
buf ( n426374 , n80158 );
not ( n80164 , n426374 );
buf ( n426376 , n80164 );
buf ( n426377 , n426376 );
nand ( n80167 , n426373 , n426377 );
buf ( n426379 , n80167 );
nand ( n80169 , n80161 , n426379 );
not ( n80170 , n80169 );
not ( n80171 , n44770 );
or ( n80172 , n80170 , n80171 );
buf ( n426384 , n392740 );
buf ( n426385 , n425923 );
nand ( n80175 , n426384 , n426385 );
buf ( n426387 , n80175 );
nand ( n80177 , n80172 , n426387 );
buf ( n426389 , n80177 );
and ( n426390 , n80157 , n426389 );
and ( n80180 , n426363 , n426367 );
or ( n80181 , n426390 , n80180 );
buf ( n426393 , n80181 );
buf ( n426394 , n426393 );
or ( n426395 , n426104 , n426394 );
xor ( n80185 , n425911 , n425936 );
xor ( n80186 , n80185 , n425962 );
buf ( n426398 , n80186 );
buf ( n426399 , n426398 );
nand ( n80189 , n426395 , n426399 );
buf ( n426401 , n80189 );
buf ( n426402 , n426401 );
buf ( n426403 , n426103 );
buf ( n426404 , n426393 );
nand ( n80194 , n426403 , n426404 );
buf ( n426406 , n80194 );
buf ( n426407 , n426406 );
nand ( n80197 , n426402 , n426407 );
buf ( n426409 , n80197 );
buf ( n426410 , n426409 );
buf ( n426411 , n395359 );
not ( n80201 , n426411 );
buf ( n426413 , n425566 );
not ( n80203 , n426413 );
or ( n80204 , n80201 , n80203 );
buf ( n426416 , n395346 );
buf ( n426417 , n47863 );
not ( n80207 , n426417 );
buf ( n426419 , n420954 );
not ( n80209 , n426419 );
or ( n426421 , n80207 , n80209 );
buf ( n426422 , n389338 );
buf ( n426423 , n419385 );
nand ( n80213 , n426422 , n426423 );
buf ( n426425 , n80213 );
buf ( n426426 , n426425 );
nand ( n80216 , n426421 , n426426 );
buf ( n426428 , n80216 );
buf ( n426429 , n426428 );
nand ( n80219 , n426416 , n426429 );
buf ( n426431 , n80219 );
buf ( n426432 , n426431 );
nand ( n80222 , n80204 , n426432 );
buf ( n426434 , n80222 );
buf ( n426435 , n426434 );
xor ( n80225 , n426410 , n426435 );
buf ( n426437 , n24116 );
not ( n80227 , n426437 );
not ( n80228 , n371751 );
not ( n80229 , n417617 );
or ( n80230 , n80228 , n80229 );
buf ( n426442 , n371751 );
buf ( n426443 , n417617 );
nor ( n80233 , n426442 , n426443 );
buf ( n426445 , n80233 );
or ( n80235 , n426445 , n402819 );
nand ( n80236 , n80230 , n80235 );
buf ( n426448 , n80236 );
nor ( n80238 , n80227 , n426448 );
buf ( n426450 , n80238 );
buf ( n426451 , n426450 );
and ( n80241 , n80225 , n426451 );
and ( n426453 , n426410 , n426435 );
or ( n426454 , n80241 , n426453 );
buf ( n426455 , n426454 );
buf ( n426456 , n426455 );
xor ( n80246 , n426079 , n426456 );
xor ( n80247 , n79218 , n425552 );
xor ( n80248 , n80247 , n425573 );
buf ( n426460 , n80248 );
and ( n80250 , n80246 , n426460 );
and ( n80251 , n426079 , n426456 );
or ( n80252 , n80250 , n80251 );
buf ( n426464 , n80252 );
buf ( n426465 , n426464 );
buf ( n426466 , n358975 );
buf ( n426467 , n41365 );
and ( n80257 , n426466 , n426467 );
not ( n426469 , n426466 );
buf ( n426470 , n410407 );
and ( n80260 , n426469 , n426470 );
nor ( n80261 , n80257 , n80260 );
buf ( n426473 , n80261 );
buf ( n426474 , n426473 );
not ( n80264 , n426474 );
buf ( n426476 , n66128 );
not ( n80266 , n426476 );
or ( n80267 , n80264 , n80266 );
buf ( n426479 , n425641 );
buf ( n426480 , n388830 );
nand ( n80270 , n426479 , n426480 );
buf ( n426482 , n80270 );
buf ( n426483 , n426482 );
nand ( n80273 , n80267 , n426483 );
buf ( n426485 , n80273 );
buf ( n426486 , n426485 );
xor ( n80276 , n426465 , n426486 );
buf ( n426488 , n59916 );
not ( n80278 , n426488 );
buf ( n426490 , n425867 );
not ( n80280 , n426490 );
or ( n80281 , n80278 , n80280 );
and ( n80282 , n47891 , n417349 );
not ( n80283 , n47891 );
and ( n80284 , n80283 , n28353 );
or ( n80285 , n80282 , n80284 );
buf ( n426497 , n80285 );
buf ( n426498 , n50579 );
nand ( n80288 , n426497 , n426498 );
buf ( n426500 , n80288 );
buf ( n426501 , n426500 );
nand ( n80291 , n80281 , n426501 );
buf ( n426503 , n80291 );
buf ( n426504 , n426503 );
and ( n80294 , n80276 , n426504 );
and ( n80295 , n426465 , n426486 );
or ( n80296 , n80294 , n80295 );
buf ( n426508 , n80296 );
buf ( n426509 , n426508 );
and ( n80299 , n79862 , n426509 );
or ( n80301 , n80299 , C0 );
buf ( n426512 , n80301 );
buf ( n426513 , n426512 );
buf ( n426514 , C0 );
buf ( n426515 , n426514 );
and ( n80326 , n426060 , n426513 );
or ( n80327 , C0 , n80326 );
buf ( n426518 , n80327 );
not ( n426519 , n426518 );
or ( n80330 , n79826 , n426519 );
not ( n80331 , n79824 );
not ( n80332 , n426518 );
not ( n426523 , n80332 );
or ( n426524 , n80331 , n426523 );
xor ( n80335 , n425436 , n425438 );
xor ( n80336 , n80335 , n425691 );
buf ( n426527 , n80336 );
nand ( n80338 , n426524 , n426527 );
nand ( n80339 , n80330 , n80338 );
nor ( n80340 , n79581 , n80339 );
and ( n80341 , n425800 , n79538 );
not ( n80342 , n425800 );
and ( n80343 , n80342 , n425769 );
or ( n80344 , n80341 , n80343 );
buf ( n80345 , n425790 );
not ( n426536 , n80345 );
and ( n426537 , n80344 , n426536 );
not ( n80348 , n80344 );
and ( n80349 , n80348 , n80345 );
nor ( n80350 , n426537 , n80349 );
or ( n426541 , n80340 , n80350 );
not ( n426542 , n79580 );
nand ( n80353 , n426542 , n80339 );
nand ( n80354 , n426541 , n80353 );
nand ( n80355 , n79578 , n80354 );
buf ( n426546 , n80355 );
not ( n80357 , n426546 );
buf ( n426548 , n79464 );
buf ( n426549 , n425812 );
nand ( n80360 , n426548 , n426549 );
buf ( n426551 , n80360 );
buf ( n426552 , n426551 );
nand ( n80363 , n80357 , n426552 );
buf ( n426554 , n80363 );
buf ( n426555 , n426554 );
nand ( n80366 , n425819 , n426555 );
buf ( n426557 , n80366 );
not ( n80368 , n426557 );
or ( n80369 , n79462 , n80368 );
buf ( n426560 , n425419 );
not ( n80371 , n426560 );
buf ( n426562 , n80371 );
buf ( n426563 , n426562 );
buf ( n426564 , n79458 );
not ( n80375 , n426564 );
buf ( n426566 , n80375 );
buf ( n426567 , n426566 );
nand ( n80378 , n426563 , n426567 );
buf ( n426569 , n80378 );
nand ( n80380 , n80369 , n426569 );
buf ( n426571 , n79066 );
buf ( n426572 , n426571 );
not ( n80383 , n426572 );
buf ( n426574 , n425382 );
not ( n80385 , n426574 );
or ( n80386 , n80383 , n80385 );
buf ( n426577 , n425382 );
buf ( n426578 , n426571 );
or ( n80389 , n426577 , n426578 );
buf ( n426580 , n425413 );
nand ( n80391 , n80389 , n426580 );
buf ( n426582 , n80391 );
buf ( n426583 , n426582 );
nand ( n80394 , n80386 , n426583 );
buf ( n426585 , n80394 );
xor ( n80396 , n422773 , n422865 );
xor ( n80397 , n80396 , n422869 );
buf ( n426588 , n80397 );
buf ( n426589 , n426588 );
not ( n80400 , n426589 );
buf ( n426591 , n80400 );
and ( n80402 , n426585 , n426591 );
not ( n80403 , n426585 );
and ( n80404 , n80403 , n426588 );
or ( n80405 , n80402 , n80404 );
buf ( n426596 , n80405 );
xor ( n80407 , n421805 , n421915 );
xor ( n80408 , n80407 , n421917 );
buf ( n426599 , n80408 );
buf ( n426600 , n426599 );
xor ( n80411 , n421603 , n421605 );
xor ( n80412 , n80411 , n421610 );
buf ( n426603 , n80412 );
buf ( n426604 , n426603 );
xor ( n80415 , n426600 , n426604 );
buf ( n426606 , n423435 );
not ( n80417 , n426606 );
buf ( n426608 , n424311 );
not ( n80419 , n426608 );
or ( n80420 , n80417 , n80419 );
buf ( n426611 , n423441 );
not ( n80422 , n426611 );
buf ( n426613 , n424314 );
not ( n80424 , n426613 );
or ( n80425 , n80422 , n80424 );
buf ( n426616 , n423431 );
nand ( n80427 , n80425 , n426616 );
buf ( n426618 , n80427 );
buf ( n426619 , n426618 );
nand ( n80430 , n80420 , n426619 );
buf ( n426621 , n80430 );
buf ( n426622 , n426621 );
xor ( n80433 , n80415 , n426622 );
buf ( n426624 , n80433 );
buf ( n426625 , n426624 );
not ( n80436 , n426625 );
buf ( n426627 , n80436 );
buf ( n426628 , n426627 );
and ( n80439 , n426596 , n426628 );
not ( n80440 , n426596 );
buf ( n426631 , n426624 );
and ( n80442 , n80440 , n426631 );
nor ( n80443 , n80439 , n80442 );
buf ( n426634 , n80443 );
xor ( n80445 , n424322 , n425375 );
and ( n80446 , n80445 , n425417 );
and ( n80447 , n424322 , n425375 );
or ( n80448 , n80446 , n80447 );
buf ( n426639 , n80448 );
nand ( n80450 , n426634 , n426639 );
nand ( n80451 , n80380 , n80450 );
buf ( n426642 , n426551 );
not ( n426643 , n426642 );
nor ( n80454 , n79578 , n80354 );
buf ( n426645 , n80454 );
nor ( n80456 , n426643 , n426645 );
buf ( n426647 , n80456 );
and ( n426648 , n426647 , n425730 );
xor ( n80459 , n425774 , n425785 );
xor ( n80460 , n80459 , n425787 );
buf ( n426651 , n80460 );
not ( n80462 , n426651 );
xor ( n80463 , n425456 , n425660 );
xor ( n80464 , n80463 , n425686 );
buf ( n426655 , n80464 );
buf ( n426656 , n426655 );
xor ( n80467 , n425582 , n425627 );
xor ( n80468 , n80467 , n425655 );
buf ( n426659 , n80468 );
buf ( n426660 , n426659 );
xor ( n426661 , n425481 , n425485 );
xor ( n80472 , n426661 , n425577 );
buf ( n426663 , n80472 );
buf ( n426664 , n426663 );
buf ( n426665 , n55055 );
not ( n80476 , n426665 );
buf ( n426667 , n62006 );
not ( n80478 , n426667 );
or ( n80479 , n80476 , n80478 );
buf ( n426670 , n24116 );
buf ( n426671 , n55054 );
nand ( n80482 , n426670 , n426671 );
buf ( n426673 , n80482 );
buf ( n426674 , n426673 );
nand ( n80485 , n80479 , n426674 );
buf ( n426676 , n80485 );
buf ( n426677 , n426676 );
not ( n80488 , n426677 );
buf ( n426679 , n73026 );
not ( n80490 , n426679 );
or ( n80491 , n80488 , n80490 );
buf ( n426682 , n426019 );
buf ( n426683 , n41664 );
nand ( n80494 , n426682 , n426683 );
buf ( n426685 , n80494 );
buf ( n426686 , n426685 );
nand ( n80497 , n80491 , n426686 );
buf ( n426688 , n80497 );
buf ( n426689 , n426688 );
buf ( n426690 , n59916 );
not ( n80501 , n426690 );
buf ( n426692 , n80285 );
not ( n80503 , n426692 );
or ( n80504 , n80501 , n80503 );
and ( n80505 , n27320 , n403668 );
not ( n80506 , n27320 );
and ( n80507 , n80506 , n47891 );
or ( n80508 , n80505 , n80507 );
buf ( n426699 , n80508 );
buf ( n426700 , n50579 );
nand ( n80511 , n426699 , n426700 );
buf ( n426702 , n80511 );
buf ( n426703 , n426702 );
nand ( n80514 , n80504 , n426703 );
buf ( n426705 , n80514 );
buf ( n426706 , n426705 );
xor ( n80517 , n426689 , n426706 );
buf ( n426708 , n400033 );
buf ( n426709 , n417617 );
and ( n80520 , n426708 , n426709 );
not ( n80521 , n426708 );
buf ( n426712 , n388751 );
and ( n80523 , n80521 , n426712 );
nor ( n426714 , n80520 , n80523 );
buf ( n426715 , n426714 );
buf ( n426716 , n426715 );
not ( n80527 , n426716 );
buf ( n426718 , n388740 );
not ( n80529 , n426718 );
or ( n80530 , n80527 , n80529 );
buf ( n426721 , n425892 );
buf ( n426722 , n388803 );
nand ( n80533 , n426721 , n426722 );
buf ( n426724 , n80533 );
buf ( n426725 , n426724 );
nand ( n80536 , n80530 , n426725 );
buf ( n426727 , n80536 );
buf ( n426728 , n426727 );
buf ( n426729 , n395359 );
not ( n80540 , n426729 );
buf ( n426731 , n426428 );
not ( n80542 , n426731 );
or ( n80543 , n80540 , n80542 );
buf ( n426734 , n47863 );
not ( n80545 , n426734 );
buf ( n426736 , n391440 );
not ( n80547 , n426736 );
or ( n80548 , n80545 , n80547 );
buf ( n426739 , n419385 );
buf ( n426740 , n420994 );
nand ( n80551 , n426739 , n426740 );
buf ( n426742 , n80551 );
buf ( n426743 , n426742 );
nand ( n80554 , n80548 , n426743 );
buf ( n426745 , n80554 );
buf ( n426746 , n426745 );
buf ( n426747 , n395346 );
nand ( n80558 , n426746 , n426747 );
buf ( n426749 , n80558 );
buf ( n426750 , n426749 );
nand ( n80561 , n80543 , n426750 );
buf ( n426752 , n80561 );
buf ( n426753 , n426752 );
buf ( n426754 , n45954 );
not ( n80565 , n426754 );
buf ( n426756 , n425954 );
not ( n426757 , n426756 );
or ( n426758 , n80565 , n426757 );
and ( n80569 , n394207 , n392217 );
not ( n80570 , n394207 );
buf ( n426761 , n392217 );
not ( n426762 , n426761 );
buf ( n426763 , n426762 );
and ( n80574 , n80570 , n426763 );
or ( n80575 , n80569 , n80574 );
nand ( n80576 , n80575 , n45949 );
buf ( n426767 , n80576 );
nand ( n80578 , n426758 , n426767 );
buf ( n426769 , n80578 );
buf ( n426770 , n426769 );
xor ( n80581 , n424647 , n424752 );
xor ( n80582 , n80581 , n78422 );
xor ( n80583 , n426294 , n426357 );
xor ( n80584 , n80582 , n80583 );
not ( n426775 , n45947 );
not ( n426776 , n426775 );
not ( n80587 , n80575 );
or ( n80588 , n426776 , n80587 );
and ( n80589 , n394814 , n392217 );
not ( n80590 , n394814 );
and ( n80591 , n80590 , n426763 );
or ( n80592 , n80589 , n80591 );
nand ( n80593 , n80592 , n45949 );
nand ( n80594 , n80588 , n80593 );
xor ( n80595 , n80584 , n80594 );
xor ( n80596 , n79909 , n79969 );
xor ( n80597 , n80596 , n426184 );
xor ( n80598 , n80121 , n426338 );
xor ( n80599 , n80597 , n80598 );
buf ( n426790 , n80599 );
xor ( n80601 , n424680 , n424693 );
xor ( n80602 , n80601 , n424710 );
xor ( n80603 , n426208 , n426257 );
xor ( n80604 , n80602 , n80603 );
buf ( n426795 , n80604 );
buf ( n426796 , n59637 );
buf ( n426797 , n14083 );
buf ( n426798 , n71681 );
and ( n80609 , n426797 , n426798 );
buf ( n426800 , n59457 );
buf ( n426801 , n418315 );
and ( n80612 , n426800 , n426801 );
nor ( n80613 , n80609 , n80612 );
buf ( n426804 , n80613 );
buf ( n426805 , n426804 );
or ( n426806 , n426796 , n426805 );
buf ( n426807 , n426134 );
buf ( n426808 , n59467 );
or ( n80619 , n426807 , n426808 );
nand ( n80620 , n426806 , n80619 );
buf ( n426811 , n80620 );
buf ( n426812 , n56045 );
buf ( n426813 , n623 );
and ( n80624 , n426812 , n426813 );
not ( n80625 , n56045 );
buf ( n426816 , n80625 );
buf ( n426817 , n422315 );
and ( n80628 , n426816 , n426817 );
buf ( n426819 , n405391 );
nor ( n80630 , n80628 , n426819 );
buf ( n426821 , n80630 );
buf ( n426822 , n426821 );
buf ( n426823 , n56041 );
nor ( n80634 , n80624 , n426822 , n426823 );
buf ( n426825 , n80634 );
xor ( n80636 , n426811 , n426825 );
buf ( n426827 , n405407 );
buf ( n426828 , n405391 );
buf ( n426829 , n74002 );
and ( n80640 , n426828 , n426829 );
buf ( n426831 , n405388 );
buf ( n426832 , n420612 );
and ( n80643 , n426831 , n426832 );
nor ( n80644 , n80640 , n80643 );
buf ( n426835 , n80644 );
buf ( n426836 , n426835 );
or ( n80647 , n426827 , n426836 );
buf ( n426838 , n426236 );
buf ( n426839 , n405378 );
or ( n80650 , n426838 , n426839 );
nand ( n80651 , n80647 , n80650 );
buf ( n426842 , n80651 );
and ( n80653 , n80636 , n426842 );
and ( n80654 , n426811 , n426825 );
or ( n80655 , n80653 , n80654 );
buf ( n426846 , n80655 );
xor ( n80657 , n426125 , n426142 );
buf ( n426848 , n80657 );
buf ( n426849 , n426848 );
xor ( n80660 , n426846 , n426849 );
buf ( n426851 , n70389 );
buf ( n426852 , n63625 );
and ( n80663 , n426851 , n426852 );
buf ( n426854 , n417024 );
buf ( n426855 , n62511 );
and ( n80666 , n426854 , n426855 );
nor ( n80667 , n80663 , n80666 );
buf ( n426858 , n80667 );
buf ( n426859 , n426858 );
buf ( n426860 , n410635 );
or ( n80671 , n426859 , n426860 );
buf ( n426862 , n426305 );
buf ( n426863 , n409504 );
or ( n426864 , n426862 , n426863 );
nand ( n426865 , n80671 , n426864 );
buf ( n426866 , n426865 );
buf ( n426867 , n426866 );
and ( n80678 , n80660 , n426867 );
and ( n426869 , n426846 , n426849 );
or ( n426870 , n80678 , n426869 );
buf ( n426871 , n426870 );
buf ( n426872 , n426871 );
xor ( n80683 , n426795 , n426872 );
xor ( n80684 , n426228 , n426245 );
xor ( n80685 , n80684 , n426253 );
buf ( n426876 , n80685 );
buf ( n426877 , n426876 );
buf ( n426878 , n405476 );
buf ( n426879 , n422315 );
nor ( n80690 , n426878 , n426879 );
buf ( n426881 , n80690 );
buf ( n426882 , n426881 );
buf ( n426883 , n59637 );
buf ( n426884 , n14083 );
buf ( n426885 , n72308 );
and ( n80696 , n426884 , n426885 );
buf ( n426887 , n59457 );
buf ( n426888 , n418942 );
and ( n80699 , n426887 , n426888 );
nor ( n80700 , n80696 , n80699 );
buf ( n426891 , n80700 );
buf ( n426892 , n426891 );
or ( n80703 , n426883 , n426892 );
buf ( n426894 , n426804 );
buf ( n426895 , n59467 );
or ( n80706 , n426894 , n426895 );
nand ( n80707 , n80703 , n80706 );
buf ( n426898 , n80707 );
buf ( n426899 , n426898 );
and ( n80710 , n426882 , n426899 );
buf ( n426901 , n80710 );
buf ( n426902 , n409429 );
buf ( n426903 , n71170 );
buf ( n426904 , n59463 );
and ( n80715 , n426903 , n426904 );
buf ( n426906 , n417804 );
buf ( n426907 , n409178 );
and ( n80718 , n426906 , n426907 );
nor ( n80719 , n80715 , n80718 );
buf ( n426910 , n80719 );
buf ( n426911 , n426910 );
or ( n80722 , n426902 , n426911 );
buf ( n426913 , n426219 );
buf ( n426914 , n409170 );
or ( n80725 , n426913 , n426914 );
nand ( n80726 , n80722 , n80725 );
buf ( n426917 , n80726 );
xor ( n80728 , n426901 , n426917 );
buf ( n426919 , n403301 );
buf ( n426920 , n623 );
or ( n80731 , n426919 , n426920 );
and ( n80732 , n56064 , n56041 , n623 );
not ( n80733 , n403309 );
nor ( n80734 , n80732 , n80733 );
buf ( n426925 , n80734 );
nand ( n80736 , n80731 , n426925 );
buf ( n426927 , n80736 );
and ( n80738 , n80728 , n426927 );
and ( n80739 , n426901 , n426917 );
or ( n80740 , n80738 , n80739 );
buf ( n426931 , n80740 );
xor ( n80742 , n426877 , n426931 );
buf ( n426933 , n70195 );
buf ( n426934 , n66411 );
and ( n80745 , n426933 , n426934 );
buf ( n426936 , n416830 );
buf ( n426937 , n62496 );
and ( n80748 , n426936 , n426937 );
nor ( n80749 , n80745 , n80748 );
buf ( n426940 , n80749 );
buf ( n426941 , n426940 );
buf ( n426942 , n410724 );
or ( n80753 , n426941 , n426942 );
buf ( n426944 , n426319 );
buf ( n426945 , n410721 );
or ( n80756 , n426944 , n426945 );
nand ( n80757 , n80753 , n80756 );
buf ( n426948 , n80757 );
buf ( n426949 , n426948 );
and ( n80760 , n80742 , n426949 );
and ( n80761 , n426877 , n426931 );
or ( n80762 , n80760 , n80761 );
buf ( n426953 , n80762 );
buf ( n426954 , n426953 );
and ( n80765 , n80683 , n426954 );
and ( n80766 , n426795 , n426872 );
or ( n80767 , n80765 , n80766 );
buf ( n426958 , n80767 );
buf ( n426959 , n426958 );
xor ( n80770 , n426790 , n426959 );
xor ( n80771 , n426846 , n426849 );
xor ( n426962 , n80771 , n426867 );
buf ( n426963 , n426962 );
buf ( n426964 , n71095 );
buf ( n426965 , n63625 );
and ( n80776 , n426964 , n426965 );
buf ( n426967 , n417729 );
buf ( n426968 , n62511 );
and ( n80779 , n426967 , n426968 );
nor ( n80780 , n80776 , n80779 );
buf ( n426971 , n80780 );
buf ( n426972 , n426971 );
buf ( n426973 , n410635 );
or ( n80784 , n426972 , n426973 );
buf ( n426975 , n426858 );
buf ( n426976 , n409504 );
or ( n80787 , n426975 , n426976 );
nand ( n80788 , n80784 , n80787 );
buf ( n426979 , n80788 );
xor ( n80790 , n426811 , n426825 );
xor ( n80791 , n80790 , n426842 );
and ( n80792 , n426979 , n80791 );
buf ( n426983 , n426835 );
buf ( n426984 , n405378 );
or ( n80795 , n426983 , n426984 );
buf ( n426986 , n405414 );
nand ( n80797 , n80795 , n426986 );
buf ( n426988 , n80797 );
buf ( n426989 , n426988 );
buf ( n426990 , n62177 );
buf ( n426991 , n71664 );
and ( n80802 , n426990 , n426991 );
buf ( n426993 , n62159 );
buf ( n426994 , n418298 );
and ( n80805 , n426993 , n426994 );
nor ( n80806 , n80802 , n80805 );
buf ( n426997 , n80806 );
buf ( n426998 , n426997 );
buf ( n426999 , n409429 );
or ( n80810 , n426998 , n426999 );
buf ( n427001 , n426910 );
buf ( n427002 , n409170 );
or ( n80813 , n427001 , n427002 );
nand ( n80814 , n80810 , n80813 );
buf ( n427005 , n80814 );
buf ( n427006 , n427005 );
xor ( n80817 , n426989 , n427006 );
buf ( n427008 , n71088 );
buf ( n427009 , n63625 );
and ( n80820 , n427008 , n427009 );
buf ( n427011 , n417722 );
buf ( n427012 , n62511 );
and ( n80823 , n427011 , n427012 );
nor ( n427014 , n80820 , n80823 );
buf ( n427015 , n427014 );
buf ( n427016 , n427015 );
buf ( n427017 , n410635 );
or ( n80828 , n427016 , n427017 );
buf ( n427019 , n426971 );
buf ( n427020 , n409504 );
or ( n80831 , n427019 , n427020 );
nand ( n80832 , n80828 , n80831 );
buf ( n427023 , n80832 );
buf ( n427024 , n427023 );
and ( n80835 , n80817 , n427024 );
and ( n80836 , n426989 , n427006 );
or ( n80837 , n80835 , n80836 );
buf ( n427028 , n80837 );
xor ( n80839 , n426811 , n426825 );
xor ( n80840 , n80839 , n426842 );
and ( n80841 , n427028 , n80840 );
and ( n80842 , n426979 , n427028 );
or ( n80843 , n80792 , n80841 , n80842 );
xor ( n80844 , n426963 , n80843 );
xor ( n80845 , n426877 , n426931 );
xor ( n80846 , n80845 , n426949 );
buf ( n427037 , n80846 );
and ( n80848 , n80844 , n427037 );
and ( n80849 , n426963 , n80843 );
or ( n80850 , n80848 , n80849 );
buf ( n427041 , n80850 );
xor ( n80852 , n426144 , n426163 );
xor ( n80853 , n80852 , n426177 );
xor ( n80854 , n426308 , n426327 );
xor ( n80855 , n80853 , n80854 );
buf ( n427046 , n80855 );
xor ( n80857 , n427041 , n427046 );
xor ( n80858 , n426795 , n426872 );
xor ( n80859 , n80858 , n426954 );
buf ( n427050 , n80859 );
buf ( n427051 , n427050 );
and ( n80862 , n80857 , n427051 );
and ( n80863 , n427041 , n427046 );
or ( n80864 , n80862 , n80863 );
buf ( n427055 , n80864 );
buf ( n427056 , n427055 );
and ( n80867 , n80770 , n427056 );
and ( n80868 , n426790 , n426959 );
or ( n80869 , n80867 , n80868 );
buf ( n427060 , n80869 );
buf ( n427061 , n427060 );
xor ( n80872 , n426344 , n426348 );
xor ( n80873 , n80872 , n426353 );
buf ( n427064 , n80873 );
buf ( n427065 , n427064 );
xor ( n80876 , n427061 , n427065 );
buf ( n427067 , n426775 );
not ( n80878 , n427067 );
buf ( n427069 , n80592 );
not ( n80880 , n427069 );
or ( n80881 , n80878 , n80880 );
buf ( n427072 , n45948 );
not ( n80883 , n427072 );
buf ( n427074 , n80883 );
buf ( n427075 , n427074 );
buf ( n427076 , n80158 );
not ( n80887 , n427076 );
buf ( n427078 , n426763 );
not ( n80889 , n427078 );
or ( n80890 , n80887 , n80889 );
buf ( n427081 , n392217 );
buf ( n427082 , n426376 );
nand ( n80893 , n427081 , n427082 );
buf ( n427084 , n80893 );
buf ( n427085 , n427084 );
nand ( n80896 , n80890 , n427085 );
buf ( n427087 , n80896 );
buf ( n427088 , n427087 );
nand ( n80899 , n427075 , n427088 );
buf ( n427090 , n80899 );
buf ( n427091 , n427090 );
nand ( n80902 , n80881 , n427091 );
buf ( n427093 , n80902 );
buf ( n427094 , n427093 );
and ( n80905 , n80876 , n427094 );
and ( n80906 , n427061 , n427065 );
or ( n80907 , n80905 , n80906 );
buf ( n427098 , n80907 );
and ( n80909 , n80595 , n427098 );
and ( n80910 , n80584 , n80594 );
or ( n80911 , n80909 , n80910 );
buf ( n427102 , n80911 );
xor ( n80913 , n426770 , n427102 );
buf ( n427104 , n395359 );
not ( n80915 , n427104 );
buf ( n427106 , n426745 );
not ( n80917 , n427106 );
or ( n80918 , n80915 , n80917 );
and ( n80919 , n372471 , n419385 );
not ( n80920 , n372471 );
and ( n80921 , n80920 , n47863 );
or ( n80922 , n80919 , n80921 );
buf ( n427113 , n80922 );
buf ( n427114 , n395346 );
nand ( n80925 , n427113 , n427114 );
buf ( n427116 , n80925 );
buf ( n427117 , n427116 );
nand ( n427118 , n80918 , n427117 );
buf ( n427119 , n427118 );
buf ( n427120 , n427119 );
and ( n80931 , n80913 , n427120 );
and ( n80932 , n426770 , n427102 );
or ( n80933 , n80931 , n80932 );
buf ( n427124 , n80933 );
buf ( n427125 , n427124 );
xor ( n80936 , n426753 , n427125 );
buf ( n427127 , n399274 );
not ( n80938 , n427127 );
buf ( n427129 , n418734 );
not ( n80940 , n427129 );
or ( n80941 , n80938 , n80940 );
buf ( n427132 , n388722 );
buf ( n427133 , n399283 );
nand ( n80944 , n427132 , n427133 );
buf ( n427135 , n80944 );
buf ( n427136 , n427135 );
nand ( n80947 , n80941 , n427136 );
buf ( n427138 , n80947 );
buf ( n427139 , n427138 );
not ( n80950 , n427139 );
buf ( n427141 , n40592 );
not ( n80952 , n427141 );
or ( n80953 , n80950 , n80952 );
buf ( n427144 , n425979 );
buf ( n427145 , n388068 );
nand ( n80956 , n427144 , n427145 );
buf ( n427147 , n80956 );
buf ( n427148 , n427147 );
nand ( n80959 , n80953 , n427148 );
buf ( n427150 , n80959 );
buf ( n427151 , n427150 );
and ( n80962 , n80936 , n427151 );
and ( n80963 , n426753 , n427125 );
or ( n80964 , n80962 , n80963 );
buf ( n427155 , n80964 );
buf ( n427156 , n427155 );
xor ( n80967 , n426728 , n427156 );
xor ( n80968 , n425967 , n425992 );
xor ( n80969 , n80968 , n425997 );
buf ( n427160 , n80969 );
buf ( n427161 , n427160 );
and ( n80972 , n80967 , n427161 );
and ( n80973 , n426728 , n427156 );
or ( n80974 , n80972 , n80973 );
buf ( n427165 , n80974 );
buf ( n427166 , n427165 );
and ( n80977 , n80517 , n427166 );
and ( n80978 , n426689 , n426706 );
or ( n80979 , n80977 , n80978 );
buf ( n427170 , n80979 );
buf ( n427171 , n427170 );
xor ( n80982 , n426664 , n427171 );
xor ( n80983 , n426007 , n426033 );
xor ( n80984 , n80983 , n426038 );
buf ( n427175 , n80984 );
buf ( n427176 , n427175 );
and ( n80987 , n80982 , n427176 );
and ( n80988 , n426664 , n427171 );
or ( n80989 , n80987 , n80988 );
buf ( n427180 , n80989 );
buf ( n427181 , n427180 );
xor ( n80992 , n426660 , n427181 );
xor ( n80993 , n425850 , n425875 );
xor ( n80994 , n80993 , n426043 );
buf ( n427185 , n80994 );
buf ( n427186 , n427185 );
and ( n427187 , n80992 , n427186 );
and ( n427188 , n426660 , n427181 );
or ( n80999 , n427187 , n427188 );
buf ( n427190 , n80999 );
buf ( n427191 , n427190 );
xor ( n81002 , n426656 , n427191 );
xor ( n81003 , n425846 , n426048 );
xor ( n81004 , n81003 , n426050 );
buf ( n427195 , n81004 );
buf ( n427196 , n427195 );
and ( n427197 , n81002 , n427196 );
and ( n81008 , n426656 , n427191 );
or ( n81009 , n427197 , n81008 );
buf ( n427200 , n81009 );
not ( n81011 , n427200 );
or ( n81012 , n80462 , n81011 );
not ( n81013 , n426651 );
not ( n81014 , n81013 );
not ( n81015 , n427200 );
not ( n81016 , n81015 );
or ( n81017 , n81014 , n81016 );
xor ( n81018 , n79824 , n426518 );
xnor ( n81019 , n81018 , n426527 );
nand ( n81020 , n81017 , n81019 );
nand ( n81021 , n81012 , n81020 );
not ( n81022 , n81021 );
not ( n81023 , n79825 );
not ( n81024 , n426518 );
or ( n81025 , n81023 , n81024 );
nand ( n81026 , n81025 , n80338 );
not ( n81027 , n81026 );
not ( n81028 , n79580 );
or ( n81029 , n81027 , n81028 );
or ( n81030 , n80339 , n79580 );
nand ( n81031 , n81029 , n81030 );
not ( n81032 , n81031 );
not ( n81033 , n80350 );
and ( n81034 , n81032 , n81033 );
and ( n81035 , n80350 , n81031 );
nor ( n81036 , n81034 , n81035 );
nand ( n81037 , n81022 , n81036 );
not ( n81038 , n81037 );
buf ( n427229 , C0 );
buf ( n427230 , n427229 );
xor ( n81056 , n426070 , n426072 );
xor ( n81057 , n81056 , n426509 );
buf ( n427233 , n81057 );
buf ( n427234 , n427233 );
xor ( n81060 , n427230 , n427234 );
xor ( n81061 , n425880 , n425905 );
xor ( n81062 , n81061 , n426002 );
buf ( n427238 , n81062 );
buf ( n427239 , n427238 );
buf ( n427240 , n59916 );
not ( n81066 , n427240 );
buf ( n427242 , n80508 );
not ( n81068 , n427242 );
or ( n81069 , n81066 , n81068 );
buf ( n427245 , n47891 );
not ( n81071 , n427245 );
buf ( n427247 , n42065 );
not ( n81073 , n427247 );
or ( n81074 , n81071 , n81073 );
buf ( n427250 , n42066 );
buf ( n427251 , n403668 );
nand ( n81077 , n427250 , n427251 );
buf ( n427253 , n81077 );
buf ( n427254 , n427253 );
nand ( n81080 , n81074 , n427254 );
buf ( n427256 , n81080 );
buf ( n427257 , n427256 );
buf ( n427258 , n50579 );
nand ( n81084 , n427257 , n427258 );
buf ( n427260 , n81084 );
buf ( n427261 , n427260 );
nand ( n81087 , n81069 , n427261 );
buf ( n427263 , n81087 );
buf ( n427264 , n427263 );
buf ( n427265 , n426393 );
buf ( n427266 , n426103 );
xor ( n81092 , n427265 , n427266 );
buf ( n427268 , n426398 );
xnor ( n81094 , n81092 , n427268 );
buf ( n427270 , n81094 );
buf ( n427271 , n427270 );
not ( n81097 , n427271 );
buf ( n427273 , n81097 );
not ( n81099 , n427273 );
not ( n81100 , n358975 );
nor ( n81101 , n81100 , n41663 );
not ( n81102 , n81101 );
or ( n81103 , n81099 , n81102 );
not ( n81104 , n427270 );
not ( n81105 , n41663 );
nand ( n81106 , n81105 , n358975 );
not ( n81107 , n81106 );
or ( n81108 , n81104 , n81107 );
xor ( n81109 , n426363 , n426367 );
xor ( n81110 , n81109 , n426389 );
buf ( n427286 , n81110 );
and ( n81112 , n55543 , n420986 );
not ( n81113 , n55543 );
and ( n81114 , n81113 , n388064 );
or ( n81115 , n81112 , n81114 );
buf ( n427291 , n81115 );
not ( n81117 , n427291 );
buf ( n427293 , n74374 );
not ( n81119 , n427293 );
or ( n81120 , n81117 , n81119 );
buf ( n427296 , n43514 );
not ( n81122 , n427296 );
buf ( n427298 , n426091 );
nand ( n81124 , n81122 , n427298 );
buf ( n427300 , n81124 );
buf ( n427301 , n427300 );
nand ( n427302 , n81120 , n427301 );
buf ( n427303 , n427302 );
xor ( n81129 , n427286 , n427303 );
not ( n81130 , n44770 );
buf ( n427306 , n397486 );
not ( n427307 , n427306 );
buf ( n427308 , n427307 );
buf ( n427309 , n427308 );
not ( n81135 , n427309 );
buf ( n427311 , n422673 );
not ( n81137 , n427311 );
or ( n81138 , n81135 , n81137 );
buf ( n427314 , n44775 );
buf ( n427315 , n397486 );
nand ( n81141 , n427314 , n427315 );
buf ( n427317 , n81141 );
buf ( n427318 , n427317 );
nand ( n81144 , n81138 , n427318 );
buf ( n427320 , n81144 );
not ( n81146 , n427320 );
or ( n81147 , n81130 , n81146 );
nand ( n81148 , n80169 , n413643 );
nand ( n81149 , n81147 , n81148 );
buf ( n427325 , n81149 );
not ( n81151 , n427325 );
buf ( n427327 , n395359 );
not ( n81153 , n427327 );
buf ( n427329 , n80922 );
not ( n81155 , n427329 );
or ( n81156 , n81153 , n81155 );
buf ( n427332 , n395346 );
buf ( n427333 , n47863 );
not ( n81159 , n427333 );
buf ( n427335 , n392878 );
not ( n81161 , n427335 );
or ( n81162 , n81159 , n81161 );
buf ( n427338 , n424808 );
buf ( n427339 , n419385 );
nand ( n81165 , n427338 , n427339 );
buf ( n427341 , n81165 );
buf ( n427342 , n427341 );
nand ( n81168 , n81162 , n427342 );
buf ( n427344 , n81168 );
buf ( n427345 , n427344 );
nand ( n81171 , n427332 , n427345 );
buf ( n427347 , n81171 );
buf ( n427348 , n427347 );
nand ( n81174 , n81156 , n427348 );
buf ( n427350 , n81174 );
buf ( n427351 , n427350 );
not ( n81177 , n427351 );
or ( n81178 , n81151 , n81177 );
buf ( n427354 , n81149 );
not ( n81180 , n427354 );
buf ( n427356 , n81180 );
buf ( n427357 , n427356 );
not ( n81183 , n427357 );
buf ( n427359 , n427350 );
not ( n81185 , n427359 );
buf ( n427361 , n81185 );
buf ( n427362 , n427361 );
not ( n81188 , n427362 );
or ( n81189 , n81183 , n81188 );
xor ( n81190 , n80584 , n80594 );
xor ( n81191 , n81190 , n427098 );
buf ( n427367 , n81191 );
nand ( n81193 , n81189 , n427367 );
buf ( n427369 , n81193 );
buf ( n427370 , n427369 );
nand ( n81196 , n81178 , n427370 );
buf ( n427372 , n81196 );
and ( n81198 , n81129 , n427372 );
and ( n81199 , n427286 , n427303 );
or ( n81200 , n81198 , n81199 );
nand ( n81201 , n81108 , n81200 );
nand ( n81202 , n81103 , n81201 );
buf ( n427378 , n81202 );
xor ( n81204 , n427264 , n427378 );
buf ( n427380 , n416762 );
not ( n81206 , n427380 );
buf ( n427382 , n358975 );
not ( n81208 , n427382 );
buf ( n427384 , n62006 );
not ( n81210 , n427384 );
or ( n81211 , n81208 , n81210 );
buf ( n427387 , n24116 );
buf ( n427388 , n402819 );
nand ( n81214 , n427387 , n427388 );
buf ( n427390 , n81214 );
buf ( n427391 , n427390 );
nand ( n81217 , n81211 , n427391 );
buf ( n427393 , n81217 );
buf ( n427394 , n427393 );
not ( n81220 , n427394 );
or ( n81221 , n81206 , n81220 );
buf ( n427397 , n426676 );
buf ( n427398 , n41664 );
nand ( n81224 , n427397 , n427398 );
buf ( n427400 , n81224 );
buf ( n427401 , n427400 );
nand ( n81227 , n81221 , n427401 );
buf ( n427403 , n81227 );
buf ( n427404 , n427403 );
and ( n81230 , n81204 , n427404 );
and ( n81231 , n427264 , n427378 );
or ( n81232 , n81230 , n81231 );
buf ( n427408 , n81232 );
buf ( n427409 , n427408 );
xor ( n81235 , n427239 , n427409 );
xor ( n81236 , n426079 , n426456 );
xor ( n81237 , n81236 , n426460 );
buf ( n427413 , n81237 );
buf ( n427414 , n427413 );
and ( n81240 , n81235 , n427414 );
and ( n81241 , n427239 , n427409 );
or ( n81242 , n81240 , n81241 );
buf ( n427418 , n81242 );
buf ( n427419 , n427418 );
xor ( n81245 , n426465 , n426486 );
xor ( n81246 , n81245 , n426504 );
buf ( n427422 , n81246 );
buf ( n427423 , n427422 );
buf ( n427424 , C0 );
buf ( n427425 , n427424 );
and ( n81276 , n427419 , n427423 );
or ( n81277 , C0 , n81276 );
buf ( n427428 , n81277 );
buf ( n427429 , n427428 );
and ( n81280 , n81060 , n427429 );
or ( n81282 , n81280 , C0 );
buf ( n427432 , n81282 );
buf ( n427433 , n427432 );
xor ( n81285 , n426060 , n426513 );
xor ( n81286 , n81285 , n426515 );
buf ( n427436 , n81286 );
buf ( n427437 , n427436 );
xor ( n81289 , n427433 , n427437 );
xor ( n81290 , n426656 , n427191 );
xor ( n81291 , n81290 , n427196 );
buf ( n427441 , n81291 );
buf ( n427442 , n427441 );
and ( n81294 , n81289 , n427442 );
and ( n81295 , n427433 , n427437 );
or ( n81296 , n81294 , n81295 );
buf ( n427446 , n81296 );
buf ( n427447 , n427446 );
xor ( n81299 , n426651 , n81015 );
xnor ( n81300 , n81299 , n81019 );
buf ( n427450 , n81300 );
xor ( n81302 , n427447 , n427450 );
xor ( n81303 , n426410 , n426435 );
xor ( n81304 , n81303 , n426451 );
buf ( n427454 , n81304 );
buf ( n427455 , n427454 );
buf ( n427456 , n51553 );
not ( n81308 , n427456 );
buf ( n427458 , n427256 );
not ( n81310 , n427458 );
or ( n81311 , n81308 , n81310 );
buf ( n427461 , n47891 );
not ( n81313 , n427461 );
buf ( n427463 , n418729 );
not ( n81315 , n427463 );
or ( n81316 , n81313 , n81315 );
buf ( n427466 , n41861 );
buf ( n427467 , n403668 );
nand ( n81319 , n427466 , n427467 );
buf ( n427469 , n81319 );
buf ( n427470 , n427469 );
nand ( n81322 , n81316 , n427470 );
buf ( n427472 , n81322 );
buf ( n427473 , n427472 );
buf ( n427474 , n50579 );
nand ( n81326 , n427473 , n427474 );
buf ( n427476 , n81326 );
buf ( n427477 , n427476 );
nand ( n81329 , n81311 , n427477 );
buf ( n427479 , n81329 );
buf ( n427480 , n427479 );
buf ( n427481 , n400033 );
not ( n81333 , n427481 );
buf ( n427483 , n388080 );
not ( n81335 , n427483 );
or ( n81336 , n81333 , n81335 );
buf ( n427486 , n388722 );
buf ( n427487 , n400042 );
nand ( n81339 , n427486 , n427487 );
buf ( n427489 , n81339 );
buf ( n427490 , n427489 );
nand ( n81342 , n81336 , n427490 );
buf ( n427492 , n81342 );
buf ( n427493 , n427492 );
not ( n81345 , n427493 );
buf ( n427495 , n67042 );
not ( n81347 , n427495 );
or ( n81348 , n81345 , n81347 );
buf ( n427498 , n40567 );
not ( n81350 , n427498 );
buf ( n427500 , n427138 );
nand ( n81352 , n81350 , n427500 );
buf ( n427502 , n81352 );
buf ( n427503 , n427502 );
nand ( n81355 , n81348 , n427503 );
buf ( n427505 , n81355 );
not ( n81357 , n427505 );
buf ( n427507 , n421646 );
buf ( n427508 , n388722 );
buf ( n427509 , n23773 );
or ( n81361 , n427508 , n427509 );
buf ( n427511 , n358975 );
nand ( n427512 , n81361 , n427511 );
buf ( n427513 , n427512 );
buf ( n427514 , n427513 );
not ( n81366 , n23774 );
nand ( n81367 , n81366 , n388722 );
buf ( n427517 , n81367 );
nand ( n81369 , n427507 , n427514 , n427517 );
buf ( n427519 , n81369 );
nand ( n81371 , n81357 , n427519 );
not ( n81372 , n81371 );
xor ( n81373 , n426770 , n427102 );
xor ( n81374 , n81373 , n427120 );
buf ( n427524 , n81374 );
not ( n81376 , n427524 );
or ( n81377 , n81372 , n81376 );
buf ( n427527 , n427519 );
not ( n81379 , n427527 );
buf ( n427529 , n81379 );
buf ( n427530 , n427529 );
buf ( n427531 , n427505 );
nand ( n81383 , n427530 , n427531 );
buf ( n427533 , n81383 );
nand ( n81385 , n81377 , n427533 );
buf ( n427535 , n81385 );
xor ( n81387 , n427480 , n427535 );
buf ( n427537 , n55055 );
not ( n81389 , n427537 );
buf ( n427539 , n371797 );
not ( n81391 , n427539 );
or ( n81392 , n81389 , n81391 );
buf ( n427542 , n421646 );
buf ( n427543 , n55054 );
nand ( n81395 , n427542 , n427543 );
buf ( n427545 , n81395 );
buf ( n427546 , n427545 );
nand ( n81398 , n81392 , n427546 );
buf ( n427548 , n81398 );
buf ( n427549 , n427548 );
not ( n81401 , n427549 );
buf ( n427551 , n388740 );
not ( n81403 , n427551 );
or ( n81404 , n81401 , n81403 );
buf ( n427554 , n426715 );
buf ( n427555 , n388803 );
nand ( n81407 , n427554 , n427555 );
buf ( n427557 , n81407 );
buf ( n427558 , n427557 );
nand ( n81410 , n81404 , n427558 );
buf ( n427560 , n81410 );
buf ( n427561 , n427560 );
and ( n81413 , n81387 , n427561 );
and ( n81414 , n427480 , n427535 );
or ( n81415 , n81413 , n81414 );
buf ( n427565 , n81415 );
buf ( n427566 , n427565 );
xor ( n81418 , n427455 , n427566 );
xor ( n81419 , n426728 , n427156 );
xor ( n81420 , n81419 , n427161 );
buf ( n427570 , n81420 );
buf ( n427571 , n427570 );
and ( n81423 , n81418 , n427571 );
and ( n81424 , n427455 , n427566 );
or ( n81425 , n81423 , n81424 );
buf ( n427575 , n81425 );
buf ( n427576 , n427575 );
xor ( n81428 , n426689 , n426706 );
xor ( n81429 , n81428 , n427166 );
buf ( n427579 , n81429 );
buf ( n427580 , n427579 );
buf ( n427581 , C0 );
buf ( n427582 , n427581 );
and ( n81448 , n427576 , n427580 );
or ( n81449 , C0 , n81448 );
buf ( n427585 , n81449 );
buf ( n427586 , n427585 );
xor ( n81452 , n426664 , n427171 );
xor ( n81453 , n81452 , n427176 );
buf ( n427589 , n81453 );
buf ( n427590 , n427589 );
buf ( n427591 , C0 );
buf ( n427592 , n427591 );
and ( n81470 , n427586 , n427590 );
or ( n81471 , C0 , n81470 );
buf ( n427595 , n81471 );
buf ( n427596 , n427595 );
xor ( n81474 , n426660 , n427181 );
xor ( n81475 , n81474 , n427186 );
buf ( n427599 , n81475 );
buf ( n427600 , n427599 );
xor ( n81478 , n427596 , n427600 );
xor ( n81479 , n427230 , n427234 );
xor ( n81480 , n81479 , n427429 );
buf ( n427604 , n81480 );
buf ( n427605 , n427604 );
and ( n81483 , n81478 , n427605 );
and ( n81484 , n427596 , n427600 );
or ( n81485 , n81483 , n81484 );
buf ( n427609 , n81485 );
buf ( n427610 , n427609 );
xor ( n81488 , n427433 , n427437 );
xor ( n81489 , n81488 , n427442 );
buf ( n427613 , n81489 );
buf ( n427614 , n427613 );
xor ( n81492 , n427610 , n427614 );
buf ( n427616 , C0 );
buf ( n427617 , n427616 );
xor ( n81507 , n427264 , n427378 );
xor ( n81508 , n81507 , n427404 );
buf ( n427620 , n81508 );
buf ( n427621 , n427620 );
or ( n81511 , n427617 , n427621 );
xor ( n81512 , n426753 , n427125 );
xor ( n81513 , n81512 , n427151 );
buf ( n427625 , n81513 );
buf ( n427626 , n427625 );
not ( n81516 , n427626 );
not ( n81517 , n51553 );
not ( n81518 , n427472 );
or ( n81519 , n81517 , n81518 );
buf ( n427631 , n47891 );
not ( n81521 , n427631 );
buf ( n427633 , n420954 );
not ( n81523 , n427633 );
or ( n81524 , n81521 , n81523 );
buf ( n427636 , n389338 );
buf ( n427637 , n403668 );
nand ( n81527 , n427636 , n427637 );
buf ( n427639 , n81527 );
buf ( n427640 , n427639 );
nand ( n81530 , n81524 , n427640 );
buf ( n427642 , n81530 );
buf ( n427643 , n427642 );
buf ( n427644 , n50579 );
nand ( n81534 , n427643 , n427644 );
buf ( n427646 , n81534 );
nand ( n81536 , n81519 , n427646 );
not ( n81537 , n81536 );
xor ( n81538 , n427286 , n427303 );
xor ( n81539 , n81538 , n427372 );
not ( n81540 , n81539 );
or ( n81541 , n81537 , n81540 );
not ( n81542 , n81536 );
not ( n81543 , n81542 );
not ( n81544 , n81539 );
not ( n81545 , n81544 );
or ( n81546 , n81543 , n81545 );
xor ( n81547 , n426790 , n426959 );
xor ( n81548 , n81547 , n427056 );
buf ( n427660 , n81548 );
buf ( n427661 , n427660 );
buf ( n427662 , n427308 );
not ( n81552 , n427662 );
buf ( n427664 , n426763 );
not ( n81554 , n427664 );
or ( n81555 , n81552 , n81554 );
buf ( n427667 , n392217 );
buf ( n427668 , n397486 );
nand ( n81558 , n427667 , n427668 );
buf ( n427670 , n81558 );
buf ( n427671 , n427670 );
nand ( n81561 , n81555 , n427671 );
buf ( n427673 , n81561 );
buf ( n427674 , n427673 );
not ( n81564 , n427674 );
buf ( n427676 , n427074 );
not ( n81566 , n427676 );
or ( n81567 , n81564 , n81566 );
buf ( n427679 , n427087 );
buf ( n427680 , n45954 );
nand ( n81570 , n427679 , n427680 );
buf ( n427682 , n81570 );
buf ( n427683 , n427682 );
nand ( n81573 , n81567 , n427683 );
buf ( n427685 , n81573 );
buf ( n427686 , n427685 );
xor ( n81576 , n427661 , n427686 );
buf ( n427688 , n395359 );
not ( n81578 , n427688 );
not ( n81579 , n23603 );
buf ( n427691 , n81579 );
not ( n81581 , n427691 );
buf ( n427693 , n394207 );
not ( n81583 , n427693 );
or ( n81584 , n81581 , n81583 );
buf ( n427696 , n81579 );
not ( n81586 , n427696 );
buf ( n427698 , n81586 );
buf ( n427699 , n427698 );
buf ( n427700 , n24828 );
nand ( n81590 , n427699 , n427700 );
buf ( n427702 , n81590 );
buf ( n427703 , n427702 );
nand ( n81593 , n81584 , n427703 );
buf ( n427705 , n81593 );
buf ( n427706 , n427705 );
not ( n81596 , n427706 );
or ( n81597 , n81578 , n81596 );
buf ( n427709 , n47863 );
buf ( n427710 , n417572 );
and ( n81600 , n427709 , n427710 );
not ( n81601 , n427709 );
buf ( n427713 , n394814 );
and ( n81603 , n81601 , n427713 );
nor ( n81604 , n81600 , n81603 );
buf ( n427716 , n81604 );
buf ( n427717 , n427716 );
buf ( n427718 , n395346 );
nand ( n81608 , n427717 , n427718 );
buf ( n427720 , n81608 );
buf ( n427721 , n427720 );
nand ( n81611 , n81597 , n427721 );
buf ( n427723 , n81611 );
buf ( n427724 , n427723 );
and ( n81614 , n81576 , n427724 );
and ( n81615 , n427661 , n427686 );
or ( n81616 , n81614 , n81615 );
buf ( n427728 , n81616 );
buf ( n427729 , n427728 );
buf ( n427730 , n59916 );
not ( n81620 , n427730 );
buf ( n427732 , n47891 );
not ( n81622 , n427732 );
buf ( n427734 , n420997 );
not ( n427735 , n427734 );
or ( n427736 , n81622 , n427735 );
buf ( n427737 , n420994 );
buf ( n427738 , n61299 );
nand ( n81628 , n427737 , n427738 );
buf ( n427740 , n81628 );
buf ( n427741 , n427740 );
nand ( n81631 , n427736 , n427741 );
buf ( n427743 , n81631 );
buf ( n427744 , n427743 );
not ( n81634 , n427744 );
or ( n81635 , n81620 , n81634 );
buf ( n427747 , n47891 );
not ( n81637 , n427747 );
buf ( n427749 , n418804 );
not ( n427750 , n427749 );
or ( n427751 , n81637 , n427750 );
buf ( n427752 , n392608 );
buf ( n427753 , n61299 );
nand ( n81643 , n427752 , n427753 );
buf ( n427755 , n81643 );
buf ( n427756 , n427755 );
nand ( n81646 , n427751 , n427756 );
buf ( n427758 , n81646 );
buf ( n427759 , n427758 );
buf ( n427760 , n50579 );
nand ( n81650 , n427759 , n427760 );
buf ( n427762 , n81650 );
buf ( n427763 , n427762 );
nand ( n81653 , n81635 , n427763 );
buf ( n427765 , n81653 );
buf ( n427766 , n427765 );
xor ( n81656 , n427729 , n427766 );
buf ( n427768 , n388076 );
not ( n81658 , n427768 );
buf ( n427770 , n81658 );
buf ( n427771 , n427770 );
buf ( n427772 , n371879 );
or ( n81662 , n427771 , n427772 );
buf ( n427774 , n358975 );
nand ( n81664 , n81662 , n427774 );
buf ( n427776 , n81664 );
buf ( n427777 , n427776 );
buf ( n427778 , n388722 );
buf ( n427779 , n427770 );
buf ( n427780 , n371879 );
nand ( n81670 , n427779 , n427780 );
buf ( n427782 , n81670 );
buf ( n427783 , n427782 );
and ( n81673 , n427777 , n427778 , n427783 );
buf ( n427785 , n81673 );
buf ( n427786 , n427785 );
and ( n81676 , n81656 , n427786 );
and ( n81677 , n427729 , n427766 );
or ( n81678 , n81676 , n81677 );
buf ( n427790 , n81678 );
not ( n81680 , n427790 );
xor ( n81681 , n427061 , n427065 );
xor ( n81682 , n81681 , n427094 );
buf ( n427794 , n81682 );
buf ( n427795 , n427794 );
buf ( n427796 , n395359 );
not ( n81686 , n427796 );
buf ( n427798 , n427344 );
not ( n81688 , n427798 );
or ( n81689 , n81686 , n81688 );
buf ( n427801 , n427705 );
buf ( n427802 , n395346 );
nand ( n81692 , n427801 , n427802 );
buf ( n427804 , n81692 );
buf ( n427805 , n427804 );
nand ( n81695 , n81689 , n427805 );
buf ( n427807 , n81695 );
buf ( n427808 , n427807 );
xor ( n81698 , n427795 , n427808 );
buf ( n427810 , n55543 );
not ( n81700 , n427810 );
buf ( n427812 , n390985 );
not ( n427813 , n427812 );
or ( n81703 , n81700 , n427813 );
buf ( n427815 , n390988 );
buf ( n427816 , n51185 );
nand ( n427817 , n427815 , n427816 );
buf ( n427818 , n427817 );
buf ( n427819 , n427818 );
nand ( n81709 , n81703 , n427819 );
buf ( n427821 , n81709 );
buf ( n427822 , n427821 );
not ( n81712 , n427822 );
buf ( n427824 , n44770 );
not ( n81714 , n427824 );
or ( n81715 , n81712 , n81714 );
buf ( n427827 , n427320 );
buf ( n427828 , n413643 );
nand ( n81718 , n427827 , n427828 );
buf ( n427830 , n81718 );
buf ( n427831 , n427830 );
nand ( n81721 , n81715 , n427831 );
buf ( n427833 , n81721 );
buf ( n427834 , n427833 );
and ( n81724 , n81698 , n427834 );
and ( n81725 , n427795 , n427808 );
or ( n81726 , n81724 , n81725 );
buf ( n427838 , n81726 );
not ( n81728 , n427838 );
buf ( n427840 , n399283 );
buf ( n427841 , n371879 );
and ( n81731 , n427840 , n427841 );
not ( n81732 , n427840 );
buf ( n427844 , n425525 );
and ( n81734 , n81732 , n427844 );
nor ( n81735 , n81731 , n81734 );
buf ( n427847 , n81735 );
buf ( n427848 , n427847 );
not ( n81738 , n427848 );
buf ( n427850 , n81738 );
buf ( n427851 , n427850 );
not ( n81741 , n427851 );
buf ( n427853 , n74375 );
not ( n81743 , n427853 );
or ( n81744 , n81741 , n81743 );
buf ( n427856 , n81115 );
buf ( n427857 , n43515 );
nand ( n81747 , n427856 , n427857 );
buf ( n427859 , n81747 );
buf ( n427860 , n427859 );
nand ( n81750 , n81744 , n427860 );
buf ( n427862 , n81750 );
not ( n81752 , n427862 );
nand ( n81753 , n81728 , n81752 );
not ( n81754 , n81753 );
or ( n81755 , n81680 , n81754 );
not ( n81756 , n81752 );
nand ( n81757 , n81756 , n427838 );
nand ( n81758 , n81755 , n81757 );
nand ( n81759 , n81546 , n81758 );
nand ( n81760 , n81541 , n81759 );
buf ( n427872 , n81760 );
not ( n81762 , n427872 );
or ( n81763 , n81516 , n81762 );
buf ( n427875 , n81760 );
buf ( n427876 , n427625 );
or ( n81766 , n427875 , n427876 );
and ( n81767 , n81200 , n427270 );
not ( n81768 , n81200 );
and ( n81769 , n81768 , n427273 );
or ( n81770 , n81767 , n81769 );
buf ( n427882 , n81770 );
buf ( n427883 , n81101 );
and ( n81773 , n427882 , n427883 );
not ( n81774 , n427882 );
buf ( n427886 , n81106 );
and ( n81776 , n81774 , n427886 );
nor ( n81777 , n81773 , n81776 );
buf ( n427889 , n81777 );
buf ( n427890 , n427889 );
nand ( n81780 , n81766 , n427890 );
buf ( n427892 , n81780 );
buf ( n427893 , n427892 );
nand ( n81783 , n81763 , n427893 );
buf ( n427895 , n81783 );
buf ( n427896 , n427895 );
nand ( n81786 , n81511 , n427896 );
buf ( n427898 , n81786 );
buf ( n427899 , n427898 );
buf ( n427900 , C1 );
buf ( n427901 , n427900 );
nand ( n81794 , n427899 , n427901 );
buf ( n427903 , n81794 );
buf ( n427904 , n427903 );
xor ( n81797 , n427239 , n427409 );
xor ( n81798 , n81797 , n427414 );
buf ( n427907 , n81798 );
buf ( n427908 , n427907 );
buf ( n427909 , C0 );
buf ( n427910 , n427909 );
and ( n81823 , n427904 , n427908 );
or ( n81824 , C0 , n81823 );
buf ( n427913 , n81824 );
buf ( n427914 , n427913 );
xor ( n81827 , n427419 , n427423 );
xor ( n81828 , n81827 , n427425 );
buf ( n427917 , n81828 );
buf ( n427918 , n427917 );
xor ( n81831 , n427914 , n427918 );
xor ( n81832 , n427586 , n427590 );
xor ( n81833 , n81832 , n427592 );
buf ( n427922 , n81833 );
buf ( n427923 , n427922 );
and ( n81836 , n81831 , n427923 );
and ( n81837 , n427914 , n427918 );
or ( n81838 , n81836 , n81837 );
buf ( n427927 , n81838 );
buf ( n427928 , n427927 );
xor ( n81841 , n427596 , n427600 );
xor ( n81842 , n81841 , n427605 );
buf ( n427931 , n81842 );
buf ( n427932 , n427931 );
xor ( n81845 , n427928 , n427932 );
xor ( n81846 , n427576 , n427580 );
xor ( n81847 , n81846 , n427582 );
buf ( n427936 , n81847 );
buf ( n427937 , n427936 );
xor ( n81850 , n427455 , n427566 );
xor ( n81851 , n81850 , n427571 );
buf ( n427940 , n81851 );
buf ( n427941 , n427940 );
buf ( n427942 , C0 );
or ( n81872 , n427941 , n427942 );
buf ( n427944 , C0 );
xor ( n81885 , n427480 , n427535 );
xor ( n81886 , n81885 , n427561 );
buf ( n427947 , n81886 );
buf ( n427948 , n427944 );
buf ( n427949 , n427947 );
or ( n81893 , n427948 , n427949 );
buf ( n427951 , n427356 );
buf ( n427952 , n427350 );
xor ( n81896 , n427951 , n427952 );
buf ( n427954 , n81191 );
xnor ( n81898 , n81896 , n427954 );
buf ( n427956 , n81898 );
buf ( n427957 , n427956 );
buf ( n427958 , n55055 );
not ( n81902 , n427958 );
buf ( n427960 , n421024 );
not ( n81904 , n427960 );
or ( n81905 , n81902 , n81904 );
buf ( n427963 , n388722 );
buf ( n427964 , n55054 );
nand ( n81908 , n427963 , n427964 );
buf ( n427966 , n81908 );
buf ( n427967 , n427966 );
nand ( n81911 , n81905 , n427967 );
buf ( n427969 , n81911 );
buf ( n427970 , n427969 );
not ( n81914 , n427970 );
buf ( n427972 , n67042 );
not ( n81916 , n427972 );
or ( n81917 , n81914 , n81916 );
buf ( n427975 , n427492 );
buf ( n427976 , n388068 );
nand ( n81920 , n427975 , n427976 );
buf ( n427978 , n81920 );
buf ( n427979 , n427978 );
nand ( n81923 , n81917 , n427979 );
buf ( n427981 , n81923 );
buf ( n427982 , n427981 );
xor ( n81926 , n427957 , n427982 );
buf ( n427984 , n388800 );
buf ( n427985 , n402819 );
nor ( n81929 , n427984 , n427985 );
buf ( n427987 , n81929 );
buf ( n427988 , n427987 );
and ( n81932 , n81926 , n427988 );
and ( n81933 , n427957 , n427982 );
or ( n81934 , n81932 , n81933 );
buf ( n427992 , n81934 );
buf ( n427993 , n427992 );
buf ( n427994 , n358975 );
buf ( n427995 , n371800 );
and ( n81939 , n427994 , n427995 );
not ( n81940 , n427994 );
buf ( n427998 , n388751 );
and ( n81942 , n81940 , n427998 );
nor ( n81943 , n81939 , n81942 );
buf ( n428001 , n81943 );
buf ( n428002 , n428001 );
not ( n81946 , n428002 );
buf ( n428004 , n388740 );
not ( n81948 , n428004 );
or ( n81949 , n81946 , n81948 );
buf ( n428007 , n427548 );
buf ( n428008 , n388803 );
nand ( n81952 , n428007 , n428008 );
buf ( n428010 , n81952 );
buf ( n428011 , n428010 );
nand ( n81955 , n81949 , n428011 );
buf ( n428013 , n81955 );
buf ( n428014 , n428013 );
xor ( n81958 , n427993 , n428014 );
buf ( n428016 , n427524 );
buf ( n428017 , n427505 );
xor ( n81961 , n428016 , n428017 );
buf ( n428019 , n427529 );
xor ( n81963 , n81961 , n428019 );
buf ( n428021 , n81963 );
buf ( n428022 , n428021 );
and ( n81966 , n81958 , n428022 );
and ( n81967 , n427993 , n428014 );
or ( n81968 , n81966 , n81967 );
buf ( n428026 , n81968 );
buf ( n428027 , n428026 );
nand ( n81971 , n81893 , n428027 );
buf ( n428029 , n81971 );
buf ( n428030 , n428029 );
nand ( n81974 , C1 , n428030 );
buf ( n428032 , n81974 );
buf ( n428033 , n428032 );
nand ( n81977 , n81872 , n428033 );
buf ( n428035 , n81977 );
buf ( n428036 , n428035 );
buf ( n428037 , C1 );
buf ( n428038 , n428037 );
nand ( n81985 , n428036 , n428038 );
buf ( n428040 , n81985 );
buf ( n428041 , n428040 );
xor ( n81988 , n427937 , n428041 );
xor ( n81989 , n427904 , n427908 );
xor ( n81990 , n81989 , n427910 );
buf ( n428045 , n81990 );
buf ( n428046 , n428045 );
and ( n81993 , n81988 , n428046 );
and ( n81994 , n427937 , n428041 );
or ( n81995 , n81993 , n81994 );
buf ( n428050 , n81995 );
buf ( n428051 , n428050 );
xor ( n81998 , n427914 , n427918 );
xor ( n81999 , n81998 , n427923 );
buf ( n428054 , n81999 );
buf ( n428055 , n428054 );
xor ( n82002 , n428051 , n428055 );
buf ( n428057 , n427895 );
buf ( n428058 , n427616 );
xor ( n82005 , n428057 , n428058 );
buf ( n428060 , n427620 );
xnor ( n82007 , n82005 , n428060 );
buf ( n428062 , n82007 );
buf ( n428063 , n428062 );
buf ( n428064 , n427625 );
buf ( n428065 , n81760 );
xor ( n82012 , n428064 , n428065 );
buf ( n428067 , n427889 );
xnor ( n82014 , n82012 , n428067 );
buf ( n428069 , n82014 );
buf ( n428070 , n428069 );
buf ( n428071 , C1 );
buf ( n428072 , n428071 );
xor ( n82040 , n81542 , n81539 );
xor ( n82041 , n82040 , n81758 );
buf ( n428075 , n82041 );
xor ( n82043 , n428072 , n428075 );
buf ( n428077 , C1 );
nand ( n82072 , n51553 , n427642 );
nand ( n82073 , n427743 , n50579 );
and ( n82074 , n82072 , n82073 );
nand ( n82077 , n428077 , n82074 );
buf ( n428082 , n43535 );
not ( n82079 , n428082 );
buf ( n428084 , n400042 );
buf ( n428085 , n388064 );
and ( n82082 , n428084 , n428085 );
not ( n82083 , n428084 );
buf ( n428088 , n425525 );
and ( n82085 , n82083 , n428088 );
nor ( n82086 , n82082 , n82085 );
buf ( n428091 , n82086 );
buf ( n428092 , n428091 );
not ( n82089 , n428092 );
and ( n82090 , n82079 , n82089 );
buf ( n428095 , n427847 );
buf ( n428096 , n43514 );
nor ( n82093 , n428095 , n428096 );
buf ( n428098 , n82093 );
buf ( n428099 , n428098 );
nor ( n82096 , n82090 , n428099 );
buf ( n428101 , n82096 );
buf ( n428102 , n428101 );
not ( n82099 , n428102 );
buf ( n428104 , n82099 );
not ( n82101 , n428104 );
buf ( n428106 , n70210 );
buf ( n428107 , n62499 );
and ( n82104 , n428106 , n428107 );
buf ( n428109 , n416845 );
buf ( n428110 , n410717 );
and ( n82107 , n428109 , n428110 );
nor ( n82108 , n82104 , n82107 );
buf ( n428113 , n82108 );
buf ( n428114 , n428113 );
buf ( n428115 , n410724 );
or ( n82112 , n428114 , n428115 );
buf ( n428117 , n426940 );
buf ( n428118 , n410721 );
or ( n82115 , n428117 , n428118 );
nand ( n82116 , n82112 , n82115 );
buf ( n428121 , n82116 );
xor ( n82118 , n426901 , n426917 );
xor ( n82119 , n82118 , n426927 );
and ( n82120 , n428121 , n82119 );
buf ( n428125 , n409429 );
buf ( n428126 , n59463 );
buf ( n428127 , n71681 );
and ( n82124 , n428126 , n428127 );
buf ( n428129 , n62159 );
buf ( n428130 , n418315 );
and ( n82127 , n428129 , n428130 );
nor ( n82128 , n82124 , n82127 );
buf ( n428133 , n82128 );
buf ( n428134 , n428133 );
or ( n82131 , n428125 , n428134 );
buf ( n428136 , n426997 );
buf ( n428137 , n409170 );
or ( n82134 , n428136 , n428137 );
nand ( n82135 , n82131 , n82134 );
buf ( n428140 , n82135 );
buf ( n428141 , n428140 );
buf ( n428142 , n58218 );
buf ( n428143 , n623 );
and ( n82140 , n428142 , n428143 );
buf ( n428145 , n13935 );
buf ( n428146 , n422315 );
and ( n82143 , n428145 , n428146 );
buf ( n428148 , n14083 );
nor ( n82145 , n82143 , n428148 );
buf ( n428150 , n82145 );
buf ( n428151 , n428150 );
buf ( n428152 , n405391 );
nor ( n82149 , n82140 , n428151 , n428152 );
buf ( n428154 , n82149 );
buf ( n428155 , n428154 );
xor ( n82152 , n428141 , n428155 );
buf ( n428157 , n59637 );
buf ( n428158 , n59628 );
buf ( n428159 , n74002 );
and ( n82156 , n428158 , n428159 );
buf ( n428161 , n59457 );
buf ( n428162 , n420612 );
and ( n82159 , n428161 , n428162 );
nor ( n82160 , n82156 , n82159 );
buf ( n428165 , n82160 );
buf ( n428166 , n428165 );
or ( n82163 , n428157 , n428166 );
buf ( n428168 , n426891 );
buf ( n428169 , n59467 );
or ( n82166 , n428168 , n428169 );
nand ( n82167 , n82163 , n82166 );
buf ( n428172 , n82167 );
buf ( n428173 , n428172 );
and ( n82170 , n82152 , n428173 );
and ( n82171 , n428141 , n428155 );
or ( n82172 , n82170 , n82171 );
buf ( n428177 , n82172 );
buf ( n428178 , n428177 );
xor ( n82175 , n426882 , n426899 );
buf ( n428180 , n82175 );
buf ( n428181 , n428180 );
xor ( n82178 , n428178 , n428181 );
buf ( n428183 , n71170 );
buf ( n428184 , n63625 );
and ( n82181 , n428183 , n428184 );
buf ( n428186 , n417804 );
buf ( n428187 , n62511 );
and ( n82184 , n428186 , n428187 );
nor ( n82185 , n82181 , n82184 );
buf ( n428190 , n82185 );
buf ( n428191 , n428190 );
buf ( n428192 , n410635 );
or ( n82189 , n428191 , n428192 );
buf ( n428194 , n427015 );
buf ( n428195 , n409504 );
or ( n428196 , n428194 , n428195 );
nand ( n82193 , n82189 , n428196 );
buf ( n428198 , n82193 );
buf ( n428199 , n428198 );
buf ( n428200 , n405384 );
buf ( n428201 , n422315 );
nor ( n82198 , n428200 , n428201 );
buf ( n428203 , n82198 );
buf ( n428204 , n428203 );
buf ( n428205 , n71664 );
buf ( n428206 , n62164 );
and ( n82203 , n428205 , n428206 );
buf ( n428208 , n418298 );
buf ( n428209 , n62511 );
and ( n82206 , n428208 , n428209 );
nor ( n82207 , n82203 , n82206 );
buf ( n428212 , n82207 );
buf ( n428213 , n428212 );
buf ( n428214 , n410635 );
or ( n82211 , n428213 , n428214 );
buf ( n428216 , n428190 );
buf ( n428217 , n409504 );
or ( n82214 , n428216 , n428217 );
nand ( n82215 , n82211 , n82214 );
buf ( n428220 , n82215 );
buf ( n428221 , n428220 );
and ( n82218 , n428204 , n428221 );
buf ( n428223 , n82218 );
buf ( n428224 , n428223 );
xor ( n82221 , n428199 , n428224 );
buf ( n428226 , n405414 );
buf ( n428227 , n623 );
or ( n82224 , n428226 , n428227 );
buf ( n428229 , n405410 );
buf ( n428230 , n405391 );
buf ( n428231 , n623 );
and ( n82228 , n428229 , n428230 , n428231 );
buf ( n428233 , n405394 );
nor ( n82230 , n82228 , n428233 );
buf ( n428235 , n82230 );
buf ( n428236 , n428235 );
nand ( n82233 , n82224 , n428236 );
buf ( n428238 , n82233 );
buf ( n428239 , n428238 );
and ( n82236 , n82221 , n428239 );
and ( n82237 , n428199 , n428224 );
or ( n82238 , n82236 , n82237 );
buf ( n428243 , n82238 );
buf ( n428244 , n428243 );
and ( n82241 , n82178 , n428244 );
and ( n82242 , n428178 , n428181 );
or ( n82243 , n82241 , n82242 );
buf ( n428248 , n82243 );
xor ( n82245 , n426901 , n426917 );
xor ( n82246 , n82245 , n426927 );
and ( n82247 , n428248 , n82246 );
and ( n82248 , n428121 , n428248 );
or ( n82249 , n82120 , n82247 , n82248 );
xor ( n82250 , n426963 , n80843 );
xor ( n82251 , n82250 , n427037 );
and ( n82252 , n82249 , n82251 );
xor ( n82253 , n426989 , n427006 );
xor ( n82254 , n82253 , n427024 );
buf ( n428259 , n82254 );
buf ( n428260 , n70389 );
buf ( n428261 , n62499 );
and ( n82258 , n428260 , n428261 );
buf ( n428263 , n417024 );
buf ( n428264 , n62496 );
and ( n82261 , n428263 , n428264 );
nor ( n82262 , n82258 , n82261 );
buf ( n428267 , n82262 );
buf ( n428268 , n428267 );
buf ( n428269 , n410724 );
or ( n82266 , n428268 , n428269 );
buf ( n428271 , n428113 );
buf ( n428272 , n410721 );
or ( n82269 , n428271 , n428272 );
nand ( n82270 , n82266 , n82269 );
buf ( n428275 , n82270 );
xor ( n82272 , n428259 , n428275 );
buf ( n428277 , n71095 );
buf ( n428278 , n62499 );
and ( n82275 , n428277 , n428278 );
buf ( n428280 , n417729 );
buf ( n428281 , n62496 );
and ( n82278 , n428280 , n428281 );
nor ( n82279 , n82275 , n82278 );
buf ( n428284 , n82279 );
buf ( n428285 , n428284 );
buf ( n428286 , n410724 );
or ( n82283 , n428285 , n428286 );
buf ( n428288 , n428267 );
buf ( n428289 , n410721 );
or ( n82286 , n428288 , n428289 );
nand ( n82287 , n82283 , n82286 );
buf ( n428292 , n82287 );
buf ( n428293 , n428292 );
xor ( n82290 , n428141 , n428155 );
xor ( n82291 , n82290 , n428173 );
buf ( n428296 , n82291 );
buf ( n428297 , n428296 );
xor ( n82294 , n428293 , n428297 );
buf ( n428299 , n428165 );
buf ( n428300 , n59467 );
or ( n82297 , n428299 , n428300 );
buf ( n428302 , n59469 );
nand ( n82299 , n82297 , n428302 );
buf ( n428304 , n82299 );
buf ( n428305 , n428304 );
buf ( n428306 , n409429 );
buf ( n428307 , n62177 );
buf ( n428308 , n72308 );
and ( n82305 , n428307 , n428308 );
buf ( n428310 , n62159 );
buf ( n428311 , n418942 );
and ( n82308 , n428310 , n428311 );
nor ( n82309 , n82305 , n82308 );
buf ( n428314 , n82309 );
buf ( n428315 , n428314 );
or ( n82312 , n428306 , n428315 );
buf ( n428317 , n428133 );
buf ( n428318 , n409170 );
or ( n82315 , n428317 , n428318 );
nand ( n82316 , n82312 , n82315 );
buf ( n428321 , n82316 );
buf ( n428322 , n428321 );
xor ( n82319 , n428305 , n428322 );
xor ( n82320 , n428204 , n428221 );
buf ( n428325 , n82320 );
buf ( n428326 , n428325 );
and ( n82323 , n82319 , n428326 );
and ( n82324 , n428305 , n428322 );
or ( n82325 , n82323 , n82324 );
buf ( n428330 , n82325 );
buf ( n428331 , n428330 );
and ( n82328 , n82294 , n428331 );
and ( n82329 , n428293 , n428297 );
or ( n82330 , n82328 , n82329 );
buf ( n428335 , n82330 );
and ( n82332 , n82272 , n428335 );
and ( n82333 , n428259 , n428275 );
or ( n82334 , n82332 , n82333 );
buf ( n428339 , n82334 );
xor ( n82336 , n426811 , n426825 );
xor ( n82337 , n82336 , n426842 );
xor ( n82338 , n426979 , n427028 );
xor ( n82339 , n82337 , n82338 );
buf ( n428344 , n82339 );
xor ( n82341 , n428339 , n428344 );
xor ( n82342 , n426901 , n426917 );
xor ( n82343 , n82342 , n426927 );
xor ( n82344 , n428121 , n428248 );
xor ( n82345 , n82343 , n82344 );
buf ( n428350 , n82345 );
and ( n82347 , n82341 , n428350 );
and ( n82348 , n428339 , n428344 );
or ( n82349 , n82347 , n82348 );
buf ( n428354 , n82349 );
xor ( n82351 , n426963 , n80843 );
xor ( n82352 , n82351 , n427037 );
and ( n82353 , n428354 , n82352 );
and ( n82354 , n82249 , n428354 );
or ( n82355 , n82252 , n82353 , n82354 );
buf ( n428360 , n82355 );
xor ( n82357 , n427041 , n427046 );
xor ( n82358 , n82357 , n427051 );
buf ( n428363 , n82358 );
buf ( n428364 , n428363 );
xor ( n82361 , n428360 , n428364 );
buf ( n428366 , n55543 );
not ( n82363 , n428366 );
buf ( n428368 , n426763 );
not ( n82365 , n428368 );
or ( n82366 , n82363 , n82365 );
buf ( n428371 , n392217 );
buf ( n428372 , n51185 );
nand ( n82369 , n428371 , n428372 );
buf ( n428374 , n82369 );
buf ( n428375 , n428374 );
nand ( n82372 , n82366 , n428375 );
buf ( n428377 , n82372 );
buf ( n428378 , n428377 );
not ( n82375 , n428378 );
buf ( n428380 , n427074 );
not ( n82377 , n428380 );
or ( n82378 , n82375 , n82377 );
buf ( n428383 , n427673 );
buf ( n428384 , n426775 );
nand ( n82381 , n428383 , n428384 );
buf ( n428386 , n82381 );
buf ( n428387 , n428386 );
nand ( n82384 , n82378 , n428387 );
buf ( n428389 , n82384 );
buf ( n428390 , n428389 );
and ( n82387 , n82361 , n428390 );
and ( n82388 , n428360 , n428364 );
or ( n82389 , n82387 , n82388 );
buf ( n428394 , n82389 );
not ( n82391 , n428394 );
buf ( n428396 , n392221 );
not ( n82393 , n428396 );
buf ( n428398 , n427821 );
not ( n82395 , n428398 );
or ( n82396 , n82393 , n82395 );
buf ( n428401 , n44770 );
buf ( n428402 , n399274 );
not ( n82399 , n428402 );
buf ( n428404 , n390985 );
not ( n82401 , n428404 );
or ( n82402 , n82399 , n82401 );
buf ( n428407 , n44775 );
buf ( n428408 , n399283 );
nand ( n82405 , n428407 , n428408 );
buf ( n428410 , n82405 );
buf ( n428411 , n428410 );
nand ( n82408 , n82402 , n428411 );
buf ( n428413 , n82408 );
buf ( n428414 , n428413 );
nand ( n82411 , n428401 , n428414 );
buf ( n428416 , n82411 );
buf ( n428417 , n428416 );
nand ( n82414 , n82396 , n428417 );
buf ( n428419 , n82414 );
buf ( n428420 , n428419 );
not ( n82417 , n428420 );
buf ( n428422 , n82417 );
nand ( n82419 , n82391 , n428422 );
not ( n82420 , n82419 );
xor ( n82421 , n427661 , n427686 );
xor ( n82422 , n82421 , n427724 );
buf ( n428427 , n82422 );
not ( n82424 , n428427 );
or ( n82425 , n82420 , n82424 );
buf ( n428430 , n428394 );
buf ( n428431 , n428419 );
nand ( n82428 , n428430 , n428431 );
buf ( n428433 , n82428 );
nand ( n82430 , n82425 , n428433 );
not ( n82431 , n82430 );
or ( n82432 , n82101 , n82431 );
buf ( n428437 , n82430 );
not ( n82434 , n428437 );
buf ( n428439 , n82434 );
not ( n82436 , n428439 );
not ( n82437 , n428101 );
or ( n82438 , n82436 , n82437 );
xor ( n82439 , n427795 , n427808 );
xor ( n82440 , n82439 , n427834 );
buf ( n428445 , n82440 );
nand ( n82442 , n82438 , n428445 );
nand ( n82443 , n82432 , n82442 );
and ( n82444 , n82077 , n82443 );
nor ( n82445 , C0 , n82444 );
buf ( n428450 , n82445 );
and ( n82447 , n82043 , n428450 );
and ( n82448 , n428072 , n428075 );
or ( n82449 , n82447 , n82448 );
buf ( n428454 , n82449 );
buf ( n428455 , n428454 );
xor ( n82452 , n428070 , n428455 );
buf ( n428457 , C1 );
buf ( n428458 , n428457 );
and ( n82466 , n82452 , n428458 );
and ( n82467 , n428070 , n428455 );
or ( n82468 , n82466 , n82467 );
buf ( n428462 , n82468 );
buf ( n428463 , n428462 );
or ( n82471 , n428063 , n428463 );
buf ( n428465 , n428032 );
buf ( n428466 , n427940 );
xor ( n82474 , n428465 , n428466 );
buf ( n428468 , C0 );
xnor ( n82476 , n82474 , n428468 );
buf ( n428470 , n82476 );
buf ( n428471 , n428470 );
buf ( n428472 , n428462 );
buf ( n428473 , n428062 );
and ( n82481 , n428472 , n428473 );
buf ( n428475 , n82481 );
buf ( n428476 , n428475 );
or ( n82484 , n428471 , n428476 );
nand ( n82485 , n82471 , n82484 );
buf ( n428479 , n82485 );
buf ( n428480 , n428479 );
xor ( n82488 , n427937 , n428041 );
xor ( n82489 , n82488 , n428046 );
buf ( n428483 , n82489 );
buf ( n428484 , n428483 );
xor ( n82492 , n428480 , n428484 );
xor ( n82493 , C1 , n427947 );
xor ( n82494 , n82493 , n428026 );
buf ( n428488 , n82494 );
not ( n82496 , n428488 );
xor ( n82497 , n428070 , n428455 );
xor ( n82498 , n82497 , n428458 );
buf ( n428492 , n82498 );
buf ( n428493 , n428492 );
not ( n82501 , n428493 );
or ( n82502 , n82496 , n82501 );
buf ( n428496 , C0 );
not ( n82518 , n427969 );
not ( n82519 , n388068 );
or ( n82520 , n82518 , n82519 );
nand ( n82521 , n421024 , n358975 );
not ( n82522 , n82521 );
buf ( n428502 , n388722 );
buf ( n428503 , n402819 );
nand ( n82525 , n428502 , n428503 );
buf ( n428505 , n82525 );
not ( n82527 , n428505 );
or ( n82528 , n82522 , n82527 );
nand ( n82529 , n82528 , n67042 );
nand ( n82530 , n82520 , n82529 );
buf ( n428510 , n82530 );
buf ( n428511 , n427716 );
not ( n82533 , n428511 );
buf ( n428513 , n395359 );
not ( n82535 , n428513 );
or ( n82536 , n82533 , n82535 );
buf ( n428516 , n81579 );
not ( n82538 , n428516 );
buf ( n428518 , n24790 );
not ( n82540 , n428518 );
buf ( n428520 , n82540 );
buf ( n428521 , n428520 );
not ( n82543 , n428521 );
or ( n82544 , n82538 , n82543 );
buf ( n428524 , n427698 );
buf ( n428525 , n24790 );
nand ( n82547 , n428524 , n428525 );
buf ( n428527 , n82547 );
buf ( n428528 , n428527 );
nand ( n82550 , n82544 , n428528 );
buf ( n428530 , n82550 );
buf ( n428531 , n428530 );
buf ( n428532 , n395346 );
nand ( n82554 , n428531 , n428532 );
buf ( n428534 , n82554 );
buf ( n428535 , n428534 );
nand ( n82557 , n82536 , n428535 );
buf ( n428537 , n82557 );
buf ( n428538 , n428537 );
xor ( n82560 , n426963 , n80843 );
xor ( n82561 , n82560 , n427037 );
xor ( n82562 , n82249 , n428354 );
xor ( n82563 , n82561 , n82562 );
buf ( n428543 , n82563 );
buf ( n428544 , n395359 );
not ( n82566 , n428544 );
buf ( n428546 , n428530 );
not ( n82568 , n428546 );
or ( n82569 , n82566 , n82568 );
buf ( n428549 , n395346 );
buf ( n428550 , n427308 );
not ( n82572 , n428550 );
buf ( n428552 , n393397 );
not ( n82574 , n428552 );
or ( n82575 , n82572 , n82574 );
buf ( n428555 , n397486 );
buf ( n428556 , n23604 );
nand ( n82578 , n428555 , n428556 );
buf ( n428558 , n82578 );
buf ( n428559 , n428558 );
nand ( n82581 , n82575 , n428559 );
buf ( n428561 , n82581 );
buf ( n428562 , n428561 );
nand ( n82584 , n428549 , n428562 );
buf ( n428564 , n82584 );
buf ( n428565 , n428564 );
nand ( n82587 , n82569 , n428565 );
buf ( n428567 , n82587 );
buf ( n428568 , n428567 );
xor ( n82590 , n428543 , n428568 );
xor ( n82591 , n428178 , n428181 );
xor ( n82592 , n82591 , n428244 );
buf ( n428572 , n82592 );
xor ( n82594 , n428259 , n428275 );
xor ( n82595 , n82594 , n428335 );
and ( n82596 , n428572 , n82595 );
buf ( n428576 , n71088 );
buf ( n428577 , n62499 );
and ( n82599 , n428576 , n428577 );
buf ( n428579 , n417722 );
buf ( n428580 , n410717 );
and ( n82602 , n428579 , n428580 );
nor ( n82603 , n82599 , n82602 );
buf ( n428583 , n82603 );
buf ( n428584 , n428583 );
buf ( n428585 , n410724 );
or ( n82607 , n428584 , n428585 );
buf ( n428587 , n428284 );
buf ( n428588 , n410721 );
or ( n82610 , n428587 , n428588 );
nand ( n82611 , n82607 , n82610 );
buf ( n428591 , n82611 );
buf ( n428592 , n59451 );
buf ( n428593 , n623 );
and ( n82615 , n428592 , n428593 );
buf ( n428595 , n406581 );
buf ( n428596 , n422315 );
and ( n82618 , n428595 , n428596 );
buf ( n428598 , n62177 );
nor ( n82620 , n82618 , n428598 );
buf ( n428600 , n82620 );
buf ( n428601 , n428600 );
buf ( n428602 , n14083 );
nor ( n82624 , n82615 , n428601 , n428602 );
buf ( n428604 , n82624 );
buf ( n428605 , n428604 );
buf ( n428606 , n410635 );
buf ( n428607 , n62164 );
buf ( n428608 , n71681 );
and ( n82630 , n428607 , n428608 );
buf ( n428610 , n418315 );
buf ( n428611 , n62511 );
and ( n82633 , n428610 , n428611 );
nor ( n82634 , n82630 , n82633 );
buf ( n428614 , n82634 );
buf ( n428615 , n428614 );
or ( n82637 , n428606 , n428615 );
buf ( n428617 , n428212 );
buf ( n428618 , n409504 );
or ( n82640 , n428617 , n428618 );
nand ( n82641 , n82637 , n82640 );
buf ( n428621 , n82641 );
buf ( n428622 , n428621 );
xor ( n82644 , n428605 , n428622 );
buf ( n428624 , n410635 );
buf ( n428625 , n62164 );
buf ( n428626 , n72308 );
and ( n82648 , n428625 , n428626 );
buf ( n428628 , n62511 );
buf ( n428629 , n418942 );
and ( n82651 , n428628 , n428629 );
nor ( n82652 , n82648 , n82651 );
buf ( n428632 , n82652 );
buf ( n428633 , n428632 );
or ( n82655 , n428624 , n428633 );
buf ( n428635 , n428614 );
buf ( n428636 , n409504 );
or ( n82658 , n428635 , n428636 );
nand ( n82659 , n82655 , n82658 );
buf ( n428639 , n82659 );
buf ( n428640 , n428639 );
buf ( n428641 , n59467 );
buf ( n428642 , n422315 );
nor ( n82664 , n428641 , n428642 );
buf ( n428644 , n82664 );
buf ( n428645 , n428644 );
and ( n82667 , n428640 , n428645 );
buf ( n428647 , n82667 );
buf ( n428648 , n428647 );
and ( n82670 , n82644 , n428648 );
and ( n82671 , n428605 , n428622 );
or ( n82672 , n82670 , n82671 );
buf ( n428652 , n82672 );
xor ( n82674 , n428591 , n428652 );
xor ( n82675 , n428305 , n428322 );
xor ( n82676 , n82675 , n428326 );
buf ( n428656 , n82676 );
and ( n82678 , n82674 , n428656 );
and ( n82679 , n428591 , n428652 );
or ( n82680 , n82678 , n82679 );
buf ( n428660 , n82680 );
xor ( n82682 , n428199 , n428224 );
xor ( n82683 , n82682 , n428239 );
buf ( n428663 , n82683 );
buf ( n428664 , n428663 );
xor ( n82686 , n428660 , n428664 );
xor ( n82687 , n428293 , n428297 );
xor ( n82688 , n82687 , n428331 );
buf ( n428668 , n82688 );
buf ( n428669 , n428668 );
and ( n82691 , n82686 , n428669 );
and ( n82692 , n428660 , n428664 );
or ( n82693 , n82691 , n82692 );
buf ( n428673 , n82693 );
xor ( n82695 , n428259 , n428275 );
xor ( n82696 , n82695 , n428335 );
and ( n82697 , n428673 , n82696 );
and ( n82698 , n428572 , n428673 );
or ( n82699 , n82596 , n82697 , n82698 );
buf ( n428679 , n82699 );
xor ( n82701 , n428339 , n428344 );
xor ( n82702 , n82701 , n428350 );
buf ( n428682 , n82702 );
buf ( n428683 , n428682 );
xor ( n82705 , n428679 , n428683 );
buf ( n428685 , n47903 );
not ( n82707 , n428685 );
nand ( n82708 , n51175 , n51178 , n51179 , n51182 );
buf ( n428688 , n82708 );
not ( n82710 , n428688 );
buf ( n428690 , n393397 );
not ( n82712 , n428690 );
or ( n82713 , n82710 , n82712 );
buf ( n428693 , n51184 );
buf ( n428694 , n23604 );
nand ( n82716 , n428693 , n428694 );
buf ( n428696 , n82716 );
buf ( n428697 , n428696 );
nand ( n82719 , n82713 , n428697 );
buf ( n428699 , n82719 );
buf ( n428700 , n428699 );
not ( n82722 , n428700 );
or ( n82723 , n82707 , n82722 );
buf ( n428703 , n428561 );
buf ( n428704 , n395359 );
nand ( n82726 , n428703 , n428704 );
buf ( n428706 , n82726 );
buf ( n428707 , n428706 );
nand ( n82729 , n82723 , n428707 );
buf ( n428709 , n82729 );
buf ( n428710 , n428709 );
and ( n82732 , n82705 , n428710 );
and ( n82733 , n428679 , n428683 );
or ( n82734 , n82732 , n82733 );
buf ( n428714 , n82734 );
buf ( n428715 , n428714 );
and ( n82737 , n82590 , n428715 );
and ( n82738 , n428543 , n428568 );
or ( n82739 , n82737 , n82738 );
buf ( n428719 , n82739 );
buf ( n428720 , n428719 );
xor ( n82742 , n428538 , n428720 );
xor ( n82743 , n428360 , n428364 );
xor ( n82744 , n82743 , n428390 );
buf ( n428724 , n82744 );
buf ( n428725 , n428724 );
and ( n82747 , n82742 , n428725 );
and ( n82748 , n428538 , n428720 );
or ( n82749 , n82747 , n82748 );
buf ( n428729 , n82749 );
buf ( n428730 , n428729 );
buf ( n428731 , n51553 );
not ( n82753 , n428731 );
buf ( n428733 , n427758 );
not ( n82755 , n428733 );
or ( n82756 , n82753 , n82755 );
buf ( n428736 , n47891 );
not ( n82758 , n428736 );
buf ( n428738 , n392878 );
not ( n82760 , n428738 );
or ( n82761 , n82758 , n82760 );
buf ( n428741 , n24841 );
buf ( n428742 , n61299 );
nand ( n82764 , n428741 , n428742 );
buf ( n428744 , n82764 );
buf ( n428745 , n428744 );
nand ( n82767 , n82761 , n428745 );
buf ( n428747 , n82767 );
buf ( n428748 , n428747 );
buf ( n428749 , n50579 );
nand ( n82771 , n428748 , n428749 );
buf ( n428751 , n82771 );
buf ( n428752 , n428751 );
nand ( n82774 , n82756 , n428752 );
buf ( n428754 , n82774 );
buf ( n428755 , n428754 );
xor ( n82777 , n428730 , n428755 );
buf ( n428757 , n40567 );
buf ( n428758 , n402819 );
nor ( n82780 , n428757 , n428758 );
buf ( n428760 , n82780 );
buf ( n428761 , n428760 );
and ( n82783 , n82777 , n428761 );
and ( n82784 , n428730 , n428755 );
or ( n82785 , n82783 , n82784 );
buf ( n428765 , n82785 );
buf ( n428766 , n428765 );
xor ( n82788 , n428510 , n428766 );
not ( n82789 , n55055 );
not ( n82790 , n420986 );
or ( n82791 , n82789 , n82790 );
buf ( n428771 , n390997 );
buf ( n428772 , n55054 );
nand ( n82794 , n428771 , n428772 );
buf ( n428774 , n82794 );
nand ( n82796 , n82791 , n428774 );
not ( n82797 , n82796 );
not ( n82798 , n74375 );
or ( n82799 , n82797 , n82798 );
buf ( n428779 , n428091 );
not ( n82801 , n428779 );
buf ( n428781 , n43515 );
nand ( n82803 , n82801 , n428781 );
buf ( n428783 , n82803 );
nand ( n82805 , n82799 , n428783 );
buf ( n428785 , n82805 );
buf ( n428786 , n51553 );
not ( n82808 , n428786 );
buf ( n428788 , n428747 );
not ( n82810 , n428788 );
or ( n82811 , n82808 , n82810 );
and ( n82812 , n394207 , n47891 );
not ( n82813 , n394207 );
and ( n82814 , n82813 , n61299 );
or ( n82815 , n82812 , n82814 );
buf ( n428795 , n82815 );
buf ( n428796 , n50579 );
nand ( n82818 , n428795 , n428796 );
buf ( n428798 , n82818 );
buf ( n428799 , n428798 );
nand ( n82821 , n82811 , n428799 );
buf ( n428801 , n82821 );
buf ( n428802 , n428801 );
buf ( n428803 , n400033 );
not ( n82825 , n428803 );
buf ( n428805 , n422673 );
not ( n82827 , n428805 );
or ( n82828 , n82825 , n82827 );
buf ( n428808 , n390988 );
buf ( n428809 , n400042 );
nand ( n82831 , n428808 , n428809 );
buf ( n428811 , n82831 );
buf ( n428812 , n428811 );
nand ( n82834 , n82828 , n428812 );
buf ( n428814 , n82834 );
buf ( n428815 , n428814 );
not ( n82837 , n428815 );
buf ( n428817 , n44770 );
not ( n82839 , n428817 );
or ( n82840 , n82837 , n82839 );
buf ( n428820 , n428413 );
buf ( n428821 , n413643 );
nand ( n82843 , n428820 , n428821 );
buf ( n428823 , n82843 );
buf ( n428824 , n428823 );
nand ( n82846 , n82840 , n428824 );
buf ( n428826 , n82846 );
buf ( n428827 , n428826 );
xor ( n82849 , n428802 , n428827 );
buf ( n428829 , n371876 );
nor ( n82851 , n44775 , n23723 );
or ( n82852 , n82851 , n402819 );
buf ( n428832 , n44775 );
buf ( n428833 , n23723 );
nand ( n82855 , n428832 , n428833 );
buf ( n428835 , n82855 );
nand ( n82857 , n82852 , n428835 );
buf ( n428837 , n82857 );
nor ( n82859 , n428829 , n428837 );
buf ( n428839 , n82859 );
buf ( n428840 , n428839 );
and ( n82862 , n82849 , n428840 );
and ( n82863 , n428802 , n428827 );
or ( n82864 , n82862 , n82863 );
buf ( n428844 , n82864 );
buf ( n428845 , n428844 );
or ( n82867 , n428785 , n428845 );
xor ( n82868 , n428394 , n428422 );
xor ( n82869 , n82868 , n428427 );
buf ( n428849 , n82869 );
not ( n82871 , n428849 );
buf ( n428851 , n82871 );
buf ( n428852 , n428851 );
nand ( n82874 , n82867 , n428852 );
buf ( n428854 , n82874 );
buf ( n428855 , n428854 );
buf ( n428856 , n82805 );
buf ( n428857 , n428844 );
nand ( n82879 , n428856 , n428857 );
buf ( n428859 , n82879 );
buf ( n428860 , n428859 );
nand ( n82882 , n428855 , n428860 );
buf ( n428862 , n82882 );
buf ( n428863 , n428862 );
and ( n82885 , n82788 , n428863 );
and ( n82886 , n428510 , n428766 );
or ( n82887 , n82885 , n82886 );
buf ( n428867 , n82887 );
not ( n82889 , n428867 );
not ( n82890 , n427838 );
not ( n82891 , n81752 );
and ( n82892 , n82890 , n82891 );
and ( n82893 , n427838 , n81752 );
nor ( n82894 , n82892 , n82893 );
not ( n82895 , n427790 );
and ( n82896 , n82894 , n82895 );
not ( n82897 , n82894 );
and ( n82898 , n82897 , n427790 );
nor ( n82899 , n82896 , n82898 );
not ( n82900 , n82899 );
nand ( n82901 , n82889 , n82900 );
not ( n82902 , n82901 );
xor ( n82903 , n427957 , n427982 );
xor ( n82904 , n82903 , n427988 );
buf ( n428884 , n82904 );
not ( n82906 , n428884 );
or ( n82907 , n82902 , n82906 );
not ( n82908 , n82900 );
nand ( n82909 , n82908 , n428867 );
nand ( n82910 , n82907 , n82909 );
buf ( n428890 , n428496 );
buf ( n428891 , n82910 );
or ( n82915 , n428890 , n428891 );
xor ( n82916 , n427993 , n428014 );
xor ( n82917 , n82916 , n428022 );
buf ( n428895 , n82917 );
buf ( n428896 , n428895 );
nand ( n82920 , n82915 , n428896 );
buf ( n428898 , n82920 );
nand ( n82922 , C1 , n428898 );
buf ( n428900 , n82922 );
nand ( n82924 , n82502 , n428900 );
buf ( n428902 , n82924 );
buf ( n428903 , n428902 );
not ( n82927 , n428492 );
buf ( n428905 , n82494 );
not ( n82929 , n428905 );
buf ( n428907 , n82929 );
nand ( n82931 , n82927 , n428907 );
buf ( n428909 , n82931 );
nand ( n82933 , n428903 , n428909 );
buf ( n428911 , n82933 );
buf ( n428912 , n428911 );
not ( n82936 , n428912 );
buf ( n428914 , n428470 );
not ( n82938 , n428914 );
xor ( n82939 , n428472 , n428473 );
buf ( n428917 , n82939 );
buf ( n428918 , n428917 );
not ( n82942 , n428918 );
and ( n82943 , n82938 , n82942 );
buf ( n428921 , n428470 );
buf ( n428922 , n428917 );
and ( n82946 , n428921 , n428922 );
nor ( n82947 , n82943 , n82946 );
buf ( n428925 , n82947 );
buf ( n428926 , n428925 );
nand ( n82950 , n82936 , n428926 );
buf ( n428928 , n82950 );
not ( n82952 , n428928 );
buf ( n428930 , n82910 );
buf ( n428931 , n428895 );
xor ( n82955 , n428930 , n428931 );
buf ( n428933 , n428496 );
xnor ( n82957 , n82955 , n428933 );
buf ( n428935 , n82957 );
buf ( n428936 , n428935 );
xor ( n82960 , n428072 , n428075 );
xor ( n82961 , n82960 , n428450 );
buf ( n428939 , n82961 );
buf ( n428940 , n428939 );
or ( n82964 , n428936 , n428940 );
buf ( n428942 , n82964 );
buf ( n428943 , n428942 );
buf ( n428944 , n428939 );
not ( n82968 , n428944 );
buf ( n428946 , n428935 );
not ( n82970 , n428946 );
or ( n82971 , n82968 , n82970 );
xor ( n82972 , n427729 , n427766 );
xor ( n82973 , n82972 , n427786 );
buf ( n428951 , n82973 );
buf ( n428952 , n428951 );
buf ( n428953 , C0 );
buf ( n428954 , n428953 );
xor ( n82990 , n428952 , n428954 );
buf ( n428956 , n82430 );
buf ( n428957 , n428445 );
xor ( n82993 , n428956 , n428957 );
buf ( n428959 , n428104 );
xor ( n82995 , n82993 , n428959 );
buf ( n428961 , n82995 );
buf ( n428962 , n428961 );
and ( n82998 , n82990 , n428962 );
or ( n83000 , n82998 , C0 );
buf ( n428965 , n83000 );
buf ( n428966 , n428965 );
not ( n83004 , n82074 );
not ( n83005 , n83004 );
not ( n83006 , n82443 );
or ( n83007 , n83005 , n83006 );
or ( n83008 , n82443 , n83004 );
nand ( n83009 , n83007 , n83008 );
not ( n83010 , n83009 );
not ( n83011 , n83010 );
or ( n83012 , C0 , n83011 );
nand ( n83014 , n83012 , C1 );
buf ( n428977 , n83014 );
buf ( n428978 , C0 );
buf ( n428979 , n428978 );
and ( n83030 , n428966 , n428977 );
or ( n83031 , C0 , n83030 );
buf ( n428982 , n83031 );
buf ( n428983 , n428982 );
nand ( n83034 , n82971 , n428983 );
buf ( n428985 , n83034 );
buf ( n428986 , n428985 );
and ( n83037 , n428943 , n428986 );
buf ( n428988 , n83037 );
buf ( n428989 , n428988 );
and ( n83040 , n82922 , n82494 );
not ( n83041 , n82922 );
and ( n83042 , n83041 , n428907 );
or ( n83043 , n83040 , n83042 );
xor ( n83044 , n83043 , n428492 );
buf ( n428995 , n83044 );
and ( n83046 , n428989 , n428995 );
buf ( n428997 , n83046 );
xnor ( n83048 , n428939 , n428982 );
xnor ( n83049 , n83048 , n428935 );
buf ( n429000 , n83049 );
buf ( n429001 , C0 );
buf ( n429002 , n429001 );
xor ( n83076 , n428538 , n428720 );
xor ( n83077 , n83076 , n428725 );
buf ( n429005 , n83077 );
buf ( n429006 , n429005 );
and ( n83080 , n399274 , n426763 );
not ( n83081 , n399274 );
and ( n83082 , n83081 , n392217 );
or ( n83083 , n83080 , n83082 );
buf ( n429011 , n83083 );
not ( n83085 , n429011 );
buf ( n429013 , n83085 );
or ( n83087 , n429013 , n45948 );
buf ( n429015 , n428377 );
not ( n83089 , n429015 );
buf ( n429017 , n83089 );
or ( n83091 , n429017 , n45947 );
nand ( n83092 , n83087 , n83091 );
buf ( n429020 , n83092 );
xor ( n83094 , n428543 , n428568 );
xor ( n83095 , n83094 , n428715 );
buf ( n429023 , n83095 );
buf ( n429024 , n429023 );
xor ( n83098 , n429020 , n429024 );
buf ( n429026 , n59916 );
not ( n83100 , n429026 );
buf ( n429028 , n82815 );
not ( n83102 , n429028 );
or ( n83103 , n83100 , n83102 );
and ( n83104 , n47891 , n394814 );
not ( n83105 , n47891 );
and ( n83106 , n83105 , n417572 );
or ( n83107 , n83104 , n83106 );
buf ( n429035 , n83107 );
buf ( n429036 , n50579 );
nand ( n83110 , n429035 , n429036 );
buf ( n429038 , n83110 );
buf ( n429039 , n429038 );
nand ( n83113 , n83103 , n429039 );
buf ( n429041 , n83113 );
buf ( n429042 , n429041 );
and ( n83116 , n83098 , n429042 );
and ( n83117 , n429020 , n429024 );
or ( n83118 , n83116 , n83117 );
buf ( n429046 , n83118 );
buf ( n429047 , n429046 );
buf ( n429048 , C0 );
buf ( n429049 , n429048 );
and ( n83148 , n429006 , n429047 );
or ( n83149 , C0 , n83148 );
buf ( n429052 , n83149 );
buf ( n429053 , n429052 );
xor ( n83152 , n429002 , n429053 );
xor ( n429055 , n428730 , n428755 );
xor ( n429056 , n429055 , n428761 );
buf ( n429057 , n429056 );
buf ( n429058 , n429057 );
and ( n429059 , n83152 , n429058 );
or ( n429060 , n429059 , C0 );
buf ( n429061 , n429060 );
buf ( n429062 , n429061 );
xor ( n429063 , n428510 , n428766 );
xor ( n429064 , n429063 , n428863 );
buf ( n429065 , n429064 );
buf ( n429066 , n429065 );
buf ( n429067 , C0 );
buf ( n429068 , n429067 );
and ( n83188 , n429062 , n429066 );
or ( n429070 , C0 , n83188 );
buf ( n429071 , n429070 );
buf ( n429072 , n429071 );
xor ( n429073 , n82899 , n82889 );
not ( n429074 , n428884 );
xor ( n83194 , n429073 , n429074 );
buf ( n429076 , n83194 );
xor ( n429077 , n429072 , n429076 );
xor ( n83197 , n428966 , n428977 );
xor ( n429079 , n83197 , n428979 );
buf ( n429080 , n429079 );
buf ( n429081 , n429080 );
and ( n429082 , n429077 , n429081 );
and ( n429083 , n429072 , n429076 );
or ( n83203 , n429082 , n429083 );
buf ( n429085 , n83203 );
buf ( n429086 , n429085 );
nor ( n83206 , n429000 , n429086 );
buf ( n429088 , n83206 );
xor ( n429089 , n428259 , n428275 );
xor ( n83209 , n429089 , n428335 );
xor ( n429091 , n428572 , n428673 );
xor ( n429092 , n83209 , n429091 );
buf ( n429093 , n429092 );
buf ( n429094 , n399271 );
not ( n429095 , n429094 );
buf ( n429096 , n393397 );
not ( n429097 , n429096 );
or ( n429098 , n429095 , n429097 );
buf ( n429099 , n81579 );
buf ( n429100 , n399271 );
not ( n429101 , n429100 );
buf ( n429102 , n429101 );
buf ( n429103 , n429102 );
nand ( n429104 , n429099 , n429103 );
buf ( n429105 , n429104 );
buf ( n429106 , n429105 );
nand ( n429107 , n429098 , n429106 );
buf ( n429108 , n429107 );
buf ( n429109 , n429108 );
not ( n429110 , n429109 );
buf ( n429111 , n47903 );
not ( n429112 , n429111 );
or ( n429113 , n429110 , n429112 );
buf ( n429114 , n428699 );
buf ( n429115 , n395359 );
nand ( n429116 , n429114 , n429115 );
buf ( n429117 , n429116 );
buf ( n429118 , n429117 );
nand ( n429119 , n429113 , n429118 );
buf ( n429120 , n429119 );
buf ( n429121 , n429120 );
xor ( n429122 , n429093 , n429121 );
buf ( n429123 , n71170 );
buf ( n429124 , n62499 );
and ( n429125 , n429123 , n429124 );
buf ( n429126 , n417804 );
buf ( n429127 , n410717 );
and ( n429128 , n429126 , n429127 );
nor ( n83248 , n429125 , n429128 );
buf ( n429130 , n83248 );
buf ( n429131 , n429130 );
buf ( n429132 , n410724 );
or ( n429133 , n429131 , n429132 );
buf ( n429134 , n428583 );
buf ( n429135 , n410721 );
or ( n429136 , n429134 , n429135 );
nand ( n429137 , n429133 , n429136 );
buf ( n429138 , n429137 );
buf ( n429139 , n429138 );
buf ( n429140 , n409429 );
buf ( n429141 , n62177 );
buf ( n429142 , n74002 );
and ( n429143 , n429141 , n429142 );
buf ( n429144 , n409178 );
buf ( n429145 , n420612 );
and ( n429146 , n429144 , n429145 );
nor ( n83266 , n429143 , n429146 );
buf ( n429148 , n83266 );
buf ( n429149 , n429148 );
or ( n83269 , n429140 , n429149 );
buf ( n429151 , n428314 );
buf ( n429152 , n409170 );
or ( n83272 , n429151 , n429152 );
nand ( n429154 , n83269 , n83272 );
buf ( n429155 , n429154 );
buf ( n429156 , n429155 );
xor ( n429157 , n429139 , n429156 );
buf ( n429158 , n59469 );
buf ( n429159 , n623 );
or ( n429160 , n429158 , n429159 );
buf ( n429161 , n59468 );
buf ( n429162 , n59628 );
buf ( n429163 , n623 );
and ( n429164 , n429161 , n429162 , n429163 );
buf ( n429165 , n406602 );
not ( n429166 , n429165 );
buf ( n429167 , n429166 );
buf ( n429168 , n429167 );
nor ( n429169 , n429164 , n429168 );
buf ( n429170 , n429169 );
buf ( n429171 , n429170 );
nand ( n429172 , n429160 , n429171 );
buf ( n429173 , n429172 );
buf ( n429174 , n429173 );
and ( n429175 , n429157 , n429174 );
and ( n429176 , n429139 , n429156 );
or ( n83296 , n429175 , n429176 );
buf ( n429178 , n83296 );
xor ( n429179 , n428591 , n428652 );
xor ( n83299 , n429179 , n428656 );
and ( n83300 , n429178 , n83299 );
buf ( n429182 , n429148 );
buf ( n429183 , n409170 );
or ( n83303 , n429182 , n429183 );
buf ( n429185 , n409181 );
nand ( n83305 , n83303 , n429185 );
buf ( n429187 , n83305 );
buf ( n429188 , n71664 );
buf ( n429189 , n62499 );
and ( n83309 , n429188 , n429189 );
buf ( n429191 , n418298 );
buf ( n429192 , n410717 );
and ( n83312 , n429191 , n429192 );
nor ( n83313 , n83309 , n83312 );
buf ( n429195 , n83313 );
buf ( n429196 , n429195 );
buf ( n429197 , n410724 );
or ( n83317 , n429196 , n429197 );
buf ( n429199 , n429130 );
buf ( n429200 , n410721 );
or ( n83320 , n429199 , n429200 );
nand ( n83321 , n83317 , n83320 );
buf ( n429203 , n83321 );
xor ( n83323 , n429187 , n429203 );
xor ( n83324 , n428640 , n428645 );
buf ( n429206 , n83324 );
and ( n83326 , n83323 , n429206 );
and ( n83327 , n429187 , n429203 );
or ( n83328 , n83326 , n83327 );
buf ( n429210 , n83328 );
xor ( n83330 , n428605 , n428622 );
xor ( n83331 , n83330 , n428648 );
buf ( n429213 , n83331 );
buf ( n429214 , n429213 );
xor ( n83334 , n429210 , n429214 );
xor ( n83335 , n429139 , n429156 );
xor ( n83336 , n83335 , n429174 );
buf ( n429218 , n83336 );
buf ( n429219 , n429218 );
and ( n83339 , n83334 , n429219 );
and ( n83340 , n429210 , n429214 );
or ( n83341 , n83339 , n83340 );
buf ( n429223 , n83341 );
xor ( n83343 , n428591 , n428652 );
xor ( n83344 , n83343 , n428656 );
and ( n83345 , n429223 , n83344 );
and ( n83346 , n429178 , n429223 );
or ( n83347 , n83300 , n83345 , n83346 );
buf ( n429229 , n83347 );
xor ( n83349 , n428660 , n428664 );
xor ( n83350 , n83349 , n428669 );
buf ( n429232 , n83350 );
buf ( n429233 , n429232 );
xor ( n83353 , n429229 , n429233 );
buf ( n429235 , n51553 );
not ( n83355 , n429235 );
buf ( n429237 , n23551 );
not ( n83357 , n429237 );
buf ( n429239 , n83357 );
and ( n83359 , n372373 , n429239 );
not ( n83360 , n372373 );
and ( n83361 , n83360 , n47891 );
or ( n83362 , n83359 , n83361 );
buf ( n429244 , n83362 );
not ( n83364 , n429244 );
or ( n83365 , n83355 , n83364 );
buf ( n429247 , n47891 );
buf ( n429248 , n82708 );
and ( n83368 , n429247 , n429248 );
not ( n83369 , n429247 );
buf ( n429251 , n82708 );
not ( n83371 , n429251 );
buf ( n429253 , n83371 );
buf ( n429254 , n429253 );
and ( n83374 , n83369 , n429254 );
nor ( n83375 , n83368 , n83374 );
buf ( n429257 , n83375 );
buf ( n429258 , n429257 );
buf ( n429259 , n50578 );
nand ( n83379 , n429258 , n429259 );
buf ( n429261 , n83379 );
buf ( n429262 , n429261 );
nand ( n83382 , n83365 , n429262 );
buf ( n429264 , n83382 );
buf ( n429265 , n429264 );
and ( n83385 , n83353 , n429265 );
and ( n83386 , n429229 , n429233 );
or ( n83387 , n83385 , n83386 );
buf ( n429269 , n83387 );
buf ( n429270 , n429269 );
xor ( n83390 , n429122 , n429270 );
buf ( n429272 , n83390 );
buf ( n429273 , n429272 );
buf ( n429274 , C0 );
buf ( n429275 , n429274 );
xor ( n83414 , n429273 , n429275 );
buf ( n429277 , n55055 );
not ( n83416 , n429277 );
buf ( n429279 , n392217 );
not ( n83418 , n429279 );
buf ( n429281 , n83418 );
buf ( n429282 , n429281 );
not ( n83421 , n429282 );
or ( n83422 , n83416 , n83421 );
buf ( n429285 , n392217 );
buf ( n429286 , n55054 );
nand ( n83425 , n429285 , n429286 );
buf ( n429288 , n83425 );
buf ( n429289 , n429288 );
nand ( n83428 , n83422 , n429289 );
buf ( n429291 , n83428 );
buf ( n429292 , n429291 );
not ( n83431 , n429292 );
buf ( n429294 , n427074 );
not ( n83433 , n429294 );
or ( n83434 , n83431 , n83433 );
buf ( n429297 , n400033 );
not ( n83436 , n429297 );
buf ( n429299 , n426763 );
not ( n83438 , n429299 );
or ( n83439 , n83436 , n83438 );
buf ( n429302 , n392217 );
buf ( n429303 , n400042 );
nand ( n83442 , n429302 , n429303 );
buf ( n429305 , n83442 );
buf ( n429306 , n429305 );
nand ( n83445 , n83439 , n429306 );
buf ( n429308 , n83445 );
buf ( n429309 , n429308 );
buf ( n429310 , n45954 );
nand ( n83449 , n429309 , n429310 );
buf ( n429312 , n83449 );
buf ( n429313 , n429312 );
nand ( n83452 , n83434 , n429313 );
buf ( n429315 , n83452 );
buf ( n429316 , n429315 );
and ( n83455 , n83414 , n429316 );
or ( n83457 , n83455 , C0 );
buf ( n429319 , n83457 );
buf ( n429320 , n429319 );
buf ( n429321 , n51553 );
not ( n83461 , n429321 );
buf ( n429323 , n83107 );
not ( n83463 , n429323 );
or ( n83464 , n83461 , n83463 );
buf ( n429326 , n50579 );
and ( n83466 , n24790 , n50584 );
not ( n83467 , n24790 );
and ( n83468 , n83467 , n47891 );
or ( n83469 , n83466 , n83468 );
buf ( n429331 , n83469 );
nand ( n83471 , n429326 , n429331 );
buf ( n429333 , n83471 );
buf ( n429334 , n429333 );
nand ( n83474 , n83464 , n429334 );
buf ( n429336 , n83474 );
buf ( n429337 , n429336 );
buf ( n429338 , n44775 );
buf ( n429339 , n392231 );
buf ( n429340 , n426763 );
nand ( n83480 , n429339 , n429340 );
buf ( n429342 , n83480 );
buf ( n429343 , n429342 );
buf ( n429344 , n358975 );
and ( n83484 , n429343 , n429344 );
and ( n83485 , n392218 , n392219 );
buf ( n429347 , n83485 );
buf ( n429348 , n429347 );
nor ( n83488 , n83484 , n429348 );
buf ( n429350 , n83488 );
buf ( n429351 , n429350 );
and ( n83491 , n429338 , n429351 );
buf ( n429353 , n83491 );
buf ( n429354 , n429353 );
xor ( n83494 , n429337 , n429354 );
buf ( n429356 , n51553 );
not ( n83496 , n429356 );
buf ( n429358 , n83469 );
not ( n83498 , n429358 );
or ( n83499 , n83496 , n83498 );
buf ( n429361 , n83362 );
buf ( n429362 , n50579 );
nand ( n83502 , n429361 , n429362 );
buf ( n429364 , n83502 );
buf ( n429365 , n429364 );
nand ( n83505 , n83499 , n429365 );
buf ( n429367 , n83505 );
buf ( n429368 , n429367 );
buf ( n429369 , n392221 );
buf ( n429370 , n358975 );
nand ( n83510 , n429369 , n429370 );
buf ( n429372 , n83510 );
buf ( n429373 , n429372 );
not ( n83513 , n429373 );
buf ( n429375 , n83513 );
buf ( n429376 , n429375 );
xor ( n83516 , n429368 , n429376 );
buf ( n429378 , n400033 );
not ( n83518 , n429378 );
buf ( n429380 , n393397 );
not ( n83520 , n429380 );
or ( n83521 , n83518 , n83520 );
buf ( n429383 , n400042 );
buf ( n429384 , n23604 );
nand ( n83524 , n429383 , n429384 );
buf ( n429386 , n83524 );
buf ( n429387 , n429386 );
nand ( n83527 , n83521 , n429387 );
buf ( n429389 , n83527 );
buf ( n429390 , n429389 );
not ( n83530 , n429390 );
buf ( n429392 , n47903 );
not ( n83532 , n429392 );
or ( n83533 , n83530 , n83532 );
buf ( n429395 , n395359 );
buf ( n429396 , n429108 );
nand ( n83536 , n429395 , n429396 );
buf ( n429398 , n83536 );
buf ( n429399 , n429398 );
nand ( n83539 , n83533 , n429399 );
buf ( n429401 , n83539 );
buf ( n429402 , n429401 );
xor ( n83542 , n429229 , n429233 );
xor ( n83543 , n83542 , n429265 );
buf ( n429405 , n83543 );
buf ( n429406 , n429405 );
xor ( n83546 , n429402 , n429406 );
buf ( n429408 , n392217 );
buf ( n429409 , n371244 );
buf ( n429410 , n81579 );
or ( n83550 , n429409 , n429410 );
buf ( n429412 , n358975 );
nand ( n83552 , n83550 , n429412 );
buf ( n429414 , n83552 );
buf ( n429415 , n429414 );
buf ( n429416 , n81579 );
buf ( n429417 , n371244 );
nand ( n83557 , n429416 , n429417 );
buf ( n429419 , n83557 );
buf ( n429420 , n429419 );
and ( n83560 , n429408 , n429415 , n429420 );
buf ( n429422 , n83560 );
buf ( n429423 , n429422 );
and ( n83563 , n83546 , n429423 );
and ( n83564 , n429402 , n429406 );
or ( n83565 , n83563 , n83564 );
buf ( n429427 , n83565 );
buf ( n429428 , n429427 );
and ( n429429 , n83516 , n429428 );
and ( n83569 , n429368 , n429376 );
or ( n429431 , n429429 , n83569 );
buf ( n429432 , n429431 );
buf ( n429433 , n429432 );
xor ( n83573 , n83494 , n429433 );
buf ( n429435 , n83573 );
buf ( n429436 , n429435 );
buf ( n429437 , C0 );
buf ( n429438 , n429437 );
and ( n429439 , n429320 , n429436 );
or ( n83591 , C0 , n429439 );
buf ( n429441 , n83591 );
buf ( n429442 , n429441 );
xor ( n429443 , n428679 , n428683 );
xor ( n83595 , n429443 , n428710 );
buf ( n429445 , n83595 );
buf ( n429446 , n429445 );
xor ( n429447 , n429093 , n429121 );
and ( n83599 , n429447 , n429270 );
and ( n429449 , n429093 , n429121 );
or ( n83601 , n83599 , n429449 );
buf ( n429451 , n83601 );
buf ( n429452 , n429451 );
xor ( n429453 , n429446 , n429452 );
buf ( n429454 , n426775 );
not ( n429455 , n429454 );
buf ( n429456 , n83083 );
not ( n429457 , n429456 );
or ( n83609 , n429455 , n429457 );
buf ( n429459 , n429308 );
buf ( n429460 , n427074 );
nand ( n429461 , n429459 , n429460 );
buf ( n429462 , n429461 );
buf ( n429463 , n429462 );
nand ( n83615 , n83609 , n429463 );
buf ( n429465 , n83615 );
buf ( n429466 , n429465 );
xor ( n429467 , n429453 , n429466 );
buf ( n429468 , n429467 );
buf ( n429469 , n429468 );
buf ( n429470 , C0 );
buf ( n429471 , n429470 );
xor ( n429472 , n429469 , n429471 );
buf ( n429473 , n413643 );
not ( n429474 , n429473 );
buf ( n429475 , n55055 );
not ( n429476 , n429475 );
buf ( n429477 , n422673 );
not ( n429478 , n429477 );
or ( n83653 , n429476 , n429478 );
buf ( n429480 , n390988 );
buf ( n429481 , n55054 );
nand ( n429482 , n429480 , n429481 );
buf ( n429483 , n429482 );
buf ( n429484 , n429483 );
nand ( n83659 , n83653 , n429484 );
buf ( n429486 , n83659 );
buf ( n429487 , n429486 );
not ( n429488 , n429487 );
or ( n83663 , n429474 , n429488 );
buf ( n429490 , n44770 );
buf ( n429491 , n358975 );
not ( n429492 , n429491 );
buf ( n429493 , n422673 );
not ( n429494 , n429493 );
or ( n83669 , n429492 , n429494 );
buf ( n429496 , n44775 );
buf ( n429497 , n402819 );
nand ( n429498 , n429496 , n429497 );
buf ( n429499 , n429498 );
buf ( n429500 , n429499 );
nand ( n83675 , n83669 , n429500 );
buf ( n429502 , n83675 );
buf ( n429503 , n429502 );
nand ( n429504 , n429490 , n429503 );
buf ( n429505 , n429504 );
buf ( n429506 , n429505 );
nand ( n83681 , n83663 , n429506 );
buf ( n429508 , n83681 );
buf ( n429509 , n429508 );
and ( n429510 , n429472 , n429509 );
or ( n429511 , n429510 , C0 );
buf ( n429512 , n429511 );
buf ( n429513 , n429512 );
xor ( n83689 , n429442 , n429513 );
xor ( n429515 , n429446 , n429452 );
and ( n83691 , n429515 , n429466 );
and ( n429517 , n429446 , n429452 );
or ( n83693 , n83691 , n429517 );
buf ( n429519 , n83693 );
buf ( n429520 , n429519 );
buf ( n429521 , n429486 );
not ( n83697 , n429521 );
buf ( n429523 , n44770 );
not ( n83699 , n429523 );
or ( n429525 , n83697 , n83699 );
buf ( n429526 , n413643 );
buf ( n429527 , n428814 );
nand ( n83703 , n429526 , n429527 );
buf ( n429529 , n83703 );
buf ( n429530 , n429529 );
nand ( n429531 , n429525 , n429530 );
buf ( n429532 , n429531 );
buf ( n429533 , n429532 );
xor ( n83709 , n429520 , n429533 );
buf ( n429535 , n43514 );
buf ( n429536 , n402819 );
nor ( n429537 , n429535 , n429536 );
buf ( n429538 , n429537 );
buf ( n429539 , n429538 );
xor ( n83715 , n83709 , n429539 );
buf ( n429541 , n83715 );
buf ( n429542 , n429541 );
and ( n429543 , n83689 , n429542 );
and ( n83719 , n429442 , n429513 );
or ( n429545 , n429543 , n83719 );
buf ( n429546 , n429545 );
buf ( n429547 , n429546 );
xor ( n83723 , n429520 , n429533 );
and ( n429549 , n83723 , n429539 );
and ( n83725 , n429520 , n429533 );
or ( n83726 , n429549 , n83725 );
buf ( n429552 , n83726 );
buf ( n429553 , n429552 );
xor ( n83729 , n428802 , n428827 );
xor ( n429555 , n83729 , n428840 );
buf ( n429556 , n429555 );
buf ( n429557 , n429556 );
xor ( n429558 , n429553 , n429557 );
buf ( n429559 , n358975 );
not ( n83735 , n429559 );
buf ( n429561 , n425525 );
not ( n83737 , n429561 );
or ( n83738 , n83735 , n83737 );
buf ( n429564 , n388064 );
buf ( n429565 , n402819 );
nand ( n83741 , n429564 , n429565 );
buf ( n429567 , n83741 );
buf ( n429568 , n429567 );
nand ( n83744 , n83738 , n429568 );
buf ( n429570 , n83744 );
buf ( n429571 , n429570 );
not ( n83747 , n429571 );
buf ( n429573 , n74375 );
not ( n83749 , n429573 );
or ( n83750 , n83747 , n83749 );
nand ( n429576 , n82796 , n43515 );
buf ( n429577 , n429576 );
nand ( n83753 , n83750 , n429577 );
buf ( n429579 , n83753 );
buf ( n429580 , n429579 );
xor ( n83756 , n429558 , n429580 );
buf ( n429582 , n83756 );
buf ( n429583 , n429582 );
xor ( n83759 , n429547 , n429583 );
xor ( n429585 , n429337 , n429354 );
and ( n83761 , n429585 , n429433 );
and ( n83762 , n429337 , n429354 );
or ( n429588 , n83761 , n83762 );
buf ( n429589 , n429588 );
buf ( n429590 , n429589 );
xor ( n429591 , n429020 , n429024 );
xor ( n83767 , n429591 , n429042 );
buf ( n429593 , n83767 );
buf ( n429594 , n429593 );
buf ( n429595 , C0 );
buf ( n429596 , n429595 );
and ( n83785 , n429590 , n429594 );
or ( n83786 , C0 , n83785 );
buf ( n429599 , n83786 );
buf ( n429600 , n429599 );
xor ( n83789 , n429006 , n429047 );
xor ( n429602 , n83789 , n429049 );
buf ( n429603 , n429602 );
buf ( n429604 , n429603 );
xor ( n429605 , n429600 , n429604 );
buf ( n429606 , C0 );
xor ( n83809 , n429605 , n429606 );
buf ( n429608 , n83809 );
buf ( n429609 , n429608 );
and ( n83812 , n83759 , n429609 );
and ( n83813 , n429547 , n429583 );
or ( n429612 , n83812 , n83813 );
buf ( n429613 , n429612 );
buf ( n429614 , n429613 );
not ( n429615 , n429614 );
xor ( n83818 , n429553 , n429557 );
and ( n83819 , n83818 , n429580 );
and ( n429618 , n429553 , n429557 );
or ( n83821 , n83819 , n429618 );
buf ( n429620 , n83821 );
buf ( n429621 , n429620 );
buf ( n429622 , n428844 );
not ( n83825 , n429622 );
buf ( n429624 , n83825 );
buf ( n429625 , n429624 );
not ( n83828 , n429625 );
buf ( n429627 , n428851 );
not ( n83830 , n429627 );
or ( n83831 , n83828 , n83830 );
buf ( n429630 , n428844 );
buf ( n429631 , n82869 );
nand ( n83834 , n429630 , n429631 );
buf ( n429633 , n83834 );
buf ( n429634 , n429633 );
nand ( n83837 , n83831 , n429634 );
buf ( n429636 , n83837 );
buf ( n429637 , n429636 );
buf ( n429638 , n82805 );
and ( n429639 , n429637 , n429638 );
not ( n83842 , n429637 );
buf ( n429641 , n82805 );
not ( n429642 , n429641 );
buf ( n429643 , n429642 );
buf ( n429644 , n429643 );
and ( n429645 , n83842 , n429644 );
nor ( n83848 , n429639 , n429645 );
buf ( n429647 , n83848 );
buf ( n429648 , n429647 );
xor ( n83851 , n429621 , n429648 );
buf ( n429650 , C0 );
buf ( n429651 , n429650 );
xor ( n83866 , n83851 , n429651 );
buf ( n429653 , n83866 );
and ( n429654 , n429600 , n429604 );
or ( n429655 , C0 , n429654 );
buf ( n429656 , n429655 );
buf ( n429657 , n429656 );
xor ( n429658 , n429002 , n429053 );
xor ( n429659 , n429658 , n429058 );
buf ( n429660 , n429659 );
buf ( n429661 , n429660 );
not ( n429662 , n429661 );
buf ( n429663 , n429662 );
buf ( n429664 , n429663 );
and ( n429665 , n429657 , n429664 );
not ( n429666 , n429657 );
buf ( n429667 , n429660 );
and ( n429668 , n429666 , n429667 );
nor ( n429669 , n429665 , n429668 );
buf ( n429670 , n429669 );
xor ( n429671 , n429653 , n429670 );
buf ( n429672 , n429671 );
nand ( n429673 , n429615 , n429672 );
buf ( n429674 , n429673 );
not ( n429675 , n429674 );
xor ( n429676 , n429273 , n429275 );
xor ( n429677 , n429676 , n429316 );
buf ( n429678 , n429677 );
buf ( n429679 , n429678 );
buf ( n429680 , n62155 );
buf ( n429681 , n623 );
and ( n429682 , n429680 , n429681 );
buf ( n429683 , n62177 );
buf ( n429684 , n409156 );
buf ( n429685 , n422315 );
and ( n83899 , n429684 , n429685 );
buf ( n429687 , n62164 );
nor ( n83901 , n83899 , n429687 );
buf ( n429689 , n83901 );
buf ( n429690 , n429689 );
nor ( n83904 , n429682 , n429683 , n429690 );
buf ( n429692 , n83904 );
buf ( n429693 , n429692 );
buf ( n429694 , n71681 );
buf ( n429695 , n62499 );
and ( n83909 , n429694 , n429695 );
buf ( n429697 , n418315 );
buf ( n429698 , n410717 );
and ( n429699 , n429697 , n429698 );
nor ( n83913 , n83909 , n429699 );
buf ( n429701 , n83913 );
buf ( n429702 , n429701 );
buf ( n429703 , n410724 );
or ( n83917 , n429702 , n429703 );
buf ( n429705 , n429195 );
buf ( n429706 , n410721 );
or ( n83920 , n429705 , n429706 );
nand ( n83921 , n83917 , n83920 );
buf ( n429709 , n83921 );
buf ( n429710 , n429709 );
xor ( n83924 , n429693 , n429710 );
buf ( n429712 , n410635 );
buf ( n429713 , n62164 );
buf ( n429714 , n74002 );
and ( n429715 , n429713 , n429714 );
buf ( n429716 , n62511 );
buf ( n429717 , n420612 );
and ( n83931 , n429716 , n429717 );
nor ( n83932 , n429715 , n83931 );
buf ( n429720 , n83932 );
buf ( n429721 , n429720 );
or ( n83935 , n429712 , n429721 );
buf ( n429723 , n428632 );
buf ( n429724 , n409504 );
or ( n83938 , n429723 , n429724 );
nand ( n83939 , n83935 , n83938 );
buf ( n429727 , n83939 );
buf ( n429728 , n429727 );
and ( n83942 , n83924 , n429728 );
and ( n83943 , n429693 , n429710 );
or ( n83944 , n83942 , n83943 );
buf ( n429732 , n83944 );
xor ( n83946 , n429187 , n429203 );
xor ( n83947 , n83946 , n429206 );
and ( n83948 , n429732 , n83947 );
buf ( n429736 , n409170 );
buf ( n429737 , n422315 );
nor ( n83951 , n429736 , n429737 );
buf ( n429739 , n83951 );
buf ( n429740 , n429739 );
buf ( n429741 , n429720 );
buf ( n429742 , n409504 );
or ( n429743 , n429741 , n429742 );
buf ( n429744 , n409512 );
nand ( n83958 , n429743 , n429744 );
buf ( n429746 , n83958 );
buf ( n429747 , n429746 );
and ( n83961 , n429740 , n429747 );
buf ( n429749 , n83961 );
buf ( n429750 , n429749 );
buf ( n429751 , n409181 );
buf ( n429752 , n623 );
or ( n83966 , n429751 , n429752 );
buf ( n429754 , n409173 );
buf ( n429755 , n62177 );
buf ( n429756 , n623 );
and ( n83970 , n429754 , n429755 , n429756 );
buf ( n429758 , n409189 );
not ( n83972 , n429758 );
buf ( n429760 , n83972 );
buf ( n429761 , n429760 );
nor ( n83975 , n83970 , n429761 );
buf ( n429763 , n83975 );
buf ( n429764 , n429763 );
nand ( n83978 , n83966 , n429764 );
buf ( n429766 , n83978 );
buf ( n429767 , n429766 );
xor ( n83981 , n429750 , n429767 );
xor ( n83982 , n429693 , n429710 );
xor ( n83983 , n83982 , n429728 );
buf ( n429771 , n83983 );
buf ( n429772 , n429771 );
and ( n83986 , n83981 , n429772 );
and ( n429774 , n429750 , n429767 );
or ( n83988 , n83986 , n429774 );
buf ( n429776 , n83988 );
xor ( n83990 , n429187 , n429203 );
xor ( n83991 , n83990 , n429206 );
and ( n83992 , n429776 , n83991 );
and ( n83993 , n429732 , n429776 );
or ( n83994 , n83948 , n83992 , n83993 );
xor ( n83995 , n429210 , n429214 );
xor ( n83996 , n83995 , n429219 );
buf ( n429784 , n83996 );
or ( n429785 , n83994 , n429784 );
not ( n83999 , n429785 );
not ( n84000 , n50578 );
not ( n84001 , n400033 );
not ( n84002 , n395333 );
or ( n84003 , n84001 , n84002 );
buf ( n429791 , n400042 );
buf ( n429792 , n47891 );
nand ( n84006 , n429791 , n429792 );
buf ( n429794 , n84006 );
nand ( n84008 , n84003 , n429794 );
not ( n84009 , n84008 );
or ( n84010 , n84000 , n84009 );
buf ( n429798 , n399271 );
buf ( n429799 , n47891 );
and ( n429800 , n429798 , n429799 );
not ( n84014 , n429798 );
buf ( n429802 , n429239 );
and ( n84016 , n84014 , n429802 );
nor ( n84017 , n429800 , n84016 );
buf ( n429805 , n84017 );
nand ( n84019 , n429805 , n51553 );
nand ( n84020 , n84010 , n84019 );
not ( n84021 , n84020 );
or ( n84022 , n83999 , n84021 );
nand ( n84023 , n83994 , n429784 );
nand ( n84024 , n84022 , n84023 );
not ( n84025 , n84024 );
buf ( n429813 , n51553 );
not ( n84027 , n429813 );
buf ( n429815 , n429257 );
not ( n84029 , n429815 );
or ( n84030 , n84027 , n84029 );
nand ( n84031 , n429805 , n50578 );
buf ( n429819 , n84031 );
nand ( n84033 , n84030 , n429819 );
buf ( n429821 , n84033 );
buf ( n429822 , n429821 );
xor ( n84036 , n428591 , n428652 );
xor ( n84037 , n84036 , n428656 );
xor ( n84038 , n429178 , n429223 );
xor ( n84039 , n84037 , n84038 );
buf ( n429827 , n84039 );
or ( n84041 , n429822 , n429827 );
buf ( n429829 , n84041 );
not ( n84043 , n429829 );
or ( n84044 , n84025 , n84043 );
buf ( n429832 , n429821 );
buf ( n429833 , n84039 );
nand ( n84047 , n429832 , n429833 );
buf ( n429835 , n84047 );
nand ( n84049 , n84044 , n429835 );
buf ( n429837 , n84049 );
not ( n84051 , n429837 );
buf ( n429839 , n358975 );
not ( n84053 , n429839 );
buf ( n429841 , n429281 );
not ( n84055 , n429841 );
or ( n84056 , n84053 , n84055 );
buf ( n429844 , n392217 );
buf ( n429845 , n402819 );
nand ( n84059 , n429844 , n429845 );
buf ( n429847 , n84059 );
buf ( n429848 , n429847 );
nand ( n84062 , n84056 , n429848 );
buf ( n429850 , n84062 );
buf ( n429851 , n429850 );
not ( n84065 , n429851 );
buf ( n429853 , n427074 );
not ( n84067 , n429853 );
or ( n84068 , n84065 , n84067 );
buf ( n429856 , n429291 );
buf ( n429857 , n426775 );
nand ( n84071 , n429856 , n429857 );
buf ( n429859 , n84071 );
buf ( n429860 , n429859 );
nand ( n84074 , n84068 , n429860 );
buf ( n429862 , n84074 );
buf ( n429863 , n429862 );
not ( n84077 , n429863 );
or ( n84078 , n84051 , n84077 );
buf ( n429866 , n84049 );
buf ( n429867 , n429862 );
or ( n84081 , n429866 , n429867 );
not ( n84082 , n47903 );
buf ( n429870 , n55054 );
buf ( n429871 , n81579 );
and ( n84085 , n429870 , n429871 );
not ( n84086 , n429870 );
buf ( n429874 , n393397 );
and ( n84088 , n84086 , n429874 );
nor ( n84089 , n84085 , n84088 );
buf ( n429877 , n84089 );
not ( n84091 , n429877 );
not ( n84092 , n84091 );
or ( n84093 , n84082 , n84092 );
nand ( n84094 , n429389 , n395359 );
nand ( n84095 , n84093 , n84094 );
not ( n84124 , n84095 );
buf ( n429884 , n84124 );
not ( n429885 , n429884 );
or ( n84129 , n429885 , C0 );
buf ( n429887 , n395325 );
buf ( n429888 , n429239 );
nand ( n84132 , n429887 , n429888 );
buf ( n429890 , n84132 );
and ( n84134 , n358975 , n429890 );
buf ( n429892 , n429239 );
not ( n84136 , n429892 );
buf ( n429894 , n84136 );
and ( n84138 , n395328 , n429894 );
nor ( n84139 , n84134 , n84138 , n393397 );
buf ( n429897 , n84139 );
xor ( n84141 , n83994 , n429784 );
and ( n84142 , n84020 , n84141 );
not ( n84143 , n84020 );
not ( n84144 , n84141 );
and ( n84145 , n84143 , n84144 );
nor ( n84146 , n84142 , n84145 );
buf ( n429904 , n84146 );
buf ( n429905 , C0 );
buf ( n429906 , n429905 );
and ( n84171 , n429897 , n429904 );
or ( n84172 , C0 , n84171 );
buf ( n429909 , n84172 );
buf ( n429910 , n429909 );
nand ( n84175 , n84129 , n429910 );
buf ( n429912 , n84175 );
buf ( n429913 , n429912 );
nand ( n84178 , C1 , n429913 );
buf ( n429915 , n84178 );
buf ( n429916 , n429915 );
nand ( n429917 , n84081 , n429916 );
buf ( n429918 , n429917 );
buf ( n429919 , n429918 );
nand ( n84184 , n84078 , n429919 );
buf ( n429921 , n84184 );
buf ( n429922 , n429921 );
not ( n84187 , n429922 );
xor ( n84188 , n429368 , n429376 );
xor ( n84189 , n84188 , n429428 );
buf ( n429926 , n84189 );
buf ( n429927 , n429926 );
not ( n84192 , n429927 );
buf ( n429929 , n84192 );
buf ( n429930 , n429929 );
nand ( n84195 , n84187 , n429930 );
buf ( n429932 , n84195 );
buf ( n429933 , n429932 );
and ( n84198 , n429679 , n429933 );
buf ( n429935 , n429921 );
not ( n84200 , n429935 );
buf ( n429937 , n429929 );
nor ( n84202 , n84200 , n429937 );
buf ( n429939 , n84202 );
buf ( n429940 , n429939 );
nor ( n84205 , n84198 , n429940 );
buf ( n429942 , n84205 );
buf ( n429943 , n429942 );
not ( n84208 , n429943 );
xor ( n84209 , n429320 , n429436 );
xor ( n84210 , n84209 , n429438 );
buf ( n429947 , n84210 );
buf ( n429948 , n429947 );
not ( n84213 , n429948 );
buf ( n429950 , n84213 );
buf ( n429951 , n429950 );
not ( n84216 , n429951 );
or ( n84217 , n84208 , n84216 );
xor ( n84218 , n429469 , n429471 );
xor ( n84219 , n84218 , n429509 );
buf ( n429956 , n84219 );
buf ( n429957 , n429956 );
nand ( n84222 , n84217 , n429957 );
buf ( n429959 , n84222 );
buf ( n429960 , n429959 );
buf ( n429961 , n429942 );
not ( n84226 , n429961 );
buf ( n429963 , n429947 );
nand ( n84228 , n84226 , n429963 );
buf ( n429965 , n84228 );
buf ( n429966 , n429965 );
nand ( n84231 , n429960 , n429966 );
buf ( n429968 , n84231 );
buf ( n429969 , n429968 );
buf ( n429970 , n84049 );
buf ( n429971 , n429862 );
xor ( n84236 , n429970 , n429971 );
buf ( n429973 , n429915 );
xnor ( n84238 , n84236 , n429973 );
buf ( n429975 , n84238 );
buf ( n429976 , n429975 );
buf ( n429977 , C1 );
buf ( n429978 , n429977 );
xor ( n84263 , n429976 , n429978 );
buf ( n429980 , C0 );
buf ( n429981 , n429980 );
xor ( n84277 , n429402 , n429406 );
xor ( n84278 , n84277 , n429423 );
buf ( n429984 , n84278 );
buf ( n429985 , n429984 );
xor ( n84281 , n429981 , n429985 );
buf ( n429987 , n402819 );
not ( n84283 , n429987 );
buf ( n429989 , n426775 );
nand ( n84285 , n84283 , n429989 );
buf ( n429991 , n84285 );
buf ( n429992 , n429991 );
buf ( n429993 , n84039 );
buf ( n429994 , n429821 );
xor ( n84290 , n429993 , n429994 );
buf ( n429996 , n84024 );
xnor ( n84292 , n84290 , n429996 );
buf ( n429998 , n84292 );
buf ( n429999 , n429998 );
nand ( n430000 , n429992 , n429999 );
buf ( n430001 , n430000 );
buf ( n430002 , n430001 );
not ( n84298 , n430002 );
xor ( n84299 , n429187 , n429203 );
xor ( n84300 , n84299 , n429206 );
xor ( n84301 , n429732 , n429776 );
xor ( n84302 , n84300 , n84301 );
buf ( n430008 , n84302 );
not ( n84304 , n430008 );
buf ( n430010 , n84304 );
buf ( n430011 , n430010 );
not ( n84307 , n430011 );
not ( n84308 , n50578 );
buf ( n430014 , n55055 );
not ( n84310 , n430014 );
buf ( n430016 , n395333 );
not ( n84312 , n430016 );
or ( n84313 , n84310 , n84312 );
buf ( n430019 , n429894 );
buf ( n430020 , n55054 );
nand ( n84316 , n430019 , n430020 );
buf ( n430022 , n84316 );
buf ( n430023 , n430022 );
nand ( n84319 , n84313 , n430023 );
buf ( n430025 , n84319 );
not ( n84321 , n430025 );
or ( n84322 , n84308 , n84321 );
nand ( n84323 , n84008 , n51553 );
nand ( n84324 , n84322 , n84323 );
buf ( n430030 , n84324 );
not ( n84326 , n430030 );
buf ( n430032 , n84326 );
buf ( n430033 , n430032 );
not ( n84329 , n430033 );
or ( n84330 , n84307 , n84329 );
buf ( n430036 , n50573 );
buf ( n430037 , C0 );
nor ( n84333 , n430036 , n430037 );
buf ( n430039 , n84333 );
buf ( n430040 , n430039 );
buf ( n430041 , n402819 );
or ( n84337 , n430040 , n430041 );
buf ( n430043 , C1 );
buf ( n430044 , n430043 );
nand ( n84343 , n84337 , n430044 );
buf ( n430046 , n84343 );
not ( n84345 , n430046 );
nand ( n84346 , n84345 , n47891 );
not ( n84347 , n84346 );
xor ( n84348 , n429740 , n429747 );
buf ( n430051 , n84348 );
buf ( n430052 , n430051 );
buf ( n430053 , n62499 );
buf ( n430054 , n72308 );
and ( n84353 , n430053 , n430054 );
buf ( n430056 , n410717 );
buf ( n430057 , n418942 );
and ( n84356 , n430056 , n430057 );
nor ( n84357 , n84353 , n84356 );
buf ( n430060 , n84357 );
buf ( n430061 , n430060 );
buf ( n430062 , n410724 );
or ( n84361 , n430061 , n430062 );
buf ( n430064 , n429701 );
buf ( n430065 , n410721 );
or ( n84364 , n430064 , n430065 );
nand ( n84365 , n84361 , n84364 );
buf ( n430068 , n84365 );
buf ( n430069 , n430068 );
xor ( n84368 , n430052 , n430069 );
buf ( n430071 , n62499 );
buf ( n430072 , n74002 );
and ( n84371 , n430071 , n430072 );
buf ( n430074 , n410717 );
buf ( n430075 , n420612 );
and ( n84374 , n430074 , n430075 );
nor ( n430077 , n84371 , n84374 );
buf ( n430078 , n430077 );
buf ( n430079 , n430078 );
buf ( n430080 , n410724 );
or ( n84379 , n430079 , n430080 );
buf ( n430082 , n430060 );
buf ( n430083 , n410721 );
or ( n84382 , n430082 , n430083 );
nand ( n84383 , n84379 , n84382 );
buf ( n430086 , n84383 );
buf ( n430087 , n430086 );
buf ( n430088 , n5744 );
buf ( n430089 , n623 );
and ( n84388 , n430088 , n430089 );
buf ( n430091 , n62164 );
buf ( n430092 , n409484 );
buf ( n430093 , n422315 );
and ( n84392 , n430092 , n430093 );
buf ( n430095 , n62499 );
nor ( n84394 , n84392 , n430095 );
buf ( n430097 , n84394 );
buf ( n430098 , n430097 );
nor ( n84397 , n84388 , n430091 , n430098 );
buf ( n430100 , n84397 );
buf ( n430101 , n430100 );
xor ( n84400 , n430087 , n430101 );
buf ( n430103 , n409512 );
buf ( n430104 , n623 );
or ( n84403 , n430103 , n430104 );
buf ( n430106 , n409507 );
buf ( n430107 , n63625 );
buf ( n430108 , n623 );
and ( n84407 , n430106 , n430107 , n430108 );
buf ( n430110 , n409520 );
not ( n84409 , n430110 );
buf ( n430112 , n84409 );
buf ( n430113 , n430112 );
nor ( n84412 , n84407 , n430113 );
buf ( n430115 , n84412 );
buf ( n430116 , n430115 );
nand ( n84415 , n84403 , n430116 );
buf ( n430118 , n84415 );
buf ( n430119 , n430118 );
and ( n84418 , n84400 , n430119 );
and ( n84419 , n430087 , n430101 );
or ( n84420 , n84418 , n84419 );
buf ( n430123 , n84420 );
buf ( n430124 , n430123 );
and ( n84423 , n84368 , n430124 );
and ( n84424 , n430052 , n430069 );
or ( n84425 , n84423 , n84424 );
buf ( n430128 , n84425 );
buf ( n430129 , n430128 );
not ( n84428 , n430129 );
buf ( n430131 , n84428 );
not ( n84430 , n430131 );
and ( n84431 , n84347 , n84430 );
buf ( n430134 , n430131 );
buf ( n430135 , n84346 );
nand ( n84434 , n430134 , n430135 );
buf ( n430137 , n84434 );
xor ( n84436 , n429750 , n429767 );
xor ( n84437 , n84436 , n429772 );
buf ( n430140 , n84437 );
and ( n84439 , n430137 , n430140 );
nor ( n84440 , n84431 , n84439 );
buf ( n430143 , n84440 );
not ( n84442 , n430143 );
buf ( n430145 , n84442 );
buf ( n430146 , n430145 );
nand ( n84445 , n84330 , n430146 );
buf ( n430148 , n84445 );
buf ( n430149 , n84324 );
buf ( n430150 , n84302 );
nand ( n84449 , n430149 , n430150 );
buf ( n430152 , n84449 );
nand ( n84451 , n430148 , n430152 );
buf ( n430154 , n402819 );
buf ( n430155 , n81579 );
xnor ( n84454 , n430154 , n430155 );
buf ( n430157 , n84454 );
not ( n84456 , n430157 );
not ( n84457 , n47903 );
or ( n84458 , n84456 , n84457 );
buf ( n430161 , n429877 );
not ( n84460 , n430161 );
buf ( n430163 , n395359 );
nand ( n84462 , n84460 , n430163 );
buf ( n430165 , n84462 );
nand ( n84464 , n84458 , n430165 );
xor ( n84465 , n84451 , n84464 );
buf ( n430168 , n395356 );
buf ( n430169 , n358975 );
nand ( n84485 , n430168 , n430169 );
buf ( n430171 , n84485 );
not ( n84492 , n84324 );
not ( n84493 , n430010 );
not ( n84494 , n430145 );
or ( n84495 , n84493 , n84494 );
buf ( n430176 , n84302 );
buf ( n430177 , n84440 );
nand ( n84498 , n430176 , n430177 );
buf ( n430179 , n84498 );
nand ( n84500 , n84495 , n430179 );
not ( n84501 , n84500 );
or ( n84502 , n84492 , n84501 );
nand ( n84503 , n430145 , n430010 );
not ( n84504 , n84324 );
nand ( n84505 , n84503 , n84504 , n430179 );
nand ( n84506 , n84502 , n84505 );
buf ( n430187 , n84506 );
not ( n84508 , n430187 );
buf ( n430189 , n84508 );
buf ( n430190 , n430189 );
buf ( n430191 , n430171 );
nand ( n430192 , C1 , n430191 );
buf ( n430193 , n430192 );
buf ( n430194 , n430193 );
nand ( n84517 , n430190 , n430194 );
buf ( n430196 , n84517 );
nand ( n84519 , C1 , n430196 );
and ( n84520 , n84465 , n84519 );
and ( n84521 , n84451 , n84464 );
or ( n84522 , n84520 , n84521 );
buf ( n430201 , n84522 );
not ( n84524 , n430201 );
or ( n84525 , n84298 , n84524 );
buf ( n430204 , n429991 );
not ( n84527 , n430204 );
buf ( n430206 , n84527 );
buf ( n430207 , n430206 );
buf ( n430208 , n429998 );
not ( n84531 , n430208 );
buf ( n430210 , n84531 );
buf ( n430211 , n430210 );
nand ( n84534 , n430207 , n430211 );
buf ( n430213 , n84534 );
buf ( n430214 , n430213 );
nand ( n84537 , n84525 , n430214 );
buf ( n430216 , n84537 );
buf ( n430217 , n430216 );
xnor ( n84540 , n84281 , n430217 );
buf ( n430219 , n84540 );
buf ( n430220 , n430219 );
xor ( n84543 , n84263 , n430220 );
buf ( n430222 , n84543 );
buf ( n430223 , n430222 );
buf ( n430224 , n84095 );
not ( n84547 , n430224 );
or ( n84550 , n84547 , C0 );
buf ( n430227 , C1 );
buf ( n430228 , n430227 );
nand ( n84556 , n84550 , n430228 );
buf ( n430230 , n84556 );
buf ( n430231 , n430230 );
buf ( n430232 , n429909 );
xnor ( n84560 , n430231 , n430232 );
buf ( n430234 , n84560 );
buf ( n430235 , n430234 );
buf ( n430236 , C1 );
buf ( n430237 , n430236 );
xor ( n84584 , n430235 , n430237 );
xor ( n84585 , n429897 , n429904 );
xor ( n84586 , n84585 , n429906 );
buf ( n430241 , n84586 );
buf ( n430242 , n430241 );
not ( n84589 , n430242 );
buf ( n430244 , C0 );
buf ( n430245 , C1 );
buf ( n430246 , n430245 );
nand ( n84613 , n84589 , n430246 );
buf ( n430248 , n84613 );
buf ( n430249 , n430248 );
xor ( n84616 , n84451 , n84464 );
xor ( n84617 , n84616 , n84519 );
buf ( n430252 , n84617 );
and ( n84619 , n430249 , n430252 );
buf ( n430254 , C0 );
buf ( n430255 , n430254 );
nor ( n84626 , n84619 , n430255 );
buf ( n430257 , n84626 );
buf ( n430258 , n430257 );
and ( n84629 , n84584 , n430258 );
and ( n84630 , n430235 , n430237 );
or ( n84631 , n84629 , n84630 );
buf ( n430262 , n84631 );
buf ( n430263 , n430262 );
or ( n84634 , n430223 , n430263 );
buf ( n430265 , n84634 );
not ( n84636 , n430265 );
xor ( n84637 , n430052 , n430069 );
xor ( n84638 , n84637 , n430124 );
buf ( n430269 , n84638 );
buf ( n430270 , n430269 );
buf ( n430271 , n409516 );
buf ( n430272 , n623 );
nand ( n84643 , n430271 , n430272 );
buf ( n430274 , n84643 );
buf ( n430275 , n430274 );
not ( n84646 , n430275 );
buf ( n430277 , n430078 );
buf ( n430278 , n410721 );
or ( n84649 , n430277 , n430278 );
buf ( n430280 , n410724 );
nand ( n84651 , n84649 , n430280 );
buf ( n430282 , n84651 );
buf ( n430283 , n430282 );
nand ( n430284 , n84646 , n430283 );
buf ( n430285 , n430284 );
buf ( n430286 , n430285 );
not ( n84657 , n430286 );
or ( n84674 , n84657 , C0 );
xor ( n84675 , n430087 , n430101 );
xor ( n84676 , n84675 , n430119 );
buf ( n430291 , n84676 );
buf ( n430292 , n430291 );
nand ( n84679 , n84674 , n430292 );
buf ( n430294 , n84679 );
buf ( n430295 , n430294 );
buf ( n430296 , C1 );
buf ( n430297 , n430296 );
nand ( n84687 , n430295 , n430297 );
buf ( n430299 , n84687 );
buf ( n430300 , n430299 );
xor ( n84690 , n430270 , n430300 );
not ( n84693 , n50533 );
and ( n84695 , n84693 , C1 );
or ( n84696 , C0 , n84695 );
and ( n84697 , n50532 , n84696 );
not ( n84698 , n50532 );
not ( n84701 , n22497 );
and ( n84703 , n84701 , C1 );
or ( n84704 , C0 , n84703 );
and ( n84705 , n84698 , n84704 );
or ( n84706 , n84697 , n84705 );
nor ( n84707 , n84706 , n402819 );
buf ( n430313 , n84707 );
and ( n84709 , n84690 , n430313 );
and ( n84710 , n430270 , n430300 );
or ( n84711 , n84709 , n84710 );
buf ( n430317 , n84711 );
buf ( n430318 , n430317 );
buf ( n430319 , C0 );
buf ( n430320 , n430319 );
xor ( n84735 , n430318 , n430320 );
not ( n84736 , n430128 );
not ( n84737 , n430140 );
or ( n84738 , n84736 , n84737 );
or ( n84739 , n430140 , n430128 );
nand ( n84740 , n84738 , n84739 );
and ( n84741 , n84346 , n84740 );
not ( n84742 , n84346 );
not ( n84743 , n84740 );
and ( n84744 , n84742 , n84743 );
nor ( n84745 , n84741 , n84744 );
buf ( n430332 , n84745 );
and ( n84747 , n84735 , n430332 );
or ( n84749 , n84747 , C0 );
buf ( n430335 , n84749 );
buf ( n430336 , n430335 );
not ( n84752 , n51553 );
not ( n84753 , n430025 );
or ( n84754 , n84752 , n84753 );
and ( n84755 , n402819 , n429239 );
not ( n84756 , n402819 );
and ( n84757 , n84756 , n47891 );
nor ( n84758 , n84755 , n84757 );
nand ( n84759 , n84758 , n50578 );
nand ( n84760 , n84754 , n84759 );
buf ( n430346 , n84760 );
buf ( n430347 , C0 );
buf ( n430348 , n430347 );
buf ( n430349 , n430282 );
not ( n84784 , n430349 );
buf ( n430351 , n430274 );
not ( n84786 , n430351 );
or ( n84787 , n84784 , n84786 );
buf ( n430354 , n430274 );
buf ( n430355 , n430282 );
or ( n84790 , n430354 , n430355 );
nand ( n84791 , n84787 , n84790 );
buf ( n430358 , n84791 );
buf ( n430359 , n430358 );
buf ( n430360 , n62499 );
buf ( n430361 , n410721 );
buf ( n430362 , n422315 );
nor ( n84797 , n430361 , n430362 );
buf ( n430364 , n84797 );
buf ( n430365 , n430364 );
nor ( n84800 , n430360 , n430365 );
buf ( n430367 , n84800 );
buf ( n430368 , n430367 );
buf ( n430369 , n410724 );
buf ( n430370 , n623 );
or ( n84805 , n430369 , n430370 );
buf ( n430372 , n410729 );
nand ( n84807 , n84805 , n430372 );
buf ( n430374 , n84807 );
buf ( n430375 , n430374 );
buf ( n430376 , C0 );
buf ( n430377 , C0 );
buf ( n430378 , n430377 );
and ( n84819 , n430368 , n430375 );
or ( n84820 , C0 , n84819 );
buf ( n430381 , n84820 );
buf ( n430382 , n430381 );
buf ( n430383 , C0 );
buf ( n430384 , n430383 );
and ( n84830 , n430359 , n430382 );
or ( n84831 , C0 , n84830 );
buf ( n430387 , n84831 );
buf ( n430388 , n430387 );
buf ( n430389 , n430285 );
not ( n84837 , n430389 );
buf ( n430391 , n430291 );
not ( n84839 , n430391 );
or ( n84840 , n84837 , n84839 );
buf ( n430394 , n430291 );
buf ( n430395 , n430285 );
or ( n84843 , n430394 , n430395 );
nand ( n84844 , n84840 , n84843 );
buf ( n430398 , n84844 );
buf ( n430399 , n430398 );
not ( n84847 , n430399 );
or ( n84848 , C0 , n84847 );
nand ( n84852 , n84848 , C1 );
buf ( n430403 , n84852 );
buf ( n430404 , n430403 );
buf ( n430405 , C0 );
buf ( n430406 , n430405 );
and ( n84874 , n430388 , n430404 );
or ( n84875 , C0 , n84874 );
buf ( n430409 , n84875 );
buf ( n430410 , n430409 );
xor ( n84878 , n430348 , n430410 );
xor ( n84879 , n430270 , n430300 );
xor ( n84880 , n84879 , n430313 );
buf ( n430414 , n84880 );
buf ( n430415 , n430414 );
and ( n84883 , n84878 , n430415 );
or ( n84885 , n84883 , C0 );
buf ( n430418 , n84885 );
buf ( n430419 , n430418 );
xor ( n84888 , n430346 , n430419 );
xor ( n84889 , n430318 , n430320 );
xor ( n84890 , n84889 , n430332 );
buf ( n430423 , n84890 );
buf ( n430424 , n430423 );
and ( n84893 , n84888 , n430424 );
and ( n84894 , n430346 , n430419 );
or ( n84895 , n84893 , n84894 );
buf ( n430428 , n84895 );
buf ( n430429 , n430428 );
xor ( n84898 , n430336 , n430429 );
buf ( n430431 , n430189 );
not ( n84900 , n430431 );
buf ( n430433 , n430171 );
and ( n84906 , C1 , n430433 );
nor ( n84907 , C0 , n84906 );
buf ( n430436 , n84907 );
buf ( n430437 , n430436 );
not ( n84910 , n430437 );
buf ( n430439 , n84910 );
buf ( n430440 , n430439 );
not ( n84913 , n430440 );
or ( n84914 , n84900 , n84913 );
buf ( n430443 , n84506 );
buf ( n430444 , n430436 );
nand ( n84917 , n430443 , n430444 );
buf ( n430446 , n84917 );
buf ( n430447 , n430446 );
nand ( n84920 , n84914 , n430447 );
buf ( n430449 , n84920 );
buf ( n430450 , n430449 );
and ( n84923 , n84898 , n430450 );
or ( n84925 , n84923 , C0 );
buf ( n430453 , n84925 );
buf ( n430454 , n430453 );
xor ( n84966 , n430388 , n430404 );
xor ( n84967 , n84966 , n430406 );
buf ( n430457 , n84967 );
buf ( n430458 , n430457 );
xor ( n84970 , n430359 , n430382 );
xor ( n84971 , n84970 , n430384 );
buf ( n430461 , n84971 );
buf ( n430462 , n430461 );
buf ( n430463 , C0 );
buf ( n430464 , n430463 );
xor ( n84976 , n430368 , n430375 );
xor ( n84977 , n84976 , n430378 );
buf ( n430467 , n84977 );
buf ( n430468 , n430467 );
buf ( n430469 , C0 );
buf ( n430470 , n430469 );
buf ( n430471 , C0 );
buf ( n430472 , n430471 );
buf ( n430473 , C0 );
buf ( n430474 , n430473 );
buf ( n430475 , C0 );
buf ( n430476 , n430475 );
buf ( n430477 , C0 );
buf ( n430478 , n430477 );
buf ( n430479 , C0 );
xor ( n85039 , n430348 , n430410 );
xor ( n85040 , n85039 , n430415 );
buf ( n430482 , n85040 );
buf ( n430483 , n430482 );
buf ( n430484 , C0 );
buf ( n430485 , n430484 );
nor ( n85060 , n430483 , n430485 );
buf ( n430487 , n85060 );
buf ( n430488 , C1 );
xor ( n85073 , n430346 , n430419 );
xor ( n85074 , n85073 , n430424 );
buf ( n430491 , n85074 );
buf ( n430492 , n430491 );
xor ( n85083 , n430336 , n430429 );
xor ( n85084 , n85083 , n430450 );
buf ( n430495 , n85084 );
buf ( n430496 , n430495 );
buf ( n430497 , C0 );
buf ( n430498 , n430497 );
xor ( n85092 , n430454 , n430498 );
buf ( n430500 , n430244 );
buf ( n430501 , n430241 );
xor ( n85095 , n430500 , n430501 );
buf ( n430503 , n84617 );
xor ( n85097 , n85095 , n430503 );
buf ( n430505 , n85097 );
buf ( n430506 , n430505 );
and ( n85100 , n85092 , n430506 );
or ( n85102 , n85100 , C0 );
buf ( n430509 , n85102 );
not ( n85104 , n430509 );
xor ( n85105 , n430235 , n430237 );
xor ( n85106 , n85105 , n430258 );
buf ( n430513 , n85106 );
buf ( n430514 , n430513 );
buf ( n430515 , n429998 );
not ( n85110 , n430515 );
buf ( n430517 , n430206 );
not ( n85112 , n430517 );
or ( n85113 , n85110 , n85112 );
buf ( n430520 , n429991 );
buf ( n430521 , n430210 );
nand ( n85116 , n430520 , n430521 );
buf ( n430523 , n85116 );
buf ( n430524 , n430523 );
nand ( n85119 , n85113 , n430524 );
buf ( n430526 , n85119 );
xnor ( n85121 , n430526 , n84522 );
buf ( n430528 , n85121 );
nand ( n85123 , n430514 , n430528 );
buf ( n430530 , n85123 );
not ( n85125 , n430530 );
or ( n85126 , n85104 , n85125 );
buf ( n430533 , n430513 );
buf ( n430534 , n85121 );
or ( n85129 , n430533 , n430534 );
buf ( n430536 , n85129 );
nand ( n85131 , n85126 , n430536 );
buf ( n430538 , n85131 );
buf ( n430539 , n430222 );
buf ( n430540 , n430262 );
nand ( n85135 , n430539 , n430540 );
buf ( n430542 , n85135 );
buf ( n430543 , n430542 );
nand ( n85138 , n430538 , n430543 );
buf ( n430545 , n85138 );
not ( n85140 , n430545 );
or ( n85141 , n84636 , n85140 );
buf ( n430548 , n429926 );
buf ( n430549 , n429921 );
xor ( n85144 , n430548 , n430549 );
buf ( n430551 , n429678 );
xor ( n85146 , n85144 , n430551 );
buf ( n430553 , n85146 );
buf ( n430554 , n430553 );
not ( n85149 , n430554 );
buf ( n430556 , n429980 );
buf ( n430557 , n429984 );
or ( n85166 , n430556 , n430557 );
buf ( n430559 , n430216 );
nand ( n85168 , n85166 , n430559 );
buf ( n430561 , n85168 );
buf ( n430562 , n430561 );
buf ( n430563 , C1 );
buf ( n430564 , n430563 );
nand ( n85176 , n430562 , n430564 );
buf ( n430566 , n85176 );
xor ( n85178 , C1 , n430566 );
buf ( n430568 , n85178 );
not ( n85180 , n430568 );
and ( n85181 , n85149 , n85180 );
buf ( n430571 , n430553 );
buf ( n430572 , n85178 );
and ( n85184 , n430571 , n430572 );
nor ( n85185 , n85181 , n85184 );
buf ( n430575 , n85185 );
xor ( n85187 , n429976 , n429978 );
and ( n85188 , n85187 , n430220 );
and ( n85189 , n429976 , n429978 );
or ( n85190 , n85188 , n85189 );
buf ( n430580 , n85190 );
nand ( n85192 , n430575 , n430580 );
nand ( n85193 , n85141 , n85192 );
buf ( n430583 , n85193 );
buf ( n430584 , n430575 );
buf ( n430585 , n430580 );
or ( n85197 , n430584 , n430585 );
buf ( n430587 , n85197 );
buf ( n430588 , n430587 );
nand ( n85200 , n430583 , n430588 );
buf ( n430590 , n85200 );
not ( n85202 , n430590 );
buf ( n430592 , n429956 );
not ( n85204 , n430592 );
buf ( n430594 , n429942 );
not ( n85206 , n430594 );
and ( n85207 , n85204 , n85206 );
buf ( n430597 , n429956 );
buf ( n430598 , n429942 );
and ( n85210 , n430597 , n430598 );
nor ( n85211 , n85207 , n85210 );
buf ( n430601 , n85211 );
buf ( n430602 , n430601 );
not ( n85214 , n430602 );
buf ( n430604 , n429947 );
not ( n85216 , n430604 );
and ( n85217 , n85214 , n85216 );
buf ( n430607 , n430601 );
buf ( n430608 , n429947 );
and ( n85220 , n430607 , n430608 );
nor ( n85221 , n85217 , n85220 );
buf ( n430611 , n85221 );
buf ( n430612 , n430611 );
buf ( n430613 , n430553 );
buf ( n430614 , n430566 );
not ( n85226 , n430614 );
buf ( n430616 , C1 );
nand ( n85228 , n85226 , n430616 );
buf ( n430618 , n85228 );
buf ( n430619 , n430618 );
nand ( n85231 , n430613 , n430619 );
buf ( n430621 , n85231 );
buf ( n430622 , n430621 );
buf ( n430623 , C1 );
buf ( n430624 , n430623 );
and ( n85240 , n430622 , n430624 );
buf ( n430626 , n85240 );
buf ( n430627 , n430626 );
nand ( n85243 , n430612 , n430627 );
buf ( n430629 , n85243 );
not ( n85245 , n430629 );
or ( n85246 , n85202 , n85245 );
buf ( n430632 , n430611 );
not ( n85248 , n430632 );
buf ( n430634 , n85248 );
buf ( n430635 , n430634 );
buf ( n430636 , n430626 );
not ( n85252 , n430636 );
buf ( n430638 , n85252 );
buf ( n430639 , n430638 );
nand ( n85255 , n430635 , n430639 );
buf ( n430641 , n85255 );
nand ( n85257 , n85246 , n430641 );
buf ( n430643 , n85257 );
xor ( n85259 , n429969 , n430643 );
buf ( n430645 , C0 );
buf ( n430646 , n430645 );
xor ( n85280 , n429590 , n429594 );
xor ( n85281 , n85280 , n429596 );
buf ( n430649 , n85281 );
buf ( n430650 , n430649 );
xor ( n85284 , n430646 , n430650 );
xor ( n85285 , n429442 , n429513 );
xor ( n85286 , n85285 , n429542 );
buf ( n430654 , n85286 );
buf ( n430655 , n430654 );
xor ( n85289 , n85284 , n430655 );
buf ( n430657 , n85289 );
buf ( n430658 , n430657 );
and ( n85292 , n85259 , n430658 );
and ( n85293 , n429969 , n430643 );
or ( n85294 , n85292 , n85293 );
buf ( n430662 , n85294 );
buf ( n430663 , n430662 );
not ( n85297 , n430663 );
buf ( n430665 , n85297 );
buf ( n430666 , n430665 );
xor ( n85300 , n429547 , n429583 );
xor ( n85301 , n85300 , n429609 );
buf ( n430669 , n85301 );
buf ( n430670 , n430669 );
xor ( n85304 , n430646 , n430650 );
and ( n85305 , n85304 , n430655 );
or ( n85307 , n85305 , C0 );
buf ( n430674 , n85307 );
buf ( n430675 , n430674 );
nor ( n85310 , n430670 , n430675 );
buf ( n430677 , n85310 );
buf ( n430678 , n430677 );
or ( n85313 , n430666 , n430678 );
buf ( n430680 , n430669 );
buf ( n430681 , n430674 );
nand ( n85316 , n430680 , n430681 );
buf ( n430683 , n85316 );
buf ( n430684 , n430683 );
nand ( n85319 , n85313 , n430684 );
buf ( n430686 , n85319 );
not ( n85321 , n430686 );
or ( n85322 , n429675 , n85321 );
buf ( n430689 , n429671 );
not ( n85324 , n430689 );
buf ( n430691 , n429613 );
nand ( n85326 , n85324 , n430691 );
buf ( n430693 , n85326 );
nand ( n85328 , n85322 , n430693 );
not ( n85329 , n85328 );
buf ( n430696 , n429656 );
not ( n85331 , n430696 );
buf ( n430698 , n429663 );
nand ( n85333 , n85331 , n430698 );
buf ( n430700 , n85333 );
buf ( n430701 , n430700 );
not ( n85336 , n430701 );
buf ( n430703 , n429653 );
not ( n85338 , n430703 );
or ( n85339 , n85336 , n85338 );
buf ( n430706 , n429660 );
buf ( n430707 , n429656 );
nand ( n85342 , n430706 , n430707 );
buf ( n430709 , n85342 );
buf ( n430710 , n430709 );
nand ( n85345 , n85339 , n430710 );
buf ( n430712 , n85345 );
buf ( n430713 , n430712 );
not ( n85348 , n430713 );
and ( n85351 , n429621 , n429648 );
or ( n85352 , C0 , n85351 );
buf ( n430717 , n85352 );
buf ( n430718 , n430717 );
xor ( n85355 , n428952 , n428954 );
xor ( n85356 , n85355 , n428962 );
buf ( n430721 , n85356 );
buf ( n430722 , n430721 );
and ( n85359 , n430718 , n430722 );
not ( n85360 , n430718 );
buf ( n430725 , n430721 );
not ( n85362 , n430725 );
buf ( n430727 , n85362 );
buf ( n430728 , n430727 );
and ( n85365 , n85360 , n430728 );
or ( n85366 , n85359 , n85365 );
buf ( n430731 , n85366 );
buf ( n430732 , n430731 );
not ( n85369 , n430732 );
xor ( n85370 , n429062 , n429066 );
xor ( n85371 , n85370 , n429068 );
buf ( n430736 , n85371 );
buf ( n430737 , n430736 );
not ( n85374 , n430737 );
and ( n85375 , n85369 , n85374 );
buf ( n430740 , n430731 );
buf ( n430741 , n430736 );
and ( n85378 , n430740 , n430741 );
nor ( n85379 , n85375 , n85378 );
buf ( n430744 , n85379 );
buf ( n430745 , n430744 );
nand ( n85382 , n85348 , n430745 );
buf ( n430747 , n85382 );
not ( n85384 , n430747 );
or ( n85385 , n85329 , n85384 );
buf ( n430750 , n430744 );
not ( n85387 , n430750 );
buf ( n430752 , n430712 );
nand ( n85389 , n85387 , n430752 );
buf ( n430754 , n85389 );
nand ( n85391 , n85385 , n430754 );
buf ( n430756 , n430721 );
not ( n85393 , n430756 );
buf ( n430758 , n430717 );
not ( n85395 , n430758 );
or ( n85396 , n85393 , n85395 );
buf ( n430761 , n430736 );
buf ( n430762 , n430717 );
not ( n85399 , n430762 );
buf ( n430764 , n430727 );
nand ( n85401 , n85399 , n430764 );
buf ( n430766 , n85401 );
buf ( n430767 , n430766 );
nand ( n85404 , n430761 , n430767 );
buf ( n430769 , n85404 );
buf ( n430770 , n430769 );
nand ( n85407 , n85396 , n430770 );
buf ( n430772 , n85407 );
not ( n85409 , n430772 );
xor ( n85410 , n429072 , n429076 );
xor ( n85411 , n85410 , n429081 );
buf ( n430776 , n85411 );
not ( n85413 , n430776 );
nand ( n85414 , n85409 , n85413 );
and ( n85415 , n85391 , n85414 );
and ( n85416 , n430776 , n430772 );
nor ( n85417 , n85415 , n85416 );
or ( n85418 , n429088 , n85417 );
buf ( n430783 , n83049 );
buf ( n430784 , n429085 );
nand ( n85421 , n430783 , n430784 );
buf ( n430786 , n85421 );
nand ( n85423 , n85418 , n430786 );
not ( n85424 , n85423 );
or ( n85425 , n428997 , n85424 );
buf ( n430790 , n83044 );
buf ( n430791 , n428988 );
or ( n85428 , n430790 , n430791 );
buf ( n430793 , n85428 );
nand ( n85430 , n85425 , n430793 );
not ( n85431 , n85430 );
or ( n85432 , n82952 , n85431 );
buf ( n430797 , n428925 );
not ( n85434 , n430797 );
buf ( n430799 , n428911 );
nand ( n85436 , n85434 , n430799 );
buf ( n430801 , n85436 );
nand ( n85438 , n85432 , n430801 );
buf ( n430803 , n85438 );
and ( n85440 , n82492 , n430803 );
and ( n85441 , n428480 , n428484 );
or ( n85442 , n85440 , n85441 );
buf ( n430807 , n85442 );
buf ( n430808 , n430807 );
and ( n85445 , n82002 , n430808 );
and ( n85446 , n428051 , n428055 );
or ( n85447 , n85445 , n85446 );
buf ( n430812 , n85447 );
buf ( n430813 , n430812 );
and ( n85450 , n81845 , n430813 );
and ( n85451 , n427928 , n427932 );
or ( n85452 , n85450 , n85451 );
buf ( n430817 , n85452 );
buf ( n430818 , n430817 );
and ( n85455 , n81492 , n430818 );
and ( n85456 , n427610 , n427614 );
or ( n85457 , n85455 , n85456 );
buf ( n430822 , n85457 );
buf ( n430823 , n430822 );
and ( n85460 , n81302 , n430823 );
and ( n85461 , n427447 , n427450 );
or ( n85462 , n85460 , n85461 );
buf ( n430827 , n85462 );
not ( n85464 , n430827 );
or ( n85465 , n81038 , n85464 );
not ( n85466 , n81036 );
nand ( n85467 , n85466 , n81021 );
nand ( n85468 , n85465 , n85467 );
nand ( n85469 , n426648 , n85468 , n80450 );
or ( n85470 , n426634 , n426639 );
nand ( n85471 , n80451 , n85469 , n85470 );
xor ( n85472 , n421599 , n421614 );
xor ( n85473 , n85472 , n421921 );
buf ( n430838 , n85473 );
buf ( n430839 , n430838 );
xor ( n85476 , n426600 , n426604 );
and ( n85477 , n85476 , n426622 );
and ( n85478 , n426600 , n426604 );
or ( n85479 , n85477 , n85478 );
buf ( n430844 , n85479 );
buf ( n430845 , n430844 );
xor ( n85482 , n430839 , n430845 );
xor ( n85483 , n422882 , n422886 );
buf ( n430848 , n85483 );
buf ( n430849 , n430848 );
buf ( n430850 , n422873 );
and ( n85487 , n430849 , n430850 );
not ( n85488 , n430849 );
buf ( n430853 , n422873 );
not ( n85490 , n430853 );
buf ( n430855 , n85490 );
buf ( n430856 , n430855 );
and ( n85493 , n85488 , n430856 );
nor ( n85494 , n85487 , n85493 );
buf ( n430859 , n85494 );
buf ( n430860 , n430859 );
xor ( n85497 , n85482 , n430860 );
buf ( n430862 , n85497 );
buf ( n430863 , n430862 );
buf ( n430864 , n426591 );
not ( n85501 , n430864 );
buf ( n430866 , n426627 );
not ( n85503 , n430866 );
or ( n85504 , n85501 , n85503 );
buf ( n430869 , n426585 );
nand ( n85506 , n85504 , n430869 );
buf ( n430871 , n85506 );
buf ( n430872 , n430871 );
buf ( n430873 , n426624 );
buf ( n430874 , n426588 );
nand ( n85511 , n430873 , n430874 );
buf ( n430876 , n85511 );
buf ( n430877 , n430876 );
nand ( n85514 , n430872 , n430877 );
buf ( n430879 , n85514 );
buf ( n430880 , n430879 );
nor ( n85517 , n430863 , n430880 );
buf ( n430882 , n85517 );
not ( n85519 , n430882 );
nand ( n85520 , n85471 , n85519 );
buf ( n430885 , n85520 );
xor ( n85522 , n430839 , n430845 );
and ( n85523 , n85522 , n430860 );
and ( n85524 , n430839 , n430845 );
or ( n85525 , n85523 , n85524 );
buf ( n430890 , n85525 );
buf ( n430891 , n430890 );
not ( n85528 , n430891 );
buf ( n430893 , n422891 );
not ( n85530 , n430893 );
buf ( n430895 , n421133 );
not ( n85532 , n430895 );
or ( n85533 , n85530 , n85532 );
buf ( n430898 , n421133 );
buf ( n430899 , n422891 );
or ( n85536 , n430898 , n430899 );
nand ( n85537 , n85533 , n85536 );
buf ( n430902 , n85537 );
xor ( n85539 , n421935 , n430902 );
buf ( n430904 , n85539 );
nand ( n85541 , n85528 , n430904 );
buf ( n430906 , n85541 );
buf ( n430907 , n430906 );
not ( n85544 , n430907 );
buf ( n430909 , n85544 );
buf ( n430910 , n430909 );
or ( n85547 , n430885 , n430910 );
buf ( n430912 , n430906 );
nand ( n85549 , n430862 , n430879 );
not ( n85550 , n85549 );
buf ( n430915 , n85550 );
and ( n85552 , n430912 , n430915 );
not ( n85553 , n430890 );
nor ( n85554 , n85553 , n85539 );
buf ( n430919 , n85554 );
nor ( n85556 , n85552 , n430919 );
buf ( n430921 , n85556 );
buf ( n430922 , n430921 );
nand ( n85559 , n85547 , n430922 );
buf ( n430924 , n85559 );
buf ( n430925 , n430924 );
and ( n85562 , n76985 , n430925 );
and ( n85563 , n422907 , n423399 );
or ( n85564 , n85562 , n85563 );
buf ( n430929 , n85564 );
buf ( n430930 , n430929 );
not ( n85567 , n430930 );
xor ( n85568 , n423157 , n423158 );
and ( n85569 , n85568 , n423165 );
or ( n85571 , n85569 , C0 );
buf ( n430935 , n85571 );
buf ( n430936 , n430935 );
buf ( n430937 , n423223 );
not ( n85575 , n430937 );
buf ( n430939 , n393544 );
not ( n85577 , n430939 );
or ( n85578 , n85575 , n85577 );
buf ( n430942 , n399274 );
buf ( n430943 , n388962 );
and ( n430944 , n430942 , n430943 );
not ( n85582 , n430942 );
buf ( n430946 , n393525 );
and ( n85584 , n85582 , n430946 );
nor ( n430948 , n430944 , n85584 );
buf ( n430949 , n430948 );
buf ( n430950 , n430949 );
buf ( n430951 , n51692 );
nand ( n430952 , n430950 , n430951 );
buf ( n430953 , n430952 );
buf ( n430954 , n430953 );
nand ( n85592 , n85578 , n430954 );
buf ( n430956 , n85592 );
buf ( n430957 , n430956 );
buf ( n430958 , n45954 );
not ( n85596 , n430958 );
buf ( n430960 , n393369 );
not ( n85598 , n430960 );
buf ( n430962 , n388409 );
not ( n85600 , n430962 );
or ( n430964 , n85598 , n85600 );
buf ( n430965 , n388406 );
buf ( n430966 , n393381 );
nand ( n85604 , n430965 , n430966 );
buf ( n430968 , n85604 );
buf ( n430969 , n430968 );
nand ( n430970 , n430964 , n430969 );
buf ( n430971 , n430970 );
buf ( n430972 , n430971 );
not ( n85610 , n430972 );
or ( n430974 , n85596 , n85610 );
buf ( n430975 , n423375 );
buf ( n430976 , n45949 );
nand ( n85614 , n430975 , n430976 );
buf ( n430978 , n85614 );
buf ( n430979 , n430978 );
nand ( n430980 , n430974 , n430979 );
buf ( n430981 , n430980 );
buf ( n430982 , n430981 );
xor ( n85620 , n430957 , n430982 );
xor ( n430984 , n423246 , n423303 );
and ( n85622 , n430984 , n423310 );
and ( n430986 , n423246 , n423303 );
or ( n85624 , n85622 , n430986 );
buf ( n430988 , n85624 );
buf ( n430989 , n430988 );
xor ( n430990 , n85620 , n430989 );
buf ( n430991 , n430990 );
buf ( n430992 , n430991 );
xor ( n85630 , n423231 , n423313 );
and ( n430994 , n85630 , n423331 );
and ( n85632 , n423231 , n423313 );
or ( n430996 , n430994 , n85632 );
buf ( n430997 , n430996 );
buf ( n430998 , n430997 );
buf ( n430999 , C1 );
buf ( n431000 , n430999 );
and ( n431001 , n430998 , n431000 );
nor ( n431002 , n431001 , C0 );
buf ( n431003 , n431002 );
buf ( n431004 , n431003 );
xor ( n431005 , n430992 , n431004 );
buf ( n431006 , n431005 );
buf ( n431007 , n431006 );
not ( n85674 , n431007 );
buf ( n431009 , n85674 );
buf ( n431010 , n431009 );
or ( n85677 , n430936 , n431010 );
xor ( n85678 , n423334 , n423338 );
and ( n85679 , n85678 , n423390 );
and ( n85680 , n423334 , n423338 );
or ( n85681 , n85679 , n85680 );
buf ( n431016 , n85681 );
buf ( n431017 , n431016 );
nand ( n85684 , n85677 , n431017 );
buf ( n431019 , n85684 );
buf ( n431020 , n431019 );
buf ( n431021 , n430935 );
buf ( n431022 , n431009 );
nand ( n85689 , n431021 , n431022 );
buf ( n431024 , n85689 );
buf ( n431025 , n431024 );
and ( n431026 , n431020 , n431025 );
buf ( n431027 , n431026 );
buf ( n431028 , n431027 );
xor ( n85695 , n422975 , n422977 );
and ( n85696 , n85695 , n422995 );
or ( n85698 , n85696 , C0 );
buf ( n431032 , n85698 );
not ( n85700 , n76935 );
not ( n85701 , n85700 );
not ( n85702 , n76944 );
or ( n85703 , n85701 , n85702 );
not ( n85704 , n76935 );
not ( n85705 , n76944 );
not ( n85706 , n85705 );
or ( n85707 , n85704 , n85706 );
nand ( n431041 , n85707 , n76966 );
nand ( n85709 , n85703 , n431041 );
buf ( n431043 , n413643 );
not ( n85711 , n431043 );
buf ( n431045 , n399986 );
not ( n85713 , n431045 );
buf ( n431047 , n45699 );
not ( n85715 , n431047 );
or ( n85716 , n85713 , n85715 );
buf ( n431050 , n27301 );
buf ( n431051 , n44776 );
nand ( n85719 , n431050 , n431051 );
buf ( n431053 , n85719 );
buf ( n431054 , n431053 );
nand ( n85722 , n85716 , n431054 );
buf ( n431056 , n85722 );
buf ( n431057 , n431056 );
not ( n85725 , n431057 );
or ( n85726 , n85711 , n85725 );
buf ( n431060 , n422921 );
buf ( n431061 , n45260 );
nand ( n85729 , n431060 , n431061 );
buf ( n431063 , n85729 );
buf ( n431064 , n431063 );
nand ( n85732 , n85726 , n431064 );
buf ( n431066 , n85732 );
not ( n85734 , n431066 );
not ( n85735 , n85734 );
not ( n85736 , n423043 );
not ( n85737 , n423059 );
or ( n85738 , n85736 , n85737 );
buf ( n431072 , n423043 );
buf ( n431073 , n423059 );
nor ( n85741 , n431072 , n431073 );
buf ( n431075 , n85741 );
or ( n85743 , n431075 , n423120 );
nand ( n85744 , n85738 , n85743 );
not ( n85745 , n85744 );
buf ( n431079 , n422949 );
not ( n85747 , n431079 );
buf ( n431081 , n396622 );
not ( n85749 , n431081 );
or ( n85750 , n85747 , n85749 );
buf ( n431084 , n394817 );
not ( n85752 , n431084 );
buf ( n431086 , n398298 );
not ( n85754 , n431086 );
or ( n431088 , n85752 , n85754 );
buf ( n431089 , n399167 );
buf ( n431090 , n394814 );
nand ( n85758 , n431089 , n431090 );
buf ( n431092 , n85758 );
buf ( n431093 , n431092 );
nand ( n85761 , n431088 , n431093 );
buf ( n431095 , n85761 );
buf ( n431096 , n431095 );
buf ( n431097 , n46921 );
nand ( n85765 , n431096 , n431097 );
buf ( n431099 , n85765 );
buf ( n431100 , n431099 );
nand ( n85768 , n85750 , n431100 );
buf ( n431102 , n85768 );
not ( n85770 , n431102 );
not ( n85771 , n85770 );
or ( n85772 , n85745 , n85771 );
not ( n85773 , n85744 );
nand ( n85774 , n431102 , n85773 );
nand ( n85775 , n85772 , n85774 );
not ( n85776 , n85775 );
or ( n85777 , n85735 , n85776 );
or ( n85778 , n85775 , n85734 );
nand ( n85779 , n85777 , n85778 );
and ( n85780 , n85709 , n85779 );
not ( n431114 , n85709 );
not ( n85782 , n85779 );
and ( n85783 , n431114 , n85782 );
nor ( n85784 , n85780 , n85783 );
xor ( n85785 , n423122 , n423147 );
and ( n85786 , n85785 , n423154 );
and ( n85787 , n423122 , n423147 );
or ( n85788 , n85786 , n85787 );
buf ( n431122 , n85788 );
and ( n85790 , n85784 , n431122 );
not ( n85791 , n85784 );
buf ( n431125 , n431122 );
not ( n85793 , n431125 );
buf ( n431127 , n85793 );
and ( n85795 , n85791 , n431127 );
nor ( n85796 , n85790 , n85795 );
xnor ( n85797 , n431032 , n85796 );
buf ( n431131 , n85797 );
xor ( n85799 , n422932 , n422957 );
and ( n85800 , n85799 , n422972 );
and ( n85801 , n422932 , n422957 );
or ( n85802 , n85800 , n85801 );
buf ( n431136 , n85802 );
buf ( n431137 , n431136 );
buf ( n431138 , n47891 );
not ( n85806 , n431138 );
buf ( n431140 , n390271 );
not ( n85808 , n431140 );
or ( n85809 , n85806 , n85808 );
buf ( n431143 , n388892 );
buf ( n431144 , n61299 );
nand ( n85812 , n431143 , n431144 );
buf ( n431146 , n85812 );
buf ( n431147 , n431146 );
nand ( n85815 , n85809 , n431147 );
buf ( n431149 , n85815 );
buf ( n431150 , n431149 );
buf ( n431151 , n61577 );
and ( n431152 , n431150 , n431151 );
buf ( n431153 , n423325 );
buf ( n431154 , n50580 );
nor ( n85822 , n431153 , n431154 );
buf ( n431156 , n85822 );
buf ( n431157 , n431156 );
nor ( n85825 , n431152 , n431157 );
buf ( n431159 , n85825 );
buf ( n431160 , n431159 );
not ( n85828 , n431160 );
buf ( n431162 , n85828 );
buf ( n431163 , n431162 );
xor ( n85831 , n431137 , n431163 );
not ( n85832 , n76501 );
not ( n85833 , n397102 );
or ( n85834 , n85832 , n85833 );
buf ( n431168 , n397489 );
not ( n85836 , n431168 );
buf ( n431170 , n49661 );
not ( n85838 , n431170 );
or ( n85839 , n85836 , n85838 );
buf ( n431173 , n49660 );
buf ( n431174 , n397492 );
nand ( n85842 , n431173 , n431174 );
buf ( n431176 , n85842 );
buf ( n431177 , n431176 );
nand ( n85845 , n85839 , n431177 );
buf ( n431179 , n85845 );
buf ( n431180 , n431179 );
not ( n85848 , n431180 );
buf ( n431182 , n85848 );
or ( n85850 , n431182 , n386474 );
nand ( n85851 , n85834 , n85850 );
buf ( n431185 , n385473 );
buf ( n431186 , n393109 );
not ( n85854 , n431186 );
buf ( n431188 , n85854 );
buf ( n431189 , n431188 );
nor ( n85857 , n431185 , n431189 );
buf ( n431191 , n85857 );
not ( n85859 , n431191 );
not ( n85860 , n402819 );
and ( n85861 , n85859 , n85860 );
not ( n85862 , n431188 );
not ( n85863 , n388962 );
or ( n85864 , n85862 , n85863 );
nand ( n85865 , n85864 , n388905 );
nor ( n85866 , n85861 , n85865 );
not ( n85867 , n76677 );
buf ( n431201 , n423078 );
buf ( n431202 , n423065 );
or ( n85870 , n431201 , n431202 );
buf ( n431204 , n85870 );
not ( n85872 , n431204 );
or ( n85873 , n85867 , n85872 );
buf ( n431207 , n423078 );
buf ( n431208 , n423065 );
nand ( n85876 , n431207 , n431208 );
buf ( n431210 , n85876 );
nand ( n431211 , n85873 , n431210 );
buf ( n431212 , n431211 );
xor ( n85880 , n417339 , n417367 );
xor ( n85881 , n85880 , n417393 );
buf ( n431215 , n85881 );
buf ( n431216 , n431215 );
xor ( n85884 , n431212 , n431216 );
buf ( n431218 , n423036 );
not ( n85886 , n431218 );
buf ( n431220 , n390429 );
not ( n85888 , n431220 );
or ( n85889 , n85886 , n85888 );
buf ( n431223 , n392884 );
not ( n85891 , n431223 );
buf ( n431225 , n24071 );
not ( n85893 , n431225 );
or ( n85894 , n85891 , n85893 );
buf ( n431228 , n53252 );
buf ( n431229 , n392887 );
nand ( n85897 , n431228 , n431229 );
buf ( n431231 , n85897 );
buf ( n431232 , n431231 );
nand ( n85900 , n85894 , n431232 );
buf ( n431234 , n85900 );
buf ( n431235 , n431234 );
buf ( n431236 , n42924 );
nand ( n85904 , n431235 , n431236 );
buf ( n431238 , n85904 );
buf ( n431239 , n431238 );
nand ( n85907 , n85889 , n431239 );
buf ( n431241 , n85907 );
buf ( n431242 , n431241 );
xor ( n85910 , n85884 , n431242 );
buf ( n431244 , n85910 );
nand ( n85912 , n85866 , n431244 );
and ( n85913 , n85851 , n85912 );
not ( n85914 , n85851 );
not ( n85915 , n431244 );
nand ( n85916 , n85866 , n85915 );
and ( n85917 , n85914 , n85916 );
or ( n85918 , n85913 , n85917 );
not ( n85919 , n85866 );
nand ( n85920 , n85919 , n85915 );
and ( n85921 , n85851 , n85920 );
not ( n85922 , n85851 );
not ( n85923 , n85866 );
nand ( n85924 , n85923 , n431244 );
and ( n85925 , n85922 , n85924 );
or ( n85926 , n85921 , n85925 );
nand ( n85927 , n85918 , n85926 );
buf ( n431261 , n85927 );
xnor ( n85929 , n85831 , n431261 );
buf ( n431263 , n85929 );
buf ( n431264 , n431263 );
and ( n85932 , n431131 , n431264 );
not ( n85933 , n431131 );
buf ( n431267 , n431263 );
not ( n431268 , n431267 );
buf ( n431269 , n431268 );
buf ( n431270 , n431269 );
and ( n85938 , n85933 , n431270 );
nor ( n85939 , n85932 , n85938 );
buf ( n431273 , n85939 );
not ( n85941 , n431273 );
buf ( n431275 , n358975 );
buf ( n431276 , n393117 );
and ( n85960 , n431275 , n431276 );
not ( n85961 , n431275 );
buf ( n431279 , n37346 );
and ( n85963 , n85961 , n431279 );
nor ( n85964 , n85960 , n85963 );
buf ( n431282 , n85964 );
not ( n85966 , n431282 );
not ( n85967 , n45662 );
or ( n85968 , n85966 , n85967 );
buf ( n431286 , n55055 );
not ( n85970 , n431286 );
buf ( n431288 , n391563 );
not ( n85972 , n431288 );
or ( n85973 , n85970 , n85972 );
buf ( n431291 , n393117 );
buf ( n431292 , n55054 );
nand ( n85976 , n431291 , n431292 );
buf ( n431294 , n85976 );
buf ( n431295 , n431294 );
nand ( n85979 , n85973 , n431295 );
buf ( n431297 , n85979 );
buf ( n431298 , n431297 );
buf ( n431299 , n37314 );
nand ( n85983 , n431298 , n431299 );
buf ( n431301 , n85983 );
nand ( n85985 , n85968 , n431301 );
buf ( n431303 , n85985 );
buf ( n431304 , n43515 );
not ( n85988 , n431304 );
buf ( n431306 , n411504 );
not ( n85990 , n431306 );
buf ( n431308 , n402836 );
not ( n85992 , n431308 );
or ( n85993 , n85990 , n85992 );
buf ( n431311 , n394666 );
buf ( n431312 , n391024 );
nand ( n85996 , n431311 , n431312 );
buf ( n431314 , n85996 );
buf ( n431315 , n431314 );
nand ( n85999 , n85993 , n431315 );
buf ( n431317 , n85999 );
buf ( n431318 , n431317 );
not ( n86002 , n431318 );
or ( n86003 , n85988 , n86002 );
buf ( n431321 , n76609 );
buf ( n431322 , n43536 );
nand ( n86006 , n431321 , n431322 );
buf ( n431324 , n86006 );
buf ( n431325 , n431324 );
nand ( n86009 , n86003 , n431325 );
buf ( n431327 , n86009 );
buf ( n431328 , n431327 );
xor ( n86012 , n423272 , n423293 );
and ( n86013 , n86012 , n423300 );
and ( n86014 , n423272 , n423293 );
or ( n86015 , n86013 , n86014 );
buf ( n431333 , n86015 );
buf ( n431334 , n431333 );
xor ( n86018 , n431328 , n431334 );
xor ( n86019 , n76651 , n423103 );
and ( n86020 , n86019 , n423116 );
and ( n86021 , n76651 , n423103 );
or ( n86022 , n86020 , n86021 );
buf ( n431340 , n86022 );
buf ( n431341 , n423285 );
not ( n86025 , n431341 );
buf ( n431343 , n406422 );
not ( n86027 , n431343 );
or ( n86028 , n86025 , n86027 );
nand ( n86029 , n70631 , n409076 );
buf ( n431347 , n86029 );
nand ( n86031 , n86028 , n431347 );
buf ( n431349 , n86031 );
buf ( n431350 , n431349 );
xor ( n86034 , n431340 , n431350 );
buf ( n431352 , n390362 );
not ( n86036 , n431352 );
buf ( n431354 , n417317 );
not ( n86038 , n431354 );
or ( n86039 , n86036 , n86038 );
buf ( n431357 , n423260 );
buf ( n431358 , n40592 );
nand ( n86042 , n431357 , n431358 );
buf ( n431360 , n86042 );
buf ( n431361 , n431360 );
nand ( n86045 , n86039 , n431361 );
buf ( n431363 , n86045 );
buf ( n431364 , n431363 );
xor ( n86048 , n86034 , n431364 );
buf ( n431366 , n86048 );
buf ( n431367 , n431366 );
xor ( n86051 , n86018 , n431367 );
buf ( n431369 , n86051 );
buf ( n431370 , n431369 );
xor ( n86054 , n431303 , n431370 );
buf ( n431372 , n395362 );
not ( n86056 , n431372 );
buf ( n431374 , n47863 );
not ( n86058 , n431374 );
buf ( n431376 , n43044 );
not ( n86060 , n431376 );
or ( n86061 , n86058 , n86060 );
buf ( n431379 , n27195 );
buf ( n431380 , n419385 );
nand ( n431381 , n431379 , n431380 );
buf ( n431382 , n431381 );
buf ( n431383 , n431382 );
nand ( n86067 , n86061 , n431383 );
buf ( n431385 , n86067 );
buf ( n431386 , n431385 );
not ( n86070 , n431386 );
or ( n86071 , n86056 , n86070 );
buf ( n431389 , n423139 );
buf ( n431390 , n395349 );
nand ( n86074 , n431389 , n431390 );
buf ( n431392 , n86074 );
buf ( n431393 , n431392 );
nand ( n86077 , n86071 , n431393 );
buf ( n431395 , n86077 );
buf ( n431396 , n431395 );
not ( n86080 , n431396 );
buf ( n431398 , n86080 );
buf ( n431399 , n431398 );
xor ( n86083 , n86054 , n431399 );
buf ( n431401 , n86083 );
buf ( n431402 , n431401 );
not ( n86086 , n431402 );
buf ( n431404 , n86086 );
not ( n86088 , n431404 );
or ( n86089 , C0 , n86088 );
buf ( n431407 , C1 );
nand ( n86097 , n86089 , n431407 );
buf ( n431409 , n76931 );
not ( n86099 , n431409 );
buf ( n431411 , n76967 );
not ( n86101 , n431411 );
buf ( n431413 , n86101 );
buf ( n431414 , n431413 );
not ( n86104 , n431414 );
or ( n86105 , n86099 , n86104 );
buf ( n431417 , n423349 );
not ( n86107 , n431417 );
buf ( n431419 , n76967 );
not ( n86109 , n431419 );
or ( n86110 , n86107 , n86109 );
buf ( n431422 , n423388 );
nand ( n86112 , n86110 , n431422 );
buf ( n431424 , n86112 );
buf ( n431425 , n431424 );
nand ( n86115 , n86105 , n431425 );
buf ( n431427 , n86115 );
buf ( n86117 , n431427 );
not ( n86118 , n86117 );
and ( n86119 , n86097 , n86118 );
not ( n86120 , n86097 );
and ( n86121 , n86120 , n86117 );
nor ( n86122 , n86119 , n86121 );
not ( n86123 , n86122 );
or ( n86124 , n85941 , n86123 );
buf ( n431436 , n422997 );
not ( n86126 , n431436 );
buf ( n431438 , n423014 );
nand ( n86128 , n86126 , n431438 );
buf ( n431440 , n86128 );
buf ( n431441 , n431440 );
not ( n431442 , n431441 );
buf ( n431443 , n423167 );
not ( n86133 , n431443 );
or ( n86134 , n431442 , n86133 );
buf ( n431446 , n423017 );
buf ( n431447 , n422997 );
nand ( n86137 , n431446 , n431447 );
buf ( n431449 , n86137 );
buf ( n431450 , n431449 );
nand ( n86140 , n86134 , n431450 );
buf ( n431452 , n86140 );
nand ( n86142 , n86124 , n431452 );
buf ( n431454 , n86142 );
not ( n86144 , n86122 );
buf ( n431456 , n431273 );
not ( n431457 , n431456 );
buf ( n431458 , n431457 );
nand ( n86148 , n86144 , n431458 );
buf ( n431460 , n86148 );
and ( n86150 , n431454 , n431460 );
buf ( n431462 , n86150 );
buf ( n431463 , n431462 );
xor ( n86153 , n431028 , n431463 );
not ( n86154 , n431263 );
not ( n86155 , n85796 );
and ( n86156 , n86154 , n86155 );
buf ( n431468 , n431263 );
buf ( n431469 , n85796 );
nand ( n86159 , n431468 , n431469 );
buf ( n431471 , n86159 );
and ( n86161 , n431471 , n431032 );
nor ( n86162 , n86156 , n86161 );
buf ( n431474 , n431122 );
not ( n86164 , n431474 );
buf ( n431476 , n85779 );
not ( n86166 , n431476 );
buf ( n431478 , n85709 );
nand ( n86168 , n86166 , n431478 );
buf ( n431480 , n86168 );
buf ( n431481 , n431480 );
not ( n86171 , n431481 );
or ( n86172 , n86164 , n86171 );
buf ( n431484 , n85709 );
not ( n86174 , n431484 );
buf ( n431486 , n85779 );
nand ( n86176 , n86174 , n431486 );
buf ( n431488 , n86176 );
buf ( n431489 , n431488 );
nand ( n86179 , n86172 , n431489 );
buf ( n431491 , n86179 );
buf ( n431492 , n431491 );
buf ( n431493 , n430991 );
not ( n86183 , n431493 );
buf ( n431495 , n86183 );
buf ( n431496 , n431495 );
not ( n86186 , n431496 );
or ( n86189 , n86186 , C0 );
buf ( n431499 , n430997 );
nand ( n86191 , n86189 , n431499 );
buf ( n431501 , n86191 );
buf ( n431502 , n431501 );
buf ( n431503 , C1 );
buf ( n431504 , n431503 );
nand ( n86199 , n431502 , n431504 );
buf ( n431506 , n86199 );
buf ( n431507 , n431506 );
xor ( n86202 , n431492 , n431507 );
buf ( n431509 , n431401 );
not ( n86206 , n431509 );
or ( n86207 , C0 , n86206 );
buf ( n431512 , n431427 );
nand ( n86209 , n86207 , n431512 );
buf ( n431514 , n86209 );
buf ( n431515 , n431514 );
buf ( n431516 , C1 );
buf ( n431517 , n431516 );
nand ( n86217 , n431515 , n431517 );
buf ( n431519 , n86217 );
buf ( n431520 , n431519 );
xor ( n86220 , n86202 , n431520 );
buf ( n431522 , n86220 );
xor ( n86222 , n86162 , n431522 );
xor ( n86223 , n430957 , n430982 );
and ( n86224 , n86223 , n430989 );
and ( n86225 , n430957 , n430982 );
or ( n86226 , n86224 , n86225 );
buf ( n431528 , n86226 );
buf ( n431529 , n431528 );
buf ( n431530 , n45954 );
not ( n86230 , n431530 );
buf ( n431532 , n393369 );
not ( n86232 , n431532 );
buf ( n431534 , n50317 );
not ( n86234 , n431534 );
or ( n86235 , n86232 , n86234 );
buf ( n431537 , n40818 );
buf ( n431538 , n393381 );
nand ( n86238 , n431537 , n431538 );
buf ( n431540 , n86238 );
buf ( n431541 , n431540 );
nand ( n86241 , n86235 , n431541 );
buf ( n431543 , n86241 );
buf ( n431544 , n431543 );
not ( n86244 , n431544 );
or ( n86245 , n86230 , n86244 );
buf ( n431547 , n430971 );
buf ( n431548 , n45949 );
nand ( n86248 , n431547 , n431548 );
buf ( n431550 , n86248 );
buf ( n431551 , n431550 );
nand ( n86251 , n86245 , n431551 );
buf ( n431553 , n86251 );
not ( n86253 , n431553 );
buf ( n431555 , n430949 );
not ( n86255 , n431555 );
buf ( n431557 , n43240 );
not ( n86257 , n431557 );
or ( n86258 , n86255 , n86257 );
buf ( n431560 , n55543 );
buf ( n431561 , n385488 );
and ( n86261 , n431560 , n431561 );
not ( n86262 , n431560 );
buf ( n431564 , n385473 );
and ( n86264 , n86262 , n431564 );
nor ( n86265 , n86261 , n86264 );
buf ( n431567 , n86265 );
buf ( n431568 , n431567 );
not ( n86268 , n431568 );
buf ( n431570 , n41447 );
nand ( n86270 , n86268 , n431570 );
buf ( n431572 , n86270 );
buf ( n431573 , n431572 );
nand ( n86273 , n86258 , n431573 );
buf ( n431575 , n86273 );
not ( n86275 , n431575 );
not ( n86276 , n86275 );
or ( n86277 , n86253 , n86276 );
not ( n86278 , n431553 );
nand ( n86279 , n86278 , n431575 );
nand ( n86280 , n86277 , n86279 );
buf ( n431582 , n43058 );
buf ( n431583 , n431297 );
not ( n86283 , n431583 );
buf ( n431585 , n86283 );
buf ( n431586 , n431585 );
or ( n86286 , n431582 , n431586 );
buf ( n431588 , n400033 );
buf ( n431589 , n388897 );
and ( n86289 , n431588 , n431589 );
not ( n86290 , n431588 );
buf ( n431592 , n393562 );
and ( n86292 , n86290 , n431592 );
nor ( n86293 , n86289 , n86292 );
buf ( n431595 , n86293 );
buf ( n431596 , n431595 );
buf ( n431597 , n398665 );
or ( n86297 , n431596 , n431597 );
nand ( n86298 , n86286 , n86297 );
buf ( n431600 , n86298 );
buf ( n86300 , n431600 );
and ( n86301 , n86280 , n86300 );
not ( n86302 , n86280 );
not ( n86303 , n86300 );
and ( n86304 , n86302 , n86303 );
nor ( n86305 , n86301 , n86304 );
buf ( n431607 , n86305 );
xor ( n86307 , n431529 , n431607 );
buf ( n431609 , C0 );
buf ( n431610 , n431609 );
xor ( n86333 , n86307 , n431610 );
buf ( n431612 , n86333 );
buf ( n431613 , n431612 );
not ( n86336 , n383904 );
nor ( n86337 , n86336 , n402819 );
xor ( n86338 , n431328 , n431334 );
and ( n86339 , n86338 , n431367 );
and ( n86340 , n431328 , n431334 );
or ( n86341 , n86339 , n86340 );
buf ( n431620 , n86341 );
xor ( n86343 , n86337 , n431620 );
buf ( n431622 , n431234 );
not ( n86345 , n431622 );
buf ( n431624 , n390429 );
not ( n86347 , n431624 );
or ( n86348 , n86345 , n86347 );
buf ( n431627 , n416220 );
buf ( n431628 , n400143 );
nand ( n86351 , n431627 , n431628 );
buf ( n431630 , n86351 );
buf ( n431631 , n431630 );
nand ( n86354 , n86348 , n431631 );
buf ( n431633 , n86354 );
buf ( n431634 , n431633 );
xor ( n86357 , n417237 , n417254 );
xor ( n86358 , n86357 , n417273 );
buf ( n431637 , n86358 );
buf ( n431638 , n431637 );
xor ( n86361 , n431634 , n431638 );
xor ( n86362 , n431340 , n431350 );
and ( n86363 , n86362 , n431364 );
and ( n86364 , n431340 , n431350 );
or ( n86365 , n86363 , n86364 );
buf ( n431644 , n86365 );
buf ( n431645 , n431644 );
xor ( n86368 , n86361 , n431645 );
buf ( n431647 , n86368 );
xor ( n86370 , n86343 , n431647 );
buf ( n431649 , n86370 );
buf ( n431650 , C0 );
buf ( n431651 , n431650 );
xor ( n86384 , n431649 , n431651 );
buf ( n431653 , n85985 );
not ( n86386 , n431653 );
buf ( n431655 , n431395 );
not ( n86388 , n431655 );
or ( n86389 , n86386 , n86388 );
buf ( n431658 , n85985 );
not ( n86391 , n431658 );
buf ( n431660 , n86391 );
buf ( n431661 , n431660 );
not ( n86394 , n431661 );
buf ( n431663 , n431398 );
not ( n86396 , n431663 );
or ( n86397 , n86394 , n86396 );
buf ( n431666 , n431369 );
nand ( n431667 , n86397 , n431666 );
buf ( n431668 , n431667 );
buf ( n431669 , n431668 );
nand ( n86402 , n86389 , n431669 );
buf ( n431671 , n86402 );
buf ( n431672 , n431671 );
xor ( n86405 , n86384 , n431672 );
buf ( n431674 , n86405 );
buf ( n431675 , n431674 );
xor ( n86408 , n431613 , n431675 );
not ( n86409 , n395349 );
not ( n86410 , n431385 );
or ( n86411 , n86409 , n86410 );
buf ( n431680 , n47863 );
not ( n86413 , n431680 );
buf ( n431682 , n40759 );
not ( n86415 , n431682 );
or ( n86416 , n86413 , n86415 );
buf ( n431685 , n40758 );
buf ( n431686 , n419385 );
nand ( n86419 , n431685 , n431686 );
buf ( n431688 , n86419 );
buf ( n431689 , n431688 );
nand ( n86422 , n86416 , n431689 );
buf ( n431691 , n86422 );
buf ( n431692 , n431691 );
buf ( n431693 , n395362 );
nand ( n86426 , n431692 , n431693 );
buf ( n431695 , n86426 );
nand ( n86428 , n86411 , n431695 );
not ( n86429 , n85744 );
not ( n86430 , n431102 );
or ( n86431 , n86429 , n86430 );
not ( n86432 , n85773 );
not ( n86433 , n85770 );
or ( n86434 , n86432 , n86433 );
nand ( n86435 , n86434 , n431066 );
nand ( n86436 , n86431 , n86435 );
xor ( n86437 , n86428 , n86436 );
not ( n86438 , n85920 );
not ( n86439 , n85851 );
or ( n86440 , n86438 , n86439 );
nand ( n86441 , n86440 , n85912 );
xor ( n86442 , n86437 , n86441 );
not ( n86443 , n431136 );
nand ( n86444 , n86443 , n431159 );
not ( n86445 , n86444 );
not ( n86446 , n85927 );
or ( n86447 , n86445 , n86446 );
buf ( n431716 , n431162 );
buf ( n431717 , n431136 );
nand ( n86450 , n431716 , n431717 );
buf ( n431719 , n86450 );
nand ( n86452 , n86447 , n431719 );
xor ( n86453 , n86442 , n86452 );
buf ( n431722 , n431095 );
not ( n86455 , n431722 );
buf ( n431724 , n396622 );
not ( n86457 , n431724 );
or ( n86458 , n86455 , n86457 );
buf ( n431727 , n394210 );
not ( n86460 , n431727 );
buf ( n431729 , n398298 );
not ( n86462 , n431729 );
or ( n86463 , n86460 , n86462 );
buf ( n431732 , n399167 );
buf ( n431733 , n394207 );
nand ( n86466 , n431732 , n431733 );
buf ( n431735 , n86466 );
buf ( n431736 , n431735 );
nand ( n86469 , n86463 , n431736 );
buf ( n431738 , n86469 );
buf ( n431739 , n431738 );
buf ( n431740 , n46921 );
nand ( n86473 , n431739 , n431740 );
buf ( n431742 , n86473 );
buf ( n431743 , n431742 );
nand ( n86476 , n86458 , n431743 );
buf ( n431745 , n86476 );
not ( n86478 , n38961 );
not ( n86479 , n431179 );
or ( n86480 , n86478 , n86479 );
buf ( n431749 , n416646 );
buf ( n431750 , n395469 );
nand ( n86483 , n431749 , n431750 );
buf ( n431752 , n86483 );
nand ( n86485 , n86480 , n431752 );
xor ( n86486 , n431745 , n86485 );
buf ( n431755 , n413643 );
not ( n86488 , n431755 );
buf ( n431757 , n64136 );
not ( n86490 , n431757 );
buf ( n431759 , n388367 );
not ( n86492 , n431759 );
or ( n86493 , n86490 , n86492 );
buf ( n431762 , n393557 );
buf ( n431763 , n44776 );
nand ( n86496 , n431762 , n431763 );
buf ( n431765 , n86496 );
buf ( n431766 , n431765 );
nand ( n86499 , n86493 , n431766 );
buf ( n431768 , n86499 );
buf ( n431769 , n431768 );
not ( n86502 , n431769 );
or ( n86503 , n86488 , n86502 );
buf ( n431772 , n431056 );
buf ( n431773 , n45260 );
nand ( n86506 , n431772 , n431773 );
buf ( n431775 , n86506 );
buf ( n431776 , n431775 );
nand ( n86509 , n86503 , n431776 );
buf ( n431778 , n86509 );
xor ( n86511 , n86486 , n431778 );
buf ( n431780 , n43515 );
not ( n86513 , n431780 );
buf ( n431782 , n416692 );
not ( n86515 , n431782 );
or ( n86516 , n86513 , n86515 );
buf ( n431785 , n431317 );
buf ( n431786 , n43536 );
nand ( n86519 , n431785 , n431786 );
buf ( n431788 , n86519 );
buf ( n431789 , n431788 );
nand ( n86522 , n86516 , n431789 );
buf ( n431791 , n86522 );
buf ( n431792 , n431791 );
xor ( n86525 , n417300 , n417325 );
xor ( n86526 , n86525 , n417398 );
buf ( n431795 , n86526 );
buf ( n431796 , n431795 );
xor ( n86529 , n431792 , n431796 );
xor ( n86530 , n431212 , n431216 );
and ( n86531 , n86530 , n431242 );
and ( n86532 , n431212 , n431216 );
or ( n86533 , n86531 , n86532 );
buf ( n431802 , n86533 );
buf ( n431803 , n431802 );
xor ( n86536 , n86529 , n431803 );
buf ( n431805 , n86536 );
xor ( n86538 , n86511 , n431805 );
not ( n86539 , n61577 );
not ( n86540 , n47891 );
not ( n86541 , n38631 );
or ( n86542 , n86540 , n86541 );
buf ( n431811 , n386179 );
not ( n86544 , n431811 );
buf ( n431813 , n61299 );
nand ( n86546 , n86544 , n431813 );
buf ( n431815 , n86546 );
nand ( n86548 , n86542 , n431815 );
not ( n86549 , n86548 );
or ( n86550 , n86539 , n86549 );
nand ( n86551 , n431149 , n50579 );
nand ( n86552 , n86550 , n86551 );
and ( n86553 , n86538 , n86552 );
not ( n86554 , n86538 );
not ( n86555 , n86552 );
and ( n86556 , n86554 , n86555 );
nor ( n86557 , n86553 , n86556 );
xor ( n86558 , n86453 , n86557 );
buf ( n431827 , n86558 );
xor ( n86560 , n86408 , n431827 );
buf ( n431829 , n86560 );
xor ( n86562 , n86222 , n431829 );
buf ( n431831 , n86562 );
xor ( n86564 , n86153 , n431831 );
buf ( n431833 , n86564 );
buf ( n431834 , n431833 );
xor ( n86567 , n430935 , n431006 );
xnor ( n86568 , n86567 , n431016 );
buf ( n431837 , n86568 );
xor ( n86570 , n423199 , n423205 );
and ( n86571 , n86570 , n423393 );
and ( n86572 , n423199 , n423205 );
or ( n86573 , n86571 , n86572 );
buf ( n431842 , n86573 );
buf ( n431843 , n431842 );
xor ( n86576 , n431837 , n431843 );
xor ( n86577 , n86122 , n431452 );
xnor ( n86578 , n86577 , n431458 );
buf ( n431847 , n86578 );
and ( n86580 , n86576 , n431847 );
and ( n86581 , n431837 , n431843 );
or ( n86582 , n86580 , n86581 );
buf ( n431851 , n86582 );
buf ( n431852 , n431851 );
not ( n86585 , n431852 );
buf ( n431854 , n86585 );
buf ( n431855 , n431854 );
nand ( n86588 , n431834 , n431855 );
buf ( n431857 , n86588 );
buf ( n431858 , n431857 );
not ( n86591 , n431858 );
xor ( n86592 , n431837 , n431843 );
xor ( n86593 , n86592 , n431847 );
buf ( n431862 , n86593 );
buf ( n431863 , n431862 );
buf ( n86596 , n431863 );
buf ( n431865 , n86596 );
buf ( n431866 , n431865 );
xor ( n86599 , n423171 , n423188 );
and ( n86600 , n86599 , n423396 );
and ( n86601 , n423171 , n423188 );
or ( n86602 , n86600 , n86601 );
buf ( n431871 , n86602 );
buf ( n431872 , n431871 );
nor ( n86605 , n431866 , n431872 );
buf ( n431874 , n86605 );
buf ( n431875 , n431874 );
nor ( n86608 , n86591 , n431875 );
buf ( n431877 , n86608 );
buf ( n431878 , n431877 );
buf ( n431879 , n413643 );
not ( n86612 , n431879 );
buf ( n431881 , n417422 );
not ( n86614 , n431881 );
or ( n86615 , n86612 , n86614 );
buf ( n431884 , n431768 );
buf ( n431885 , n45260 );
nand ( n86618 , n431884 , n431885 );
buf ( n431887 , n86618 );
buf ( n431888 , n431887 );
nand ( n86621 , n86615 , n431888 );
buf ( n431890 , n86621 );
not ( n86623 , n431890 );
xor ( n86624 , n431634 , n431638 );
and ( n86625 , n86624 , n431645 );
and ( n86626 , n431634 , n431638 );
or ( n86627 , n86625 , n86626 );
buf ( n431896 , n86627 );
not ( n86629 , n431896 );
not ( n86630 , n86629 );
or ( n86631 , n86623 , n86630 );
not ( n86632 , n431890 );
nand ( n86633 , n431896 , n86632 );
nand ( n86634 , n86631 , n86633 );
xor ( n86635 , n417278 , n417295 );
xor ( n86636 , n86635 , n417403 );
buf ( n431905 , n86636 );
and ( n86638 , n86634 , n431905 );
not ( n86639 , n86634 );
not ( n86640 , n431905 );
and ( n86641 , n86639 , n86640 );
nor ( n86642 , n86638 , n86641 );
buf ( n431911 , n86642 );
xor ( n86644 , n86428 , n86436 );
and ( n86645 , n86644 , n86441 );
and ( n86646 , n86428 , n86436 );
or ( n86647 , n86645 , n86646 );
buf ( n431916 , n86647 );
xor ( n86649 , n431911 , n431916 );
or ( n86650 , n86511 , n431805 );
not ( n86651 , n86650 );
not ( n86652 , n86552 );
or ( n86653 , n86651 , n86652 );
nand ( n86654 , n86511 , n431805 );
nand ( n86655 , n86653 , n86654 );
buf ( n431924 , n86655 );
xor ( n86657 , n86649 , n431924 );
buf ( n431926 , n86657 );
buf ( n431927 , n431926 );
buf ( n431928 , n43058 );
not ( n86661 , n431928 );
buf ( n431930 , n431595 );
not ( n86663 , n431930 );
and ( n86664 , n86661 , n86663 );
buf ( n431933 , n417445 );
buf ( n431934 , n37315 );
nor ( n86667 , n431933 , n431934 );
buf ( n431936 , n86667 );
buf ( n431937 , n431936 );
nor ( n86670 , n86664 , n431937 );
buf ( n431939 , n86670 );
not ( n86672 , n431939 );
not ( n86673 , n44077 );
not ( n86674 , n431567 );
and ( n86675 , n86673 , n86674 );
and ( n86676 , n416560 , n49166 );
nor ( n86677 , n86675 , n86676 );
not ( n86678 , n86677 );
xor ( n86679 , n431792 , n431796 );
and ( n86680 , n86679 , n431803 );
and ( n86681 , n431792 , n431796 );
or ( n86682 , n86680 , n86681 );
buf ( n431951 , n86682 );
xnor ( n86684 , n86678 , n431951 );
not ( n86685 , n86684 );
or ( n86686 , n86672 , n86685 );
or ( n86687 , n86684 , n431939 );
nand ( n86688 , n86686 , n86687 );
buf ( n431957 , n86688 );
buf ( n431958 , C1 );
buf ( n431959 , n431958 );
xor ( n86714 , n431957 , n431959 );
xor ( n86715 , n431745 , n86485 );
and ( n86716 , n86715 , n431778 );
and ( n86717 , n431745 , n86485 );
or ( n86718 , n86716 , n86717 );
and ( n86719 , n45949 , n431543 );
and ( n86720 , n27195 , n393384 );
not ( n86721 , n27195 );
and ( n86722 , n86721 , n393369 );
or ( n86723 , n86720 , n86722 );
and ( n86724 , n86723 , n45954 );
nor ( n86725 , n86719 , n86724 );
buf ( n431972 , n86725 );
not ( n86727 , n431972 );
buf ( n431974 , n86727 );
xor ( n86729 , n86718 , n431974 );
not ( n86730 , n395362 );
not ( n86731 , n70093 );
or ( n86732 , n86730 , n86731 );
buf ( n431979 , n431691 );
not ( n86734 , n431979 );
buf ( n431981 , n395352 );
nor ( n86736 , n86734 , n431981 );
buf ( n431983 , n86736 );
not ( n86738 , n431983 );
nand ( n86739 , n86732 , n86738 );
xnor ( n86740 , n86729 , n86739 );
buf ( n431987 , n86740 );
xor ( n86742 , n86714 , n431987 );
buf ( n431989 , n86742 );
buf ( n431990 , n431989 );
xor ( n86745 , n431927 , n431990 );
xor ( n86746 , n431492 , n431507 );
and ( n86747 , n86746 , n431520 );
and ( n86748 , n431492 , n431507 );
or ( n86749 , n86747 , n86748 );
buf ( n431996 , n86749 );
buf ( n431997 , n431996 );
xnor ( n86752 , n86745 , n431997 );
buf ( n431999 , n86752 );
buf ( n432000 , n431999 );
buf ( n432001 , n431522 );
not ( n86756 , n432001 );
buf ( n432003 , n86162 );
nand ( n86758 , n86756 , n432003 );
buf ( n432005 , n86758 );
buf ( n432006 , n432005 );
not ( n86761 , n432006 );
buf ( n432008 , n431829 );
not ( n86763 , n432008 );
or ( n86764 , n86761 , n86763 );
buf ( n432011 , n86162 );
not ( n86766 , n432011 );
buf ( n432013 , n431522 );
nand ( n86768 , n86766 , n432013 );
buf ( n432015 , n86768 );
buf ( n432016 , n432015 );
nand ( n86771 , n86764 , n432016 );
buf ( n432018 , n86771 );
buf ( n432019 , n432018 );
xor ( n86774 , n432000 , n432019 );
xor ( n86775 , n68388 , n68368 );
xnor ( n86776 , n86775 , n68414 );
buf ( n432023 , n86776 );
buf ( n432024 , n431738 );
not ( n86779 , n432024 );
buf ( n432026 , n389122 );
not ( n86781 , n432026 );
or ( n86782 , n86779 , n86781 );
buf ( n432029 , n416190 );
buf ( n432030 , n41563 );
nand ( n86785 , n432029 , n432030 );
buf ( n432032 , n86785 );
buf ( n432033 , n432032 );
nand ( n86788 , n86782 , n432033 );
buf ( n432035 , n86788 );
buf ( n432036 , n432035 );
xor ( n86791 , n432023 , n432036 );
buf ( n432038 , n416322 );
buf ( n432039 , n416252 );
xor ( n86794 , n432038 , n432039 );
buf ( n432041 , n416232 );
xnor ( n86796 , n86794 , n432041 );
buf ( n432043 , n86796 );
buf ( n432044 , n432043 );
xor ( n86799 , n86791 , n432044 );
buf ( n432046 , n86799 );
buf ( n432047 , n432046 );
buf ( n432048 , n416661 );
not ( n86803 , n432048 );
buf ( n432050 , n416699 );
not ( n86805 , n432050 );
or ( n86806 , n86803 , n86805 );
buf ( n432053 , n416699 );
buf ( n432054 , n416661 );
or ( n86809 , n432053 , n432054 );
nand ( n86810 , n86806 , n86809 );
buf ( n432057 , n86810 );
xnor ( n86812 , n70040 , n432057 );
buf ( n432059 , n86812 );
xor ( n86814 , n432047 , n432059 );
buf ( n432061 , n50357 );
buf ( n432062 , n402819 );
buf ( n432063 , n40791 );
and ( n86818 , n432062 , n432063 );
not ( n86819 , n432062 );
buf ( n432066 , n391764 );
and ( n86821 , n86819 , n432066 );
nor ( n86822 , n86818 , n86821 );
buf ( n432069 , n86822 );
buf ( n432070 , n432069 );
or ( n86825 , n432061 , n432070 );
buf ( n432072 , n55054 );
buf ( n432073 , n389928 );
and ( n86828 , n432072 , n432073 );
not ( n86829 , n432072 );
buf ( n432076 , n388266 );
and ( n86831 , n86829 , n432076 );
nor ( n86832 , n86828 , n86831 );
buf ( n432079 , n86832 );
buf ( n432080 , n432079 );
buf ( n432081 , n383910 );
or ( n86836 , n432080 , n432081 );
nand ( n86837 , n86825 , n86836 );
buf ( n432084 , n86837 );
buf ( n432085 , n432084 );
xor ( n86840 , n86814 , n432085 );
buf ( n432087 , n86840 );
buf ( n432088 , n432087 );
buf ( n432089 , C0 );
buf ( n432090 , n432089 );
xor ( n86863 , n432088 , n432090 );
and ( n86866 , n431529 , n431607 );
or ( n86867 , C0 , n86866 );
buf ( n432094 , n86867 );
buf ( n432095 , n432094 );
xor ( n86870 , n86863 , n432095 );
buf ( n432097 , n86870 );
buf ( n432098 , n432097 );
not ( n86873 , n86337 );
not ( n86874 , n431647 );
or ( n86875 , n86873 , n86874 );
nor ( n86876 , n86337 , n431647 );
not ( n86877 , n431620 );
or ( n86878 , n86876 , n86877 );
nand ( n86879 , n86875 , n86878 );
nand ( n86880 , n86275 , n86278 );
not ( n86881 , n86880 );
not ( n86882 , n86300 );
or ( n86883 , n86881 , n86882 );
nand ( n86884 , n431553 , n431575 );
nand ( n86885 , n86883 , n86884 );
xor ( n86886 , n86879 , n86885 );
not ( n86887 , n61577 );
buf ( n432114 , n47891 );
not ( n86889 , n432114 );
buf ( n432116 , n385345 );
not ( n86891 , n432116 );
or ( n86892 , n86889 , n86891 );
not ( n86893 , n44007 );
nand ( n86894 , n86893 , n61299 );
buf ( n432121 , n86894 );
nand ( n86896 , n86892 , n432121 );
buf ( n432123 , n86896 );
not ( n86898 , n432123 );
or ( n86899 , n86887 , n86898 );
nand ( n86900 , n86548 , n50579 );
nand ( n86901 , n86899 , n86900 );
xor ( n86902 , n86886 , n86901 );
buf ( n432129 , n86902 );
xor ( n86904 , n431649 , n431651 );
and ( n86905 , n86904 , n431672 );
or ( n86907 , n86905 , C0 );
buf ( n432133 , n86907 );
buf ( n432134 , n432133 );
xor ( n86910 , n432129 , n432134 );
xor ( n86911 , n86442 , n86452 );
and ( n86912 , n86911 , n86557 );
and ( n86913 , n86442 , n86452 );
or ( n86914 , n86912 , n86913 );
buf ( n432140 , n86914 );
xor ( n86916 , n86910 , n432140 );
buf ( n432142 , n86916 );
buf ( n432143 , n432142 );
xor ( n86919 , n432098 , n432143 );
xor ( n86920 , n431613 , n431675 );
and ( n86921 , n86920 , n431827 );
and ( n86922 , n431613 , n431675 );
or ( n86923 , n86921 , n86922 );
buf ( n432149 , n86923 );
buf ( n432150 , n432149 );
xor ( n86926 , n86919 , n432150 );
buf ( n432152 , n86926 );
buf ( n432153 , n432152 );
xnor ( n86929 , n86774 , n432153 );
buf ( n432155 , n86929 );
buf ( n432156 , n432155 );
xor ( n86932 , n431028 , n431463 );
and ( n86933 , n86932 , n431831 );
and ( n86934 , n431028 , n431463 );
or ( n86935 , n86933 , n86934 );
buf ( n432161 , n86935 );
buf ( n432162 , n432161 );
nand ( n86938 , n432156 , n432162 );
buf ( n432164 , n86938 );
buf ( n432165 , n432164 );
and ( n86941 , n431878 , n432165 );
buf ( n432167 , n86941 );
buf ( n432168 , n432167 );
not ( n86944 , n432168 );
or ( n86945 , n85567 , n86944 );
not ( n86946 , n431857 );
and ( n86947 , n431862 , n431871 );
not ( n86948 , n86947 );
or ( n86949 , n86946 , n86948 );
buf ( n432175 , n431833 );
buf ( n432176 , n431854 );
or ( n86952 , n432175 , n432176 );
buf ( n432178 , n86952 );
nand ( n86954 , n86949 , n432178 );
not ( n86955 , n86954 );
not ( n86956 , n432164 );
or ( n86957 , n86955 , n86956 );
buf ( n432183 , n432155 );
buf ( n432184 , n432161 );
or ( n86960 , n432183 , n432184 );
buf ( n432186 , n86960 );
nand ( n86962 , n86957 , n432186 );
buf ( n432188 , n86962 );
not ( n86964 , n432188 );
buf ( n432190 , n86964 );
buf ( n432191 , n432190 );
nand ( n86967 , n86945 , n432191 );
buf ( n432193 , n86967 );
buf ( n432194 , n432193 );
buf ( n432195 , n416202 );
buf ( n432196 , n416177 );
xor ( n86972 , n432195 , n432196 );
buf ( n432198 , n416333 );
xnor ( n86974 , n86972 , n432198 );
buf ( n432200 , n86974 );
buf ( n432201 , n432200 );
nand ( n86977 , n86629 , n86632 );
not ( n86978 , n86977 );
not ( n86979 , n431905 );
or ( n86980 , n86978 , n86979 );
nand ( n86981 , n431896 , n431890 );
nand ( n86982 , n86980 , n86981 );
buf ( n432208 , n86982 );
xor ( n86984 , n432201 , n432208 );
buf ( n432210 , n86678 );
not ( n86986 , n432210 );
buf ( n432212 , n431939 );
not ( n86988 , n432212 );
buf ( n432214 , n86988 );
buf ( n432215 , n432214 );
not ( n86991 , n432215 );
or ( n86992 , n86986 , n86991 );
buf ( n432218 , n86677 );
not ( n86994 , n432218 );
buf ( n432220 , n431939 );
not ( n86996 , n432220 );
or ( n86997 , n86994 , n86996 );
buf ( n432223 , n431951 );
nand ( n86999 , n86997 , n432223 );
buf ( n432225 , n86999 );
buf ( n432226 , n432225 );
nand ( n87002 , n86992 , n432226 );
buf ( n432228 , n87002 );
buf ( n432229 , n432228 );
and ( n87005 , n86984 , n432229 );
and ( n87006 , n432201 , n432208 );
or ( n87007 , n87005 , n87006 );
buf ( n432233 , n87007 );
buf ( n432234 , n432233 );
not ( n87010 , n70093 );
not ( n87011 , n395362 );
or ( n87012 , n87010 , n87011 );
not ( n87013 , n86725 );
nor ( n87014 , n87013 , n431983 );
nand ( n87015 , n87012 , n87014 );
not ( n87016 , n87015 );
not ( n87017 , n86718 );
or ( n87018 , n87016 , n87017 );
nand ( n87019 , n431974 , n86739 );
nand ( n87020 , n87018 , n87019 );
buf ( n432246 , n87020 );
buf ( n432247 , C0 );
buf ( n432248 , n432247 );
or ( n87047 , n432246 , n432248 );
xor ( n87048 , n432047 , n432059 );
and ( n87049 , n87048 , n432085 );
and ( n87050 , n432047 , n432059 );
or ( n87051 , n87049 , n87050 );
buf ( n432254 , n87051 );
buf ( n432255 , n432254 );
nand ( n87054 , n87047 , n432255 );
buf ( n432257 , n87054 );
buf ( n432258 , n432257 );
buf ( n432259 , C1 );
buf ( n432260 , n432259 );
and ( n87062 , n432258 , n432260 );
buf ( n432262 , n87062 );
buf ( n432263 , n432262 );
not ( n87065 , n432263 );
buf ( n432265 , n87065 );
buf ( n432266 , n432265 );
xor ( n87068 , n432234 , n432266 );
buf ( n432268 , n416632 );
buf ( n432269 , n417460 );
xor ( n87071 , n432268 , n432269 );
buf ( n432271 , n416737 );
xnor ( n87073 , n87071 , n432271 );
buf ( n432273 , n87073 );
buf ( n432274 , n432273 );
not ( n87076 , n432274 );
buf ( n432276 , n87076 );
buf ( n432277 , n432276 );
xnor ( n87079 , n87068 , n432277 );
buf ( n432279 , n87079 );
buf ( n432280 , n432279 );
not ( n87082 , n432280 );
buf ( n432282 , n87082 );
buf ( n432283 , n432282 );
not ( n87085 , n432283 );
buf ( n432285 , n415928 );
buf ( n432286 , n415959 );
xor ( n87088 , n432285 , n432286 );
buf ( n432288 , n416012 );
xnor ( n87090 , n87088 , n432288 );
buf ( n432290 , n87090 );
buf ( n432291 , n432290 );
not ( n87093 , n432291 );
buf ( n432293 , n87093 );
buf ( n432294 , n432293 );
not ( n87096 , n432294 );
buf ( n432296 , n69726 );
buf ( n432297 , n61577 );
and ( n87099 , n432296 , n432297 );
buf ( n432299 , n47891 );
not ( n87101 , n432299 );
buf ( n432301 , n41904 );
not ( n87103 , n432301 );
or ( n87104 , n87101 , n87103 );
buf ( n432304 , n388952 );
buf ( n432305 , n61299 );
nand ( n87107 , n432304 , n432305 );
buf ( n432307 , n87107 );
buf ( n432308 , n432307 );
nand ( n87110 , n87104 , n432308 );
buf ( n432310 , n87110 );
buf ( n432311 , n432310 );
not ( n87113 , n432311 );
buf ( n432313 , n50580 );
nor ( n87115 , n87113 , n432313 );
buf ( n432315 , n87115 );
buf ( n432316 , n432315 );
nor ( n87118 , n87099 , n432316 );
buf ( n432318 , n87118 );
buf ( n432319 , n432318 );
not ( n87121 , n432319 );
or ( n87122 , n87096 , n87121 );
buf ( n432322 , n432318 );
not ( n87124 , n432322 );
buf ( n432324 , n87124 );
buf ( n432325 , n432324 );
buf ( n432326 , n432290 );
nand ( n87128 , n432325 , n432326 );
buf ( n432328 , n87128 );
buf ( n432329 , n432328 );
nand ( n87131 , n87122 , n432329 );
buf ( n432331 , n87131 );
xor ( n87133 , n416336 , n416361 );
xor ( n87134 , n87133 , n416387 );
buf ( n432334 , n87134 );
xor ( n87136 , n432331 , n432334 );
buf ( n432336 , n87136 );
buf ( n432337 , C0 );
xor ( n87150 , n432023 , n432036 );
and ( n87151 , n87150 , n432044 );
and ( n87152 , n432023 , n432036 );
or ( n87153 , n87151 , n87152 );
buf ( n432342 , n87153 );
buf ( n432343 , n432342 );
buf ( n432344 , n45949 );
not ( n87157 , n432344 );
buf ( n432346 , n86723 );
not ( n87159 , n432346 );
or ( n87160 , n87157 , n87159 );
buf ( n432349 , n416118 );
not ( n87162 , n432349 );
buf ( n432351 , n45954 );
nand ( n87164 , n87162 , n432351 );
buf ( n432353 , n87164 );
buf ( n432354 , n432353 );
nand ( n87167 , n87160 , n432354 );
buf ( n432356 , n87167 );
buf ( n432357 , n432356 );
xor ( n87170 , n432343 , n432357 );
buf ( n432359 , n432079 );
not ( n87172 , n432359 );
buf ( n432361 , n87172 );
buf ( n432362 , n432361 );
not ( n87175 , n432362 );
buf ( n432364 , n383894 );
not ( n87177 , n432364 );
or ( n87178 , n87175 , n87177 );
buf ( n432367 , n416374 );
buf ( n432368 , n383907 );
nand ( n87181 , n432367 , n432368 );
buf ( n432370 , n87181 );
buf ( n432371 , n432370 );
nand ( n87184 , n87178 , n432371 );
buf ( n432373 , n87184 );
buf ( n432374 , n432373 );
and ( n87187 , n87170 , n432374 );
and ( n87188 , n432343 , n432357 );
or ( n87189 , n87187 , n87188 );
buf ( n432378 , n87189 );
xor ( n87191 , n432337 , n432378 );
not ( n87192 , n416151 );
not ( n87193 , n69432 );
or ( n87194 , n87192 , n87193 );
nand ( n87195 , n69456 , n416127 );
nand ( n87196 , n87194 , n87195 );
not ( n87197 , n416109 );
and ( n87198 , n87196 , n87197 );
not ( n87199 , n87196 );
and ( n87200 , n87199 , n416109 );
nor ( n87201 , n87198 , n87200 );
not ( n87202 , n87201 );
xor ( n87203 , n87191 , n87202 );
buf ( n432392 , n87203 );
xor ( n87205 , n432336 , n432392 );
xor ( n87206 , n416712 , n416719 );
xor ( n87207 , n87206 , n416733 );
buf ( n432396 , n87207 );
buf ( n432397 , C0 );
buf ( n432398 , n432397 );
buf ( n432399 , n432396 );
or ( n87237 , n432398 , n432399 );
xor ( n87238 , n432343 , n432357 );
xor ( n87239 , n87238 , n432374 );
buf ( n432403 , n87239 );
buf ( n432404 , n432403 );
nand ( n87242 , n87237 , n432404 );
buf ( n432406 , n87242 );
buf ( n432407 , n432406 );
nand ( n87245 , C1 , n432407 );
buf ( n432409 , n87245 );
buf ( n432410 , n432409 );
xor ( n87248 , n87205 , n432410 );
buf ( n432412 , n87248 );
buf ( n432413 , n432412 );
not ( n87251 , n432413 );
or ( n87252 , n87085 , n87251 );
buf ( n432416 , n432412 );
buf ( n432417 , n432282 );
or ( n87255 , n432416 , n432417 );
buf ( n432419 , n432403 );
buf ( n432420 , n432396 );
xor ( n87258 , n432419 , n432420 );
xor ( n87261 , n87258 , C1 );
buf ( n432423 , n87261 );
buf ( n432424 , n432423 );
not ( n87264 , n432424 );
buf ( n432426 , n87264 );
not ( n87266 , n432426 );
xor ( n87267 , n432088 , n432090 );
and ( n87268 , n87267 , n432095 );
or ( n87270 , n87268 , C0 );
buf ( n432431 , n87270 );
not ( n87272 , n432431 );
or ( n87273 , n87266 , n87272 );
buf ( n432434 , n432431 );
not ( n87275 , n432434 );
buf ( n432436 , n87275 );
not ( n87277 , n432436 );
not ( n87278 , n432423 );
or ( n87279 , n87277 , n87278 );
not ( n87280 , n86885 );
not ( n87281 , n86901 );
or ( n87282 , n87280 , n87281 );
or ( n87283 , n86901 , n86885 );
nand ( n87284 , n87283 , n86879 );
nand ( n87285 , n87282 , n87284 );
buf ( n432446 , n87285 );
xor ( n87287 , n432201 , n432208 );
xor ( n87288 , n87287 , n432229 );
buf ( n432449 , n87288 );
buf ( n432450 , n432449 );
xor ( n87291 , n432446 , n432450 );
buf ( n432452 , n87291 );
buf ( n432453 , n432452 );
buf ( n432454 , n416547 );
not ( n87295 , n432454 );
not ( n87296 , n416572 );
not ( n87297 , n68419 );
not ( n87298 , n69922 );
or ( n87299 , n87297 , n87298 );
or ( n87300 , n68419 , n69928 );
nand ( n87301 , n87299 , n87300 );
not ( n87302 , n87301 );
or ( n87303 , n87296 , n87302 );
or ( n87304 , n416572 , n69930 );
nand ( n87305 , n87303 , n87304 );
buf ( n432466 , n87305 );
not ( n87307 , n432466 );
or ( n87308 , n87295 , n87307 );
buf ( n432469 , n87305 );
buf ( n432470 , n416547 );
or ( n87311 , n432469 , n432470 );
nand ( n87312 , n87308 , n87311 );
buf ( n432473 , n87312 );
buf ( n432474 , n432473 );
buf ( n432475 , n50579 );
not ( n87316 , n432475 );
buf ( n432477 , n432123 );
not ( n87318 , n432477 );
or ( n87319 , n87316 , n87318 );
buf ( n432480 , n432310 );
buf ( n432481 , n61577 );
nand ( n87322 , n432480 , n432481 );
buf ( n432483 , n87322 );
buf ( n432484 , n432483 );
nand ( n87325 , n87319 , n432484 );
buf ( n432486 , n87325 );
buf ( n432487 , n432486 );
xor ( n87328 , n432474 , n432487 );
xor ( n87329 , n417408 , n417433 );
xor ( n87330 , n87329 , n417456 );
buf ( n432491 , n87330 );
buf ( n432492 , n432491 );
xor ( n87333 , n87328 , n432492 );
buf ( n432494 , n87333 );
buf ( n432495 , n432494 );
and ( n87336 , n432453 , n432495 );
not ( n87337 , n432453 );
buf ( n432498 , n432494 );
not ( n87339 , n432498 );
buf ( n432500 , n87339 );
buf ( n432501 , n432500 );
and ( n87342 , n87337 , n432501 );
nor ( n87343 , n87336 , n87342 );
buf ( n432504 , n87343 );
nand ( n87345 , n87279 , n432504 );
nand ( n87346 , n87273 , n87345 );
buf ( n432507 , n87346 );
nand ( n87348 , n87255 , n432507 );
buf ( n432509 , n87348 );
buf ( n432510 , n432509 );
nand ( n87351 , n87252 , n432510 );
buf ( n432512 , n87351 );
buf ( n432513 , n432512 );
xor ( n87354 , n416624 , n416628 );
xor ( n87355 , n87354 , n417467 );
buf ( n432516 , n87355 );
buf ( n432517 , n432516 );
buf ( n432518 , n416605 );
not ( n87359 , n432518 );
buf ( n432520 , n87359 );
not ( n87364 , n432520 );
and ( n87365 , n87364 , n69844 );
nor ( n87366 , C0 , n87365 );
nand ( n87368 , C1 , n69843 );
and ( n87369 , n432520 , n87368 );
not ( n87370 , n432520 );
and ( n87371 , n87370 , C1 );
or ( n87372 , n87369 , n87371 );
nand ( n87373 , n87366 , n87372 );
buf ( n432530 , n87373 );
xor ( n87375 , n432517 , n432530 );
xor ( n87376 , n432336 , n432392 );
and ( n87377 , n87376 , n432410 );
and ( n87378 , n432336 , n432392 );
or ( n87379 , n87377 , n87378 );
buf ( n432536 , n87379 );
buf ( n432537 , n432536 );
xor ( n87382 , n87375 , n432537 );
buf ( n432539 , n87382 );
buf ( n432540 , n432539 );
and ( n87385 , n432513 , n432540 );
not ( n87386 , n432513 );
buf ( n432543 , n432539 );
not ( n87388 , n432543 );
buf ( n432545 , n87388 );
buf ( n432546 , n432545 );
and ( n87391 , n87386 , n432546 );
nor ( n87392 , n87385 , n87391 );
buf ( n432549 , n87392 );
buf ( n432550 , n432549 );
buf ( n432551 , n432293 );
not ( n87396 , n432551 );
buf ( n432553 , n432324 );
not ( n87398 , n432553 );
or ( n87399 , n87396 , n87398 );
buf ( n432556 , n432290 );
not ( n87401 , n432556 );
buf ( n432558 , n432318 );
not ( n87403 , n432558 );
or ( n87404 , n87401 , n87403 );
buf ( n432561 , n432334 );
nand ( n87406 , n87404 , n432561 );
buf ( n432563 , n87406 );
buf ( n432564 , n432563 );
nand ( n87409 , n87399 , n432564 );
buf ( n432566 , n87409 );
buf ( n432567 , n432566 );
xor ( n87412 , n69728 , n69737 );
xor ( n87413 , n87412 , n69748 );
buf ( n432570 , n87413 );
xor ( n87415 , n432567 , n432570 );
xor ( n87416 , n69461 , n416391 );
xor ( n87417 , n87416 , n416395 );
buf ( n432574 , n87417 );
xnor ( n87419 , n87415 , n432574 );
buf ( n432576 , n87419 );
buf ( n432577 , n432576 );
not ( n87422 , n432265 );
not ( n87423 , n432276 );
or ( n87424 , n87422 , n87423 );
not ( n87425 , n432273 );
not ( n87426 , n432262 );
or ( n87427 , n87425 , n87426 );
nand ( n87428 , n87427 , n432233 );
nand ( n87429 , n87424 , n87428 );
not ( n87430 , n87429 );
not ( n87431 , n87202 );
or ( n87435 , n87431 , C1 );
not ( n87437 , n87201 );
or ( n87438 , C0 , n87437 );
nand ( n87439 , n87438 , n432378 );
nand ( n87440 , n87435 , n87439 );
not ( n87441 , n87440 );
not ( n87442 , n87441 );
buf ( n432595 , n69934 );
not ( n87458 , n432595 );
buf ( n432597 , n416520 );
not ( n87460 , n432597 );
or ( n87461 , n87458 , n87460 );
buf ( n432600 , n69934 );
not ( n87463 , n432600 );
buf ( n432602 , n416517 );
nand ( n87465 , n87463 , n432602 );
buf ( n432604 , n87465 );
buf ( n432605 , n432604 );
nand ( n87468 , n87461 , n432605 );
buf ( n432607 , n87468 );
buf ( n432608 , n432607 );
buf ( n432609 , n416540 );
and ( n87472 , n432608 , n432609 );
not ( n87473 , n432608 );
buf ( n432612 , n416598 );
and ( n87475 , n87473 , n432612 );
nor ( n87476 , n87472 , n87475 );
buf ( n432615 , n87476 );
buf ( n432616 , n432615 );
not ( n87479 , n432616 );
or ( n87480 , C0 , n87479 );
xor ( n87481 , n432474 , n432487 );
and ( n87482 , n87481 , n432492 );
and ( n87483 , n432474 , n432487 );
or ( n87484 , n87482 , n87483 );
buf ( n432623 , n87484 );
buf ( n432624 , n432623 );
nand ( n87487 , n87480 , n432624 );
buf ( n432626 , n87487 );
buf ( n432627 , n432615 );
not ( n87490 , n432627 );
buf ( n432629 , n87490 );
buf ( n432630 , C1 );
nand ( n87499 , n432626 , n432630 );
not ( n87500 , n87499 );
or ( n87501 , n87442 , n87500 );
or ( n87502 , n87499 , n87441 );
nand ( n87503 , n87501 , n87502 );
not ( n87504 , n87503 );
or ( n87505 , n87430 , n87504 );
not ( n87506 , n87429 );
not ( n87507 , n87506 );
or ( n87508 , n87507 , n87503 );
nand ( n87509 , n87505 , n87508 );
buf ( n432642 , n87509 );
xor ( n87511 , n432577 , n432642 );
buf ( n432644 , n432449 );
buf ( n432645 , n87285 );
or ( n87514 , n432644 , n432645 );
buf ( n432647 , n87514 );
buf ( n432648 , n432647 );
buf ( n432649 , n432494 );
and ( n87518 , n432648 , n432649 );
and ( n87519 , n432446 , n432450 );
buf ( n432652 , n87519 );
buf ( n432653 , n432652 );
nor ( n87522 , n87518 , n432653 );
buf ( n432655 , n87522 );
buf ( n432656 , n432655 );
and ( n87525 , n432623 , C1 );
or ( n432658 , n87525 , C0 );
buf ( n432659 , n432658 );
buf ( n432660 , n432629 );
xnor ( n87531 , n432659 , n432660 );
buf ( n432662 , n87531 );
buf ( n432663 , n432662 );
xor ( n432664 , n432656 , n432663 );
and ( n87535 , n86647 , n86642 );
or ( n432666 , n86655 , n87535 );
or ( n87537 , n86647 , n86642 );
nand ( n432668 , n432666 , n87537 );
buf ( n432669 , n432668 );
xor ( n432670 , n431957 , n431959 );
and ( n87541 , n432670 , n431987 );
and ( n432672 , n431957 , n431959 );
or ( n87543 , n87541 , n432672 );
buf ( n432674 , n87543 );
buf ( n432675 , n432674 );
xor ( n432676 , n432669 , n432675 );
xor ( n87547 , n87020 , n432247 );
xnor ( n432678 , n87547 , n432254 );
buf ( n432679 , n432678 );
and ( n432680 , n432676 , n432679 );
and ( n87551 , n432669 , n432675 );
or ( n432682 , n432680 , n87551 );
buf ( n432683 , n432682 );
buf ( n432684 , n432683 );
and ( n87555 , n432664 , n432684 );
and ( n432686 , n432656 , n432663 );
or ( n87557 , n87555 , n432686 );
buf ( n432688 , n87557 );
buf ( n432689 , n432688 );
xor ( n432690 , n87511 , n432689 );
buf ( n432691 , n432690 );
buf ( n432692 , n432691 );
and ( n87563 , n432550 , n432692 );
not ( n432694 , n432550 );
buf ( n432695 , n432691 );
not ( n432696 , n432695 );
buf ( n432697 , n432696 );
buf ( n432698 , n432697 );
and ( n87569 , n432694 , n432698 );
nor ( n432700 , n87563 , n87569 );
buf ( n432701 , n432700 );
buf ( n432702 , n432701 );
xor ( n87573 , n432656 , n432663 );
xor ( n432704 , n87573 , n432684 );
buf ( n432705 , n432704 );
buf ( n432706 , n432705 );
not ( n87577 , n431989 );
buf ( n432708 , n431926 );
not ( n87579 , n432708 );
buf ( n432710 , n87579 );
not ( n87581 , n432710 );
and ( n432712 , n87577 , n87581 );
buf ( n432713 , n431989 );
buf ( n432714 , n432710 );
nand ( n87585 , n432713 , n432714 );
buf ( n432716 , n87585 );
and ( n87587 , n432716 , n431996 );
nor ( n432718 , n432712 , n87587 );
buf ( n432719 , n432718 );
not ( n432720 , n432719 );
xor ( n432721 , n432669 , n432675 );
xor ( n432722 , n432721 , n432679 );
buf ( n432723 , n432722 );
buf ( n432724 , n432723 );
not ( n432725 , n432724 );
or ( n432726 , n432720 , n432725 );
xor ( n432727 , n432129 , n432134 );
and ( n432728 , n432727 , n432140 );
and ( n432729 , n432129 , n432134 );
or ( n432730 , n432728 , n432729 );
buf ( n432731 , n432730 );
buf ( n432732 , n432731 );
nand ( n432733 , n432726 , n432732 );
buf ( n432734 , n432733 );
buf ( n432735 , n432734 );
buf ( n432736 , n432718 );
not ( n432737 , n432736 );
buf ( n432738 , n432723 );
not ( n432739 , n432738 );
buf ( n432740 , n432739 );
buf ( n432741 , n432740 );
nand ( n432742 , n432737 , n432741 );
buf ( n432743 , n432742 );
buf ( n432744 , n432743 );
and ( n432745 , n432735 , n432744 );
buf ( n432746 , n432745 );
buf ( n432747 , n432746 );
xor ( n432748 , n432706 , n432747 );
buf ( n432749 , n432279 );
buf ( n432750 , n432412 );
xor ( n432751 , n432749 , n432750 );
buf ( n432752 , n87346 );
xor ( n432753 , n432751 , n432752 );
buf ( n432754 , n432753 );
buf ( n432755 , n432754 );
and ( n432756 , n432748 , n432755 );
and ( n432757 , n432706 , n432747 );
or ( n432758 , n432756 , n432757 );
buf ( n432759 , n432758 );
buf ( n432760 , n432759 );
nand ( n432761 , n432702 , n432760 );
buf ( n432762 , n432761 );
buf ( n432763 , n432762 );
buf ( n432764 , n432431 );
not ( n432765 , n432764 );
buf ( n432766 , n432423 );
not ( n432767 , n432766 );
or ( n432768 , n432765 , n432767 );
buf ( n432769 , n432426 );
buf ( n432770 , n432436 );
nand ( n432771 , n432769 , n432770 );
buf ( n432772 , n432771 );
buf ( n432773 , n432772 );
nand ( n432774 , n432768 , n432773 );
buf ( n432775 , n432774 );
buf ( n432776 , n432775 );
buf ( n432777 , n432504 );
xor ( n432778 , n432776 , n432777 );
buf ( n432779 , n432778 );
buf ( n432780 , n432779 );
xor ( n432781 , n432098 , n432143 );
and ( n432782 , n432781 , n432150 );
and ( n432783 , n432098 , n432143 );
or ( n432784 , n432782 , n432783 );
buf ( n432785 , n432784 );
buf ( n432786 , n432785 );
xor ( n432787 , n432780 , n432786 );
buf ( n432788 , n432731 );
buf ( n432789 , n432718 );
xor ( n432790 , n432788 , n432789 );
buf ( n432791 , n432740 );
xnor ( n432792 , n432790 , n432791 );
buf ( n432793 , n432792 );
buf ( n432794 , n432793 );
and ( n432795 , n432787 , n432794 );
and ( n432796 , n432780 , n432786 );
or ( n432797 , n432795 , n432796 );
buf ( n432798 , n432797 );
buf ( n432799 , n432798 );
not ( n432800 , n432799 );
xor ( n432801 , n432706 , n432747 );
xor ( n432802 , n432801 , n432755 );
buf ( n432803 , n432802 );
buf ( n432804 , n432803 );
nand ( n432805 , n432800 , n432804 );
buf ( n432806 , n432805 );
buf ( n432807 , n432806 );
not ( n432808 , n432807 );
xor ( n432809 , n432780 , n432786 );
xor ( n432810 , n432809 , n432794 );
buf ( n432811 , n432810 );
buf ( n432812 , n432811 );
buf ( n432813 , n431999 );
not ( n432814 , n432813 );
buf ( n432815 , n432018 );
not ( n432816 , n432815 );
or ( n432817 , n432814 , n432816 );
or ( n432818 , n431999 , n432018 );
nand ( n432819 , n432818 , n432152 );
buf ( n432820 , n432819 );
nand ( n432821 , n432817 , n432820 );
buf ( n432822 , n432821 );
buf ( n432823 , n432822 );
nor ( n432824 , n432812 , n432823 );
buf ( n432825 , n432824 );
buf ( n432826 , n432825 );
nor ( n432827 , n432808 , n432826 );
buf ( n432828 , n432827 );
buf ( n432829 , n432828 );
nand ( n432830 , n432194 , n432763 , n432829 );
buf ( n432831 , n432830 );
buf ( n432832 , n432831 );
not ( n432833 , n432806 );
buf ( n432834 , n432822 );
buf ( n432835 , n432811 );
and ( n432836 , n432834 , n432835 );
buf ( n432837 , n432836 );
not ( n432838 , n432837 );
or ( n432839 , n432833 , n432838 );
buf ( n432840 , n432803 );
not ( n432841 , n432840 );
buf ( n432842 , n432798 );
nand ( n432843 , n432841 , n432842 );
buf ( n432844 , n432843 );
nand ( n432845 , n432839 , n432844 );
buf ( n432846 , n432845 );
buf ( n432847 , n432762 );
nand ( n432848 , n432846 , n432847 );
buf ( n432849 , n432848 );
buf ( n432850 , n432849 );
buf ( n432851 , n432701 );
buf ( n432852 , n432759 );
or ( n432853 , n432851 , n432852 );
buf ( n432854 , n432853 );
buf ( n432855 , n432854 );
nand ( n432856 , n432832 , n432850 , n432855 );
buf ( n432857 , n432856 );
buf ( n432858 , n432857 );
xor ( n432859 , n69144 , n416056 );
xor ( n432860 , n432859 , n416458 );
buf ( n432861 , n432860 );
buf ( n432862 , n416030 );
buf ( n432863 , n416035 );
xor ( n432864 , n432862 , n432863 );
buf ( n432865 , n416050 );
xnor ( n432866 , n432864 , n432865 );
buf ( n432867 , n432866 );
buf ( n432868 , n432867 );
not ( n432869 , n432868 );
xor ( n432870 , n416404 , n416407 );
xor ( n432871 , n432870 , n416454 );
buf ( n432872 , n432871 );
buf ( n432873 , n432872 );
not ( n432874 , n432873 );
buf ( n432875 , n432874 );
buf ( n432876 , n432875 );
not ( n432877 , n432876 );
or ( n432878 , n432869 , n432877 );
not ( n432879 , n432566 );
not ( n432880 , n87417 );
or ( n432881 , n432879 , n432880 );
buf ( n432882 , n87417 );
buf ( n432883 , n432566 );
or ( n432884 , n432882 , n432883 );
buf ( n432885 , n87413 );
nand ( n432886 , n432884 , n432885 );
buf ( n432887 , n432886 );
nand ( n432888 , n432881 , n432887 );
xor ( n432889 , n416411 , n416444 );
xor ( n432890 , n432889 , n416449 );
buf ( n432891 , n432890 );
xor ( n432892 , n432888 , n432891 );
xor ( n432893 , n416485 , n416488 );
xor ( n432894 , n432893 , n416609 );
buf ( n432895 , n432894 );
and ( n432896 , n432892 , n432895 );
and ( n432897 , n432888 , n432891 );
or ( n432898 , n432896 , n432897 );
buf ( n432899 , n432898 );
nand ( n432900 , n432878 , n432899 );
buf ( n432901 , n432900 );
buf ( n432902 , n432901 );
buf ( n432903 , n432867 );
not ( n432904 , n432903 );
buf ( n432905 , n432872 );
nand ( n432906 , n432904 , n432905 );
buf ( n432907 , n432906 );
buf ( n432908 , n432907 );
nand ( n432909 , n432902 , n432908 );
buf ( n432910 , n432909 );
buf ( n432911 , n432910 );
xor ( n432912 , n432861 , n432911 );
xor ( n432913 , n416469 , n416473 );
xor ( n432914 , n432913 , n417486 );
buf ( n432915 , n432914 );
buf ( n432916 , n432915 );
xor ( n432917 , n432912 , n432916 );
buf ( n432918 , n432917 );
buf ( n432919 , n432918 );
not ( n432920 , n432919 );
buf ( n432921 , n432920 );
buf ( n432922 , n432921 );
xor ( n432923 , n416613 , n416617 );
xor ( n432924 , n432923 , n417481 );
buf ( n432925 , n432924 );
not ( n432926 , n432925 );
buf ( n432927 , n432926 );
not ( n432928 , n432927 );
buf ( n432929 , n432867 );
buf ( n432930 , n432898 );
xor ( n432931 , n432929 , n432930 );
buf ( n432932 , n432872 );
xor ( n432933 , n432931 , n432932 );
buf ( n432934 , n432933 );
buf ( n432935 , n432934 );
not ( n432936 , n432935 );
or ( n432937 , n432928 , n432936 );
xor ( n432938 , n416622 , n417471 );
xor ( n432939 , n432938 , n417476 );
buf ( n432940 , n432939 );
buf ( n432941 , n432940 );
not ( n432942 , n87440 );
not ( n432943 , n87429 );
or ( n432944 , n432942 , n432943 );
not ( n432945 , n87441 );
not ( n432946 , n87506 );
or ( n432947 , n432945 , n432946 );
nand ( n432948 , n432947 , n87499 );
nand ( n432949 , n432944 , n432948 );
buf ( n432950 , n432949 );
or ( n432951 , n432941 , n432950 );
buf ( n432952 , n432951 );
buf ( n432953 , n432952 );
xor ( n432954 , n432517 , n432530 );
and ( n432955 , n432954 , n432537 );
and ( n432956 , n432517 , n432530 );
or ( n432957 , n432955 , n432956 );
buf ( n432958 , n432957 );
buf ( n432959 , n432958 );
and ( n432960 , n432953 , n432959 );
buf ( n432961 , n432940 );
buf ( n432962 , n432949 );
and ( n432963 , n432961 , n432962 );
buf ( n432964 , n432963 );
buf ( n432965 , n432964 );
nor ( n432966 , n432960 , n432965 );
buf ( n432967 , n432966 );
not ( n432968 , n432967 );
buf ( n432969 , n432968 );
nand ( n432970 , n432937 , n432969 );
buf ( n432971 , n432970 );
buf ( n432972 , n432971 );
buf ( n432973 , n432934 );
not ( n432974 , n432973 );
buf ( n432975 , n432974 );
buf ( n432976 , n432975 );
buf ( n432977 , n432925 );
nand ( n432978 , n432976 , n432977 );
buf ( n432979 , n432978 );
buf ( n432980 , n432979 );
nand ( n432981 , n432972 , n432980 );
buf ( n432982 , n432981 );
buf ( n432983 , n432982 );
not ( n432984 , n432983 );
buf ( n432985 , n432984 );
buf ( n432986 , n432985 );
nand ( n432987 , n432922 , n432986 );
buf ( n432988 , n432987 );
buf ( n432989 , n432988 );
not ( n432990 , n432989 );
xor ( n432991 , n417496 , n417497 );
buf ( n432992 , n432991 );
buf ( n432993 , n432992 );
buf ( n432994 , n69132 );
and ( n432995 , n432993 , n432994 );
not ( n432996 , n432993 );
buf ( n432997 , n69132 );
not ( n432998 , n432997 );
buf ( n432999 , n432998 );
buf ( n433000 , n432999 );
and ( n433001 , n432996 , n433000 );
nor ( n433002 , n432995 , n433001 );
buf ( n433003 , n433002 );
buf ( n433004 , n433003 );
xor ( n433005 , n432861 , n432911 );
and ( n433006 , n433005 , n432916 );
and ( n433007 , n432861 , n432911 );
or ( n433008 , n433006 , n433007 );
buf ( n433009 , n433008 );
buf ( n433010 , n433009 );
nor ( n433011 , n433004 , n433010 );
buf ( n433012 , n433011 );
buf ( n433013 , n433012 );
nor ( n433014 , n432990 , n433013 );
buf ( n433015 , n433014 );
buf ( n433016 , n433015 );
buf ( n433017 , n432545 );
not ( n433018 , n433017 );
buf ( n433019 , n432691 );
not ( n433020 , n433019 );
or ( n433021 , n433018 , n433020 );
buf ( n433022 , n432512 );
nand ( n433023 , n433021 , n433022 );
buf ( n433024 , n433023 );
buf ( n433025 , n433024 );
buf ( n433026 , n432697 );
buf ( n433027 , n432539 );
nand ( n433028 , n433026 , n433027 );
buf ( n433029 , n433028 );
buf ( n433030 , n433029 );
nand ( n433031 , n433025 , n433030 );
buf ( n433032 , n433031 );
buf ( n433033 , n433032 );
xor ( n433034 , n432961 , n432962 );
buf ( n433035 , n433034 );
buf ( n433036 , n433035 );
buf ( n433037 , n432958 );
not ( n433038 , n433037 );
buf ( n433039 , n433038 );
buf ( n433040 , n433039 );
and ( n433041 , n433036 , n433040 );
not ( n433042 , n433036 );
buf ( n433043 , n432958 );
and ( n433044 , n433042 , n433043 );
nor ( n433045 , n433041 , n433044 );
buf ( n433046 , n433045 );
xor ( n433047 , n432888 , n432891 );
xor ( n433048 , n433047 , n432895 );
buf ( n433049 , n433048 );
not ( n433050 , n433049 );
buf ( n433051 , n433050 );
buf ( n433052 , n433051 );
not ( n433053 , n433052 );
xor ( n433054 , n432577 , n432642 );
and ( n433055 , n433054 , n432689 );
and ( n433056 , n432577 , n432642 );
or ( n433057 , n433055 , n433056 );
buf ( n433058 , n433057 );
buf ( n433059 , n433058 );
not ( n433060 , n433059 );
buf ( n433061 , n433060 );
buf ( n433062 , n433061 );
not ( n433063 , n433062 );
or ( n433064 , n433053 , n433063 );
buf ( n433065 , n433058 );
buf ( n433066 , n433048 );
nand ( n433067 , n433065 , n433066 );
buf ( n433068 , n433067 );
buf ( n433069 , n433068 );
nand ( n433070 , n433064 , n433069 );
buf ( n433071 , n433070 );
xnor ( n433072 , n433046 , n433071 );
buf ( n433073 , n433072 );
or ( n433074 , n433033 , n433073 );
buf ( n433075 , n433074 );
buf ( n433076 , n433075 );
not ( n433077 , n432926 );
not ( n433078 , n432967 );
or ( n433079 , n433077 , n433078 );
nand ( n433080 , n432968 , n432925 );
nand ( n433081 , n433079 , n433080 );
and ( n433082 , n433081 , n432975 );
not ( n433083 , n433081 );
not ( n433084 , n432975 );
and ( n433085 , n433083 , n433084 );
nor ( n433086 , n433082 , n433085 );
buf ( n433087 , n433086 );
not ( n433088 , n433046 );
not ( n433089 , n433051 );
and ( n433090 , n433088 , n433089 );
buf ( n433091 , n433046 );
buf ( n433092 , n433051 );
nand ( n433093 , n433091 , n433092 );
buf ( n433094 , n433093 );
and ( n433095 , n433094 , n433061 );
nor ( n433096 , n433090 , n433095 );
buf ( n433097 , n433096 );
nand ( n433098 , n433087 , n433097 );
buf ( n433099 , n433098 );
buf ( n433100 , n433099 );
and ( n433101 , n433076 , n433100 );
buf ( n433102 , n433101 );
buf ( n433103 , n433102 );
nand ( n433104 , n432858 , n433016 , n433103 );
buf ( n433105 , n433104 );
buf ( n433106 , n433105 );
not ( n433107 , n432988 );
not ( n433108 , n433099 );
buf ( n433109 , n433072 );
buf ( n433110 , n433032 );
and ( n433111 , n433109 , n433110 );
buf ( n433112 , n433111 );
not ( n433113 , n433112 );
or ( n433114 , n433108 , n433113 );
buf ( n433115 , n433086 );
not ( n433116 , n433115 );
buf ( n433117 , n433116 );
buf ( n433118 , n433117 );
buf ( n433119 , n433096 );
not ( n433120 , n433119 );
buf ( n433121 , n433120 );
buf ( n433122 , n433121 );
nand ( n433123 , n433118 , n433122 );
buf ( n433124 , n433123 );
nand ( n433125 , n433114 , n433124 );
not ( n433126 , n433125 );
or ( n433127 , n433107 , n433126 );
buf ( n433128 , n433003 );
buf ( n433129 , n433009 );
nand ( n433130 , n433128 , n433129 );
buf ( n433131 , n433130 );
buf ( n433132 , n433131 );
buf ( n433133 , n432918 );
buf ( n433134 , n432982 );
nand ( n433135 , n433133 , n433134 );
buf ( n433136 , n433135 );
buf ( n433137 , n433136 );
and ( n433138 , n433132 , n433137 );
buf ( n433139 , n433138 );
nand ( n433140 , n433127 , n433139 );
buf ( n433141 , n433012 );
not ( n433142 , n433141 );
buf ( n433143 , n433142 );
nand ( n433144 , n433140 , n433143 );
buf ( n433145 , n433144 );
nand ( n433146 , n433106 , n433145 );
buf ( n433147 , n433146 );
not ( n433148 , n433147 );
or ( n433149 , n70878 , n433148 );
not ( n433150 , n415844 );
buf ( n433151 , n415848 );
buf ( n433152 , n417502 );
nor ( n433153 , n433151 , n433152 );
buf ( n433154 , n433153 );
not ( n433155 , n433154 );
or ( n433156 , n433150 , n433155 );
buf ( n433157 , n415768 );
not ( n433158 , n433157 );
buf ( n433159 , n433158 );
buf ( n433160 , n433159 );
buf ( n433161 , n415841 );
not ( n433162 , n433161 );
buf ( n433163 , n433162 );
buf ( n433164 , n433163 );
nand ( n433165 , n433160 , n433164 );
buf ( n433166 , n433165 );
nand ( n433167 , n433156 , n433166 );
and ( n433168 , n433167 , n69045 );
nor ( n433169 , n414401 , n415763 );
nor ( n433170 , n433168 , n433169 );
nand ( n433171 , n433149 , n433170 );
not ( n433172 , n412499 );
not ( n433173 , n412404 );
and ( n433174 , n433172 , n433173 );
nor ( n433175 , n67615 , n412627 );
nor ( n433176 , n433174 , n433175 );
nand ( n433177 , n433176 , n414370 , n67622 );
not ( n433178 , n433177 );
nand ( n433179 , n433171 , n433178 , n67642 );
not ( n433180 , n414379 );
not ( n433181 , n414384 );
nand ( n433182 , n433180 , n433181 );
nand ( n433183 , n67643 , n433179 , n433182 );
nand ( n433184 , n52628 , n405627 , n63019 , n433183 );
not ( n433185 , n433184 );
buf ( n433186 , n48197 );
not ( n433187 , n433186 );
buf ( n433188 , n48741 );
not ( n433189 , n433188 );
or ( n433190 , n433187 , n433189 );
buf ( n433191 , n48741 );
buf ( n433192 , n48197 );
or ( n433193 , n433191 , n433192 );
buf ( n433194 , n48207 );
nand ( n433195 , n433193 , n433194 );
buf ( n433196 , n433195 );
buf ( n433197 , n433196 );
nand ( n433198 , n433190 , n433197 );
buf ( n433199 , n433198 );
buf ( n433200 , n433199 );
not ( n433201 , n433200 );
buf ( n433202 , n433201 );
buf ( n433203 , n433202 );
buf ( n433204 , n388806 );
not ( n433205 , n433204 );
buf ( n433206 , n388743 );
not ( n433207 , n433206 );
or ( n433208 , n433205 , n433207 );
buf ( n433209 , n48524 );
nand ( n433210 , n433208 , n433209 );
buf ( n433211 , n433210 );
buf ( n433212 , n433211 );
buf ( n433213 , n386480 );
not ( n433214 , n433213 );
buf ( n433215 , n38972 );
not ( n433216 , n433215 );
buf ( n433217 , n383762 );
not ( n433218 , n433217 );
or ( n433219 , n433216 , n433218 );
buf ( n433220 , n42152 );
buf ( n433221 , n38971 );
nand ( n433222 , n433220 , n433221 );
buf ( n433223 , n433222 );
buf ( n433224 , n433223 );
nand ( n433225 , n433219 , n433224 );
buf ( n433226 , n433225 );
buf ( n433227 , n433226 );
not ( n433228 , n433227 );
or ( n433229 , n433214 , n433228 );
buf ( n433230 , n395680 );
buf ( n433231 , n386496 );
nand ( n433232 , n433230 , n433231 );
buf ( n433233 , n433232 );
buf ( n433234 , n433233 );
nand ( n433235 , n433229 , n433234 );
buf ( n433236 , n433235 );
buf ( n433237 , n433236 );
xor ( n433238 , n433212 , n433237 );
buf ( n433239 , n389162 );
not ( n433240 , n433239 );
buf ( n433241 , n41671 );
not ( n433242 , n433241 );
buf ( n433243 , n382535 );
not ( n433244 , n433243 );
or ( n433245 , n433242 , n433244 );
buf ( n433246 , n382548 );
not ( n433247 , n433246 );
buf ( n433248 , n41670 );
nand ( n433249 , n433247 , n433248 );
buf ( n433250 , n433249 );
buf ( n433251 , n433250 );
nand ( n433252 , n433245 , n433251 );
buf ( n433253 , n433252 );
buf ( n433254 , n433253 );
not ( n433255 , n433254 );
or ( n433256 , n433240 , n433255 );
buf ( n433257 , n48423 );
buf ( n433258 , n41711 );
nand ( n433259 , n433257 , n433258 );
buf ( n433260 , n433259 );
buf ( n433261 , n433260 );
nand ( n433262 , n433256 , n433261 );
buf ( n433263 , n433262 );
buf ( n433264 , n433263 );
xor ( n433265 , n433238 , n433264 );
buf ( n433266 , n433265 );
buf ( n433267 , n433266 );
xor ( n433268 , n395851 , n395868 );
and ( n433269 , n433268 , n395940 );
and ( n433270 , n395851 , n395868 );
or ( n433271 , n433269 , n433270 );
buf ( n433272 , n433271 );
buf ( n433273 , n433272 );
xor ( n433274 , n433267 , n433273 );
xor ( n433275 , n396053 , n396064 );
and ( n433276 , n433275 , n396087 );
and ( n433277 , n396053 , n396064 );
or ( n433278 , n433276 , n433277 );
buf ( n433279 , n433278 );
buf ( n433280 , n433279 );
xor ( n433281 , n433274 , n433280 );
buf ( n433282 , n433281 );
buf ( n433283 , n433282 );
not ( n433284 , n396089 );
not ( n433285 , n396106 );
xor ( n433286 , n396164 , n396148 );
not ( n433287 , n433286 );
nand ( n433288 , n433287 , n396170 );
not ( n433289 , n396170 );
nand ( n433290 , n433289 , n433286 );
nand ( n433291 , n433285 , n433288 , n433290 );
not ( n433292 , n433291 );
or ( n433293 , n433284 , n433292 );
nand ( n433294 , n396106 , n48734 );
nand ( n433295 , n433293 , n433294 );
buf ( n433296 , n433295 );
xor ( n433297 , n433283 , n433296 );
xor ( n433298 , n396114 , n396139 );
and ( n433299 , n433298 , n396146 );
and ( n433300 , n396114 , n396139 );
or ( n433301 , n433299 , n433300 );
buf ( n433302 , n433301 );
buf ( n433303 , n433302 );
buf ( n433304 , n390403 );
not ( n433305 , n433304 );
buf ( n433306 , n24074 );
buf ( n433307 , n37370 );
and ( n433308 , n433306 , n433307 );
not ( n433309 , n433306 );
buf ( n433310 , n49933 );
and ( n433311 , n433309 , n433310 );
nor ( n433312 , n433308 , n433311 );
buf ( n433313 , n433312 );
buf ( n433314 , n433313 );
not ( n433315 , n433314 );
or ( n433316 , n433305 , n433315 );
buf ( n433317 , n396005 );
buf ( n433318 , n391080 );
nand ( n433319 , n433317 , n433318 );
buf ( n433320 , n433319 );
buf ( n433321 , n433320 );
nand ( n433322 , n433316 , n433321 );
buf ( n433323 , n433322 );
buf ( n433324 , n433323 );
xor ( n433325 , n433303 , n433324 );
xor ( n433326 , n395691 , n395697 );
and ( n433327 , n433326 , n395769 );
and ( n433328 , n395691 , n395697 );
or ( n433329 , n433327 , n433328 );
buf ( n433330 , n433329 );
buf ( n433331 , n433330 );
xor ( n433332 , n433325 , n433331 );
buf ( n433333 , n433332 );
buf ( n433334 , n433333 );
buf ( n433335 , n37695 );
not ( n433336 , n433335 );
buf ( n433337 , n391895 );
not ( n433338 , n433337 );
buf ( n433339 , n433338 );
buf ( n433340 , n433339 );
not ( n433341 , n433340 );
buf ( n433342 , n389467 );
not ( n433343 , n433342 );
or ( n433344 , n433341 , n433343 );
buf ( n433345 , n384974 );
buf ( n433346 , n37346 );
nand ( n433347 , n433345 , n433346 );
buf ( n433348 , n433347 );
buf ( n433349 , n433348 );
nand ( n433350 , n433344 , n433349 );
buf ( n433351 , n433350 );
buf ( n433352 , n433351 );
not ( n433353 , n433352 );
or ( n433354 , n433336 , n433353 );
buf ( n433355 , n395840 );
buf ( n433356 , n385269 );
nand ( n433357 , n433355 , n433356 );
buf ( n433358 , n433357 );
buf ( n433359 , n433358 );
nand ( n433360 , n433354 , n433359 );
buf ( n433361 , n433360 );
buf ( n433362 , n433361 );
buf ( n433363 , n395735 );
not ( n433364 , n433363 );
buf ( n433365 , n48275 );
not ( n433366 , n433365 );
or ( n433367 , n433364 , n433366 );
buf ( n433368 , n395763 );
nand ( n433369 , n433367 , n433368 );
buf ( n433370 , n433369 );
not ( n433371 , n48275 );
nand ( n433372 , n433371 , n395738 );
nand ( n433373 , n433370 , n433372 );
buf ( n433374 , n433373 );
xor ( n433375 , n433362 , n433374 );
buf ( n433376 , n38324 );
not ( n433377 , n433376 );
buf ( n433378 , n385494 );
not ( n433379 , n433378 );
buf ( n433380 , n385734 );
not ( n433381 , n433380 );
or ( n433382 , n433379 , n433381 );
buf ( n433383 , n384186 );
buf ( n433384 , n385491 );
nand ( n433385 , n433383 , n433384 );
buf ( n433386 , n433385 );
buf ( n433387 , n433386 );
nand ( n433388 , n433382 , n433387 );
buf ( n433389 , n433388 );
buf ( n433390 , n433389 );
not ( n433391 , n433390 );
or ( n433392 , n433377 , n433391 );
buf ( n433393 , n396131 );
buf ( n433394 , n385479 );
nand ( n433395 , n433393 , n433394 );
buf ( n433396 , n433395 );
buf ( n433397 , n433396 );
nand ( n433398 , n433392 , n433397 );
buf ( n433399 , n433398 );
buf ( n433400 , n433399 );
xor ( n433401 , n433375 , n433400 );
buf ( n433402 , n433401 );
buf ( n433403 , n433402 );
not ( n433404 , n388141 );
not ( n433405 , n35301 );
not ( n433406 , n388157 );
or ( n433407 , n433405 , n433406 );
nand ( n433408 , n388160 , n386385 );
nand ( n433409 , n433407 , n433408 );
not ( n433410 , n433409 );
or ( n433411 , n433404 , n433410 );
buf ( n433412 , n396076 );
buf ( n433413 , n40701 );
nand ( n433414 , n433412 , n433413 );
buf ( n433415 , n433414 );
nand ( n433416 , n433411 , n433415 );
buf ( n433417 , n433416 );
xor ( n433418 , n433403 , n433417 );
buf ( n433419 , n388833 );
not ( n433420 , n433419 );
and ( n433421 , n383059 , n41342 );
not ( n433422 , n383059 );
and ( n433423 , n433422 , n41349 );
or ( n433424 , n433421 , n433423 );
buf ( n433425 , n433424 );
not ( n433426 , n433425 );
or ( n433427 , n433420 , n433426 );
buf ( n433428 , n48717 );
buf ( n433429 , n388872 );
nand ( n433430 , n433428 , n433429 );
buf ( n433431 , n433430 );
buf ( n433432 , n433431 );
nand ( n433433 , n433427 , n433432 );
buf ( n433434 , n433433 );
buf ( n433435 , n433434 );
xor ( n433436 , n433418 , n433435 );
buf ( n433437 , n433436 );
buf ( n433438 , n433437 );
xor ( n433439 , n433334 , n433438 );
buf ( n433440 , n396148 );
buf ( n433441 , n433440 );
not ( n433442 , n433441 );
buf ( n433443 , n396164 );
not ( n433444 , n433443 );
or ( n433445 , n433442 , n433444 );
buf ( n433446 , n433440 );
buf ( n433447 , n396164 );
or ( n433448 , n433446 , n433447 );
buf ( n433449 , n396170 );
nand ( n433450 , n433448 , n433449 );
buf ( n433451 , n433450 );
buf ( n433452 , n433451 );
nand ( n433453 , n433445 , n433452 );
buf ( n433454 , n433453 );
buf ( n433455 , n433454 );
xor ( n433456 , n433439 , n433455 );
buf ( n433457 , n433456 );
buf ( n433458 , n433457 );
xor ( n433459 , n433297 , n433458 );
buf ( n433460 , n433459 );
not ( n433461 , n433460 );
not ( n433462 , n48213 );
nand ( n433463 , n48585 , n433462 );
not ( n433464 , n433463 );
not ( n433465 , n396177 );
or ( n433466 , n433464 , n433465 );
nand ( n433467 , n396021 , n48213 );
nand ( n433468 , n433466 , n433467 );
xor ( n433469 , n433461 , n433468 );
xor ( n433470 , n395658 , n395946 );
and ( n433471 , n433470 , n396019 );
and ( n433472 , n395658 , n395946 );
or ( n433473 , n433471 , n433472 );
buf ( n433474 , n433473 );
buf ( n433475 , n433474 );
xor ( n433476 , n395664 , n395772 );
and ( n433477 , n433476 , n395943 );
and ( n433478 , n395664 , n395772 );
or ( n433479 , n433477 , n433478 );
buf ( n433480 , n433479 );
buf ( n433481 , n433480 );
xor ( n433482 , n395953 , n396009 );
and ( n433483 , n433482 , n396016 );
and ( n433484 , n395953 , n396009 );
or ( n433485 , n433483 , n433484 );
buf ( n433486 , n433485 );
buf ( n433487 , n433486 );
xor ( n433488 , n433481 , n433487 );
buf ( n433489 , n395815 );
buf ( n433490 , n395757 );
not ( n433491 , n433490 );
buf ( n433492 , n389744 );
not ( n433493 , n433492 );
or ( n433494 , n433491 , n433493 );
buf ( n433495 , n379463 );
buf ( n433496 , n388646 );
not ( n433497 , n433496 );
buf ( n433498 , n382994 );
not ( n433499 , n433498 );
or ( n433500 , n433497 , n433499 );
buf ( n433501 , n385975 );
buf ( n433502 , n388654 );
nand ( n433503 , n433501 , n433502 );
buf ( n433504 , n433503 );
buf ( n433505 , n433504 );
nand ( n433506 , n433500 , n433505 );
buf ( n433507 , n433506 );
buf ( n433508 , n433507 );
nand ( n433509 , n433495 , n433508 );
buf ( n433510 , n433509 );
buf ( n433511 , n433510 );
nand ( n433512 , n433494 , n433511 );
buf ( n433513 , n433512 );
buf ( n433514 , n433513 );
xor ( n433515 , n433489 , n433514 );
buf ( n433516 , n395929 );
not ( n433517 , n433516 );
buf ( n433518 , n391270 );
not ( n433519 , n433518 );
or ( n433520 , n433517 , n433519 );
buf ( n433521 , n391173 );
not ( n433522 , n44399 );
not ( n433523 , n389598 );
or ( n433524 , n433522 , n433523 );
buf ( n433525 , n383423 );
buf ( n433526 , n41195 );
nand ( n433527 , n433525 , n433526 );
buf ( n433528 , n433527 );
nand ( n433529 , n433524 , n433528 );
buf ( n433530 , n433529 );
nand ( n433531 , n433521 , n433530 );
buf ( n433532 , n433531 );
buf ( n433533 , n433532 );
nand ( n433534 , n433520 , n433533 );
buf ( n433535 , n433534 );
buf ( n433536 , n433535 );
xor ( n433537 , n433515 , n433536 );
buf ( n433538 , n433537 );
buf ( n433539 , n433538 );
xor ( n433540 , n395895 , n395909 );
and ( n433541 , n433540 , n395937 );
and ( n433542 , n395895 , n395909 );
or ( n433543 , n433541 , n433542 );
buf ( n433544 , n433543 );
buf ( n433545 , n433544 );
xor ( n433546 , n433539 , n433545 );
buf ( n433547 , n384644 );
not ( n433548 , n433547 );
buf ( n433549 , n389928 );
not ( n433550 , n433549 );
buf ( n433551 , n38159 );
not ( n433552 , n433551 );
or ( n433553 , n433550 , n433552 );
buf ( n433554 , n36564 );
buf ( n433555 , n36252 );
nand ( n433556 , n433554 , n433555 );
buf ( n433557 , n433556 );
buf ( n433558 , n433557 );
nand ( n433559 , n433553 , n433558 );
buf ( n433560 , n433559 );
buf ( n433561 , n433560 );
not ( n433562 , n433561 );
or ( n433563 , n433548 , n433562 );
buf ( n433564 , n395787 );
buf ( n433565 , n383897 );
nand ( n433566 , n433564 , n433565 );
buf ( n433567 , n433566 );
buf ( n433568 , n433567 );
nand ( n433569 , n433563 , n433568 );
buf ( n433570 , n433569 );
buf ( n433571 , n433570 );
buf ( n433572 , n395889 );
not ( n433573 , n433572 );
buf ( n433574 , n433573 );
buf ( n433575 , n433574 );
not ( n433576 , n433575 );
buf ( n433577 , n384627 );
not ( n433578 , n433577 );
or ( n433579 , n433576 , n433578 );
and ( n433580 , n27196 , n42390 );
not ( n433581 , n27196 );
and ( n433582 , n433581 , n395885 );
or ( n433583 , n433580 , n433582 );
buf ( n433584 , n433583 );
buf ( n433585 , n384557 );
nand ( n433586 , n433584 , n433585 );
buf ( n433587 , n433586 );
buf ( n433588 , n433587 );
nand ( n433589 , n433579 , n433588 );
buf ( n433590 , n433589 );
buf ( n433591 , n433590 );
xor ( n433592 , n433571 , n433591 );
buf ( n433593 , n48469 );
not ( n433594 , n433593 );
buf ( n433595 , n383017 );
not ( n433596 , n433595 );
or ( n433597 , n433594 , n433596 );
buf ( n433598 , n383137 );
buf ( n433599 , n390490 );
not ( n433600 , n433599 );
buf ( n433601 , n398740 );
not ( n433602 , n433601 );
or ( n433603 , n433600 , n433602 );
buf ( n433604 , n40714 );
not ( n433605 , n433604 );
buf ( n433606 , n433605 );
buf ( n433607 , n433606 );
buf ( n433608 , n388569 );
nand ( n433609 , n433607 , n433608 );
buf ( n433610 , n433609 );
buf ( n433611 , n433610 );
nand ( n433612 , n433603 , n433611 );
buf ( n433613 , n433612 );
buf ( n433614 , n433613 );
nand ( n433615 , n433598 , n433614 );
buf ( n433616 , n433615 );
buf ( n433617 , n433616 );
nand ( n433618 , n433597 , n433617 );
buf ( n433619 , n433618 );
buf ( n433620 , n433619 );
xor ( n433621 , n433592 , n433620 );
buf ( n433622 , n433621 );
buf ( n433623 , n433622 );
xor ( n433624 , n433546 , n433623 );
buf ( n433625 , n433624 );
not ( n433626 , n41565 );
buf ( n433627 , n24050 );
not ( n433628 , n433627 );
buf ( n433629 , n38357 );
not ( n433630 , n433629 );
or ( n433631 , n433628 , n433630 );
buf ( n433632 , n51163 );
buf ( n433633 , n389075 );
nand ( n433634 , n433632 , n433633 );
buf ( n433635 , n433634 );
buf ( n433636 , n433635 );
nand ( n433637 , n433631 , n433636 );
buf ( n433638 , n433637 );
not ( n433639 , n433638 );
or ( n433640 , n433626 , n433639 );
nand ( n433641 , n395983 , n389125 );
nand ( n433642 , n433640 , n433641 );
not ( n433643 , n433642 );
xor ( n433644 , n395798 , n395819 );
and ( n433645 , n433644 , n395848 );
and ( n433646 , n395798 , n395819 );
or ( n433647 , n433645 , n433646 );
buf ( n433648 , n433647 );
not ( n433649 , n433648 );
not ( n433650 , n433649 );
or ( n433651 , n433643 , n433650 );
not ( n433652 , n433642 );
nand ( n433653 , n433648 , n433652 );
nand ( n433654 , n433651 , n433653 );
buf ( n433655 , n40972 );
not ( n433656 , n433655 );
buf ( n433657 , n385356 );
not ( n433658 , n433657 );
or ( n433659 , n433656 , n433658 );
buf ( n433660 , n385342 );
buf ( n433661 , n36395 );
nand ( n433662 , n433660 , n433661 );
buf ( n433663 , n433662 );
buf ( n433664 , n433663 );
nand ( n433665 , n433659 , n433664 );
buf ( n433666 , n433665 );
not ( n433667 , n433666 );
not ( n433668 , n43272 );
or ( n433669 , n433667 , n433668 );
nand ( n433670 , n40840 , n388928 );
or ( n433671 , n40840 , n388928 );
nand ( n433672 , n433670 , n433671 , n64851 );
nand ( n433673 , n433669 , n433672 );
not ( n433674 , n433673 );
buf ( n433675 , n395729 );
not ( n433676 , n433675 );
buf ( n433677 , n433676 );
not ( n433678 , n433677 );
not ( n433679 , n36801 );
or ( n433680 , n433678 , n433679 );
buf ( n433681 , n392111 );
buf ( n433682 , n40886 );
buf ( n433683 , n390271 );
and ( n433684 , n433682 , n433683 );
not ( n433685 , n433682 );
buf ( n433686 , n375784 );
and ( n433687 , n433685 , n433686 );
nor ( n433688 , n433684 , n433687 );
buf ( n433689 , n433688 );
buf ( n433690 , n433689 );
nand ( n433691 , n433681 , n433690 );
buf ( n433692 , n433691 );
nand ( n433693 , n433680 , n433692 );
xor ( n433694 , n433674 , n433693 );
buf ( n433695 , n389348 );
buf ( n433696 , n389602 );
buf ( n433697 , n384143 );
and ( n433698 , n433696 , n433697 );
not ( n433699 , n433696 );
buf ( n433700 , n382857 );
and ( n433701 , n433699 , n433700 );
nor ( n433702 , n433698 , n433701 );
buf ( n433703 , n433702 );
buf ( n433704 , n433703 );
or ( n433705 , n433695 , n433704 );
nand ( n433706 , C1 , n433705 );
buf ( n433707 , n433706 );
xnor ( n433708 , n433694 , n433707 );
not ( n433709 , n433708 );
xor ( n433710 , n433654 , n433709 );
or ( n433711 , n48551 , n48570 );
nand ( n433712 , n433711 , n48531 );
nand ( n433713 , n48570 , n48551 );
nand ( n433714 , n433712 , n433713 );
not ( n433715 , n433714 );
nand ( n433716 , n433710 , n433715 );
nand ( n433717 , n433625 , n433716 );
not ( n433718 , n433717 );
nor ( n433719 , n433716 , n433625 );
nor ( n433720 , n433710 , n433715 );
nor ( n433721 , n433719 , n433720 );
not ( n433722 , n433721 );
or ( n433723 , n433718 , n433722 );
not ( n433724 , n433710 );
nand ( n433725 , n433724 , n433625 , n433714 );
nand ( n433726 , n433723 , n433725 );
buf ( n433727 , n433726 );
xor ( n433728 , n433488 , n433727 );
buf ( n433729 , n433728 );
buf ( n433730 , n433729 );
xor ( n433731 , n433475 , n433730 );
xor ( n433732 , n396029 , n396035 );
and ( n433733 , n433732 , n396175 );
and ( n433734 , n396029 , n396035 );
or ( n433735 , n433733 , n433734 );
buf ( n433736 , n433735 );
buf ( n433737 , n433736 );
xor ( n433738 , n433731 , n433737 );
buf ( n433739 , n433738 );
xnor ( n433740 , n433469 , n433739 );
buf ( n433741 , n433740 );
not ( n433742 , n433741 );
buf ( n433743 , n433742 );
buf ( n433744 , n433743 );
nand ( n433745 , n433203 , n433744 );
buf ( n433746 , n433745 );
buf ( n433747 , n433746 );
xor ( n433748 , n433212 , n433237 );
and ( n433749 , n433748 , n433264 );
and ( n433750 , n433212 , n433237 );
or ( n433751 , n433749 , n433750 );
buf ( n433752 , n433751 );
buf ( n433753 , n433752 );
buf ( n433754 , n386496 );
not ( n433755 , n433754 );
buf ( n433756 , n433226 );
not ( n433757 , n433756 );
or ( n433758 , n433755 , n433757 );
buf ( n433759 , n386480 );
buf ( n433760 , n38972 );
buf ( n433761 , n37173 );
and ( n433762 , n433760 , n433761 );
not ( n433763 , n433760 );
buf ( n433764 , n389525 );
and ( n433765 , n433763 , n433764 );
nor ( n433766 , n433762 , n433765 );
buf ( n433767 , n433766 );
buf ( n433768 , n433767 );
nand ( n433769 , n433759 , n433768 );
buf ( n433770 , n433769 );
buf ( n433771 , n433770 );
nand ( n433772 , n433758 , n433771 );
buf ( n433773 , n433772 );
buf ( n433774 , n41711 );
not ( n433775 , n433774 );
buf ( n433776 , n433253 );
not ( n433777 , n433776 );
or ( n433778 , n433775 , n433777 );
not ( n433779 , n24117 );
not ( n433780 , n399653 );
or ( n433781 , n433779 , n433780 );
nand ( n433782 , n41671 , n388113 );
nand ( n433783 , n433781 , n433782 );
nand ( n433784 , n433783 , n389162 );
buf ( n433785 , n433784 );
nand ( n433786 , n433778 , n433785 );
buf ( n433787 , n433786 );
xor ( n433788 , n433773 , n433787 );
xor ( n433789 , n433571 , n433591 );
and ( n433790 , n433789 , n433620 );
and ( n433791 , n433571 , n433591 );
or ( n433792 , n433790 , n433791 );
buf ( n433793 , n433792 );
xor ( n433794 , n433788 , n433793 );
buf ( n433795 , n433794 );
xor ( n433796 , n433753 , n433795 );
buf ( n433797 , n388872 );
not ( n433798 , n433797 );
buf ( n433799 , n433424 );
not ( n433800 , n433799 );
or ( n433801 , n433798 , n433800 );
buf ( n433802 , n41349 );
buf ( n433803 , n35519 );
and ( n433804 , n433802 , n433803 );
not ( n433805 , n433802 );
buf ( n433806 , n392144 );
and ( n433807 , n433805 , n433806 );
nor ( n433808 , n433804 , n433807 );
buf ( n433809 , n433808 );
buf ( n433810 , n433809 );
not ( n433811 , n433810 );
buf ( n433812 , n388833 );
nand ( n433813 , n433811 , n433812 );
buf ( n433814 , n433813 );
buf ( n433815 , n433814 );
nand ( n433816 , n433801 , n433815 );
buf ( n433817 , n433816 );
buf ( n433818 , n433817 );
xor ( n433819 , n433362 , n433374 );
and ( n433820 , n433819 , n433400 );
and ( n433821 , n433362 , n433374 );
or ( n433822 , n433820 , n433821 );
buf ( n433823 , n433822 );
buf ( n433824 , n433823 );
xor ( n433825 , n433818 , n433824 );
buf ( n433826 , n391080 );
not ( n433827 , n433826 );
buf ( n433828 , n433313 );
not ( n433829 , n433828 );
or ( n433830 , n433827 , n433829 );
buf ( n433831 , n24074 );
not ( n433832 , n433831 );
buf ( n433833 , n37027 );
not ( n433834 , n433833 );
or ( n433835 , n433832 , n433834 );
nand ( n433836 , n39051 , n24073 );
buf ( n433837 , n433836 );
nand ( n433838 , n433835 , n433837 );
buf ( n433839 , n433838 );
buf ( n433840 , n433839 );
buf ( n433841 , n390403 );
nand ( n433842 , n433840 , n433841 );
buf ( n433843 , n433842 );
buf ( n433844 , n433843 );
nand ( n433845 , n433830 , n433844 );
buf ( n433846 , n433845 );
buf ( n433847 , n433846 );
xnor ( n433848 , n433825 , n433847 );
buf ( n433849 , n433848 );
buf ( n433850 , n433849 );
xnor ( n433851 , n433796 , n433850 );
buf ( n433852 , n433851 );
buf ( n433853 , n433852 );
xor ( n433854 , n433334 , n433438 );
and ( n433855 , n433854 , n433455 );
and ( n433856 , n433334 , n433438 );
or ( n433857 , n433855 , n433856 );
buf ( n433858 , n433857 );
buf ( n433859 , n433858 );
xor ( n433860 , n433853 , n433859 );
xor ( n433861 , n433403 , n433417 );
and ( n433862 , n433861 , n433435 );
and ( n433863 , n433403 , n433417 );
or ( n433864 , n433862 , n433863 );
buf ( n433865 , n433864 );
buf ( n433866 , n433865 );
not ( n433867 , n433866 );
buf ( n433868 , n433867 );
xor ( n433869 , n433303 , n433324 );
and ( n433870 , n433869 , n433331 );
and ( n433871 , n433303 , n433324 );
or ( n433872 , n433870 , n433871 );
buf ( n433873 , n433872 );
not ( n433874 , n433873 );
and ( n433875 , n433868 , n433874 );
not ( n433876 , n433868 );
and ( n433877 , n433876 , n433873 );
or ( n433878 , n433875 , n433877 );
buf ( n433879 , n433642 );
not ( n433880 , n433879 );
buf ( n433881 , n433708 );
not ( n433882 , n433881 );
or ( n433883 , n433880 , n433882 );
not ( n433884 , n433652 );
not ( n433885 , n433709 );
or ( n433886 , n433884 , n433885 );
nand ( n433887 , n433886 , n433648 );
buf ( n433888 , n433887 );
nand ( n433889 , n433883 , n433888 );
buf ( n433890 , n433889 );
not ( n433891 , n40701 );
not ( n433892 , n433409 );
or ( n433893 , n433891 , n433892 );
xor ( n433894 , n388160 , n382921 );
nand ( n433895 , n433894 , n388141 );
nand ( n433896 , n433893 , n433895 );
not ( n433897 , n433896 );
buf ( n433898 , n433613 );
not ( n433899 , n433898 );
buf ( n433900 , n396868 );
not ( n433901 , n433900 );
or ( n433902 , n433899 , n433901 );
buf ( n433903 , n383137 );
buf ( n433904 , n389862 );
not ( n433905 , n433904 );
buf ( n433906 , n398740 );
not ( n433907 , n433906 );
or ( n433908 , n433905 , n433907 );
buf ( n433909 , n386223 );
buf ( n433910 , n389859 );
nand ( n433911 , n433909 , n433910 );
buf ( n433912 , n433911 );
buf ( n433913 , n433912 );
nand ( n433914 , n433908 , n433913 );
buf ( n433915 , n433914 );
buf ( n433916 , n433915 );
nand ( n433917 , n433903 , n433916 );
buf ( n433918 , n433917 );
buf ( n433919 , n433918 );
nand ( n433920 , n433902 , n433919 );
buf ( n433921 , n433920 );
buf ( n433922 , n433921 );
buf ( n433923 , n433529 );
not ( n433924 , n433923 );
buf ( n433925 , n391164 );
not ( n433926 , n433925 );
buf ( n433927 , n433926 );
buf ( n433928 , n433927 );
not ( n433929 , n433928 );
or ( n433930 , n433924 , n433929 );
buf ( n433931 , n383423 );
not ( n433932 , n433931 );
buf ( n433933 , n388445 );
not ( n433934 , n433933 );
and ( n433935 , n433932 , n433934 );
buf ( n433936 , n389589 );
buf ( n433937 , n388445 );
and ( n433938 , n433936 , n433937 );
nor ( n433939 , n433935 , n433938 );
buf ( n433940 , n433939 );
buf ( n433941 , n433940 );
not ( n433942 , n433941 );
buf ( n433943 , n383406 );
nand ( n433944 , n433942 , n433943 );
buf ( n433945 , n433944 );
buf ( n433946 , n433945 );
nand ( n433947 , n433930 , n433946 );
buf ( n433948 , n433947 );
buf ( n433949 , n433948 );
xor ( n433950 , n433922 , n433949 );
buf ( n433951 , n433674 );
not ( n433952 , n433951 );
not ( n433953 , n433693 );
buf ( n433954 , n433953 );
not ( n433955 , n433954 );
or ( n433956 , n433952 , n433955 );
buf ( n433957 , n433707 );
nand ( n433958 , n433956 , n433957 );
buf ( n433959 , n433958 );
buf ( n433960 , n433959 );
buf ( n433961 , n433693 );
buf ( n433962 , n433673 );
nand ( n433963 , n433961 , n433962 );
buf ( n433964 , n433963 );
buf ( n433965 , n433964 );
nand ( n433966 , n433960 , n433965 );
buf ( n433967 , n433966 );
buf ( n433968 , n433967 );
xor ( n433969 , n433950 , n433968 );
buf ( n433970 , n433969 );
not ( n433971 , n433970 );
xor ( n433972 , n433897 , n433971 );
xnor ( n433973 , n433890 , n433972 );
buf ( n433974 , n433973 );
and ( n433975 , n433878 , n433974 );
not ( n433976 , n433878 );
not ( n433977 , n433974 );
and ( n433978 , n433976 , n433977 );
nor ( n433979 , n433975 , n433978 );
buf ( n433980 , n433979 );
xor ( n433981 , n433860 , n433980 );
buf ( n433982 , n433981 );
xor ( n433983 , n433475 , n433730 );
and ( n433984 , n433983 , n433737 );
and ( n433985 , n433475 , n433730 );
or ( n433986 , n433984 , n433985 );
buf ( n433987 , n433986 );
xor ( n433988 , n433982 , n433987 );
not ( n433989 , n433716 );
not ( n433990 , n433625 );
or ( n433991 , n433989 , n433990 );
not ( n433992 , n433720 );
nand ( n433993 , n433991 , n433992 );
buf ( n433994 , n433993 );
xor ( n433995 , n433267 , n433273 );
and ( n433996 , n433995 , n433280 );
and ( n433997 , n433267 , n433273 );
or ( n433998 , n433996 , n433997 );
buf ( n433999 , n433998 );
buf ( n434000 , n433999 );
xor ( n434001 , n433994 , n434000 );
buf ( n434002 , n385269 );
not ( n434003 , n434002 );
buf ( n434004 , n433351 );
not ( n434005 , n434004 );
or ( n434006 , n434003 , n434005 );
buf ( n434007 , n433339 );
not ( n434008 , n434007 );
buf ( n434009 , n384239 );
not ( n434010 , n434009 );
or ( n434011 , n434008 , n434010 );
buf ( n434012 , n389692 );
buf ( n434013 , n37346 );
nand ( n434014 , n434012 , n434013 );
buf ( n434015 , n434014 );
buf ( n434016 , n434015 );
nand ( n434017 , n434011 , n434016 );
buf ( n434018 , n434017 );
buf ( n434019 , n434018 );
buf ( n434020 , n37695 );
nand ( n434021 , n434019 , n434020 );
buf ( n434022 , n434021 );
buf ( n434023 , n434022 );
nand ( n434024 , n434006 , n434023 );
buf ( n434025 , n434024 );
buf ( n434026 , n434025 );
buf ( n434027 , n385479 );
not ( n434028 , n434027 );
buf ( n434029 , n433389 );
not ( n434030 , n434029 );
or ( n434031 , n434028 , n434030 );
buf ( n434032 , n385494 );
not ( n434033 , n434032 );
buf ( n434034 , n48233 );
not ( n434035 , n434034 );
or ( n434036 , n434033 , n434035 );
buf ( n434037 , n69799 );
buf ( n434038 , n385491 );
nand ( n434039 , n434037 , n434038 );
buf ( n434040 , n434039 );
buf ( n434041 , n434040 );
nand ( n434042 , n434036 , n434041 );
buf ( n434043 , n434042 );
buf ( n434044 , n434043 );
buf ( n434045 , n41447 );
nand ( n434046 , n434044 , n434045 );
buf ( n434047 , n434046 );
buf ( n434048 , n434047 );
nand ( n434049 , n434031 , n434048 );
buf ( n434050 , n434049 );
buf ( n434051 , n434050 );
xor ( n434052 , n434026 , n434051 );
xor ( n434053 , n433489 , n433514 );
and ( n434054 , n434053 , n433536 );
and ( n434055 , n433489 , n433514 );
or ( n434056 , n434054 , n434055 );
buf ( n434057 , n434056 );
buf ( n434058 , n434057 );
xor ( n434059 , n434052 , n434058 );
buf ( n434060 , n434059 );
buf ( n434061 , n434060 );
xor ( n434062 , n433539 , n433545 );
and ( n434063 , n434062 , n433623 );
and ( n434064 , n433539 , n433545 );
or ( n434065 , n434063 , n434064 );
buf ( n434066 , n434065 );
buf ( n434067 , n434066 );
xor ( n434068 , n434061 , n434067 );
buf ( n434069 , n384644 );
not ( n434070 , n434069 );
buf ( n434071 , n389928 );
not ( n434072 , n434071 );
buf ( n434073 , n395830 );
not ( n434074 , n434073 );
or ( n434075 , n434072 , n434074 );
buf ( n434076 , n390657 );
buf ( n434077 , n36252 );
nand ( n434078 , n434076 , n434077 );
buf ( n434079 , n434078 );
buf ( n434080 , n434079 );
nand ( n434081 , n434075 , n434080 );
buf ( n434082 , n434081 );
buf ( n434083 , n434082 );
not ( n434084 , n434083 );
or ( n434085 , n434070 , n434084 );
buf ( n434086 , n433560 );
buf ( n434087 , n383897 );
nand ( n434088 , n434086 , n434087 );
buf ( n434089 , n434088 );
buf ( n434090 , n434089 );
nand ( n434091 , n434085 , n434090 );
buf ( n434092 , n434091 );
and ( n434093 , n433583 , n389883 );
buf ( n434094 , n40758 );
not ( n434095 , n434094 );
buf ( n434096 , n42390 );
not ( n434097 , n434096 );
or ( n434098 , n434095 , n434097 );
buf ( n434099 , n37037 );
buf ( n434100 , n40971 );
nand ( n434101 , n434099 , n434100 );
buf ( n434102 , n434101 );
buf ( n434103 , n434102 );
nand ( n434104 , n434098 , n434103 );
buf ( n434105 , n434104 );
and ( n434106 , n434105 , n384554 );
nor ( n434107 , n434093 , n434106 );
xor ( n434108 , n434092 , n434107 );
not ( n434109 , n40901 );
not ( n434110 , n40890 );
not ( n434111 , n421471 );
or ( n434112 , n434110 , n434111 );
nand ( n434113 , n38630 , n40891 );
nand ( n434114 , n434112 , n434113 );
not ( n434115 , n434114 );
or ( n434116 , n434109 , n434115 );
nand ( n434117 , n433689 , n40858 );
nand ( n434118 , n434116 , n434117 );
buf ( n434119 , n434118 );
not ( n434120 , n434119 );
buf ( n434121 , n434120 );
and ( n434122 , n434108 , n434121 );
not ( n434123 , n434108 );
and ( n434124 , n434123 , n434118 );
nor ( n434125 , n434122 , n434124 );
buf ( n434126 , n433666 );
not ( n434127 , n434126 );
buf ( n434128 , n390260 );
not ( n434129 , n434128 );
or ( n434130 , n434127 , n434129 );
buf ( n434131 , n40972 );
not ( n434132 , n434131 );
buf ( n434133 , n41904 );
not ( n434134 , n434133 );
or ( n434135 , n434132 , n434134 );
buf ( n434136 , n388952 );
buf ( n434137 , n42799 );
nand ( n434138 , n434136 , n434137 );
buf ( n434139 , n434138 );
buf ( n434140 , n434139 );
nand ( n434141 , n434135 , n434140 );
buf ( n434142 , n434141 );
buf ( n434143 , n434142 );
buf ( n434144 , n388346 );
nand ( n434145 , n434143 , n434144 );
buf ( n434146 , n434145 );
buf ( n434147 , n434146 );
nand ( n434148 , n434130 , n434147 );
buf ( n434149 , n434148 );
buf ( n434150 , n434149 );
buf ( n434151 , n388549 );
not ( n434152 , n434151 );
buf ( n434153 , n384143 );
not ( n434154 , n434153 );
or ( n434155 , n434152 , n434154 );
buf ( n434156 , n385328 );
buf ( n434157 , n388546 );
nand ( n434158 , n434156 , n434157 );
buf ( n434159 , n434158 );
buf ( n434160 , n434159 );
nand ( n434161 , n434155 , n434160 );
buf ( n434162 , n434161 );
buf ( n434163 , n434162 );
not ( n434164 , n434163 );
buf ( n434165 , n434164 );
buf ( n434166 , n434165 );
buf ( n434167 , n389348 );
or ( n434168 , n434166 , n434167 );
nand ( n434169 , C1 , n434168 );
buf ( n434170 , n434169 );
buf ( n434171 , n434170 );
xor ( n434172 , n434150 , n434171 );
buf ( n434173 , n391782 );
not ( n434174 , n434173 );
buf ( n434175 , n434174 );
buf ( n434176 , n434175 );
buf ( n434177 , n433507 );
not ( n434178 , n434177 );
buf ( n434179 , n434178 );
buf ( n434180 , n434179 );
or ( n434181 , n434176 , n434180 );
buf ( n434182 , n389024 );
not ( n434183 , n434182 );
buf ( n434184 , n434183 );
buf ( n434185 , n434184 );
buf ( n434186 , n388376 );
not ( n434187 , n434186 );
buf ( n434188 , n385987 );
not ( n434189 , n434188 );
or ( n434190 , n434187 , n434189 );
buf ( n434191 , n397524 );
buf ( n434192 , n388373 );
nand ( n434193 , n434191 , n434192 );
buf ( n434194 , n434193 );
buf ( n434195 , n434194 );
nand ( n434196 , n434190 , n434195 );
buf ( n434197 , n434196 );
buf ( n434198 , n434197 );
not ( n434199 , n434198 );
buf ( n434200 , n434199 );
buf ( n434201 , n434200 );
or ( n434202 , n434185 , n434201 );
nand ( n434203 , n434181 , n434202 );
buf ( n434204 , n434203 );
buf ( n434205 , n434204 );
xor ( n434206 , n434172 , n434205 );
buf ( n434207 , n434206 );
buf ( n434208 , n434207 );
buf ( n434209 , n41565 );
not ( n434210 , n434209 );
buf ( n434211 , n24050 );
not ( n434212 , n434211 );
buf ( n434213 , n36900 );
not ( n434214 , n434213 );
or ( n434215 , n434212 , n434214 );
buf ( n434216 , n37381 );
buf ( n434217 , n389075 );
nand ( n434218 , n434216 , n434217 );
buf ( n434219 , n434218 );
buf ( n434220 , n434219 );
nand ( n434221 , n434215 , n434220 );
buf ( n434222 , n434221 );
buf ( n434223 , n434222 );
not ( n434224 , n434223 );
or ( n434225 , n434210 , n434224 );
buf ( n434226 , n433638 );
buf ( n434227 , n389125 );
nand ( n434228 , n434226 , n434227 );
buf ( n434229 , n434228 );
buf ( n434230 , n434229 );
nand ( n434231 , n434225 , n434230 );
buf ( n434232 , n434231 );
buf ( n434233 , n434232 );
xor ( n434234 , n434208 , n434233 );
buf ( n434235 , n434234 );
xor ( n434236 , n434125 , n434235 );
buf ( n434237 , n434236 );
not ( n434238 , n434237 );
buf ( n434239 , n434238 );
buf ( n434240 , n434239 );
xor ( n434241 , n434068 , n434240 );
buf ( n434242 , n434241 );
buf ( n434243 , n434242 );
xor ( n434244 , n434001 , n434243 );
buf ( n434245 , n434244 );
buf ( n434246 , n434245 );
xor ( n434247 , n433481 , n433487 );
and ( n434248 , n434247 , n433727 );
and ( n434249 , n433481 , n433487 );
or ( n434250 , n434248 , n434249 );
buf ( n434251 , n434250 );
buf ( n434252 , n434251 );
xor ( n434253 , n434246 , n434252 );
xor ( n434254 , n433283 , n433296 );
and ( n434255 , n434254 , n433458 );
and ( n434256 , n433283 , n433296 );
or ( n434257 , n434255 , n434256 );
buf ( n434258 , n434257 );
buf ( n434259 , n434258 );
xor ( n434260 , n434253 , n434259 );
buf ( n434261 , n434260 );
xnor ( n434262 , n433988 , n434261 );
not ( n434263 , n433739 );
nand ( n434264 , n434263 , n433461 );
buf ( n434265 , n433468 );
and ( n434266 , n434264 , n434265 );
not ( n434267 , n433739 );
nor ( n434268 , n434267 , n433461 );
nor ( n434269 , n434266 , n434268 );
nand ( n434270 , n434262 , n434269 );
buf ( n434271 , n434270 );
and ( n434272 , n433747 , n434271 );
buf ( n434273 , n434272 );
not ( n434274 , n433982 );
not ( n434275 , n434274 );
not ( n434276 , n433987 );
not ( n434277 , n434276 );
or ( n434278 , n434275 , n434277 );
nand ( n434279 , n434278 , n434261 );
nand ( n434280 , n433982 , n433987 );
nand ( n434281 , n434279 , n434280 );
xor ( n434282 , n433773 , n433787 );
and ( n434283 , n434282 , n433793 );
and ( n434284 , n433773 , n433787 );
or ( n434285 , n434283 , n434284 );
buf ( n434286 , n389162 );
not ( n434287 , n434286 );
buf ( n434288 , n434287 );
not ( n434289 , n434288 );
not ( n434290 , n41710 );
or ( n434291 , n434289 , n434290 );
nand ( n434292 , n434291 , n433783 );
not ( n434293 , n433809 );
not ( n434294 , n41374 );
and ( n434295 , n434293 , n434294 );
buf ( n434296 , n41342 );
not ( n434297 , n434296 );
buf ( n434298 , n382548 );
not ( n434299 , n434298 );
or ( n434300 , n434297 , n434299 );
buf ( n434301 , n398938 );
buf ( n434302 , n41349 );
nand ( n434303 , n434301 , n434302 );
buf ( n434304 , n434303 );
buf ( n434305 , n434304 );
nand ( n434306 , n434300 , n434305 );
buf ( n434307 , n434306 );
and ( n434308 , n434307 , n388833 );
nor ( n434309 , n434295 , n434308 );
and ( n434310 , n434292 , n434309 );
not ( n434311 , n434292 );
buf ( n434312 , n434309 );
not ( n434313 , n434312 );
buf ( n434314 , n434313 );
and ( n434315 , n434311 , n434314 );
or ( n434316 , n434310 , n434315 );
not ( n434317 , n38324 );
not ( n434318 , n385494 );
not ( n434319 , n383762 );
or ( n434320 , n434318 , n434319 );
buf ( n434321 , n42152 );
buf ( n434322 , n385491 );
nand ( n434323 , n434321 , n434322 );
buf ( n434324 , n434323 );
nand ( n434325 , n434320 , n434324 );
not ( n434326 , n434325 );
or ( n434327 , n434317 , n434326 );
not ( n434328 , n385482 );
nand ( n434329 , n434328 , n434043 );
nand ( n434330 , n434327 , n434329 );
and ( n434331 , n434316 , n434330 );
not ( n434332 , n434316 );
not ( n434333 , n434330 );
and ( n434334 , n434332 , n434333 );
nor ( n434335 , n434331 , n434334 );
xor ( n434336 , n434285 , n434335 );
not ( n434337 , n433846 );
not ( n434338 , n433817 );
or ( n434339 , n434337 , n434338 );
or ( n434340 , n433817 , n433846 );
nand ( n434341 , n434340 , n433823 );
nand ( n434342 , n434339 , n434341 );
xor ( n434343 , n434336 , n434342 );
buf ( n434344 , n434343 );
not ( n434345 , n433868 );
not ( n434346 , n433973 );
or ( n434347 , n434345 , n434346 );
nand ( n434348 , n434347 , n433873 );
buf ( n434349 , n434348 );
not ( n434350 , n433973 );
nand ( n434351 , n434350 , n433865 );
buf ( n434352 , n434351 );
nand ( n434353 , n434349 , n434352 );
buf ( n434354 , n434353 );
buf ( n434355 , n434354 );
xor ( n434356 , n434344 , n434355 );
xor ( n434357 , n433922 , n433949 );
and ( n434358 , n434357 , n433968 );
and ( n434359 , n433922 , n433949 );
or ( n434360 , n434358 , n434359 );
buf ( n434361 , n434360 );
buf ( n434362 , n434361 );
buf ( n434363 , n41565 );
not ( n434364 , n434363 );
buf ( n434365 , n24050 );
not ( n434366 , n434365 );
buf ( n434367 , n37369 );
not ( n434368 , n434367 );
or ( n434369 , n434366 , n434368 );
buf ( n434370 , n37370 );
buf ( n434371 , n389075 );
nand ( n434372 , n434370 , n434371 );
buf ( n434373 , n434372 );
buf ( n434374 , n434373 );
nand ( n434375 , n434369 , n434374 );
buf ( n434376 , n434375 );
buf ( n434377 , n434376 );
not ( n434378 , n434377 );
or ( n434379 , n434364 , n434378 );
buf ( n434380 , n434222 );
buf ( n434381 , n389125 );
nand ( n434382 , n434380 , n434381 );
buf ( n434383 , n434382 );
buf ( n434384 , n434383 );
nand ( n434385 , n434379 , n434384 );
buf ( n434386 , n434385 );
buf ( n434387 , n434386 );
xor ( n434388 , n434362 , n434387 );
buf ( n434389 , n433915 );
not ( n434390 , n434389 );
buf ( n434391 , n383017 );
not ( n434392 , n434391 );
or ( n434393 , n434390 , n434392 );
buf ( n434394 , n390635 );
buf ( n434395 , n388646 );
not ( n434396 , n434395 );
buf ( n434397 , n398740 );
not ( n434398 , n434397 );
or ( n434399 , n434396 , n434398 );
buf ( n434400 , n433606 );
buf ( n434401 , n388654 );
nand ( n434402 , n434400 , n434401 );
buf ( n434403 , n434402 );
buf ( n434404 , n434403 );
nand ( n434405 , n434399 , n434404 );
buf ( n434406 , n434405 );
buf ( n434407 , n434406 );
nand ( n434408 , n434394 , n434407 );
buf ( n434409 , n434408 );
buf ( n434410 , n434409 );
nand ( n434411 , n434393 , n434410 );
buf ( n434412 , n434411 );
buf ( n434413 , n434105 );
not ( n434414 , n434413 );
buf ( n434415 , n384627 );
not ( n434416 , n434415 );
or ( n434417 , n434414 , n434416 );
buf ( n434418 , n390271 );
buf ( n434419 , n390498 );
and ( n434420 , n434418 , n434419 );
not ( n434421 , n434418 );
buf ( n434422 , n391129 );
and ( n434423 , n434421 , n434422 );
nor ( n434424 , n434420 , n434423 );
buf ( n434425 , n434424 );
buf ( n434426 , n434425 );
not ( n434427 , n434426 );
buf ( n434428 , n389908 );
nand ( n434429 , n434427 , n434428 );
buf ( n434430 , n434429 );
buf ( n434431 , n434430 );
nand ( n434432 , n434417 , n434431 );
buf ( n434433 , n434432 );
not ( n434434 , n434433 );
xor ( n434435 , n434412 , n434434 );
buf ( n434436 , n37695 );
not ( n434437 , n434436 );
buf ( n434438 , n37347 );
not ( n434439 , n434438 );
buf ( n434440 , n385734 );
not ( n434441 , n434440 );
or ( n434442 , n434439 , n434441 );
buf ( n434443 , n384186 );
buf ( n434444 , n391895 );
nand ( n434445 , n434443 , n434444 );
buf ( n434446 , n434445 );
buf ( n434447 , n434446 );
nand ( n434448 , n434442 , n434447 );
buf ( n434449 , n434448 );
buf ( n434450 , n434449 );
not ( n434451 , n434450 );
or ( n434452 , n434437 , n434451 );
buf ( n434453 , n434018 );
buf ( n434454 , n385269 );
nand ( n434455 , n434453 , n434454 );
buf ( n434456 , n434455 );
buf ( n434457 , n434456 );
nand ( n434458 , n434452 , n434457 );
buf ( n434459 , n434458 );
xnor ( n434460 , n434435 , n434459 );
buf ( n434461 , n434460 );
xor ( n434462 , n434388 , n434461 );
buf ( n434463 , n434462 );
buf ( n434464 , n434463 );
xor ( n434465 , n434026 , n434051 );
and ( n434466 , n434465 , n434058 );
and ( n434467 , n434026 , n434051 );
or ( n434468 , n434466 , n434467 );
buf ( n434469 , n434468 );
not ( n434470 , n434469 );
not ( n434471 , n434470 );
buf ( n434472 , n390403 );
not ( n434473 , n434472 );
and ( n434474 , n35301 , n24073 );
not ( n434475 , n35301 );
and ( n434476 , n434475 , n24074 );
or ( n434477 , n434474 , n434476 );
buf ( n434478 , n434477 );
not ( n434479 , n434478 );
or ( n434480 , n434473 , n434479 );
buf ( n434481 , n433839 );
buf ( n434482 , n391080 );
nand ( n434483 , n434481 , n434482 );
buf ( n434484 , n434483 );
buf ( n434485 , n434484 );
nand ( n434486 , n434480 , n434485 );
buf ( n434487 , n434486 );
not ( n434488 , n434487 );
or ( n434489 , n434471 , n434488 );
not ( n434490 , n434487 );
nand ( n434491 , n434490 , n434469 );
nand ( n434492 , n434489 , n434491 );
buf ( n434493 , n40701 );
not ( n434494 , n434493 );
buf ( n434495 , n433894 );
not ( n434496 , n434495 );
or ( n434497 , n434494 , n434496 );
not ( n434498 , n388160 );
not ( n434499 , n386424 );
or ( n434500 , n434498 , n434499 );
not ( n434501 , n388771 );
nand ( n434502 , n434501 , n388157 );
nand ( n434503 , n434500 , n434502 );
buf ( n434504 , n434503 );
buf ( n434505 , n388141 );
nand ( n434506 , n434504 , n434505 );
buf ( n434507 , n434506 );
buf ( n434508 , n434507 );
nand ( n434509 , n434497 , n434508 );
buf ( n434510 , n434509 );
and ( n434511 , n434492 , n434510 );
not ( n434512 , n434492 );
not ( n434513 , n434510 );
and ( n434514 , n434512 , n434513 );
nor ( n434515 , n434511 , n434514 );
buf ( n434516 , n434515 );
xor ( n434517 , n434464 , n434516 );
not ( n434518 , n433896 );
not ( n434519 , n433970 );
or ( n434520 , n434518 , n434519 );
not ( n434521 , n433890 );
and ( n434522 , n433897 , n433971 );
or ( n434523 , n434521 , n434522 );
nand ( n434524 , n434520 , n434523 );
buf ( n434525 , n434524 );
xor ( n434526 , n434517 , n434525 );
buf ( n434527 , n434526 );
buf ( n434528 , n434527 );
xor ( n434529 , n434356 , n434528 );
buf ( n434530 , n434529 );
xor ( n434531 , n434246 , n434252 );
and ( n434532 , n434531 , n434259 );
and ( n434533 , n434246 , n434252 );
or ( n434534 , n434532 , n434533 );
buf ( n434535 , n434534 );
xor ( n434536 , n434530 , n434535 );
xor ( n434537 , n433994 , n434000 );
and ( n434538 , n434537 , n434243 );
and ( n434539 , n433994 , n434000 );
or ( n434540 , n434538 , n434539 );
buf ( n434541 , n434540 );
not ( n434542 , n434541 );
buf ( n434543 , n434060 );
not ( n434544 , n434543 );
buf ( n434545 , n434544 );
buf ( n434546 , n434545 );
not ( n434547 , n434546 );
buf ( n434548 , n434236 );
not ( n434549 , n434548 );
or ( n434550 , n434547 , n434549 );
buf ( n434551 , n434066 );
nand ( n434552 , n434550 , n434551 );
buf ( n434553 , n434552 );
buf ( n434554 , n434553 );
buf ( n434555 , n434239 );
buf ( n434556 , n434060 );
nand ( n434557 , n434555 , n434556 );
buf ( n434558 , n434557 );
buf ( n434559 , n434558 );
nand ( n434560 , n434554 , n434559 );
buf ( n434561 , n434560 );
buf ( n434562 , n434561 );
buf ( n434563 , n433849 );
buf ( n434564 , n433794 );
buf ( n434565 , n433752 );
nor ( n434566 , n434564 , n434565 );
buf ( n434567 , n434566 );
buf ( n434568 , n434567 );
or ( n434569 , n434563 , n434568 );
buf ( n434570 , n433794 );
buf ( n434571 , n433752 );
nand ( n434572 , n434570 , n434571 );
buf ( n434573 , n434572 );
buf ( n434574 , n434573 );
nand ( n434575 , n434569 , n434574 );
buf ( n434576 , n434575 );
buf ( n434577 , n434576 );
xor ( n434578 , n434562 , n434577 );
buf ( n434579 , n384644 );
not ( n434580 , n434579 );
buf ( n434581 , n36252 );
not ( n434582 , n434581 );
buf ( n434583 , n434582 );
buf ( n434584 , n434583 );
not ( n434585 , n434584 );
buf ( n434586 , n390172 );
not ( n434587 , n434586 );
or ( n434588 , n434585 , n434587 );
buf ( n434589 , n384974 );
buf ( n434590 , n36252 );
nand ( n434591 , n434589 , n434590 );
buf ( n434592 , n434591 );
buf ( n434593 , n434592 );
nand ( n434594 , n434588 , n434593 );
buf ( n434595 , n434594 );
buf ( n434596 , n434595 );
not ( n434597 , n434596 );
or ( n434598 , n434580 , n434597 );
buf ( n434599 , n434082 );
buf ( n434600 , n383897 );
nand ( n434601 , n434599 , n434600 );
buf ( n434602 , n434601 );
buf ( n434603 , n434602 );
nand ( n434604 , n434598 , n434603 );
buf ( n434605 , n434604 );
xor ( n434606 , n434150 , n434171 );
and ( n434607 , n434606 , n434205 );
and ( n434608 , n434150 , n434171 );
or ( n434609 , n434607 , n434608 );
buf ( n434610 , n434609 );
xor ( n434611 , n434605 , n434610 );
not ( n434612 , n434092 );
not ( n434613 , n434121 );
or ( n434614 , n434612 , n434613 );
buf ( n434615 , n434092 );
buf ( n434616 , n434121 );
nor ( n434617 , n434615 , n434616 );
buf ( n434618 , n434617 );
or ( n434619 , n434618 , n434107 );
nand ( n434620 , n434614 , n434619 );
xor ( n434621 , n434611 , n434620 );
buf ( n434622 , n434125 );
not ( n434623 , n434622 );
buf ( n434624 , n434623 );
not ( n434625 , n434624 );
buf ( n434626 , n434207 );
buf ( n434627 , n434232 );
or ( n434628 , n434626 , n434627 );
buf ( n434629 , n434628 );
not ( n434630 , n434629 );
or ( n434631 , n434625 , n434630 );
and ( n434632 , n434208 , n434233 );
buf ( n434633 , n434632 );
not ( n434634 , n434633 );
nand ( n434635 , n434631 , n434634 );
xor ( n434636 , n434621 , n434635 );
buf ( n434637 , n40840 );
buf ( n434638 , n434637 );
not ( n434639 , n434638 );
buf ( n434640 , n41896 );
not ( n434641 , n434640 );
or ( n434642 , n434639 , n434641 );
buf ( n434643 , n38155 );
buf ( n434644 , n40835 );
nand ( n434645 , n434643 , n434644 );
buf ( n434646 , n434645 );
buf ( n434647 , n434646 );
nand ( n434648 , n434642 , n434647 );
buf ( n434649 , n434648 );
buf ( n434650 , n434649 );
buf ( n434651 , n383946 );
and ( n434652 , n434650 , n434651 );
buf ( n434653 , n388460 );
buf ( n434654 , n434142 );
and ( n434655 , n434653 , n434654 );
buf ( n434656 , n434655 );
buf ( n434657 , n434656 );
nor ( n434658 , n434652 , n434657 );
buf ( n434659 , n434658 );
buf ( n434660 , n434659 );
not ( n434661 , n434660 );
buf ( n434662 , n434661 );
xor ( n434663 , n434121 , n434662 );
buf ( n434664 , n391164 );
buf ( n434665 , n433940 );
or ( n434666 , n434664 , n434665 );
buf ( n434667 , n391176 );
buf ( n434668 , n27196 );
buf ( n434669 , n389598 );
and ( n434670 , n434668 , n434669 );
not ( n434671 , n434668 );
buf ( n434672 , n388556 );
and ( n434673 , n434671 , n434672 );
nor ( n434674 , n434670 , n434673 );
buf ( n434675 , n434674 );
buf ( n434676 , n434675 );
or ( n434677 , n434667 , n434676 );
nand ( n434678 , n434666 , n434677 );
buf ( n434679 , n434678 );
not ( n434680 , n434679 );
xnor ( n434681 , n434663 , n434680 );
not ( n434682 , n434681 );
not ( n434683 , n386480 );
buf ( n434684 , n38972 );
not ( n434685 , n434684 );
buf ( n434686 , n37147 );
not ( n434687 , n434686 );
or ( n434688 , n434685 , n434687 );
buf ( n434689 , n394463 );
buf ( n434690 , n38971 );
nand ( n434691 , n434689 , n434690 );
buf ( n434692 , n434691 );
buf ( n434693 , n434692 );
nand ( n434694 , n434688 , n434693 );
buf ( n434695 , n434694 );
not ( n434696 , n434695 );
or ( n434697 , n434683 , n434696 );
buf ( n434698 , n433767 );
buf ( n434699 , n386496 );
nand ( n434700 , n434698 , n434699 );
buf ( n434701 , n434700 );
nand ( n434702 , n434697 , n434701 );
not ( n434703 , n434702 );
not ( n434704 , n434703 );
buf ( n434705 , n434197 );
not ( n434706 , n434705 );
buf ( n434707 , n391782 );
not ( n434708 , n434707 );
or ( n434709 , n434706 , n434708 );
not ( n434710 , n44399 );
not ( n434711 , n382994 );
or ( n434712 , n434710 , n434711 );
buf ( n434713 , n389759 );
buf ( n434714 , n41195 );
nand ( n434715 , n434713 , n434714 );
buf ( n434716 , n434715 );
nand ( n434717 , n434712 , n434716 );
nand ( n434718 , n379463 , n434717 );
buf ( n434719 , n434718 );
nand ( n434720 , n434709 , n434719 );
buf ( n434721 , n434720 );
not ( n434722 , n40858 );
not ( n434723 , n434114 );
or ( n434724 , n434722 , n434723 );
not ( n434725 , n385342 );
not ( n434726 , n40890 );
or ( n434727 , n434725 , n434726 );
nand ( n434728 , n385356 , n40891 );
nand ( n434729 , n434727 , n434728 );
buf ( n434730 , n434729 );
buf ( n434731 , n384413 );
nand ( n434732 , n434730 , n434731 );
buf ( n434733 , n434732 );
nand ( n434734 , n434724 , n434733 );
buf ( n434735 , n434734 );
xor ( n434736 , n434721 , n434735 );
buf ( n434737 , n389547 );
buf ( n434738 , n390490 );
not ( n434739 , n434738 );
buf ( n434740 , n384096 );
not ( n434741 , n434740 );
or ( n434742 , n434739 , n434741 );
buf ( n434743 , n385292 );
buf ( n434744 , n388569 );
nand ( n434745 , n434743 , n434744 );
buf ( n434746 , n434745 );
buf ( n434747 , n434746 );
nand ( n434748 , n434742 , n434747 );
buf ( n434749 , n434748 );
buf ( n434750 , n434749 );
nand ( n434751 , n434737 , n434750 );
buf ( n434752 , n434751 );
buf ( n434753 , n434752 );
nand ( n434754 , C1 , n434753 );
buf ( n434755 , n434754 );
buf ( n434756 , n434755 );
xor ( n434757 , n434736 , n434756 );
not ( n434758 , n434757 );
or ( n434759 , n434704 , n434758 );
buf ( n434760 , n434721 );
not ( n434761 , n434760 );
xnor ( n434762 , n434735 , n434756 );
not ( n434763 , n434762 );
or ( n434764 , n434761 , n434763 );
or ( n434765 , n434760 , n434762 );
nand ( n434766 , n434764 , n434765 );
or ( n434767 , n434766 , n434703 );
nand ( n434768 , n434759 , n434767 );
not ( n434769 , n434768 );
or ( n434770 , n434682 , n434769 );
and ( n434771 , n434118 , n434659 );
not ( n434772 , n434118 );
and ( n434773 , n434772 , n434662 );
nor ( n434774 , n434771 , n434773 );
not ( n434775 , n434680 );
and ( n434776 , n434774 , n434775 );
not ( n434777 , n434774 );
and ( n434778 , n434777 , n434680 );
nor ( n434779 , n434776 , n434778 );
or ( n434780 , n434779 , n434768 );
nand ( n434781 , n434770 , n434780 );
not ( n434782 , n434781 );
xnor ( n434783 , n434636 , n434782 );
buf ( n434784 , n434783 );
xor ( n434785 , n434578 , n434784 );
buf ( n434786 , n434785 );
not ( n434787 , n434786 );
not ( n434788 , n434787 );
or ( n434789 , n434542 , n434788 );
not ( n434790 , n434541 );
nand ( n434791 , n434786 , n434790 );
nand ( n434792 , n434789 , n434791 );
xor ( n434793 , n433853 , n433859 );
and ( n434794 , n434793 , n433980 );
and ( n434795 , n433853 , n433859 );
or ( n434796 , n434794 , n434795 );
buf ( n434797 , n434796 );
and ( n434798 , n434792 , n434797 );
not ( n434799 , n434792 );
not ( n434800 , n434797 );
and ( n434801 , n434799 , n434800 );
nor ( n434802 , n434798 , n434801 );
xor ( n434803 , n434536 , n434802 );
nor ( n434804 , n434281 , n434803 );
buf ( n434805 , n434729 );
not ( n434806 , n434805 );
buf ( n434807 , n36801 );
not ( n434808 , n434807 );
or ( n434809 , n434806 , n434808 );
buf ( n434810 , n390929 );
buf ( n434811 , n385324 );
and ( n434812 , n434810 , n434811 );
not ( n434813 , n434810 );
buf ( n434814 , n389964 );
and ( n434815 , n434813 , n434814 );
nor ( n434816 , n434812 , n434815 );
buf ( n434817 , n434816 );
buf ( n434818 , n434817 );
buf ( n434819 , n392111 );
nand ( n434820 , n434818 , n434819 );
buf ( n434821 , n434820 );
buf ( n434822 , n434821 );
nand ( n434823 , n434809 , n434822 );
buf ( n434824 , n434823 );
not ( n434825 , n40840 );
nand ( n434826 , n434825 , n390651 );
nand ( n434827 , n40840 , n36509 );
nand ( n434828 , n434826 , n434827 );
buf ( n434829 , n434828 );
not ( n434830 , n434829 );
buf ( n434831 , n388349 );
not ( n434832 , n434831 );
and ( n434833 , n434830 , n434832 );
buf ( n434834 , n434649 );
buf ( n434835 , n388460 );
and ( n434836 , n434834 , n434835 );
nor ( n434837 , n434833 , n434836 );
buf ( n434838 , n434837 );
buf ( n434839 , n434838 );
not ( n434840 , n434839 );
buf ( n434841 , n434840 );
xor ( n434842 , n434824 , n434841 );
not ( n434843 , n389024 );
buf ( n434844 , n40819 );
not ( n434845 , n434844 );
buf ( n434846 , n385972 );
not ( n434847 , n434846 );
or ( n434848 , n434845 , n434847 );
buf ( n434849 , n388445 );
buf ( n434850 , n397524 );
nand ( n434851 , n434849 , n434850 );
buf ( n434852 , n434851 );
buf ( n434853 , n434852 );
nand ( n434854 , n434848 , n434853 );
buf ( n434855 , n434854 );
not ( n434856 , n434855 );
or ( n434857 , n434843 , n434856 );
nand ( n434858 , n382598 , n434717 );
nand ( n434859 , n434857 , n434858 );
xnor ( n434860 , n434842 , n434859 );
not ( n434861 , n434860 );
not ( n434862 , n434861 );
buf ( n434863 , n388872 );
not ( n434864 , n434863 );
buf ( n434865 , n434307 );
not ( n434866 , n434865 );
or ( n434867 , n434864 , n434866 );
buf ( n434868 , n388833 );
not ( n434869 , n434868 );
buf ( n434870 , n434869 );
buf ( n434871 , n434870 );
not ( n434872 , n434871 );
buf ( n434873 , n41342 );
not ( n434874 , n434873 );
buf ( n434875 , n385502 );
not ( n434876 , n434875 );
or ( n434877 , n434874 , n434876 );
buf ( n434878 , n385499 );
buf ( n434879 , n41349 );
nand ( n434880 , n434878 , n434879 );
buf ( n434881 , n434880 );
buf ( n434882 , n434881 );
nand ( n434883 , n434877 , n434882 );
buf ( n434884 , n434883 );
buf ( n434885 , n434884 );
nand ( n434886 , n434872 , n434885 );
buf ( n434887 , n434886 );
buf ( n434888 , n434887 );
nand ( n434889 , n434867 , n434888 );
buf ( n434890 , n434889 );
buf ( n434891 , n434890 );
not ( n434892 , n434891 );
buf ( n434893 , n434892 );
not ( n434894 , n434893 );
or ( n434895 , n434862 , n434894 );
buf ( n434896 , n434890 );
buf ( n434897 , n434860 );
nand ( n434898 , n434896 , n434897 );
buf ( n434899 , n434898 );
nand ( n434900 , n434895 , n434899 );
buf ( n434901 , n384621 );
buf ( n434902 , n434425 );
or ( n434903 , n434901 , n434902 );
buf ( n434904 , n391635 );
buf ( n434905 , n395885 );
not ( n434906 , n434905 );
buf ( n434907 , n38631 );
not ( n434908 , n434907 );
and ( n434909 , n434906 , n434908 );
buf ( n434910 , n390498 );
buf ( n434911 , n386182 );
and ( n434912 , n434910 , n434911 );
nor ( n434913 , n434909 , n434912 );
buf ( n434914 , n434913 );
buf ( n434915 , n434914 );
or ( n434916 , n434904 , n434915 );
nand ( n434917 , n434903 , n434916 );
buf ( n434918 , n434917 );
buf ( n434919 , n434406 );
not ( n434920 , n434919 );
buf ( n434921 , n396868 );
not ( n434922 , n434921 );
or ( n434923 , n434920 , n434922 );
buf ( n434924 , n390476 );
buf ( n434925 , n388376 );
not ( n434926 , n434925 );
buf ( n434927 , n37402 );
not ( n434928 , n434927 );
or ( n434929 , n434926 , n434928 );
buf ( n434930 , n35435 );
buf ( n434931 , n388373 );
nand ( n434932 , n434930 , n434931 );
buf ( n434933 , n434932 );
buf ( n434934 , n434933 );
nand ( n434935 , n434929 , n434934 );
buf ( n434936 , n434935 );
buf ( n434937 , n434936 );
nand ( n434938 , n434924 , n434937 );
buf ( n434939 , n434938 );
buf ( n434940 , n434939 );
nand ( n434941 , n434923 , n434940 );
buf ( n434942 , n434941 );
xor ( n434943 , n434918 , n434942 );
not ( n434944 , n434675 );
not ( n434945 , n434944 );
not ( n434946 , n391652 );
or ( n434947 , n434945 , n434946 );
buf ( n434948 , n40971 );
buf ( n434949 , n395919 );
not ( n434950 , n434949 );
buf ( n434951 , n434950 );
buf ( n434952 , n434951 );
and ( n434953 , n434948 , n434952 );
not ( n434954 , n434948 );
buf ( n434955 , n385633 );
and ( n434956 , n434954 , n434955 );
nor ( n434957 , n434953 , n434956 );
buf ( n434958 , n434957 );
or ( n434959 , n383403 , n434958 );
nand ( n434960 , n434947 , n434959 );
xor ( n434961 , n434943 , n434960 );
and ( n434962 , n434900 , n434961 );
not ( n434963 , n434900 );
buf ( n434964 , n434961 );
not ( n434965 , n434964 );
buf ( n434966 , n434965 );
and ( n434967 , n434963 , n434966 );
nor ( n434968 , n434962 , n434967 );
buf ( n434969 , n434118 );
not ( n434970 , n434969 );
buf ( n434971 , n434662 );
not ( n434972 , n434971 );
or ( n434973 , n434970 , n434972 );
buf ( n434974 , n434121 );
not ( n434975 , n434974 );
buf ( n434976 , n434659 );
not ( n434977 , n434976 );
or ( n434978 , n434975 , n434977 );
buf ( n434979 , n434679 );
nand ( n434980 , n434978 , n434979 );
buf ( n434981 , n434980 );
buf ( n434982 , n434981 );
nand ( n434983 , n434973 , n434982 );
buf ( n434984 , n434983 );
buf ( n434985 , n434984 );
buf ( n434986 , n37695 );
not ( n434987 , n434986 );
and ( n434988 , n36216 , n391895 );
not ( n434989 , n36216 );
and ( n434990 , n434989 , n37347 );
or ( n434991 , n434988 , n434990 );
buf ( n434992 , n434991 );
not ( n434993 , n434992 );
or ( n434994 , n434987 , n434993 );
buf ( n434995 , n434449 );
buf ( n434996 , n385269 );
nand ( n434997 , n434995 , n434996 );
buf ( n434998 , n434997 );
buf ( n434999 , n434998 );
nand ( n435000 , n434994 , n434999 );
buf ( n435001 , n435000 );
buf ( n435002 , n435001 );
not ( n435003 , n435002 );
buf ( n435004 , n435003 );
buf ( n435005 , n435004 );
and ( n435006 , n434985 , n435005 );
not ( n435007 , n434985 );
buf ( n435008 , n435001 );
and ( n435009 , n435007 , n435008 );
nor ( n435010 , n435006 , n435009 );
buf ( n435011 , n435010 );
buf ( n435012 , n386496 );
not ( n435013 , n435012 );
buf ( n435014 , n434695 );
not ( n435015 , n435014 );
or ( n435016 , n435013 , n435015 );
buf ( n435017 , n38972 );
not ( n435018 , n435017 );
buf ( n435019 , n403567 );
not ( n435020 , n435019 );
or ( n435021 , n435018 , n435020 );
buf ( n435022 , n396298 );
buf ( n435023 , n38971 );
nand ( n435024 , n435022 , n435023 );
buf ( n435025 , n435024 );
buf ( n435026 , n435025 );
nand ( n435027 , n435021 , n435026 );
buf ( n435028 , n435027 );
buf ( n435029 , n435028 );
buf ( n435030 , n386480 );
nand ( n435031 , n435029 , n435030 );
buf ( n435032 , n435031 );
buf ( n435033 , n435032 );
nand ( n435034 , n435016 , n435033 );
buf ( n435035 , n435034 );
and ( n435036 , n435011 , n435035 );
not ( n435037 , n435011 );
buf ( n435038 , n435035 );
not ( n435039 , n435038 );
buf ( n435040 , n435039 );
and ( n435041 , n435037 , n435040 );
or ( n435042 , n435036 , n435041 );
not ( n435043 , n435042 );
xor ( n435044 , n434968 , n435043 );
xor ( n435045 , n434362 , n434387 );
and ( n435046 , n435045 , n434461 );
and ( n435047 , n434362 , n434387 );
or ( n435048 , n435046 , n435047 );
buf ( n435049 , n435048 );
not ( n435050 , n435049 );
xor ( n435051 , n435044 , n435050 );
xor ( n435052 , n434464 , n434516 );
and ( n435053 , n435052 , n434525 );
and ( n435054 , n434464 , n434516 );
or ( n435055 , n435053 , n435054 );
buf ( n435056 , n435055 );
not ( n435057 , n435056 );
xor ( n435058 , n435051 , n435057 );
not ( n435059 , n385889 );
not ( n435060 , n434325 );
or ( n435061 , n435059 , n435060 );
buf ( n435062 , n385494 );
not ( n435063 , n435062 );
buf ( n435064 , n389525 );
not ( n435065 , n435064 );
or ( n435066 , n435063 , n435065 );
nand ( n435067 , n37173 , n385491 );
buf ( n435068 , n435067 );
nand ( n435069 , n435066 , n435068 );
buf ( n435070 , n435069 );
buf ( n435071 , n435070 );
buf ( n435072 , n38324 );
nand ( n435073 , n435071 , n435072 );
buf ( n435074 , n435073 );
nand ( n435075 , n435061 , n435074 );
not ( n435076 , n435075 );
not ( n435077 , n434412 );
nand ( n435078 , n435077 , n434434 );
not ( n435079 , n435078 );
not ( n435080 , n434459 );
or ( n435081 , n435079 , n435080 );
nand ( n435082 , n434433 , n434412 );
nand ( n435083 , n435081 , n435082 );
xor ( n435084 , n435076 , n435083 );
not ( n435085 , n434376 );
not ( n435086 , n389125 );
or ( n435087 , n435085 , n435086 );
buf ( n435088 , n24050 );
not ( n435089 , n435088 );
buf ( n435090 , n383575 );
not ( n435091 , n435090 );
or ( n435092 , n435089 , n435091 );
buf ( n435093 , n385834 );
buf ( n435094 , n389075 );
nand ( n435095 , n435093 , n435094 );
buf ( n435096 , n435095 );
buf ( n435097 , n435096 );
nand ( n435098 , n435092 , n435097 );
buf ( n435099 , n435098 );
buf ( n435100 , n435099 );
buf ( n435101 , n41565 );
nand ( n435102 , n435100 , n435101 );
buf ( n435103 , n435102 );
nand ( n435104 , n435087 , n435103 );
xnor ( n435105 , n435084 , n435104 );
not ( n435106 , n435105 );
not ( n435107 , n435106 );
not ( n435108 , n434510 );
not ( n435109 , n434469 );
nand ( n435110 , n435109 , n434490 );
not ( n435111 , n435110 );
or ( n435112 , n435108 , n435111 );
not ( n435113 , n434470 );
nand ( n435114 , n435113 , n434487 );
nand ( n435115 , n435112 , n435114 );
not ( n435116 , n435115 );
not ( n435117 , n435116 );
or ( n435118 , n435107 , n435117 );
or ( n435119 , n435116 , n435106 );
nand ( n435120 , n435118 , n435119 );
not ( n435121 , n435120 );
buf ( n435122 , n434781 );
buf ( n435123 , n434621 );
buf ( n435124 , n435123 );
or ( n435125 , n435122 , n435124 );
buf ( n435126 , n434635 );
nand ( n435127 , n435125 , n435126 );
buf ( n435128 , n435127 );
buf ( n435129 , n434781 );
buf ( n435130 , n435123 );
nand ( n435131 , n435129 , n435130 );
buf ( n435132 , n435131 );
nand ( n435133 , n435128 , n435132 );
buf ( n435134 , n435133 );
not ( n435135 , n435134 );
or ( n435136 , n435121 , n435135 );
or ( n435137 , n435134 , n435120 );
nand ( n435138 , n435136 , n435137 );
xnor ( n435139 , n435058 , n435138 );
buf ( n435140 , n435139 );
xor ( n435141 , n434562 , n434577 );
and ( n435142 , n435141 , n434784 );
and ( n435143 , n434562 , n434577 );
or ( n435144 , n435142 , n435143 );
buf ( n435145 , n435144 );
buf ( n435146 , n435145 );
buf ( n435147 , n40701 );
not ( n435148 , n435147 );
buf ( n435149 , n434503 );
not ( n435150 , n435149 );
or ( n435151 , n435148 , n435150 );
buf ( n435152 , n388160 );
not ( n435153 , n435152 );
buf ( n435154 , n38532 );
not ( n435155 , n435154 );
or ( n435156 , n435153 , n435155 );
buf ( n435157 , n35519 );
buf ( n435158 , n388157 );
nand ( n435159 , n435157 , n435158 );
buf ( n435160 , n435159 );
buf ( n435161 , n435160 );
nand ( n435162 , n435156 , n435161 );
buf ( n435163 , n435162 );
buf ( n435164 , n435163 );
buf ( n435165 , n388141 );
nand ( n435166 , n435164 , n435165 );
buf ( n435167 , n435166 );
buf ( n435168 , n435167 );
nand ( n435169 , n435151 , n435168 );
buf ( n435170 , n435169 );
buf ( n435171 , n391080 );
not ( n435172 , n435171 );
buf ( n435173 , n434477 );
not ( n435174 , n435173 );
or ( n435175 , n435172 , n435174 );
and ( n435176 , n382921 , n24073 );
not ( n435177 , n382921 );
and ( n435178 , n435177 , n24074 );
or ( n435179 , n435176 , n435178 );
buf ( n435180 , n435179 );
buf ( n435181 , n390403 );
nand ( n435182 , n435180 , n435181 );
buf ( n435183 , n435182 );
buf ( n435184 , n435183 );
nand ( n435185 , n435175 , n435184 );
buf ( n435186 , n435185 );
not ( n435187 , n435186 );
xor ( n435188 , n435170 , n435187 );
xor ( n435189 , n434605 , n434610 );
and ( n435190 , n435189 , n434620 );
and ( n435191 , n434605 , n434610 );
or ( n435192 , n435190 , n435191 );
not ( n435193 , n435192 );
xor ( n435194 , n435188 , n435193 );
buf ( n435195 , n435194 );
buf ( n435196 , n385292 );
not ( n435197 , n435196 );
buf ( n435198 , n389859 );
not ( n435199 , n435198 );
and ( n435200 , n435197 , n435199 );
buf ( n435201 , n382854 );
buf ( n435202 , n389859 );
and ( n435203 , n435201 , n435202 );
nor ( n435204 , n435200 , n435203 );
buf ( n435205 , n435204 );
not ( n435206 , n435205 );
and ( n435207 , n382947 , n435206 );
nor ( n435208 , C0 , n435207 );
buf ( n435209 , n435208 );
buf ( n435210 , n383897 );
not ( n435211 , n435210 );
buf ( n435212 , n434595 );
not ( n435213 , n435212 );
or ( n435214 , n435211 , n435213 );
not ( n435215 , n434583 );
not ( n435216 , n397419 );
or ( n435217 , n435215 , n435216 );
buf ( n435218 , n389928 );
not ( n435219 , n435218 );
buf ( n435220 , n38472 );
nand ( n435221 , n435219 , n435220 );
buf ( n435222 , n435221 );
nand ( n435223 , n435217 , n435222 );
nand ( n435224 , n435223 , n384644 );
buf ( n435225 , n435224 );
nand ( n435226 , n435214 , n435225 );
buf ( n435227 , n435226 );
buf ( n435228 , n435227 );
xor ( n435229 , n435209 , n435228 );
buf ( n435230 , n434734 );
not ( n435231 , n435230 );
buf ( n435232 , n434755 );
not ( n435233 , n435232 );
or ( n435234 , n435231 , n435233 );
buf ( n435235 , n434755 );
buf ( n435236 , n434734 );
or ( n435237 , n435235 , n435236 );
buf ( n435238 , n434721 );
nand ( n435239 , n435237 , n435238 );
buf ( n435240 , n435239 );
buf ( n435241 , n435240 );
nand ( n435242 , n435234 , n435241 );
buf ( n435243 , n435242 );
buf ( n435244 , n435243 );
xor ( n435245 , n435229 , n435244 );
buf ( n435246 , n435245 );
buf ( n435247 , n434333 );
not ( n435248 , n435247 );
buf ( n435249 , n434309 );
not ( n435250 , n435249 );
or ( n435251 , n435248 , n435250 );
buf ( n435252 , n434292 );
nand ( n435253 , n435251 , n435252 );
buf ( n435254 , n435253 );
buf ( n435255 , n435254 );
buf ( n435256 , n434314 );
buf ( n435257 , n434330 );
nand ( n435258 , n435256 , n435257 );
buf ( n435259 , n435258 );
buf ( n435260 , n435259 );
nand ( n435261 , n435255 , n435260 );
buf ( n435262 , n435261 );
xor ( n435263 , n435246 , n435262 );
buf ( n435264 , n435263 );
nand ( n435265 , n434779 , n434703 );
and ( n435266 , n435265 , n434766 );
nor ( n435267 , n434779 , n434703 );
nor ( n435268 , n435266 , n435267 );
buf ( n435269 , n435268 );
xnor ( n435270 , n435264 , n435269 );
buf ( n435271 , n435270 );
buf ( n435272 , n435271 );
xor ( n435273 , n435195 , n435272 );
xor ( n435274 , n434285 , n434335 );
and ( n435275 , n435274 , n434342 );
and ( n435276 , n434285 , n434335 );
or ( n435277 , n435275 , n435276 );
buf ( n435278 , n435277 );
xor ( n435279 , n435273 , n435278 );
buf ( n435280 , n435279 );
buf ( n435281 , n435280 );
xor ( n435282 , n435146 , n435281 );
xor ( n435283 , n434344 , n434355 );
and ( n435284 , n435283 , n434528 );
and ( n435285 , n434344 , n434355 );
or ( n435286 , n435284 , n435285 );
buf ( n435287 , n435286 );
buf ( n435288 , n435287 );
xor ( n435289 , n435282 , n435288 );
buf ( n435290 , n435289 );
buf ( n435291 , n435290 );
xor ( n435292 , n435140 , n435291 );
nand ( n435293 , n434787 , n434790 );
not ( n435294 , n435293 );
not ( n435295 , n434797 );
or ( n435296 , n435294 , n435295 );
nand ( n435297 , n434786 , n434541 );
nand ( n435298 , n435296 , n435297 );
buf ( n435299 , n435298 );
xor ( n435300 , n435292 , n435299 );
buf ( n435301 , n435300 );
buf ( n435302 , n435301 );
xor ( n435303 , n434530 , n434535 );
and ( n435304 , n435303 , n434802 );
and ( n435305 , n434530 , n434535 );
or ( n435306 , n435304 , n435305 );
buf ( n435307 , n435306 );
nor ( n435308 , n435302 , n435307 );
buf ( n435309 , n435308 );
nor ( n435310 , n434804 , n435309 );
nand ( n435311 , n434273 , n435310 );
not ( n435312 , n435311 );
buf ( n435313 , n386480 );
not ( n435314 , n435313 );
buf ( n435315 , n22982 );
not ( n435316 , n435315 );
buf ( n435317 , n38823 );
not ( n435318 , n435317 );
or ( n435319 , n435316 , n435318 );
buf ( n435320 , n49938 );
buf ( n435321 , n38971 );
nand ( n435322 , n435320 , n435321 );
buf ( n435323 , n435322 );
buf ( n435324 , n435323 );
nand ( n435325 , n435319 , n435324 );
buf ( n435326 , n435325 );
buf ( n435327 , n435326 );
not ( n435328 , n435327 );
or ( n435329 , n435314 , n435328 );
buf ( n435330 , n435028 );
buf ( n435331 , n386496 );
nand ( n435332 , n435330 , n435331 );
buf ( n435333 , n435332 );
buf ( n435334 , n435333 );
nand ( n435335 , n435329 , n435334 );
buf ( n435336 , n435335 );
buf ( n435337 , n435336 );
buf ( n435338 , n41565 );
not ( n435339 , n435338 );
buf ( n435340 , n24050 );
not ( n435341 , n435340 );
buf ( n435342 , n42616 );
not ( n435343 , n435342 );
or ( n435344 , n435341 , n435343 );
buf ( n435345 , n35301 );
buf ( n435346 , n389075 );
nand ( n435347 , n435345 , n435346 );
buf ( n435348 , n435347 );
buf ( n435349 , n435348 );
nand ( n435350 , n435344 , n435349 );
buf ( n435351 , n435350 );
buf ( n435352 , n435351 );
not ( n435353 , n435352 );
or ( n435354 , n435339 , n435353 );
buf ( n435355 , n435099 );
buf ( n435356 , n389125 );
nand ( n435357 , n435355 , n435356 );
buf ( n435358 , n435357 );
buf ( n435359 , n435358 );
nand ( n435360 , n435354 , n435359 );
buf ( n435361 , n435360 );
buf ( n435362 , n435361 );
xor ( n435363 , n435337 , n435362 );
buf ( n435364 , n390213 );
buf ( n435365 , n434936 );
not ( n435366 , n435365 );
buf ( n435367 , n435366 );
buf ( n435368 , n435367 );
or ( n435369 , n435364 , n435368 );
buf ( n435370 , n386307 );
and ( n435371 , n44399 , n398740 );
not ( n435372 , n44399 );
and ( n435373 , n435372 , n384965 );
nor ( n435374 , n435371 , n435373 );
buf ( n435375 , n435374 );
or ( n435376 , n435370 , n435375 );
nand ( n435377 , n435369 , n435376 );
buf ( n435378 , n435377 );
buf ( n435379 , n435378 );
buf ( n435380 , n383946 );
not ( n435381 , n435380 );
buf ( n435382 , n434637 );
not ( n435383 , n435382 );
buf ( n435384 , n384280 );
not ( n435385 , n435384 );
or ( n435386 , n435383 , n435385 );
buf ( n435387 , n58546 );
buf ( n435388 , n36398 );
nand ( n435389 , n435387 , n435388 );
buf ( n435390 , n435389 );
buf ( n435391 , n435390 );
nand ( n435392 , n435386 , n435391 );
buf ( n435393 , n435392 );
buf ( n435394 , n435393 );
not ( n435395 , n435394 );
or ( n435396 , n435381 , n435395 );
buf ( n435397 , n434828 );
not ( n435398 , n435397 );
buf ( n435399 , n398406 );
nand ( n435400 , n435398 , n435399 );
buf ( n435401 , n435400 );
buf ( n435402 , n435401 );
nand ( n435403 , n435396 , n435402 );
buf ( n435404 , n435403 );
buf ( n435405 , n435404 );
xor ( n435406 , n435379 , n435405 );
buf ( n435407 , n384644 );
not ( n435408 , n435407 );
buf ( n435409 , n434583 );
not ( n435410 , n435409 );
buf ( n435411 , n405715 );
not ( n435412 , n435411 );
or ( n435413 , n435410 , n435412 );
buf ( n435414 , n385740 );
buf ( n435415 , n36252 );
nand ( n435416 , n435414 , n435415 );
buf ( n435417 , n435416 );
buf ( n435418 , n435417 );
nand ( n435419 , n435413 , n435418 );
buf ( n435420 , n435419 );
buf ( n435421 , n435420 );
not ( n435422 , n435421 );
or ( n435423 , n435408 , n435422 );
nand ( n435424 , n435223 , n383897 );
buf ( n435425 , n435424 );
nand ( n435426 , n435423 , n435425 );
buf ( n435427 , n435426 );
buf ( n435428 , n435427 );
xor ( n435429 , n435406 , n435428 );
buf ( n435430 , n435429 );
buf ( n435431 , n435430 );
xor ( n435432 , n435363 , n435431 );
buf ( n435433 , n435432 );
not ( n435434 , n435433 );
or ( n435435 , n435104 , n435075 );
nand ( n435436 , n435435 , n435083 );
nand ( n435437 , n435104 , n435075 );
nand ( n435438 , n435436 , n435437 );
not ( n435439 , n435438 );
nand ( n435440 , n435434 , n435439 );
not ( n435441 , n435440 );
not ( n435442 , n435170 );
not ( n435443 , n435442 );
not ( n435444 , n435187 );
or ( n435445 , n435443 , n435444 );
nand ( n435446 , n435445 , n435192 );
nand ( n435447 , n435186 , n435170 );
nand ( n435448 , n435446 , n435447 );
not ( n435449 , n435448 );
or ( n435450 , n435441 , n435449 );
nand ( n435451 , n435438 , n435433 );
nand ( n435452 , n435450 , n435451 );
buf ( n435453 , n434870 );
not ( n435454 , n435453 );
buf ( n435455 , n41374 );
not ( n435456 , n435455 );
or ( n435457 , n435454 , n435456 );
buf ( n435458 , n434884 );
nand ( n435459 , n435457 , n435458 );
buf ( n435460 , n435459 );
buf ( n435461 , n435460 );
buf ( n435462 , n37695 );
not ( n435463 , n435462 );
buf ( n435464 , n37347 );
not ( n435465 , n435464 );
buf ( n435466 , n390373 );
not ( n435467 , n435466 );
or ( n435468 , n435465 , n435467 );
buf ( n435469 , n390379 );
buf ( n435470 , n37354 );
nand ( n435471 , n435469 , n435470 );
buf ( n435472 , n435471 );
buf ( n435473 , n435472 );
nand ( n435474 , n435468 , n435473 );
buf ( n435475 , n435474 );
buf ( n435476 , n435475 );
not ( n435477 , n435476 );
or ( n435478 , n435463 , n435477 );
buf ( n435479 , n434991 );
buf ( n435480 , n385269 );
nand ( n435481 , n435479 , n435480 );
buf ( n435482 , n435481 );
buf ( n435483 , n435482 );
nand ( n435484 , n435478 , n435483 );
buf ( n435485 , n435484 );
buf ( n435486 , n435485 );
xor ( n435487 , n435461 , n435486 );
xor ( n435488 , n435209 , n435228 );
and ( n435489 , n435488 , n435244 );
and ( n435490 , n435209 , n435228 );
or ( n435491 , n435489 , n435490 );
buf ( n435492 , n435491 );
buf ( n435493 , n435492 );
and ( n435494 , n435487 , n435493 );
and ( n435495 , n435461 , n435486 );
or ( n435496 , n435494 , n435495 );
buf ( n435497 , n435496 );
not ( n435498 , n386480 );
not ( n435499 , n22982 );
not ( n435500 , n383575 );
or ( n435501 , n435499 , n435500 );
not ( n435502 , n22982 );
nand ( n435503 , n435502 , n39051 );
nand ( n435504 , n435501 , n435503 );
not ( n435505 , n435504 );
or ( n435506 , n435498 , n435505 );
buf ( n435507 , n435326 );
buf ( n435508 , n386496 );
nand ( n435509 , n435507 , n435508 );
buf ( n435510 , n435509 );
nand ( n435511 , n435506 , n435510 );
not ( n435512 , n435511 );
not ( n435513 , n391080 );
buf ( n435514 , n24074 );
not ( n435515 , n435514 );
buf ( n435516 , n386421 );
not ( n435517 , n435516 );
or ( n435518 , n435515 , n435517 );
buf ( n435519 , n383056 );
buf ( n435520 , n24073 );
nand ( n435521 , n435519 , n435520 );
buf ( n435522 , n435521 );
buf ( n435523 , n435522 );
nand ( n435524 , n435518 , n435523 );
buf ( n435525 , n435524 );
not ( n435526 , n435525 );
or ( n435527 , n435513 , n435526 );
buf ( n435528 , n24074 );
not ( n435529 , n435528 );
buf ( n435530 , n383108 );
not ( n435531 , n435530 );
or ( n435532 , n435529 , n435531 );
buf ( n435533 , n383111 );
buf ( n435534 , n24073 );
nand ( n435535 , n435533 , n435534 );
buf ( n435536 , n435535 );
buf ( n435537 , n435536 );
nand ( n435538 , n435532 , n435537 );
buf ( n435539 , n435538 );
nand ( n435540 , n390403 , n435539 );
nand ( n435541 , n435527 , n435540 );
not ( n435542 , n435541 );
not ( n435543 , n389547 );
buf ( n435544 , n388376 );
not ( n435545 , n435544 );
buf ( n435546 , n384096 );
not ( n435547 , n435546 );
or ( n435548 , n435545 , n435547 );
buf ( n435549 , n382854 );
buf ( n435550 , n388373 );
nand ( n435551 , n435549 , n435550 );
buf ( n435552 , n435551 );
buf ( n435553 , n435552 );
nand ( n435554 , n435548 , n435553 );
buf ( n435555 , n435554 );
not ( n435556 , n435555 );
or ( n435557 , n435543 , n435556 );
and ( n435558 , n385292 , n388646 );
not ( n435559 , n385292 );
and ( n435560 , n435559 , n388654 );
nor ( n435561 , n435558 , n435560 );
nand ( n435562 , n435557 , C1 );
buf ( n435563 , n435562 );
buf ( n435564 , n385359 );
not ( n435565 , n435564 );
buf ( n435566 , n394392 );
not ( n435567 , n435566 );
or ( n435568 , n435565 , n435567 );
buf ( n435569 , n44007 );
buf ( n435570 , n395885 );
nand ( n435571 , n435569 , n435570 );
buf ( n435572 , n435571 );
buf ( n435573 , n435572 );
nand ( n435574 , n435568 , n435573 );
buf ( n435575 , n435574 );
buf ( n435576 , n435575 );
not ( n435577 , n435576 );
buf ( n435578 , n390485 );
not ( n435579 , n435578 );
or ( n435580 , n435577 , n435579 );
buf ( n435581 , n385324 );
not ( n435582 , n435581 );
buf ( n435583 , n384562 );
not ( n435584 , n435583 );
or ( n435585 , n435582 , n435584 );
buf ( n435586 , n395885 );
buf ( n435587 , n386236 );
nand ( n435588 , n435586 , n435587 );
buf ( n435589 , n435588 );
buf ( n435590 , n435589 );
nand ( n435591 , n435585 , n435590 );
buf ( n435592 , n435591 );
buf ( n435593 , n435592 );
buf ( n435594 , n384554 );
nand ( n435595 , n435593 , n435594 );
buf ( n435596 , n435595 );
buf ( n435597 , n435596 );
nand ( n435598 , n435580 , n435597 );
buf ( n435599 , n435598 );
buf ( n435600 , n435599 );
xor ( n435601 , n435563 , n435600 );
buf ( n435602 , n390213 );
buf ( n435603 , n435374 );
or ( n435604 , n435602 , n435603 );
buf ( n435605 , n386307 );
buf ( n435606 , n388445 );
buf ( n435607 , n35435 );
and ( n435608 , n435606 , n435607 );
not ( n435609 , n435606 );
buf ( n435610 , n38685 );
and ( n435611 , n435609 , n435610 );
nor ( n435612 , n435608 , n435611 );
buf ( n435613 , n435612 );
buf ( n435614 , n435613 );
or ( n435615 , n435605 , n435614 );
nand ( n435616 , n435604 , n435615 );
buf ( n435617 , n435616 );
buf ( n435618 , n435617 );
xor ( n435619 , n435601 , n435618 );
buf ( n435620 , n435619 );
buf ( n435621 , n435620 );
not ( n435622 , n435621 );
buf ( n435623 , n435622 );
and ( n435624 , n435542 , n435623 );
not ( n435625 , n435542 );
and ( n435626 , n435625 , n435620 );
nor ( n435627 , n435624 , n435626 );
not ( n435628 , n435627 );
or ( n435629 , n435512 , n435628 );
not ( n435630 , n435623 );
nand ( n435631 , n435630 , n435542 );
not ( n435632 , n435620 );
nand ( n435633 , n435632 , n435541 );
not ( n435634 , n435511 );
nand ( n435635 , n435631 , n435633 , n435634 );
nand ( n435636 , n435629 , n435635 );
xor ( n435637 , n435497 , n435636 );
xor ( n435638 , n435337 , n435362 );
and ( n435639 , n435638 , n435431 );
and ( n435640 , n435337 , n435362 );
or ( n435641 , n435639 , n435640 );
buf ( n435642 , n435641 );
xnor ( n435643 , n435637 , n435642 );
not ( n435644 , n435208 );
not ( n435645 , n435644 );
not ( n435646 , n390485 );
not ( n435647 , n390498 );
not ( n435648 , n386182 );
or ( n435649 , n435647 , n435648 );
or ( n435650 , n395885 , n38631 );
nand ( n435651 , n435649 , n435650 );
not ( n435652 , n435651 );
or ( n435653 , n435646 , n435652 );
buf ( n435654 , n435575 );
buf ( n435655 , n389908 );
nand ( n435656 , n435654 , n435655 );
buf ( n435657 , n435656 );
nand ( n435658 , n435653 , n435657 );
not ( n435659 , n435658 );
or ( n435660 , n435645 , n435659 );
not ( n435661 , n435208 );
buf ( n435662 , n435658 );
not ( n435663 , n435662 );
buf ( n435664 , n435663 );
not ( n435665 , n435664 );
or ( n435666 , n435661 , n435665 );
buf ( n435667 , n391920 );
buf ( n435668 , n434958 );
or ( n435669 , n435667 , n435668 );
buf ( n435670 , n383403 );
buf ( n435671 , n386150 );
buf ( n435672 , n389589 );
and ( n435673 , n435671 , n435672 );
not ( n435674 , n435671 );
buf ( n435675 , n391183 );
and ( n435676 , n435674 , n435675 );
nor ( n435677 , n435673 , n435676 );
buf ( n435678 , n435677 );
buf ( n435679 , n435678 );
or ( n435680 , n435670 , n435679 );
nand ( n435681 , n435669 , n435680 );
buf ( n435682 , n435681 );
nand ( n435683 , n435666 , n435682 );
nand ( n435684 , n435660 , n435683 );
not ( n435685 , n435684 );
not ( n435686 , n435685 );
buf ( n435687 , n388141 );
not ( n435688 , n435687 );
buf ( n435689 , n388160 );
not ( n435690 , n435689 );
buf ( n435691 , n34861 );
not ( n435692 , n435691 );
or ( n435693 , n435690 , n435692 );
buf ( n435694 , n399653 );
buf ( n435695 , n388157 );
nand ( n435696 , n435694 , n435695 );
buf ( n435697 , n435696 );
buf ( n435698 , n435697 );
nand ( n435699 , n435693 , n435698 );
buf ( n435700 , n435699 );
buf ( n435701 , n435700 );
not ( n435702 , n435701 );
or ( n435703 , n435688 , n435702 );
buf ( n435704 , n388160 );
not ( n435705 , n435704 );
buf ( n435706 , n382548 );
not ( n435707 , n435706 );
or ( n435708 , n435705 , n435707 );
buf ( n435709 , n391212 );
buf ( n435710 , n388157 );
nand ( n435711 , n435709 , n435710 );
buf ( n435712 , n435711 );
buf ( n435713 , n435712 );
nand ( n435714 , n435708 , n435713 );
buf ( n435715 , n435714 );
buf ( n435716 , n435715 );
buf ( n435717 , n40701 );
nand ( n435718 , n435716 , n435717 );
buf ( n435719 , n435718 );
buf ( n435720 , n435719 );
nand ( n435721 , n435703 , n435720 );
buf ( n435722 , n435721 );
not ( n435723 , n435722 );
or ( n435724 , n435686 , n435723 );
not ( n435725 , n435722 );
nand ( n435726 , n435725 , n435684 );
nand ( n435727 , n435724 , n435726 );
not ( n435728 , n385889 );
buf ( n435729 , n385494 );
not ( n435730 , n435729 );
buf ( n435731 , n38357 );
not ( n435732 , n435731 );
or ( n435733 , n435730 , n435732 );
buf ( n435734 , n389435 );
buf ( n435735 , n385491 );
nand ( n435736 , n435734 , n435735 );
buf ( n435737 , n435736 );
buf ( n435738 , n435737 );
nand ( n435739 , n435733 , n435738 );
buf ( n435740 , n435739 );
not ( n435741 , n435740 );
or ( n435742 , n435728 , n435741 );
buf ( n435743 , n385494 );
not ( n435744 , n435743 );
buf ( n435745 , n385774 );
not ( n435746 , n435745 );
or ( n435747 , n435744 , n435746 );
buf ( n435748 , n38227 );
buf ( n435749 , n385491 );
nand ( n435750 , n435748 , n435749 );
buf ( n435751 , n435750 );
buf ( n435752 , n435751 );
nand ( n435753 , n435747 , n435752 );
buf ( n435754 , n435753 );
buf ( n435755 , n435754 );
buf ( n435756 , n38324 );
nand ( n435757 , n435755 , n435756 );
buf ( n435758 , n435757 );
nand ( n435759 , n435742 , n435758 );
not ( n435760 , n435759 );
and ( n435761 , n435727 , n435760 );
not ( n435762 , n435727 );
and ( n435763 , n435762 , n435759 );
nor ( n435764 , n435761 , n435763 );
buf ( n435765 , n388141 );
not ( n435766 , n435765 );
buf ( n435767 , n435715 );
not ( n435768 , n435767 );
or ( n435769 , n435766 , n435768 );
buf ( n435770 , n40701 );
buf ( n435771 , n435163 );
nand ( n435772 , n435770 , n435771 );
buf ( n435773 , n435772 );
buf ( n435774 , n435773 );
nand ( n435775 , n435769 , n435774 );
buf ( n435776 , n435775 );
buf ( n435777 , n435776 );
xor ( n435778 , n434918 , n434942 );
and ( n435779 , n435778 , n434960 );
and ( n435780 , n434918 , n434942 );
or ( n435781 , n435779 , n435780 );
buf ( n435782 , n435781 );
xor ( n435783 , n435777 , n435782 );
buf ( n435784 , n435658 );
buf ( n435785 , n435208 );
xor ( n435786 , n435784 , n435785 );
buf ( n435787 , n435682 );
not ( n435788 , n435787 );
xor ( n435789 , n435786 , n435788 );
buf ( n435790 , n435789 );
buf ( n435791 , n435790 );
and ( n435792 , n435783 , n435791 );
and ( n435793 , n435777 , n435782 );
or ( n435794 , n435792 , n435793 );
buf ( n435795 , n435794 );
and ( n435796 , n435764 , n435795 );
not ( n435797 , n435764 );
not ( n435798 , n435795 );
and ( n435799 , n435797 , n435798 );
nor ( n435800 , n435796 , n435799 );
xor ( n435801 , n435379 , n435405 );
and ( n435802 , n435801 , n435428 );
and ( n435803 , n435379 , n435405 );
or ( n435804 , n435802 , n435803 );
buf ( n435805 , n435804 );
not ( n435806 , n435805 );
not ( n435807 , n435806 );
buf ( n435808 , n385269 );
not ( n435809 , n435808 );
buf ( n435810 , n435475 );
not ( n435811 , n435810 );
or ( n435812 , n435809 , n435811 );
buf ( n435813 , n37347 );
not ( n435814 , n435813 );
buf ( n435815 , n389525 );
not ( n435816 , n435815 );
or ( n435817 , n435814 , n435816 );
buf ( n435818 , n384741 );
buf ( n435819 , n37354 );
nand ( n435820 , n435818 , n435819 );
buf ( n435821 , n435820 );
buf ( n435822 , n435821 );
nand ( n435823 , n435817 , n435822 );
buf ( n435824 , n435823 );
buf ( n435825 , n435824 );
buf ( n435826 , n37695 );
nand ( n435827 , n435825 , n435826 );
buf ( n435828 , n435827 );
buf ( n435829 , n435828 );
nand ( n435830 , n435812 , n435829 );
buf ( n435831 , n435830 );
not ( n435832 , n435831 );
not ( n435833 , n435832 );
buf ( n435834 , n42825 );
not ( n435835 , n435834 );
buf ( n435836 , n385972 );
not ( n435837 , n435836 );
or ( n435838 , n435835 , n435837 );
buf ( n435839 , n31964 );
buf ( n435840 , n74955 );
nand ( n435841 , n435839 , n435840 );
buf ( n435842 , n435841 );
buf ( n435843 , n435842 );
nand ( n435844 , n435838 , n435843 );
buf ( n435845 , n435844 );
buf ( n435846 , n435845 );
not ( n435847 , n435846 );
buf ( n435848 , n398431 );
not ( n435849 , n435848 );
or ( n435850 , n435847 , n435849 );
buf ( n435851 , n379463 );
buf ( n435852 , n27613 );
not ( n435853 , n435852 );
buf ( n435854 , n385987 );
not ( n435855 , n435854 );
or ( n435856 , n435853 , n435855 );
buf ( n435857 , n397524 );
buf ( n435858 , n40971 );
nand ( n435859 , n435857 , n435858 );
buf ( n435860 , n435859 );
buf ( n435861 , n435860 );
nand ( n435862 , n435856 , n435861 );
buf ( n435863 , n435862 );
buf ( n435864 , n435863 );
nand ( n435865 , n435851 , n435864 );
buf ( n435866 , n435865 );
buf ( n435867 , n435866 );
nand ( n435868 , n435850 , n435867 );
buf ( n435869 , n435868 );
buf ( n435870 , n435869 );
not ( n435871 , n435870 );
buf ( n435872 , n384413 );
not ( n435873 , n435872 );
buf ( n435874 , n40943 );
not ( n435875 , n435874 );
buf ( n435876 , n384083 );
not ( n435877 , n435876 );
or ( n435878 , n435875 , n435877 );
buf ( n435879 , n385983 );
buf ( n435880 , n388419 );
nand ( n435881 , n435879 , n435880 );
buf ( n435882 , n435881 );
buf ( n435883 , n435882 );
nand ( n435884 , n435878 , n435883 );
buf ( n435885 , n435884 );
buf ( n435886 , n435885 );
not ( n435887 , n435886 );
or ( n435888 , n435873 , n435887 );
buf ( n435889 , n36801 );
and ( n435890 , n41896 , n388419 );
not ( n435891 , n41896 );
and ( n435892 , n435891 , n36808 );
nor ( n435893 , n435890 , n435892 );
buf ( n435894 , n435893 );
nand ( n435895 , n435889 , n435894 );
buf ( n435896 , n435895 );
buf ( n435897 , n435896 );
nand ( n435898 , n435888 , n435897 );
buf ( n435899 , n435898 );
buf ( n435900 , n435899 );
not ( n435901 , n435900 );
buf ( n435902 , n435901 );
buf ( n435903 , n435902 );
not ( n435904 , n435903 );
or ( n435905 , n435871 , n435904 );
buf ( n435906 , n435899 );
buf ( n435907 , n435869 );
not ( n435908 , n435907 );
buf ( n435909 , n435908 );
buf ( n435910 , n435909 );
nand ( n435911 , n435906 , n435910 );
buf ( n435912 , n435911 );
buf ( n435913 , n435912 );
nand ( n435914 , n435905 , n435913 );
buf ( n435915 , n435914 );
not ( n435916 , n391173 );
buf ( n435917 , n386182 );
not ( n435918 , n435917 );
buf ( n435919 , n435918 );
buf ( n435920 , n435919 );
not ( n435921 , n435920 );
buf ( n435922 , n383426 );
not ( n435923 , n435922 );
or ( n435924 , n435921 , n435923 );
buf ( n435925 , n388556 );
buf ( n435926 , n386182 );
nand ( n435927 , n435925 , n435926 );
buf ( n435928 , n435927 );
buf ( n435929 , n435928 );
nand ( n435930 , n435924 , n435929 );
buf ( n435931 , n435930 );
not ( n435932 , n435931 );
or ( n435933 , n435916 , n435932 );
not ( n435934 , n435678 );
nand ( n435935 , n435934 , n391652 );
nand ( n435936 , n435933 , n435935 );
buf ( n435937 , n435936 );
not ( n435938 , n435937 );
buf ( n435939 , n435938 );
and ( n435940 , n435915 , n435939 );
not ( n435941 , n435915 );
and ( n435942 , n435941 , n435936 );
nor ( n435943 , n435940 , n435942 );
not ( n435944 , n435943 );
not ( n435945 , n435944 );
or ( n435946 , n435833 , n435945 );
or ( n435947 , n435944 , n435832 );
nand ( n435948 , n435946 , n435947 );
not ( n435949 , n435948 );
or ( n435950 , n435807 , n435949 );
or ( n435951 , n435948 , n435806 );
nand ( n435952 , n435950 , n435951 );
xor ( n435953 , n435800 , n435952 );
not ( n435954 , n435953 );
nor ( n435955 , n435452 , n435643 , n435954 );
not ( n435956 , n435955 );
not ( n435957 , n435643 );
nand ( n435958 , n435452 , n435957 , n435954 );
not ( n435959 , n435452 );
buf ( n435960 , n435643 );
nand ( n435961 , n435959 , n435960 , n435954 );
nand ( n435962 , n435960 , n435452 , n435953 );
nand ( n435963 , n435956 , n435958 , n435961 , n435962 );
not ( n435964 , n435963 );
not ( n435965 , n434824 );
nand ( n435966 , n435965 , n434838 );
not ( n435967 , n435966 );
not ( n435968 , n434859 );
or ( n435969 , n435967 , n435968 );
buf ( n435970 , n434841 );
buf ( n435971 , n434824 );
nand ( n435972 , n435970 , n435971 );
buf ( n435973 , n435972 );
nand ( n435974 , n435969 , n435973 );
buf ( n435975 , n435974 );
buf ( n435976 , n434855 );
not ( n435977 , n435976 );
buf ( n435978 , n389015 );
not ( n435979 , n435978 );
or ( n435980 , n435977 , n435979 );
buf ( n435981 , n389024 );
buf ( n435982 , n435845 );
nand ( n435983 , n435981 , n435982 );
buf ( n435984 , n435983 );
buf ( n435985 , n435984 );
nand ( n435986 , n435980 , n435985 );
buf ( n435987 , n435986 );
buf ( n435988 , n435987 );
not ( n435989 , n435893 );
not ( n435990 , n40901 );
or ( n435991 , n435989 , n435990 );
buf ( n435992 , n36801 );
buf ( n435993 , n434817 );
nand ( n435994 , n435992 , n435993 );
buf ( n435995 , n435994 );
nand ( n435996 , n435991 , n435995 );
buf ( n435997 , n435996 );
xor ( n435998 , n435988 , n435997 );
not ( n435999 , n388498 );
nand ( n436000 , n435999 , n435561 );
nand ( n436001 , C1 , n436000 );
buf ( n436002 , n436001 );
xor ( n436003 , n435998 , n436002 );
buf ( n436004 , n436003 );
buf ( n436005 , n436004 );
xor ( n436006 , n435975 , n436005 );
buf ( n436007 , n38324 );
not ( n436008 , n436007 );
buf ( n436009 , n435740 );
not ( n436010 , n436009 );
or ( n436011 , n436008 , n436010 );
buf ( n436012 , n435070 );
buf ( n436013 , n385889 );
nand ( n436014 , n436012 , n436013 );
buf ( n436015 , n436014 );
buf ( n436016 , n436015 );
nand ( n436017 , n436011 , n436016 );
buf ( n436018 , n436017 );
buf ( n436019 , n436018 );
xor ( n436020 , n436006 , n436019 );
buf ( n436021 , n436020 );
buf ( n436022 , n436021 );
xor ( n436023 , n435461 , n435486 );
xor ( n436024 , n436023 , n435493 );
buf ( n436025 , n436024 );
buf ( n436026 , n436025 );
xor ( n436027 , n436022 , n436026 );
xor ( n436028 , n435777 , n435782 );
xor ( n436029 , n436028 , n435791 );
buf ( n436030 , n436029 );
buf ( n436031 , n436030 );
xor ( n436032 , n436027 , n436031 );
buf ( n436033 , n436032 );
buf ( n436034 , n436033 );
buf ( n436035 , n435106 );
not ( n436036 , n436035 );
buf ( n436037 , n435116 );
not ( n436038 , n436037 );
or ( n436039 , n436036 , n436038 );
buf ( n436040 , n435133 );
nand ( n436041 , n436039 , n436040 );
buf ( n436042 , n436041 );
buf ( n436043 , n436042 );
buf ( n436044 , n435115 );
buf ( n436045 , n435105 );
nand ( n436046 , n436044 , n436045 );
buf ( n436047 , n436046 );
buf ( n436048 , n436047 );
nand ( n436049 , n436043 , n436048 );
buf ( n436050 , n436049 );
buf ( n436051 , n436050 );
xor ( n436052 , n436034 , n436051 );
nand ( n436053 , n435434 , n435438 );
nand ( n436054 , n435433 , n435439 );
nand ( n436055 , n436053 , n436054 );
xor ( n436056 , n436055 , n435448 );
buf ( n436057 , n436056 );
and ( n436058 , n436052 , n436057 );
and ( n436059 , n436034 , n436051 );
or ( n436060 , n436058 , n436059 );
buf ( n436061 , n436060 );
buf ( n436062 , n436061 );
buf ( n436063 , n435262 );
buf ( n436064 , n435246 );
nor ( n436065 , n436063 , n436064 );
buf ( n436066 , n436065 );
buf ( n436067 , n436066 );
buf ( n436068 , n435268 );
or ( n436069 , n436067 , n436068 );
buf ( n436070 , n435262 );
buf ( n436071 , n435246 );
nand ( n436072 , n436070 , n436071 );
buf ( n436073 , n436072 );
buf ( n436074 , n436073 );
nand ( n436075 , n436069 , n436074 );
buf ( n436076 , n436075 );
buf ( n436077 , n436076 );
not ( n436078 , n434890 );
nand ( n436079 , n436078 , n434860 );
not ( n436080 , n436079 );
not ( n436081 , n434961 );
or ( n436082 , n436080 , n436081 );
not ( n436083 , n434860 );
nand ( n436084 , n436083 , n434890 );
nand ( n436085 , n436082 , n436084 );
buf ( n436086 , n435040 );
buf ( n436087 , n435004 );
nand ( n436088 , n436086 , n436087 );
buf ( n436089 , n436088 );
buf ( n436090 , n436089 );
buf ( n436091 , n434984 );
and ( n436092 , n436090 , n436091 );
buf ( n436093 , n435035 );
buf ( n436094 , n435001 );
and ( n436095 , n436093 , n436094 );
buf ( n436096 , n436095 );
buf ( n436097 , n436096 );
nor ( n436098 , n436092 , n436097 );
buf ( n436099 , n436098 );
buf ( n436100 , n436099 );
not ( n436101 , n436100 );
buf ( n436102 , n436101 );
buf ( n436103 , n436102 );
not ( n436104 , n436103 );
buf ( n436105 , n435179 );
buf ( n436106 , n391080 );
and ( n436107 , n436105 , n436106 );
buf ( n436108 , n435525 );
not ( n436109 , n436108 );
buf ( n436110 , n42925 );
nor ( n436111 , n436109 , n436110 );
buf ( n436112 , n436111 );
buf ( n436113 , n436112 );
nor ( n436114 , n436107 , n436113 );
buf ( n436115 , n436114 );
buf ( n436116 , n436115 );
not ( n436117 , n436116 );
or ( n436118 , n436104 , n436117 );
buf ( n436119 , n436115 );
not ( n436120 , n436119 );
buf ( n436121 , n436120 );
buf ( n436122 , n436121 );
buf ( n436123 , n436099 );
nand ( n436124 , n436122 , n436123 );
buf ( n436125 , n436124 );
buf ( n436126 , n436125 );
nand ( n436127 , n436118 , n436126 );
buf ( n436128 , n436127 );
xor ( n436129 , n436085 , n436128 );
buf ( n436130 , n436129 );
xor ( n436131 , n436077 , n436130 );
not ( n436132 , n435049 );
not ( n436133 , n434968 );
buf ( n436134 , n436133 );
buf ( n436135 , n435043 );
nand ( n436136 , n436134 , n436135 );
buf ( n436137 , n436136 );
not ( n436138 , n436137 );
or ( n436139 , n436132 , n436138 );
not ( n436140 , n436133 );
nand ( n436141 , n436140 , n435042 );
nand ( n436142 , n436139 , n436141 );
buf ( n436143 , n436142 );
and ( n436144 , n436131 , n436143 );
and ( n436145 , n436077 , n436130 );
or ( n436146 , n436144 , n436145 );
buf ( n436147 , n436146 );
buf ( n436148 , n436147 );
not ( n436149 , n436102 );
not ( n436150 , n436121 );
or ( n436151 , n436149 , n436150 );
not ( n436152 , n436099 );
not ( n436153 , n436115 );
or ( n436154 , n436152 , n436153 );
nand ( n436155 , n436154 , n436085 );
nand ( n436156 , n436151 , n436155 );
buf ( n436157 , n41565 );
not ( n436158 , n436157 );
buf ( n436159 , n24050 );
not ( n436160 , n436159 );
buf ( n436161 , n386561 );
not ( n436162 , n436161 );
or ( n436163 , n436160 , n436162 );
buf ( n436164 , n382921 );
buf ( n436165 , n389075 );
nand ( n436166 , n436164 , n436165 );
buf ( n436167 , n436166 );
buf ( n436168 , n436167 );
nand ( n436169 , n436163 , n436168 );
buf ( n436170 , n436169 );
buf ( n436171 , n436170 );
not ( n436172 , n436171 );
or ( n436173 , n436158 , n436172 );
buf ( n436174 , n435351 );
buf ( n436175 , n389125 );
nand ( n436176 , n436174 , n436175 );
buf ( n436177 , n436176 );
buf ( n436178 , n436177 );
nand ( n436179 , n436173 , n436178 );
buf ( n436180 , n436179 );
buf ( n436181 , n398406 );
not ( n436182 , n436181 );
buf ( n436183 , n435393 );
not ( n436184 , n436183 );
or ( n436185 , n436182 , n436184 );
buf ( n436186 , n434637 );
not ( n436187 , n436186 );
buf ( n436188 , n390810 );
not ( n436189 , n436188 );
or ( n436190 , n436187 , n436189 );
buf ( n436191 , n38472 );
buf ( n436192 , n36398 );
nand ( n436193 , n436191 , n436192 );
buf ( n436194 , n436193 );
buf ( n436195 , n436194 );
nand ( n436196 , n436190 , n436195 );
buf ( n436197 , n436196 );
buf ( n436198 , n436197 );
buf ( n436199 , n383946 );
nand ( n436200 , n436198 , n436199 );
buf ( n436201 , n436200 );
buf ( n436202 , n436201 );
nand ( n436203 , n436185 , n436202 );
buf ( n436204 , n436203 );
buf ( n436205 , n436204 );
buf ( n436206 , n383897 );
not ( n436207 , n436206 );
buf ( n436208 , n435420 );
not ( n436209 , n436208 );
or ( n436210 , n436207 , n436209 );
buf ( n436211 , n434583 );
not ( n436212 , n436211 );
buf ( n436213 , n36218 );
not ( n436214 , n436213 );
or ( n436215 , n436212 , n436214 );
buf ( n436216 , n48234 );
buf ( n436217 , n36252 );
nand ( n436218 , n436216 , n436217 );
buf ( n436219 , n436218 );
buf ( n436220 , n436219 );
nand ( n436221 , n436215 , n436220 );
buf ( n436222 , n436221 );
buf ( n436223 , n436222 );
buf ( n436224 , n384644 );
nand ( n436225 , n436223 , n436224 );
buf ( n436226 , n436225 );
buf ( n436227 , n436226 );
nand ( n436228 , n436210 , n436227 );
buf ( n436229 , n436228 );
buf ( n436230 , n436229 );
xor ( n436231 , n436205 , n436230 );
xor ( n436232 , n435988 , n435997 );
and ( n436233 , n436232 , n436002 );
and ( n436234 , n435988 , n435997 );
or ( n436235 , n436233 , n436234 );
buf ( n436236 , n436235 );
buf ( n436237 , n436236 );
xor ( n436238 , n436231 , n436237 );
buf ( n436239 , n436238 );
xor ( n436240 , n436180 , n436239 );
xor ( n436241 , n435975 , n436005 );
and ( n436242 , n436241 , n436019 );
and ( n436243 , n435975 , n436005 );
or ( n436244 , n436242 , n436243 );
buf ( n436245 , n436244 );
xor ( n436246 , n436240 , n436245 );
xor ( n436247 , n436156 , n436246 );
xor ( n436248 , n436022 , n436026 );
and ( n436249 , n436248 , n436031 );
and ( n436250 , n436022 , n436026 );
or ( n436251 , n436249 , n436250 );
buf ( n436252 , n436251 );
xor ( n436253 , n436247 , n436252 );
buf ( n436254 , n436253 );
not ( n436255 , n436254 );
buf ( n436256 , n436255 );
buf ( n436257 , n436256 );
and ( n436258 , n436148 , n436257 );
not ( n436259 , n436148 );
buf ( n436260 , n436253 );
and ( n436261 , n436259 , n436260 );
nor ( n436262 , n436258 , n436261 );
buf ( n436263 , n436262 );
buf ( n436264 , n436263 );
and ( n436265 , n436062 , n436264 );
not ( n436266 , n436062 );
buf ( n436267 , n436263 );
not ( n436268 , n436267 );
buf ( n436269 , n436268 );
buf ( n436270 , n436269 );
and ( n436271 , n436266 , n436270 );
nor ( n436272 , n436265 , n436271 );
buf ( n436273 , n436272 );
not ( n436274 , n436273 );
not ( n436275 , n436274 );
or ( n436276 , n435964 , n436275 );
not ( n436277 , n435963 );
nand ( n436278 , n436273 , n436277 );
nand ( n436279 , n436276 , n436278 );
xor ( n436280 , n436077 , n436130 );
xor ( n436281 , n436280 , n436143 );
buf ( n436282 , n436281 );
not ( n436283 , n436282 );
xor ( n436284 , n435195 , n435272 );
and ( n436285 , n436284 , n435278 );
and ( n436286 , n435195 , n435272 );
or ( n436287 , n436285 , n436286 );
buf ( n436288 , n436287 );
not ( n436289 , n436288 );
nand ( n436290 , n436283 , n436289 );
not ( n436291 , n436290 );
not ( n436292 , n435138 );
not ( n436293 , n435051 );
nand ( n436294 , n435057 , n436293 );
not ( n436295 , n436294 );
or ( n436296 , n436292 , n436295 );
nand ( n436297 , n435056 , n435051 );
nand ( n436298 , n436296 , n436297 );
not ( n436299 , n436298 );
or ( n436300 , n436291 , n436299 );
nand ( n436301 , n436282 , n436288 );
nand ( n436302 , n436300 , n436301 );
buf ( n436303 , n436302 );
not ( n436304 , n436303 );
buf ( n436305 , n436304 );
and ( n436306 , n436279 , n436305 );
not ( n436307 , n436279 );
and ( n436308 , n436307 , n436302 );
nor ( n436309 , n436306 , n436308 );
xor ( n436310 , n436034 , n436051 );
xor ( n436311 , n436310 , n436057 );
buf ( n436312 , n436311 );
buf ( n436313 , n436312 );
xor ( n436314 , n435146 , n435281 );
and ( n436315 , n436314 , n435288 );
and ( n436316 , n435146 , n435281 );
or ( n436317 , n436315 , n436316 );
buf ( n436318 , n436317 );
buf ( n436319 , n436318 );
xor ( n436320 , n436313 , n436319 );
not ( n436321 , n436288 );
not ( n436322 , n436282 );
not ( n436323 , n436322 );
or ( n436324 , n436321 , n436323 );
nand ( n436325 , n436289 , n436282 );
nand ( n436326 , n436324 , n436325 );
and ( n436327 , n436326 , n436298 );
not ( n436328 , n436326 );
not ( n436329 , n436298 );
and ( n436330 , n436328 , n436329 );
nor ( n436331 , n436327 , n436330 );
buf ( n436332 , n436331 );
and ( n436333 , n436320 , n436332 );
and ( n436334 , n436313 , n436319 );
or ( n436335 , n436333 , n436334 );
buf ( n436336 , n436335 );
nor ( n436337 , n436309 , n436336 );
buf ( n436338 , n436337 );
not ( n436339 , n436338 );
buf ( n436340 , n436339 );
xor ( n436341 , n436313 , n436319 );
xor ( n436342 , n436341 , n436332 );
buf ( n436343 , n436342 );
xor ( n436344 , n435140 , n435291 );
and ( n436345 , n436344 , n435299 );
and ( n436346 , n435140 , n435291 );
or ( n436347 , n436345 , n436346 );
buf ( n436348 , n436347 );
or ( n436349 , n436343 , n436348 );
nand ( n436350 , n436340 , n436349 );
not ( n436351 , n40640 );
not ( n436352 , n40700 );
or ( n436353 , n436351 , n436352 );
nand ( n436354 , n436353 , n435700 );
not ( n436355 , n436222 );
not ( n436356 , n383897 );
or ( n436357 , n436355 , n436356 );
not ( n436358 , n383910 );
not ( n436359 , n42153 );
not ( n436360 , n36253 );
or ( n436361 , n436359 , n436360 );
buf ( n436362 , n383765 );
buf ( n436363 , n36252 );
nand ( n436364 , n436362 , n436363 );
buf ( n436365 , n436364 );
nand ( n436366 , n436361 , n436365 );
nand ( n436367 , n436358 , n436366 );
nand ( n436368 , n436357 , n436367 );
xor ( n436369 , n436354 , n436368 );
buf ( n436370 , n435562 );
not ( n436371 , n436370 );
buf ( n436372 , n435617 );
not ( n436373 , n436372 );
buf ( n436374 , n436373 );
buf ( n436375 , n436374 );
not ( n436376 , n436375 );
or ( n436377 , n436371 , n436376 );
buf ( n436378 , n435599 );
nand ( n436379 , n436377 , n436378 );
buf ( n436380 , n436379 );
not ( n436381 , n435562 );
nand ( n436382 , n435617 , n436381 );
nand ( n436383 , n436380 , n436382 );
and ( n436384 , n436369 , n436383 );
and ( n436385 , n436354 , n436368 );
or ( n436386 , n436384 , n436385 );
buf ( n436387 , n435869 );
not ( n436388 , n436387 );
buf ( n436389 , n435899 );
not ( n436390 , n436389 );
or ( n436391 , n436388 , n436390 );
buf ( n436392 , n435936 );
buf ( n436393 , n435902 );
buf ( n436394 , n435909 );
nand ( n436395 , n436393 , n436394 );
buf ( n436396 , n436395 );
buf ( n436397 , n436396 );
nand ( n436398 , n436392 , n436397 );
buf ( n436399 , n436398 );
buf ( n436400 , n436399 );
nand ( n436401 , n436391 , n436400 );
buf ( n436402 , n436401 );
not ( n436403 , n436402 );
buf ( n436404 , n390403 );
not ( n436405 , n436404 );
buf ( n436406 , n24074 );
not ( n436407 , n436406 );
buf ( n436408 , n382548 );
not ( n436409 , n436408 );
or ( n436410 , n436407 , n436409 );
buf ( n436411 , n390345 );
buf ( n436412 , n24073 );
nand ( n436413 , n436411 , n436412 );
buf ( n436414 , n436413 );
buf ( n436415 , n436414 );
nand ( n436416 , n436410 , n436415 );
buf ( n436417 , n436416 );
buf ( n436418 , n436417 );
not ( n436419 , n436418 );
or ( n436420 , n436405 , n436419 );
buf ( n436421 , n435539 );
buf ( n436422 , n391080 );
nand ( n436423 , n436421 , n436422 );
buf ( n436424 , n436423 );
buf ( n436425 , n436424 );
nand ( n436426 , n436420 , n436425 );
buf ( n436427 , n436426 );
not ( n436428 , n436427 );
or ( n436429 , n436403 , n436428 );
not ( n436430 , n436402 );
not ( n436431 , n436430 );
not ( n436432 , n436427 );
not ( n436433 , n436432 );
or ( n436434 , n436431 , n436433 );
buf ( n436435 , n389348 );
buf ( n436436 , n41195 );
buf ( n436437 , n382857 );
and ( n436438 , n436436 , n436437 );
not ( n436439 , n436436 );
buf ( n436440 , n385331 );
and ( n436441 , n436439 , n436440 );
nor ( n436442 , n436438 , n436441 );
buf ( n436443 , n436442 );
buf ( n436444 , n436443 );
or ( n436445 , n436435 , n436444 );
nand ( n436446 , C1 , n436445 );
buf ( n436447 , n436446 );
buf ( n436448 , n436447 );
buf ( n436449 , n435863 );
not ( n436450 , n436449 );
buf ( n436451 , n382598 );
not ( n436452 , n436451 );
or ( n436453 , n436450 , n436452 );
buf ( n436454 , n375784 );
buf ( n436455 , n31964 );
and ( n436456 , n436454 , n436455 );
not ( n436457 , n436454 );
buf ( n436458 , n385972 );
and ( n436459 , n436457 , n436458 );
or ( n436460 , n436456 , n436459 );
buf ( n436461 , n436460 );
buf ( n436462 , n436461 );
not ( n436463 , n436462 );
buf ( n436464 , n379466 );
nand ( n436465 , n436463 , n436464 );
buf ( n436466 , n436465 );
buf ( n436467 , n436466 );
nand ( n436468 , n436453 , n436467 );
buf ( n436469 , n436468 );
buf ( n436470 , n436469 );
xor ( n436471 , n436448 , n436470 );
buf ( n436472 , n383479 );
buf ( n436473 , n435931 );
not ( n436474 , n436473 );
buf ( n436475 , n436474 );
buf ( n436476 , n436475 );
or ( n436477 , n436472 , n436476 );
buf ( n436478 , n383499 );
buf ( n436479 , n385345 );
buf ( n436480 , n385729 );
and ( n436481 , n436479 , n436480 );
not ( n436482 , n436479 );
buf ( n436483 , n383426 );
and ( n436484 , n436482 , n436483 );
nor ( n436485 , n436481 , n436484 );
buf ( n436486 , n436485 );
buf ( n436487 , n436486 );
or ( n436488 , n436478 , n436487 );
nand ( n436489 , n436477 , n436488 );
buf ( n436490 , n436489 );
buf ( n436491 , n436490 );
xor ( n436492 , n436471 , n436491 );
buf ( n436493 , n436492 );
nand ( n436494 , n436434 , n436493 );
nand ( n436495 , n436429 , n436494 );
xor ( n436496 , n436386 , n436495 );
buf ( n436497 , n384369 );
not ( n436498 , n436497 );
buf ( n436499 , n36821 );
not ( n436500 , n436499 );
buf ( n436501 , n384280 );
not ( n436502 , n436501 );
or ( n436503 , n436500 , n436502 );
buf ( n436504 , n384286 );
buf ( n436505 , n40886 );
nand ( n436506 , n436504 , n436505 );
buf ( n436507 , n436506 );
buf ( n436508 , n436507 );
nand ( n436509 , n436503 , n436508 );
buf ( n436510 , n436509 );
buf ( n436511 , n436510 );
not ( n436512 , n436511 );
or ( n436513 , n436498 , n436512 );
buf ( n436514 , n36821 );
not ( n436515 , n436514 );
buf ( n436516 , n41596 );
not ( n436517 , n436516 );
or ( n436518 , n436515 , n436517 );
buf ( n436519 , n397419 );
not ( n436520 , n436519 );
buf ( n436521 , n40886 );
nand ( n436522 , n436520 , n436521 );
buf ( n436523 , n436522 );
buf ( n436524 , n436523 );
nand ( n436525 , n436518 , n436524 );
buf ( n436526 , n436525 );
buf ( n436527 , n436526 );
buf ( n436528 , n384416 );
nand ( n436529 , n436527 , n436528 );
buf ( n436530 , n436529 );
buf ( n436531 , n436530 );
nand ( n436532 , n436513 , n436531 );
buf ( n436533 , n436532 );
buf ( n436534 , n436533 );
buf ( n436535 , n385269 );
not ( n436536 , n436535 );
buf ( n436537 , n37347 );
not ( n436538 , n436537 );
buf ( n436539 , n384715 );
not ( n436540 , n436539 );
or ( n436541 , n436538 , n436540 );
buf ( n436542 , n389435 );
buf ( n436543 , n37354 );
nand ( n436544 , n436542 , n436543 );
buf ( n436545 , n436544 );
buf ( n436546 , n436545 );
nand ( n436547 , n436541 , n436546 );
buf ( n436548 , n436547 );
buf ( n436549 , n436548 );
not ( n436550 , n436549 );
or ( n436551 , n436536 , n436550 );
not ( n436552 , n37347 );
not ( n436553 , n36899 );
or ( n436554 , n436552 , n436553 );
nand ( n436555 , n389423 , n37354 );
nand ( n436556 , n436554 , n436555 );
nand ( n436557 , n436556 , n37695 );
buf ( n436558 , n436557 );
nand ( n436559 , n436551 , n436558 );
buf ( n436560 , n436559 );
buf ( n436561 , n436560 );
xor ( n436562 , n436534 , n436561 );
xor ( n436563 , n436448 , n436470 );
and ( n436564 , n436563 , n436491 );
and ( n436565 , n436448 , n436470 );
or ( n436566 , n436564 , n436565 );
buf ( n436567 , n436566 );
buf ( n436568 , n436567 );
xor ( n436569 , n436562 , n436568 );
buf ( n436570 , n436569 );
xor ( n436571 , n436496 , n436570 );
buf ( n436572 , n436571 );
buf ( n436573 , n435511 );
buf ( n436574 , n435541 );
or ( n436575 , n436573 , n436574 );
buf ( n436576 , n435623 );
nand ( n436577 , n436575 , n436576 );
buf ( n436578 , n436577 );
buf ( n436579 , n436578 );
buf ( n436580 , n435511 );
buf ( n436581 , n435541 );
nand ( n436582 , n436580 , n436581 );
buf ( n436583 , n436582 );
buf ( n436584 , n436583 );
and ( n436585 , n436579 , n436584 );
buf ( n436586 , n436585 );
buf ( n436587 , n436586 );
not ( n436588 , n436587 );
buf ( n436589 , n436588 );
buf ( n436590 , n436589 );
not ( n436591 , n436590 );
xor ( n436592 , n436354 , n436368 );
xor ( n436593 , n436592 , n436383 );
buf ( n436594 , n436593 );
not ( n436595 , n436594 );
or ( n436596 , n436591 , n436595 );
buf ( n436597 , n38324 );
not ( n436598 , n436597 );
buf ( n436599 , n385494 );
not ( n436600 , n436599 );
buf ( n436601 , n41359 );
not ( n436602 , n436601 );
or ( n436603 , n436600 , n436602 );
buf ( n436604 , n49938 );
buf ( n436605 , n385491 );
nand ( n436606 , n436604 , n436605 );
buf ( n436607 , n436606 );
buf ( n436608 , n436607 );
nand ( n436609 , n436603 , n436608 );
buf ( n436610 , n436609 );
buf ( n436611 , n436610 );
not ( n436612 , n436611 );
or ( n436613 , n436598 , n436612 );
buf ( n436614 , n435754 );
buf ( n436615 , n385889 );
nand ( n436616 , n436614 , n436615 );
buf ( n436617 , n436616 );
buf ( n436618 , n436617 );
nand ( n436619 , n436613 , n436618 );
buf ( n436620 , n436619 );
buf ( n436621 , n435562 );
buf ( n436622 , n435592 );
not ( n436623 , n436622 );
buf ( n436624 , n389883 );
not ( n436625 , n436624 );
or ( n436626 , n436623 , n436625 );
buf ( n436627 , n389894 );
not ( n436628 , n436627 );
buf ( n436629 , n44423 );
not ( n436630 , n436629 );
or ( n436631 , n436628 , n436630 );
buf ( n436632 , n38155 );
buf ( n436633 , n42390 );
nand ( n436634 , n436632 , n436633 );
buf ( n436635 , n436634 );
buf ( n436636 , n436635 );
nand ( n436637 , n436631 , n436636 );
buf ( n436638 , n436637 );
buf ( n436639 , n436638 );
buf ( n436640 , n389908 );
nand ( n436641 , n436639 , n436640 );
buf ( n436642 , n436641 );
buf ( n436643 , n436642 );
nand ( n436644 , n436626 , n436643 );
buf ( n436645 , n436644 );
buf ( n436646 , n436645 );
xor ( n436647 , n436621 , n436646 );
and ( n436648 , n27196 , n59976 );
not ( n436649 , n27196 );
and ( n436650 , n436649 , n383027 );
or ( n436651 , n436648 , n436650 );
not ( n436652 , n436651 );
not ( n436653 , n386310 );
or ( n436654 , n436652 , n436653 );
not ( n436655 , n435613 );
nand ( n436656 , n436655 , n386300 );
nand ( n436657 , n436654 , n436656 );
buf ( n436658 , n436657 );
not ( n436659 , n436658 );
buf ( n436660 , n436659 );
buf ( n436661 , n436660 );
xor ( n436662 , n436647 , n436661 );
buf ( n436663 , n436662 );
xor ( n436664 , n436620 , n436663 );
xor ( n436665 , n436205 , n436230 );
and ( n436666 , n436665 , n436237 );
and ( n436667 , n436205 , n436230 );
or ( n436668 , n436666 , n436667 );
buf ( n436669 , n436668 );
xnor ( n436670 , n436664 , n436669 );
buf ( n436671 , n436670 );
buf ( n436672 , n436593 );
not ( n436673 , n436672 );
buf ( n436674 , n436586 );
nand ( n436675 , n436673 , n436674 );
buf ( n436676 , n436675 );
buf ( n436677 , n436676 );
nand ( n436678 , n436671 , n436677 );
buf ( n436679 , n436678 );
buf ( n436680 , n436679 );
nand ( n436681 , n436596 , n436680 );
buf ( n436682 , n436681 );
buf ( n436683 , n436682 );
xor ( n436684 , n436572 , n436683 );
buf ( n436685 , n383897 );
not ( n436686 , n436685 );
buf ( n436687 , n436366 );
not ( n436688 , n436687 );
or ( n436689 , n436686 , n436688 );
buf ( n436690 , n36253 );
not ( n436691 , n436690 );
buf ( n436692 , n399538 );
not ( n436693 , n436692 );
or ( n436694 , n436691 , n436693 );
buf ( n436695 , n384741 );
buf ( n436696 , n36252 );
nand ( n436697 , n436695 , n436696 );
buf ( n436698 , n436697 );
buf ( n436699 , n436698 );
nand ( n436700 , n436694 , n436699 );
buf ( n436701 , n436700 );
buf ( n436702 , n436701 );
buf ( n436703 , n384644 );
nand ( n436704 , n436702 , n436703 );
buf ( n436705 , n436704 );
buf ( n436706 , n436705 );
nand ( n436707 , n436689 , n436706 );
buf ( n436708 , n436707 );
buf ( n436709 , n385889 );
not ( n436710 , n436709 );
buf ( n436711 , n436610 );
not ( n436712 , n436711 );
or ( n436713 , n436710 , n436712 );
buf ( n436714 , n385494 );
not ( n436715 , n436714 );
buf ( n436716 , n37027 );
not ( n436717 , n436716 );
or ( n436718 , n436715 , n436717 );
buf ( n436719 , n385834 );
buf ( n436720 , n385491 );
nand ( n436721 , n436719 , n436720 );
buf ( n436722 , n436721 );
buf ( n436723 , n436722 );
nand ( n436724 , n436718 , n436723 );
buf ( n436725 , n436724 );
buf ( n436726 , n436725 );
buf ( n436727 , n38324 );
nand ( n436728 , n436726 , n436727 );
buf ( n436729 , n436728 );
buf ( n436730 , n436729 );
nand ( n436731 , n436713 , n436730 );
buf ( n436732 , n436731 );
not ( n436733 , n436732 );
xor ( n436734 , n436708 , n436733 );
buf ( n436735 , n389777 );
buf ( n436736 , n385292 );
not ( n436737 , n436736 );
buf ( n436738 , n388445 );
not ( n436739 , n436738 );
and ( n436740 , n436737 , n436739 );
buf ( n436741 , n385328 );
buf ( n436742 , n388445 );
and ( n436743 , n436741 , n436742 );
nor ( n436744 , n436740 , n436743 );
buf ( n436745 , n436744 );
buf ( n436746 , n436745 );
or ( n436747 , n436735 , n436746 );
nand ( n436748 , C1 , n436747 );
buf ( n436749 , n436748 );
not ( n436750 , n436749 );
buf ( n436751 , n436750 );
buf ( n436752 , n436651 );
not ( n436753 , n436752 );
buf ( n436754 , n386300 );
not ( n436755 , n436754 );
or ( n436756 , n436753 , n436755 );
buf ( n436757 , n386310 );
buf ( n436758 , n27613 );
not ( n436759 , n436758 );
buf ( n436760 , n59976 );
not ( n436761 , n436760 );
or ( n436762 , n436759 , n436761 );
buf ( n436763 , n386223 );
not ( n436764 , n27613 );
buf ( n436765 , n436764 );
nand ( n436766 , n436763 , n436765 );
buf ( n436767 , n436766 );
buf ( n436768 , n436767 );
nand ( n436769 , n436762 , n436768 );
buf ( n436770 , n436769 );
buf ( n436771 , n436770 );
nand ( n436772 , n436757 , n436771 );
buf ( n436773 , n436772 );
buf ( n436774 , n436773 );
nand ( n436775 , n436756 , n436774 );
buf ( n436776 , n436775 );
buf ( n436777 , n436776 );
xor ( n436778 , n436751 , n436777 );
not ( n436779 , n398406 );
buf ( n436780 , n434637 );
buf ( n436781 , n384186 );
and ( n436782 , n436780 , n436781 );
not ( n436783 , n436780 );
buf ( n436784 , n384211 );
and ( n436785 , n436783 , n436784 );
nor ( n436786 , n436782 , n436785 );
buf ( n436787 , n436786 );
not ( n436788 , n436787 );
or ( n436789 , n436779 , n436788 );
buf ( n436790 , n36399 );
not ( n436791 , n436790 );
buf ( n436792 , n48233 );
not ( n436793 , n436792 );
or ( n436794 , n436791 , n436793 );
buf ( n436795 , n37216 );
buf ( n436796 , n36398 );
nand ( n436797 , n436795 , n436796 );
buf ( n436798 , n436797 );
buf ( n436799 , n436798 );
nand ( n436800 , n436794 , n436799 );
buf ( n436801 , n436800 );
nand ( n436802 , n383946 , n436801 );
nand ( n436803 , n436789 , n436802 );
buf ( n436804 , n436803 );
xor ( n436805 , n436778 , n436804 );
buf ( n436806 , n436805 );
xnor ( n436807 , n436734 , n436806 );
not ( n436808 , n390403 );
buf ( n436809 , n24074 );
buf ( n436810 , n385499 );
and ( n436811 , n436809 , n436810 );
not ( n436812 , n436809 );
buf ( n436813 , n34861 );
and ( n436814 , n436812 , n436813 );
nor ( n436815 , n436811 , n436814 );
buf ( n436816 , n436815 );
not ( n436817 , n436816 );
or ( n436818 , n436808 , n436817 );
buf ( n436819 , n436417 );
buf ( n436820 , n391080 );
nand ( n436821 , n436819 , n436820 );
buf ( n436822 , n436821 );
nand ( n436823 , n436818 , n436822 );
not ( n436824 , n436381 );
not ( n436825 , n436660 );
or ( n436826 , n436824 , n436825 );
nand ( n436827 , n436826 , n436645 );
buf ( n436828 , n436657 );
buf ( n436829 , n435562 );
nand ( n436830 , n436828 , n436829 );
buf ( n436831 , n436830 );
nand ( n436832 , n436827 , n436831 );
xor ( n436833 , n436823 , n436832 );
buf ( n436834 , n383479 );
buf ( n436835 , n436486 );
or ( n436836 , n436834 , n436835 );
buf ( n436837 , n383499 );
buf ( n436838 , n388556 );
buf ( n436839 , n386236 );
and ( n436840 , n436838 , n436839 );
not ( n436841 , n436838 );
buf ( n436842 , n385318 );
not ( n436843 , n436842 );
buf ( n436844 , n436843 );
buf ( n436845 , n436844 );
and ( n436846 , n436841 , n436845 );
nor ( n436847 , n436840 , n436846 );
buf ( n436848 , n436847 );
buf ( n436849 , n436848 );
or ( n436850 , n436837 , n436849 );
nand ( n436851 , n436836 , n436850 );
buf ( n436852 , n436851 );
buf ( n436853 , n436638 );
not ( n436854 , n436853 );
buf ( n436855 , n389883 );
not ( n436856 , n436855 );
or ( n436857 , n436854 , n436856 );
buf ( n436858 , n389894 );
not ( n436859 , n436858 );
buf ( n436860 , n384083 );
not ( n436861 , n436860 );
or ( n436862 , n436859 , n436861 );
buf ( n436863 , n385983 );
buf ( n436864 , n391129 );
nand ( n436865 , n436863 , n436864 );
buf ( n436866 , n436865 );
buf ( n436867 , n436866 );
nand ( n436868 , n436862 , n436867 );
buf ( n436869 , n436868 );
buf ( n436870 , n436869 );
buf ( n436871 , n384554 );
nand ( n436872 , n436870 , n436871 );
buf ( n436873 , n436872 );
buf ( n436874 , n436873 );
nand ( n436875 , n436857 , n436874 );
buf ( n436876 , n436875 );
buf ( n436877 , n436876 );
buf ( n436878 , n382598 );
not ( n436879 , n436878 );
buf ( n436880 , n436879 );
buf ( n436881 , n436880 );
buf ( n436882 , n436461 );
or ( n436883 , n436881 , n436882 );
buf ( n436884 , n379460 );
buf ( n436885 , n436884 );
buf ( n436886 , n386182 );
not ( n436887 , n436886 );
buf ( n436888 , n31964 );
not ( n436889 , n436888 );
and ( n436890 , n436887 , n436889 );
buf ( n436891 , n389997 );
buf ( n436892 , n386182 );
and ( n436893 , n436891 , n436892 );
nor ( n436894 , n436890 , n436893 );
buf ( n436895 , n436894 );
buf ( n436896 , n436895 );
or ( n436897 , n436885 , n436896 );
nand ( n436898 , n436883 , n436897 );
buf ( n436899 , n436898 );
buf ( n436900 , n436899 );
and ( n436901 , n436877 , n436900 );
not ( n436902 , n436877 );
buf ( n436903 , n436899 );
not ( n436904 , n436903 );
buf ( n436905 , n436904 );
buf ( n436906 , n436905 );
and ( n436907 , n436902 , n436906 );
nor ( n436908 , n436901 , n436907 );
buf ( n436909 , n436908 );
xor ( n436910 , n436852 , n436909 );
xor ( n436911 , n436833 , n436910 );
xor ( n436912 , n436807 , n436911 );
buf ( n436913 , n384416 );
not ( n436914 , n436913 );
buf ( n436915 , n436510 );
not ( n436916 , n436915 );
or ( n436917 , n436914 , n436916 );
buf ( n436918 , n435885 );
buf ( n436919 , n384369 );
nand ( n436920 , n436918 , n436919 );
buf ( n436921 , n436920 );
buf ( n436922 , n436921 );
nand ( n436923 , n436917 , n436922 );
buf ( n436924 , n436923 );
not ( n436925 , n436924 );
not ( n436926 , n383946 );
not ( n436927 , n436787 );
or ( n436928 , n436926 , n436927 );
nand ( n436929 , n436197 , n384011 );
nand ( n436930 , n436928 , n436929 );
not ( n436931 , n436930 );
not ( n436932 , n436931 );
or ( n436933 , n436925 , n436932 );
not ( n436934 , n436924 );
nand ( n436935 , n436934 , n436930 );
nand ( n436936 , n436933 , n436935 );
not ( n436937 , n37316 );
not ( n436938 , n436548 );
or ( n436939 , n436937 , n436938 );
buf ( n436940 , n435824 );
buf ( n436941 , n385269 );
nand ( n436942 , n436940 , n436941 );
buf ( n436943 , n436942 );
nand ( n436944 , n436939 , n436943 );
and ( n436945 , n436936 , n436944 );
not ( n436946 , n436936 );
not ( n436947 , n436944 );
and ( n436948 , n436946 , n436947 );
nor ( n436949 , n436945 , n436948 );
not ( n436950 , n436949 );
buf ( n436951 , n386480 );
not ( n436952 , n436951 );
buf ( n436953 , n22982 );
not ( n436954 , n436953 );
buf ( n436955 , n386391 );
not ( n436956 , n436955 );
or ( n436957 , n436954 , n436956 );
buf ( n436958 , n402307 );
buf ( n436959 , n38971 );
nand ( n436960 , n436958 , n436959 );
buf ( n436961 , n436960 );
buf ( n436962 , n436961 );
nand ( n436963 , n436957 , n436962 );
buf ( n436964 , n436963 );
buf ( n436965 , n436964 );
not ( n436966 , n436965 );
or ( n436967 , n436952 , n436966 );
buf ( n436968 , n435504 );
buf ( n436969 , n386496 );
nand ( n436970 , n436968 , n436969 );
buf ( n436971 , n436970 );
buf ( n436972 , n436971 );
nand ( n436973 , n436967 , n436972 );
buf ( n436974 , n436973 );
buf ( n436975 , n436974 );
buf ( n436976 , n389125 );
not ( n436977 , n436976 );
buf ( n436978 , n436170 );
not ( n436979 , n436978 );
or ( n436980 , n436977 , n436979 );
buf ( n436981 , n24050 );
not ( n436982 , n436981 );
buf ( n436983 , n388771 );
not ( n436984 , n436983 );
or ( n436985 , n436982 , n436984 );
buf ( n436986 , n388774 );
buf ( n436987 , n389075 );
nand ( n436988 , n436986 , n436987 );
buf ( n436989 , n436988 );
buf ( n436990 , n436989 );
nand ( n436991 , n436985 , n436990 );
buf ( n436992 , n436991 );
buf ( n436993 , n436992 );
buf ( n436994 , n41565 );
nand ( n436995 , n436993 , n436994 );
buf ( n436996 , n436995 );
buf ( n436997 , n436996 );
nand ( n436998 , n436980 , n436997 );
buf ( n436999 , n436998 );
buf ( n437000 , n436999 );
or ( n437001 , n436975 , n437000 );
buf ( n437002 , n437001 );
not ( n437003 , n437002 );
or ( n437004 , n436950 , n437003 );
buf ( n437005 , n436999 );
buf ( n437006 , n436974 );
and ( n437007 , n437005 , n437006 );
buf ( n437008 , n437007 );
not ( n437009 , n437008 );
nand ( n437010 , n437004 , n437009 );
xor ( n437011 , n436912 , n437010 );
buf ( n437012 , n437011 );
xor ( n437013 , n436684 , n437012 );
buf ( n437014 , n437013 );
buf ( n437015 , n437014 );
not ( n437016 , n435957 );
not ( n437017 , n435954 );
or ( n437018 , n437016 , n437017 );
not ( n437019 , n435953 );
not ( n437020 , n435643 );
or ( n437021 , n437019 , n437020 );
nand ( n437022 , n437021 , n435452 );
nand ( n437023 , n437018 , n437022 );
buf ( n437024 , n437023 );
not ( n437025 , n437024 );
xor ( n437026 , n436156 , n436246 );
and ( n437027 , n437026 , n436252 );
and ( n437028 , n436156 , n436246 );
or ( n437029 , n437027 , n437028 );
buf ( n437030 , n437029 );
not ( n437031 , n437030 );
buf ( n437032 , n437031 );
xor ( n437033 , n437005 , n437006 );
buf ( n437034 , n437033 );
not ( n437035 , n436949 );
and ( n437036 , n437034 , n437035 );
not ( n437037 , n437034 );
and ( n437038 , n437037 , n436949 );
nor ( n437039 , n437036 , n437038 );
xor ( n437040 , n436180 , n436239 );
and ( n437041 , n437040 , n436245 );
and ( n437042 , n436180 , n436239 );
or ( n437043 , n437041 , n437042 );
and ( n437044 , n437039 , n437043 );
not ( n437045 , n437039 );
not ( n437046 , n437043 );
and ( n437047 , n437045 , n437046 );
or ( n437048 , n437044 , n437047 );
not ( n437049 , n435952 );
nand ( n437050 , n435764 , n435798 );
not ( n437051 , n437050 );
or ( n437052 , n437049 , n437051 );
not ( n437053 , n435764 );
nand ( n437054 , n437053 , n435795 );
nand ( n437055 , n437052 , n437054 );
not ( n437056 , n437055 );
and ( n437057 , n437048 , n437056 );
not ( n437058 , n437048 );
and ( n437059 , n437058 , n437055 );
nor ( n437060 , n437057 , n437059 );
nand ( n437061 , n437032 , n437060 );
buf ( n437062 , n437061 );
not ( n437063 , n437062 );
or ( n437064 , n437025 , n437063 );
not ( n437065 , n437060 );
buf ( n437066 , n437065 );
buf ( n437067 , n437029 );
nand ( n437068 , n437066 , n437067 );
buf ( n437069 , n437068 );
buf ( n437070 , n437069 );
nand ( n437071 , n437064 , n437070 );
buf ( n437072 , n437071 );
buf ( n437073 , n437072 );
xor ( n437074 , n437015 , n437073 );
buf ( n437075 , n436669 );
buf ( n437076 , n436620 );
or ( n437077 , n437075 , n437076 );
buf ( n437078 , n436663 );
not ( n437079 , n437078 );
buf ( n437080 , n437079 );
buf ( n437081 , n437080 );
nand ( n437082 , n437077 , n437081 );
buf ( n437083 , n437082 );
buf ( n437084 , n437083 );
buf ( n437085 , n436669 );
buf ( n437086 , n436620 );
nand ( n437087 , n437085 , n437086 );
buf ( n437088 , n437087 );
buf ( n437089 , n437088 );
and ( n437090 , n437084 , n437089 );
buf ( n437091 , n437090 );
buf ( n437092 , n437091 );
not ( n437093 , n436944 );
nand ( n437094 , n436931 , n436934 );
not ( n437095 , n437094 );
or ( n437096 , n437093 , n437095 );
nand ( n437097 , n436924 , n436930 );
nand ( n437098 , n437096 , n437097 );
not ( n437099 , n386496 );
not ( n437100 , n436964 );
or ( n437101 , n437099 , n437100 );
buf ( n437102 , n38972 );
not ( n437103 , n437102 );
buf ( n437104 , n386561 );
not ( n437105 , n437104 );
or ( n437106 , n437103 , n437105 );
buf ( n437107 , n382921 );
buf ( n437108 , n38971 );
nand ( n437109 , n437107 , n437108 );
buf ( n437110 , n437109 );
buf ( n437111 , n437110 );
nand ( n437112 , n437106 , n437111 );
buf ( n437113 , n437112 );
buf ( n437114 , n437113 );
buf ( n437115 , n386480 );
nand ( n437116 , n437114 , n437115 );
buf ( n437117 , n437116 );
nand ( n437118 , n437101 , n437117 );
not ( n437119 , n437118 );
not ( n437120 , n389125 );
not ( n437121 , n436992 );
or ( n437122 , n437120 , n437121 );
buf ( n437123 , n24050 );
not ( n437124 , n437123 );
buf ( n437125 , n38532 );
not ( n437126 , n437125 );
or ( n437127 , n437124 , n437126 );
buf ( n437128 , n35519 );
buf ( n437129 , n389075 );
nand ( n437130 , n437128 , n437129 );
buf ( n437131 , n437130 );
buf ( n437132 , n437131 );
nand ( n437133 , n437127 , n437132 );
buf ( n437134 , n437133 );
buf ( n437135 , n437134 );
buf ( n437136 , n41565 );
nand ( n437137 , n437135 , n437136 );
buf ( n437138 , n437137 );
nand ( n437139 , n437122 , n437138 );
and ( n437140 , n437098 , n437119 , n437139 );
not ( n437141 , n437140 );
not ( n437142 , n437139 );
and ( n437143 , n437098 , n437118 , n437142 );
not ( n437144 , n437098 );
nor ( n437145 , n437118 , n437139 );
and ( n437146 , n437144 , n437145 );
nor ( n437147 , n437143 , n437146 );
nand ( n437148 , n437118 , n437139 , n437144 );
nand ( n437149 , n437141 , n437147 , n437148 );
buf ( n437150 , n437149 );
xor ( n437151 , n437092 , n437150 );
not ( n437152 , n435944 );
not ( n437153 , n435831 );
or ( n437154 , n437152 , n437153 );
not ( n437155 , n435832 );
not ( n437156 , n435943 );
or ( n437157 , n437155 , n437156 );
nand ( n437158 , n437157 , n435805 );
nand ( n437159 , n437154 , n437158 );
not ( n437160 , n437159 );
not ( n437161 , n437160 );
not ( n437162 , n435684 );
not ( n437163 , n435722 );
or ( n437164 , n437162 , n437163 );
not ( n437165 , n435685 );
not ( n437166 , n435725 );
or ( n437167 , n437165 , n437166 );
nand ( n437168 , n437167 , n435759 );
nand ( n437169 , n437164 , n437168 );
buf ( n437170 , n437169 );
not ( n437171 , n437170 );
buf ( n437172 , n437171 );
not ( n437173 , n437172 );
and ( n437174 , n437161 , n437173 );
not ( n437175 , n436493 );
and ( n437176 , n436402 , n436427 );
not ( n437177 , n436402 );
and ( n437178 , n437177 , n436432 );
nor ( n437179 , n437176 , n437178 );
not ( n437180 , n437179 );
not ( n437181 , n437180 );
or ( n437182 , n437175 , n437181 );
not ( n437183 , n436493 );
nand ( n437184 , n437183 , n437179 );
nand ( n437185 , n437182 , n437184 );
or ( n437186 , n437159 , n437169 );
and ( n437187 , n437185 , n437186 );
nor ( n437188 , n437174 , n437187 );
buf ( n437189 , n437188 );
xor ( n437190 , n437151 , n437189 );
buf ( n437191 , n437190 );
buf ( n437192 , n437191 );
not ( n437193 , n437046 );
not ( n437194 , n437039 );
and ( n437195 , n437193 , n437194 );
nand ( n437196 , n437046 , n437039 );
and ( n437197 , n437055 , n437196 );
nor ( n437198 , n437195 , n437197 );
buf ( n437199 , n437198 );
and ( n437200 , n437192 , n437199 );
not ( n437201 , n437192 );
buf ( n437202 , n437198 );
not ( n437203 , n437202 );
buf ( n437204 , n437203 );
buf ( n437205 , n437204 );
and ( n437206 , n437201 , n437205 );
nor ( n437207 , n437200 , n437206 );
buf ( n437208 , n437207 );
buf ( n437209 , n437208 );
buf ( n437210 , n437169 );
not ( n437211 , n437210 );
buf ( n437212 , n437160 );
not ( n437213 , n437212 );
or ( n437214 , n437211 , n437213 );
buf ( n437215 , n437159 );
buf ( n437216 , n437172 );
nand ( n437217 , n437215 , n437216 );
buf ( n437218 , n437217 );
buf ( n437219 , n437218 );
nand ( n437220 , n437214 , n437219 );
buf ( n437221 , n437220 );
not ( n437222 , n437185 );
and ( n437223 , n437221 , n437222 );
not ( n437224 , n437221 );
and ( n437225 , n437224 , n437185 );
nor ( n437226 , n437223 , n437225 );
buf ( n437227 , n437226 );
not ( n437228 , n437227 );
xor ( n437229 , n436593 , n436586 );
xor ( n437230 , n437229 , n436670 );
buf ( n437231 , n437230 );
not ( n437232 , n437231 );
or ( n437233 , n437228 , n437232 );
not ( n437234 , n435497 );
buf ( n437235 , n435636 );
not ( n437236 , n437235 );
or ( n437237 , n437234 , n437236 );
or ( n437238 , n437235 , n435497 );
nand ( n437239 , n437238 , n435642 );
nand ( n437240 , n437237 , n437239 );
buf ( n437241 , n437240 );
nand ( n437242 , n437233 , n437241 );
buf ( n437243 , n437242 );
buf ( n437244 , n437243 );
buf ( n437245 , n437226 );
not ( n437246 , n437245 );
buf ( n437247 , n437230 );
not ( n437248 , n437247 );
buf ( n437249 , n437248 );
buf ( n437250 , n437249 );
nand ( n437251 , n437246 , n437250 );
buf ( n437252 , n437251 );
buf ( n437253 , n437252 );
nand ( n437254 , n437244 , n437253 );
buf ( n437255 , n437254 );
buf ( n437256 , n437255 );
xor ( n437257 , n437209 , n437256 );
buf ( n437258 , n437257 );
buf ( n437259 , n437258 );
xor ( n437260 , n437074 , n437259 );
buf ( n437261 , n437260 );
not ( n437262 , n437261 );
not ( n437263 , n437240 );
and ( n437264 , n437226 , n437263 );
not ( n437265 , n437226 );
and ( n437266 , n437265 , n437240 );
nor ( n437267 , n437264 , n437266 );
and ( n437268 , n437267 , n437230 );
not ( n437269 , n437267 );
and ( n437270 , n437269 , n437249 );
nor ( n437271 , n437268 , n437270 );
not ( n437272 , n437029 );
not ( n437273 , n437060 );
or ( n437274 , n437272 , n437273 );
buf ( n437275 , n437065 );
buf ( n437276 , n437032 );
nand ( n437277 , n437275 , n437276 );
buf ( n437278 , n437277 );
nand ( n437279 , n437274 , n437278 );
not ( n437280 , n437023 );
and ( n437281 , n437279 , n437280 );
not ( n437282 , n437279 );
and ( n437283 , n437282 , n437023 );
nor ( n437284 , n437281 , n437283 );
xor ( n437285 , n437271 , n437284 );
buf ( n437286 , n436061 );
buf ( n437287 , n436147 );
not ( n437288 , n437287 );
buf ( n437289 , n436256 );
nand ( n437290 , n437288 , n437289 );
buf ( n437291 , n437290 );
buf ( n437292 , n437291 );
and ( n437293 , n437286 , n437292 );
buf ( n437294 , n436147 );
not ( n437295 , n437294 );
buf ( n437296 , n436256 );
nor ( n437297 , n437295 , n437296 );
buf ( n437298 , n437297 );
buf ( n437299 , n437298 );
nor ( n437300 , n437293 , n437299 );
buf ( n437301 , n437300 );
and ( n437302 , n437285 , n437301 );
and ( n437303 , n437271 , n437284 );
or ( n437304 , n437302 , n437303 );
nand ( n437305 , n437262 , n437304 );
not ( n437306 , n437305 );
not ( n437307 , n436305 );
buf ( n437308 , n435963 );
not ( n437309 , n437308 );
buf ( n437310 , n437309 );
not ( n437311 , n437310 );
and ( n437312 , n437307 , n437311 );
buf ( n437313 , n436305 );
buf ( n437314 , n437310 );
nand ( n437315 , n437313 , n437314 );
buf ( n437316 , n437315 );
buf ( n437317 , n436273 );
not ( n437318 , n437317 );
buf ( n437319 , n437318 );
and ( n437320 , n437316 , n437319 );
nor ( n437321 , n437312 , n437320 );
xor ( n437322 , n437271 , n437284 );
xor ( n437323 , n437322 , n437301 );
nand ( n437324 , n437321 , n437323 );
not ( n437325 , n437324 );
nor ( n437326 , n436350 , n437306 , n437325 );
xor ( n437327 , n437015 , n437073 );
and ( n437328 , n437327 , n437259 );
and ( n437329 , n437015 , n437073 );
or ( n437330 , n437328 , n437329 );
buf ( n437331 , n437330 );
not ( n437332 , n437331 );
xor ( n437333 , n436534 , n436561 );
and ( n437334 , n437333 , n436568 );
and ( n437335 , n436534 , n436561 );
or ( n437336 , n437334 , n437335 );
buf ( n437337 , n437336 );
buf ( n437338 , n437337 );
not ( n437339 , n437338 );
buf ( n437340 , n437339 );
buf ( n437341 , n437340 );
not ( n437342 , n437341 );
buf ( n437343 , n384557 );
not ( n437344 , n437343 );
buf ( n437345 , n42390 );
buf ( n437346 , n390172 );
and ( n437347 , n437345 , n437346 );
not ( n437348 , n437345 );
buf ( n437349 , n398327 );
and ( n437350 , n437348 , n437349 );
nor ( n437351 , n437347 , n437350 );
buf ( n437352 , n437351 );
buf ( n437353 , n437352 );
not ( n437354 , n437353 );
or ( n437355 , n437344 , n437354 );
buf ( n437356 , n384627 );
buf ( n437357 , n436869 );
nand ( n437358 , n437356 , n437357 );
buf ( n437359 , n437358 );
buf ( n437360 , n437359 );
nand ( n437361 , n437355 , n437360 );
buf ( n437362 , n437361 );
not ( n437363 , n383897 );
not ( n437364 , n436701 );
or ( n437365 , n437363 , n437364 );
buf ( n437366 , n36253 );
not ( n437367 , n437366 );
buf ( n437368 , n38357 );
not ( n437369 , n437368 );
or ( n437370 , n437367 , n437369 );
buf ( n437371 , n51163 );
buf ( n437372 , n36252 );
nand ( n437373 , n437371 , n437372 );
buf ( n437374 , n437373 );
buf ( n437375 , n437374 );
nand ( n437376 , n437370 , n437375 );
buf ( n437377 , n437376 );
nand ( n437378 , n437377 , n384644 );
nand ( n437379 , n437365 , n437378 );
xor ( n437380 , n437362 , n437379 );
buf ( n437381 , n436899 );
not ( n437382 , n437381 );
buf ( n437383 , n436876 );
not ( n437384 , n437383 );
or ( n437385 , n437382 , n437384 );
buf ( n437386 , n436905 );
not ( n437387 , n437386 );
buf ( n437388 , n436876 );
not ( n437389 , n437388 );
buf ( n437390 , n437389 );
buf ( n437391 , n437390 );
not ( n437392 , n437391 );
or ( n437393 , n437387 , n437392 );
buf ( n437394 , n436852 );
nand ( n437395 , n437393 , n437394 );
buf ( n437396 , n437395 );
buf ( n437397 , n437396 );
nand ( n437398 , n437385 , n437397 );
buf ( n437399 , n437398 );
xnor ( n437400 , n437380 , n437399 );
buf ( n437401 , n437400 );
not ( n437402 , n437401 );
buf ( n437403 , n437402 );
buf ( n437404 , n437403 );
not ( n437405 , n437404 );
or ( n437406 , n437342 , n437405 );
buf ( n437407 , n437400 );
buf ( n437408 , n437337 );
nand ( n437409 , n437407 , n437408 );
buf ( n437410 , n437409 );
buf ( n437411 , n437410 );
nand ( n437412 , n437406 , n437411 );
buf ( n437413 , n437412 );
xor ( n437414 , n436823 , n436832 );
and ( n437415 , n437414 , n436910 );
and ( n437416 , n436823 , n436832 );
or ( n437417 , n437415 , n437416 );
and ( n437418 , n437413 , n437417 );
not ( n437419 , n437413 );
not ( n437420 , n437417 );
and ( n437421 , n437419 , n437420 );
nor ( n437422 , n437418 , n437421 );
buf ( n437423 , n437422 );
buf ( n437424 , n41565 );
not ( n437425 , n437424 );
buf ( n437426 , n24050 );
not ( n437427 , n437426 );
buf ( n437428 , n390351 );
not ( n437429 , n437428 );
or ( n437430 , n437427 , n437429 );
buf ( n437431 , n382532 );
buf ( n437432 , n389075 );
nand ( n437433 , n437431 , n437432 );
buf ( n437434 , n437433 );
buf ( n437435 , n437434 );
nand ( n437436 , n437430 , n437435 );
buf ( n437437 , n437436 );
buf ( n437438 , n437437 );
not ( n437439 , n437438 );
or ( n437440 , n437425 , n437439 );
buf ( n437441 , n437134 );
buf ( n437442 , n389125 );
nand ( n437443 , n437441 , n437442 );
buf ( n437444 , n437443 );
buf ( n437445 , n437444 );
nand ( n437446 , n437440 , n437445 );
buf ( n437447 , n437446 );
buf ( n437448 , n437447 );
buf ( n437449 , n383946 );
not ( n437450 , n437449 );
buf ( n437451 , n434637 );
not ( n437452 , n437451 );
buf ( n437453 , n383762 );
not ( n437454 , n437453 );
or ( n437455 , n437452 , n437454 );
buf ( n437456 , n42152 );
buf ( n437457 , n36398 );
nand ( n437458 , n437456 , n437457 );
buf ( n437459 , n437458 );
buf ( n437460 , n437459 );
nand ( n437461 , n437455 , n437460 );
buf ( n437462 , n437461 );
buf ( n437463 , n437462 );
not ( n437464 , n437463 );
or ( n437465 , n437450 , n437464 );
buf ( n437466 , n436801 );
buf ( n437467 , n384011 );
nand ( n437468 , n437466 , n437467 );
buf ( n437469 , n437468 );
buf ( n437470 , n437469 );
nand ( n437471 , n437465 , n437470 );
buf ( n437472 , n437471 );
buf ( n437473 , n437472 );
xor ( n437474 , n437448 , n437473 );
buf ( n437475 , n389547 );
buf ( n437476 , n42825 );
not ( n437477 , n437476 );
buf ( n437478 , n384143 );
not ( n437479 , n437478 );
or ( n437480 , n437477 , n437479 );
buf ( n437481 , n385292 );
buf ( n437482 , n74955 );
nand ( n437483 , n437481 , n437482 );
buf ( n437484 , n437483 );
buf ( n437485 , n437484 );
nand ( n437486 , n437480 , n437485 );
buf ( n437487 , n437486 );
buf ( n437488 , n437487 );
nand ( n437489 , n437475 , n437488 );
buf ( n437490 , n437489 );
buf ( n437491 , n437490 );
nand ( n437492 , C1 , n437491 );
buf ( n437493 , n437492 );
buf ( n437494 , n437493 );
not ( n437495 , n389024 );
buf ( n437496 , n31964 );
not ( n437497 , n437496 );
buf ( n437498 , n385345 );
not ( n437499 , n437498 );
or ( n437500 , n437497 , n437499 );
buf ( n437501 , n385359 );
buf ( n437502 , n385972 );
nand ( n437503 , n437501 , n437502 );
buf ( n437504 , n437503 );
buf ( n437505 , n437504 );
nand ( n437506 , n437500 , n437505 );
buf ( n437507 , n437506 );
not ( n437508 , n437507 );
or ( n437509 , n437495 , n437508 );
not ( n437510 , n436895 );
nand ( n437511 , n437510 , n382598 );
nand ( n437512 , n437509 , n437511 );
buf ( n437513 , n437512 );
xor ( n437514 , n437494 , n437513 );
buf ( n437515 , n391920 );
buf ( n437516 , n436848 );
or ( n437517 , n437515 , n437516 );
and ( n437518 , n38159 , n434951 );
not ( n437519 , n38159 );
and ( n437520 , n437519 , n388576 );
nor ( n437521 , n437518 , n437520 );
buf ( n437522 , n437521 );
buf ( n437523 , n391176 );
or ( n437524 , n437522 , n437523 );
nand ( n437525 , n437517 , n437524 );
buf ( n437526 , n437525 );
buf ( n437527 , n437526 );
xor ( n437528 , n437514 , n437527 );
buf ( n437529 , n437528 );
buf ( n437530 , n437529 );
xor ( n437531 , n437474 , n437530 );
buf ( n437532 , n437531 );
buf ( n437533 , n437532 );
not ( n437534 , n436806 );
not ( n437535 , n436708 );
nand ( n437536 , n437535 , n436733 );
not ( n437537 , n437536 );
or ( n437538 , n437534 , n437537 );
nand ( n437539 , n436732 , n436708 );
nand ( n437540 , n437538 , n437539 );
buf ( n437541 , n437540 );
and ( n437542 , n437533 , n437541 );
not ( n437543 , n437533 );
buf ( n437544 , n437540 );
not ( n437545 , n437544 );
buf ( n437546 , n437545 );
buf ( n437547 , n437546 );
and ( n437548 , n437543 , n437547 );
nor ( n437549 , n437542 , n437548 );
buf ( n437550 , n437549 );
buf ( n437551 , n437550 );
buf ( n437552 , n42925 );
not ( n437553 , n437552 );
buf ( n437554 , n390435 );
not ( n437555 , n437554 );
or ( n437556 , n437553 , n437555 );
buf ( n437557 , n436816 );
nand ( n437558 , n437556 , n437557 );
buf ( n437559 , n437558 );
xor ( n437560 , n436751 , n436777 );
and ( n437561 , n437560 , n436804 );
and ( n437562 , n436751 , n436777 );
or ( n437563 , n437561 , n437562 );
buf ( n437564 , n437563 );
xor ( n437565 , n437559 , n437564 );
buf ( n437566 , n436770 );
not ( n437567 , n437566 );
buf ( n437568 , n396868 );
not ( n437569 , n437568 );
or ( n437570 , n437567 , n437569 );
buf ( n437571 , n386310 );
and ( n437572 , n390271 , n386223 );
not ( n437573 , n390271 );
and ( n437574 , n437573 , n398740 );
or ( n437575 , n437572 , n437574 );
buf ( n437576 , n437575 );
nand ( n437577 , n437571 , n437576 );
buf ( n437578 , n437577 );
buf ( n437579 , n437578 );
nand ( n437580 , n437570 , n437579 );
buf ( n437581 , n437580 );
xor ( n437582 , n437581 , n436750 );
buf ( n437583 , n36821 );
buf ( n437584 , n384211 );
and ( n437585 , n437583 , n437584 );
not ( n437586 , n437583 );
buf ( n437587 , n385740 );
and ( n437588 , n437586 , n437587 );
nor ( n437589 , n437585 , n437588 );
buf ( n437590 , n437589 );
buf ( n437591 , n437590 );
buf ( n437592 , n386770 );
or ( n437593 , n437591 , n437592 );
buf ( n437594 , n436526 );
buf ( n437595 , n384369 );
nand ( n437596 , n437594 , n437595 );
buf ( n437597 , n437596 );
buf ( n437598 , n437597 );
nand ( n437599 , n437593 , n437598 );
buf ( n437600 , n437599 );
xnor ( n437601 , n437582 , n437600 );
xor ( n437602 , n437565 , n437601 );
buf ( n437603 , n437602 );
not ( n437604 , n437603 );
buf ( n437605 , n437604 );
buf ( n437606 , n437605 );
and ( n437607 , n437551 , n437606 );
not ( n437608 , n437551 );
buf ( n437609 , n437602 );
and ( n437610 , n437608 , n437609 );
nor ( n437611 , n437607 , n437610 );
buf ( n437612 , n437611 );
buf ( n437613 , n437612 );
xor ( n437614 , n437423 , n437613 );
not ( n437615 , n436807 );
not ( n437616 , n436911 );
nor ( n437617 , n437615 , n437616 );
or ( n437618 , n437617 , n437010 );
not ( n437619 , n436911 );
nand ( n437620 , n437619 , n437615 );
nand ( n437621 , n437618 , n437620 );
buf ( n437622 , n437621 );
xnor ( n437623 , n437614 , n437622 );
buf ( n437624 , n437623 );
buf ( n437625 , n437624 );
buf ( n437626 , n437198 );
not ( n437627 , n437626 );
buf ( n437628 , n437191 );
not ( n437629 , n437628 );
or ( n437630 , n437627 , n437629 );
buf ( n437631 , n437255 );
nand ( n437632 , n437630 , n437631 );
buf ( n437633 , n437632 );
buf ( n437634 , n437633 );
buf ( n437635 , n437191 );
not ( n437636 , n437635 );
buf ( n437637 , n437204 );
nand ( n437638 , n437636 , n437637 );
buf ( n437639 , n437638 );
buf ( n437640 , n437639 );
and ( n437641 , n437634 , n437640 );
buf ( n437642 , n437641 );
buf ( n437643 , n437642 );
xor ( n437644 , n437625 , n437643 );
buf ( n437645 , n37316 );
not ( n437646 , n437645 );
buf ( n437647 , n37347 );
not ( n437648 , n437647 );
buf ( n437649 , n41359 );
not ( n437650 , n437649 );
or ( n437651 , n437648 , n437650 );
nand ( n437652 , n37370 , n37354 );
buf ( n437653 , n437652 );
nand ( n437654 , n437651 , n437653 );
buf ( n437655 , n437654 );
buf ( n437656 , n437655 );
not ( n437657 , n437656 );
or ( n437658 , n437646 , n437657 );
buf ( n437659 , n436556 );
buf ( n437660 , n385269 );
nand ( n437661 , n437659 , n437660 );
buf ( n437662 , n437661 );
buf ( n437663 , n437662 );
nand ( n437664 , n437658 , n437663 );
buf ( n437665 , n437664 );
buf ( n437666 , n437665 );
buf ( n437667 , n38324 );
not ( n437668 , n437667 );
buf ( n437669 , n385494 );
not ( n437670 , n437669 );
buf ( n437671 , n386385 );
not ( n437672 , n437671 );
or ( n437673 , n437670 , n437672 );
buf ( n437674 , n35301 );
buf ( n437675 , n385491 );
nand ( n437676 , n437674 , n437675 );
buf ( n437677 , n437676 );
buf ( n437678 , n437677 );
nand ( n437679 , n437673 , n437678 );
buf ( n437680 , n437679 );
buf ( n437681 , n437680 );
not ( n437682 , n437681 );
or ( n437683 , n437668 , n437682 );
buf ( n437684 , n436725 );
buf ( n437685 , n385889 );
nand ( n437686 , n437684 , n437685 );
buf ( n437687 , n437686 );
buf ( n437688 , n437687 );
nand ( n437689 , n437683 , n437688 );
buf ( n437690 , n437689 );
buf ( n437691 , n437690 );
xor ( n437692 , n437666 , n437691 );
buf ( n437693 , n437113 );
buf ( n437694 , n386496 );
and ( n437695 , n437693 , n437694 );
buf ( n437696 , n22982 );
not ( n437697 , n437696 );
buf ( n437698 , n386421 );
not ( n437699 , n437698 );
or ( n437700 , n437697 , n437699 );
buf ( n437701 , n386418 );
buf ( n437702 , n38971 );
nand ( n437703 , n437701 , n437702 );
buf ( n437704 , n437703 );
buf ( n437705 , n437704 );
nand ( n437706 , n437700 , n437705 );
buf ( n437707 , n437706 );
buf ( n437708 , n437707 );
not ( n437709 , n437708 );
buf ( n437710 , n386483 );
nor ( n437711 , n437709 , n437710 );
buf ( n437712 , n437711 );
buf ( n437713 , n437712 );
nor ( n437714 , n437695 , n437713 );
buf ( n437715 , n437714 );
buf ( n437716 , n437715 );
not ( n437717 , n437716 );
buf ( n437718 , n437717 );
buf ( n437719 , n437718 );
xnor ( n437720 , n437692 , n437719 );
buf ( n437721 , n437720 );
buf ( n437722 , n437721 );
not ( n437723 , n437722 );
buf ( n437724 , n437723 );
buf ( n437725 , n437724 );
not ( n437726 , n437725 );
or ( n437727 , n437144 , n437145 );
nand ( n437728 , n437118 , n437139 );
nand ( n437729 , n437727 , n437728 );
buf ( n437730 , n437729 );
not ( n437731 , n437730 );
buf ( n437732 , n437731 );
buf ( n437733 , n437732 );
not ( n437734 , n437733 );
or ( n437735 , n437726 , n437734 );
buf ( n437736 , n437721 );
buf ( n437737 , n437729 );
nand ( n437738 , n437736 , n437737 );
buf ( n437739 , n437738 );
buf ( n437740 , n437739 );
nand ( n437741 , n437735 , n437740 );
buf ( n437742 , n437741 );
buf ( n437743 , n437742 );
xor ( n437744 , n436386 , n436495 );
and ( n437745 , n437744 , n436570 );
and ( n437746 , n436386 , n436495 );
or ( n437747 , n437745 , n437746 );
buf ( n437748 , n437747 );
and ( n437749 , n437743 , n437748 );
not ( n437750 , n437743 );
buf ( n437751 , n437747 );
not ( n437752 , n437751 );
buf ( n437753 , n437752 );
buf ( n437754 , n437753 );
and ( n437755 , n437750 , n437754 );
nor ( n437756 , n437749 , n437755 );
buf ( n437757 , n437756 );
xor ( n437758 , n437092 , n437150 );
and ( n437759 , n437758 , n437189 );
and ( n437760 , n437092 , n437150 );
or ( n437761 , n437759 , n437760 );
buf ( n437762 , n437761 );
xor ( n437763 , n437757 , n437762 );
xor ( n437764 , n436572 , n436683 );
and ( n437765 , n437764 , n437012 );
and ( n437766 , n436572 , n436683 );
or ( n437767 , n437765 , n437766 );
buf ( n437768 , n437767 );
xor ( n437769 , n437763 , n437768 );
buf ( n437770 , n437769 );
xor ( n437771 , n437644 , n437770 );
buf ( n437772 , n437771 );
nand ( n437773 , n437332 , n437772 );
buf ( n437774 , n385494 );
buf ( n437775 , n386561 );
and ( n437776 , n437774 , n437775 );
not ( n437777 , n437774 );
buf ( n437778 , n382921 );
and ( n437779 , n437777 , n437778 );
nor ( n437780 , n437776 , n437779 );
buf ( n437781 , n437780 );
buf ( n437782 , n437781 );
not ( n437783 , n437782 );
buf ( n437784 , n37924 );
not ( n437785 , n437784 );
and ( n437786 , n437783 , n437785 );
buf ( n437787 , n437680 );
buf ( n437788 , n385889 );
and ( n437789 , n437787 , n437788 );
nor ( n437790 , n437786 , n437789 );
buf ( n437791 , n437790 );
not ( n437792 , n437362 );
not ( n437793 , n437792 );
not ( n437794 , n437379 );
not ( n437795 , n437794 );
or ( n437796 , n437793 , n437795 );
nand ( n437797 , n437796 , n437399 );
nand ( n437798 , n437362 , n437379 );
nand ( n437799 , n437797 , n437798 );
xor ( n437800 , n437791 , n437799 );
xor ( n437801 , n437448 , n437473 );
and ( n437802 , n437801 , n437530 );
and ( n437803 , n437448 , n437473 );
or ( n437804 , n437802 , n437803 );
buf ( n437805 , n437804 );
xnor ( n437806 , n437800 , n437805 );
buf ( n437807 , n437532 );
not ( n437808 , n437807 );
buf ( n437809 , n437540 );
not ( n437810 , n437809 );
or ( n437811 , n437808 , n437810 );
buf ( n437812 , n437540 );
buf ( n437813 , n437532 );
or ( n437814 , n437812 , n437813 );
buf ( n437815 , n437602 );
nand ( n437816 , n437814 , n437815 );
buf ( n437817 , n437816 );
buf ( n437818 , n437817 );
nand ( n437819 , n437811 , n437818 );
buf ( n437820 , n437819 );
xor ( n437821 , n437806 , n437820 );
xor ( n437822 , n437494 , n437513 );
and ( n437823 , n437822 , n437527 );
and ( n437824 , n437494 , n437513 );
or ( n437825 , n437823 , n437824 );
buf ( n437826 , n437825 );
buf ( n437827 , n437826 );
buf ( n437828 , n389125 );
not ( n437829 , n437828 );
buf ( n437830 , n437437 );
not ( n437831 , n437830 );
or ( n437832 , n437829 , n437831 );
buf ( n437833 , n24050 );
not ( n437834 , n437833 );
buf ( n437835 , n385502 );
not ( n437836 , n437835 );
or ( n437837 , n437834 , n437836 );
buf ( n437838 , n388113 );
not ( n437839 , n437838 );
buf ( n437840 , n389075 );
nand ( n437841 , n437839 , n437840 );
buf ( n437842 , n437841 );
buf ( n437843 , n437842 );
nand ( n437844 , n437837 , n437843 );
buf ( n437845 , n437844 );
buf ( n437846 , n437845 );
buf ( n437847 , n41565 );
nand ( n437848 , n437846 , n437847 );
buf ( n437849 , n437848 );
buf ( n437850 , n437849 );
nand ( n437851 , n437832 , n437850 );
buf ( n437852 , n437851 );
buf ( n437853 , n437852 );
xor ( n437854 , n437827 , n437853 );
buf ( n437855 , n383897 );
not ( n437856 , n437855 );
buf ( n437857 , n437377 );
not ( n437858 , n437857 );
or ( n437859 , n437856 , n437858 );
buf ( n437860 , n36253 );
not ( n437861 , n437860 );
buf ( n437862 , n36900 );
not ( n437863 , n437862 );
or ( n437864 , n437861 , n437863 );
buf ( n437865 , n38227 );
buf ( n437866 , n36252 );
nand ( n437867 , n437865 , n437866 );
buf ( n437868 , n437867 );
buf ( n437869 , n437868 );
nand ( n437870 , n437864 , n437869 );
buf ( n437871 , n437870 );
buf ( n437872 , n437871 );
buf ( n437873 , n384644 );
nand ( n437874 , n437872 , n437873 );
buf ( n437875 , n437874 );
buf ( n437876 , n437875 );
nand ( n437877 , n437859 , n437876 );
buf ( n437878 , n437877 );
buf ( n437879 , n437878 );
xor ( n437880 , n437854 , n437879 );
buf ( n437881 , n437880 );
buf ( n437882 , n437881 );
buf ( n437883 , n384011 );
not ( n437884 , n437883 );
buf ( n437885 , n437462 );
not ( n437886 , n437885 );
or ( n437887 , n437884 , n437886 );
buf ( n437888 , n434637 );
not ( n437889 , n437888 );
buf ( n437890 , n389525 );
not ( n437891 , n437890 );
or ( n437892 , n437889 , n437891 );
buf ( n437893 , n384741 );
buf ( n437894 , n36398 );
nand ( n437895 , n437893 , n437894 );
buf ( n437896 , n437895 );
buf ( n437897 , n437896 );
nand ( n437898 , n437892 , n437897 );
buf ( n437899 , n437898 );
buf ( n437900 , n437899 );
buf ( n437901 , n383946 );
nand ( n437902 , n437900 , n437901 );
buf ( n437903 , n437902 );
buf ( n437904 , n437903 );
nand ( n437905 , n437887 , n437904 );
buf ( n437906 , n437905 );
buf ( n437907 , n437906 );
buf ( n437908 , n386496 );
not ( n437909 , n437908 );
buf ( n437910 , n437707 );
not ( n437911 , n437910 );
or ( n437912 , n437909 , n437911 );
buf ( n437913 , n38972 );
not ( n437914 , n437913 );
buf ( n437915 , n38532 );
not ( n437916 , n437915 );
or ( n437917 , n437914 , n437916 );
buf ( n437918 , n383111 );
buf ( n437919 , n38971 );
nand ( n437920 , n437918 , n437919 );
buf ( n437921 , n437920 );
buf ( n437922 , n437921 );
nand ( n437923 , n437917 , n437922 );
buf ( n437924 , n437923 );
buf ( n437925 , n437924 );
buf ( n437926 , n386480 );
nand ( n437927 , n437925 , n437926 );
buf ( n437928 , n437927 );
buf ( n437929 , n437928 );
nand ( n437930 , n437912 , n437929 );
buf ( n437931 , n437930 );
buf ( n437932 , n437931 );
xor ( n437933 , n437907 , n437932 );
buf ( n437934 , n437507 );
not ( n437935 , n437934 );
buf ( n437936 , n382598 );
not ( n437937 , n437936 );
or ( n437938 , n437935 , n437937 );
buf ( n437939 , n385975 );
buf ( n437940 , n386236 );
and ( n437941 , n437939 , n437940 );
not ( n437942 , n437939 );
buf ( n437943 , n385324 );
and ( n437944 , n437942 , n437943 );
nor ( n437945 , n437941 , n437944 );
buf ( n437946 , n437945 );
buf ( n437947 , n437946 );
not ( n437948 , n437947 );
buf ( n437949 , n379466 );
nand ( n437950 , n437948 , n437949 );
buf ( n437951 , n437950 );
buf ( n437952 , n437951 );
nand ( n437953 , n437938 , n437952 );
buf ( n437954 , n437953 );
buf ( n437955 , n437954 );
not ( n437956 , n59976 );
not ( n437957 , n435919 );
or ( n437958 , n437956 , n437957 );
buf ( n437959 , n384965 );
buf ( n437960 , n386182 );
nand ( n437961 , n437959 , n437960 );
buf ( n437962 , n437961 );
nand ( n437963 , n437958 , n437962 );
not ( n437964 , n437963 );
not ( n437965 , n386310 );
or ( n437966 , n437964 , n437965 );
nand ( n437967 , n386300 , n437575 );
nand ( n437968 , n437966 , n437967 );
buf ( n437969 , n437968 );
xor ( n437970 , n437955 , n437969 );
buf ( n437971 , n383479 );
buf ( n437972 , n437521 );
or ( n437973 , n437971 , n437972 );
buf ( n437974 , n383426 );
buf ( n437975 , n384092 );
and ( n437976 , n437974 , n437975 );
not ( n437977 , n437974 );
buf ( n437978 , n389485 );
and ( n437979 , n437977 , n437978 );
nor ( n437980 , n437976 , n437979 );
buf ( n437981 , n437980 );
buf ( n437982 , n437981 );
buf ( n437983 , n383403 );
or ( n437984 , n437982 , n437983 );
nand ( n437985 , n437973 , n437984 );
buf ( n437986 , n437985 );
buf ( n437987 , n437986 );
xor ( n437988 , n437970 , n437987 );
buf ( n437989 , n437988 );
buf ( n437990 , n437989 );
xor ( n437991 , n437933 , n437990 );
buf ( n437992 , n437991 );
buf ( n437993 , n437992 );
xor ( n437994 , n437882 , n437993 );
xor ( n437995 , n437559 , n437564 );
and ( n437996 , n437995 , n437601 );
and ( n437997 , n437559 , n437564 );
or ( n437998 , n437996 , n437997 );
buf ( n437999 , n437998 );
xor ( n438000 , n437994 , n437999 );
buf ( n438001 , n438000 );
xnor ( n438002 , n437821 , n438001 );
buf ( n438003 , n438002 );
not ( n438004 , n437724 );
not ( n438005 , n437729 );
or ( n438006 , n438004 , n438005 );
not ( n438007 , n437721 );
not ( n438008 , n437732 );
or ( n438009 , n438007 , n438008 );
nand ( n438010 , n438009 , n437747 );
nand ( n438011 , n438006 , n438010 );
not ( n438012 , n437581 );
nand ( n438013 , n436750 , n438012 );
and ( n438014 , n437600 , n438013 );
nor ( n438015 , n436750 , n438012 );
nor ( n438016 , n438014 , n438015 );
not ( n438017 , n438016 );
buf ( n438018 , n385269 );
not ( n438019 , n438018 );
buf ( n438020 , n437655 );
not ( n438021 , n438020 );
or ( n438022 , n438019 , n438021 );
buf ( n438023 , n37347 );
not ( n438024 , n438023 );
buf ( n438025 , n37027 );
not ( n438026 , n438025 );
or ( n438027 , n438024 , n438026 );
buf ( n438028 , n385834 );
buf ( n438029 , n37354 );
nand ( n438030 , n438028 , n438029 );
buf ( n438031 , n438030 );
buf ( n438032 , n438031 );
nand ( n438033 , n438027 , n438032 );
buf ( n438034 , n438033 );
buf ( n438035 , n438034 );
buf ( n438036 , n37695 );
nand ( n438037 , n438035 , n438036 );
buf ( n438038 , n438037 );
buf ( n438039 , n438038 );
nand ( n438040 , n438022 , n438039 );
buf ( n438041 , n438040 );
and ( n438042 , n438017 , n438041 );
not ( n438043 , n438017 );
not ( n438044 , n438041 );
and ( n438045 , n438043 , n438044 );
nor ( n438046 , n438042 , n438045 );
not ( n438047 , n382944 );
buf ( n438048 , n382857 );
not ( n438049 , n438048 );
buf ( n438050 , n436764 );
not ( n438051 , n438050 );
and ( n438052 , n438049 , n438051 );
buf ( n438053 , n382854 );
buf ( n438054 , n40971 );
and ( n438055 , n438053 , n438054 );
nor ( n438056 , n438052 , n438055 );
buf ( n438057 , n438056 );
not ( n438058 , n438057 );
and ( n438059 , n438047 , n438058 );
nor ( n438060 , n438059 , C0 );
buf ( n438061 , n384627 );
not ( n438062 , n438061 );
buf ( n438063 , n437352 );
not ( n438064 , n438063 );
or ( n438065 , n438062 , n438064 );
buf ( n438066 , n384568 );
not ( n438067 , n438066 );
buf ( n438068 , n386012 );
not ( n438069 , n438068 );
or ( n438070 , n438067 , n438069 );
buf ( n438071 , n41595 );
buf ( n438072 , n42390 );
nand ( n438073 , n438071 , n438072 );
buf ( n438074 , n438073 );
buf ( n438075 , n438074 );
nand ( n438076 , n438070 , n438075 );
buf ( n438077 , n438076 );
buf ( n438078 , n438077 );
buf ( n438079 , n384557 );
nand ( n438080 , n438078 , n438079 );
buf ( n438081 , n438080 );
buf ( n438082 , n438081 );
nand ( n438083 , n438065 , n438082 );
buf ( n438084 , n438083 );
xor ( n438085 , n438060 , n438084 );
buf ( n438086 , n384416 );
not ( n438087 , n438086 );
buf ( n438088 , n36821 );
not ( n438089 , n438088 );
buf ( n438090 , n48233 );
not ( n438091 , n438090 );
or ( n438092 , n438089 , n438091 );
buf ( n438093 , n48234 );
buf ( n438094 , n40886 );
nand ( n438095 , n438093 , n438094 );
buf ( n438096 , n438095 );
buf ( n438097 , n438096 );
nand ( n438098 , n438092 , n438097 );
buf ( n438099 , n438098 );
buf ( n438100 , n438099 );
not ( n438101 , n438100 );
or ( n438102 , n438087 , n438101 );
buf ( n438103 , n437590 );
not ( n438104 , n438103 );
buf ( n438105 , n384369 );
nand ( n438106 , n438104 , n438105 );
buf ( n438107 , n438106 );
buf ( n438108 , n438107 );
nand ( n438109 , n438102 , n438108 );
buf ( n438110 , n438109 );
xor ( n438111 , n438085 , n438110 );
not ( n438112 , n438111 );
and ( n438113 , n438046 , n438112 );
not ( n438114 , n438046 );
and ( n438115 , n438114 , n438111 );
nor ( n438116 , n438113 , n438115 );
not ( n438117 , n437718 );
not ( n438118 , n437665 );
or ( n438119 , n438117 , n438118 );
buf ( n438120 , n437665 );
not ( n438121 , n438120 );
buf ( n438122 , n438121 );
not ( n438123 , n438122 );
not ( n438124 , n437715 );
or ( n438125 , n438123 , n438124 );
nand ( n438126 , n438125 , n437690 );
nand ( n438127 , n438119 , n438126 );
and ( n438128 , n438116 , n438127 );
not ( n438129 , n438116 );
buf ( n438130 , n438127 );
not ( n438131 , n438130 );
buf ( n438132 , n438131 );
and ( n438133 , n438129 , n438132 );
nor ( n438134 , n438128 , n438133 );
buf ( n438135 , n437337 );
not ( n438136 , n438135 );
buf ( n438137 , n437403 );
not ( n438138 , n438137 );
or ( n438139 , n438136 , n438138 );
not ( n438140 , n437340 );
not ( n438141 , n437400 );
or ( n438142 , n438140 , n438141 );
nand ( n438143 , n438142 , n437417 );
buf ( n438144 , n438143 );
nand ( n438145 , n438139 , n438144 );
buf ( n438146 , n438145 );
xor ( n438147 , n438134 , n438146 );
xor ( n438148 , n438011 , n438147 );
not ( n438149 , n437612 );
not ( n438150 , n437621 );
and ( n438151 , n438149 , n438150 );
nand ( n438152 , n437612 , n437621 );
buf ( n438153 , n437413 );
and ( n438154 , n438153 , n437417 );
not ( n438155 , n438153 );
and ( n438156 , n438155 , n437420 );
nor ( n438157 , n438154 , n438156 );
and ( n438158 , n438152 , n438157 );
nor ( n438159 , n438151 , n438158 );
xnor ( n438160 , n438148 , n438159 );
buf ( n438161 , n438160 );
xor ( n438162 , n438003 , n438161 );
buf ( n438163 , n437768 );
buf ( n438164 , n437757 );
not ( n438165 , n438164 );
buf ( n438166 , n437762 );
nand ( n438167 , n438165 , n438166 );
buf ( n438168 , n438167 );
buf ( n438169 , n438168 );
nand ( n438170 , n438163 , n438169 );
buf ( n438171 , n438170 );
buf ( n438172 , n438171 );
buf ( n438173 , n437762 );
not ( n438174 , n438173 );
buf ( n438175 , n437757 );
nand ( n438176 , n438174 , n438175 );
buf ( n438177 , n438176 );
buf ( n438178 , n438177 );
and ( n438179 , n438172 , n438178 );
buf ( n438180 , n438179 );
buf ( n438181 , n438180 );
xor ( n438182 , n438162 , n438181 );
buf ( n438183 , n438182 );
xor ( n438184 , n437625 , n437643 );
and ( n438185 , n438184 , n437770 );
and ( n438186 , n437625 , n437643 );
or ( n438187 , n438185 , n438186 );
buf ( n438188 , n438187 );
nand ( n438189 , n438183 , n438188 );
nand ( n438190 , n437773 , n438189 );
not ( n438191 , n438190 );
xor ( n438192 , n437882 , n437993 );
and ( n438193 , n438192 , n437999 );
and ( n438194 , n437882 , n437993 );
or ( n438195 , n438193 , n438194 );
buf ( n438196 , n438195 );
buf ( n438197 , n438196 );
buf ( n438198 , n385491 );
buf ( n438199 , n388774 );
and ( n438200 , n438198 , n438199 );
not ( n438201 , n438198 );
buf ( n438202 , n388771 );
and ( n438203 , n438201 , n438202 );
nor ( n438204 , n438200 , n438203 );
buf ( n438205 , n438204 );
not ( n438206 , n438205 );
not ( n438207 , n37924 );
and ( n438208 , n438206 , n438207 );
buf ( n438209 , n437781 );
not ( n438210 , n438209 );
buf ( n438211 , n438210 );
and ( n438212 , n438211 , n385889 );
nor ( n438213 , n438208 , n438212 );
buf ( n438214 , n438213 );
buf ( n438215 , n37354 );
not ( n438216 , n438215 );
buf ( n438217 , n382893 );
not ( n438218 , n438217 );
or ( n438219 , n438216 , n438218 );
buf ( n438220 , n402307 );
not ( n438221 , n438220 );
buf ( n438222 , n37347 );
nand ( n438223 , n438221 , n438222 );
buf ( n438224 , n438223 );
buf ( n438225 , n438224 );
nand ( n438226 , n438219 , n438225 );
buf ( n438227 , n438226 );
buf ( n438228 , n438227 );
buf ( n438229 , n37695 );
and ( n438230 , n438228 , n438229 );
buf ( n438231 , n438034 );
not ( n438232 , n438231 );
buf ( n438233 , n384901 );
nor ( n438234 , n438232 , n438233 );
buf ( n438235 , n438234 );
buf ( n438236 , n438235 );
nor ( n438237 , n438230 , n438236 );
buf ( n438238 , n438237 );
buf ( n438239 , n438238 );
xor ( n438240 , n438214 , n438239 );
buf ( n438241 , n438240 );
buf ( n438242 , n438241 );
xor ( n438243 , n437827 , n437853 );
and ( n438244 , n438243 , n437879 );
and ( n438245 , n437827 , n437853 );
or ( n438246 , n438244 , n438245 );
buf ( n438247 , n438246 );
buf ( n438248 , n438247 );
xnor ( n438249 , n438242 , n438248 );
buf ( n438250 , n438249 );
buf ( n438251 , n438250 );
not ( n438252 , n438251 );
buf ( n438253 , n438252 );
buf ( n438254 , n438253 );
and ( n438255 , n438197 , n438254 );
not ( n438256 , n438197 );
buf ( n438257 , n438250 );
and ( n438258 , n438256 , n438257 );
nor ( n438259 , n438255 , n438258 );
buf ( n438260 , n438259 );
buf ( n438261 , n438260 );
xor ( n438262 , n437907 , n437932 );
and ( n438263 , n438262 , n437990 );
and ( n438264 , n437907 , n437932 );
or ( n438265 , n438263 , n438264 );
buf ( n438266 , n438265 );
buf ( n438267 , n384416 );
not ( n438268 , n438267 );
not ( n438269 , n36821 );
not ( n438270 , n46361 );
or ( n438271 , n438269 , n438270 );
nand ( n438272 , n383765 , n37597 );
nand ( n438273 , n438271 , n438272 );
buf ( n438274 , n438273 );
not ( n438275 , n438274 );
or ( n438276 , n438268 , n438275 );
buf ( n438277 , n438099 );
buf ( n438278 , n384369 );
nand ( n438279 , n438277 , n438278 );
buf ( n438280 , n438279 );
buf ( n438281 , n438280 );
nand ( n438282 , n438276 , n438281 );
buf ( n438283 , n438282 );
buf ( n438284 , n438283 );
buf ( n438285 , n41564 );
not ( n438286 , n438285 );
buf ( n438287 , n389125 );
not ( n438288 , n438287 );
buf ( n438289 , n438288 );
buf ( n438290 , n438289 );
not ( n438291 , n438290 );
or ( n438292 , n438286 , n438291 );
buf ( n438293 , n437845 );
nand ( n438294 , n438292 , n438293 );
buf ( n438295 , n438294 );
buf ( n438296 , n438295 );
not ( n438297 , n438296 );
buf ( n438298 , n438297 );
buf ( n438299 , n438298 );
and ( n438300 , n438284 , n438299 );
not ( n438301 , n438284 );
buf ( n438302 , n438295 );
and ( n438303 , n438301 , n438302 );
nor ( n438304 , n438300 , n438303 );
buf ( n438305 , n438304 );
xor ( n438306 , n437955 , n437969 );
and ( n438307 , n438306 , n437987 );
and ( n438308 , n437955 , n437969 );
or ( n438309 , n438307 , n438308 );
buf ( n438310 , n438309 );
xor ( n438311 , n438305 , n438310 );
and ( n438312 , n438266 , n438311 );
not ( n438313 , n438266 );
buf ( n438314 , n438311 );
not ( n438315 , n438314 );
buf ( n438316 , n438315 );
and ( n438317 , n438313 , n438316 );
or ( n438318 , n438312 , n438317 );
buf ( n438319 , n438318 );
buf ( n438320 , n383946 );
not ( n438321 , n438320 );
buf ( n438322 , n36399 );
not ( n438323 , n438322 );
buf ( n438324 , n38357 );
not ( n438325 , n438324 );
or ( n438326 , n438323 , n438325 );
buf ( n438327 , n389435 );
buf ( n438328 , n36398 );
nand ( n438329 , n438327 , n438328 );
buf ( n438330 , n438329 );
buf ( n438331 , n438330 );
nand ( n438332 , n438326 , n438331 );
buf ( n438333 , n438332 );
buf ( n438334 , n438333 );
not ( n438335 , n438334 );
or ( n438336 , n438321 , n438335 );
buf ( n438337 , n437899 );
buf ( n438338 , n384011 );
nand ( n438339 , n438337 , n438338 );
buf ( n438340 , n438339 );
buf ( n438341 , n438340 );
nand ( n438342 , n438336 , n438341 );
buf ( n438343 , n438342 );
buf ( n438344 , n438343 );
buf ( n438345 , n386480 );
not ( n438346 , n438345 );
buf ( n438347 , n38972 );
not ( n438348 , n438347 );
buf ( n438349 , n382535 );
not ( n438350 , n438349 );
or ( n438351 , n438348 , n438350 );
buf ( n438352 , n382532 );
buf ( n438353 , n38971 );
nand ( n438354 , n438352 , n438353 );
buf ( n438355 , n438354 );
buf ( n438356 , n438355 );
nand ( n438357 , n438351 , n438356 );
buf ( n438358 , n438357 );
buf ( n438359 , n438358 );
not ( n438360 , n438359 );
or ( n438361 , n438346 , n438360 );
buf ( n438362 , n437924 );
buf ( n438363 , n386496 );
nand ( n438364 , n438362 , n438363 );
buf ( n438365 , n438364 );
buf ( n438366 , n438365 );
nand ( n438367 , n438361 , n438366 );
buf ( n438368 , n438367 );
buf ( n438369 , n438368 );
xor ( n438370 , n438344 , n438369 );
buf ( n438371 , n434175 );
not ( n438372 , n438371 );
buf ( n438373 , n437946 );
not ( n438374 , n438373 );
and ( n438375 , n438372 , n438374 );
buf ( n438376 , n38667 );
buf ( n438377 , n389024 );
and ( n438378 , n438376 , n438377 );
nor ( n438379 , n438375 , n438378 );
buf ( n438380 , n438379 );
not ( n438381 , n438380 );
not ( n438382 , n438381 );
buf ( n438383 , n389777 );
buf ( n438384 , n386158 );
nor ( n438385 , n438383 , n438384 );
buf ( n438386 , n438385 );
buf ( n438387 , n438386 );
nor ( n438388 , C0 , n438387 );
buf ( n438389 , n438388 );
not ( n438390 , n438389 );
or ( n438391 , n438382 , n438390 );
buf ( n438392 , n438389 );
not ( n438393 , n438392 );
buf ( n438394 , n438393 );
nand ( n438395 , n438394 , n438380 );
nand ( n438396 , n438391 , n438395 );
buf ( n438397 , n438060 );
not ( n438398 , n438397 );
buf ( n438399 , n438398 );
buf ( n438400 , n438399 );
not ( n438401 , n438400 );
buf ( n438402 , n438401 );
xnor ( n438403 , n438396 , n438402 );
buf ( n438404 , n438403 );
xor ( n438405 , n438370 , n438404 );
buf ( n438406 , n438405 );
buf ( n438407 , n438406 );
not ( n438408 , n438407 );
buf ( n438409 , n438408 );
buf ( n438410 , n438409 );
and ( n438411 , n438319 , n438410 );
not ( n438412 , n438319 );
buf ( n438413 , n438406 );
and ( n438414 , n438412 , n438413 );
nor ( n438415 , n438411 , n438414 );
buf ( n438416 , n438415 );
buf ( n438417 , n438416 );
buf ( n438418 , n438417 );
buf ( n438419 , n438418 );
buf ( n438420 , n438419 );
xor ( n438421 , n438261 , n438420 );
buf ( n438422 , n438421 );
buf ( n438423 , n438422 );
not ( n438424 , n438423 );
buf ( n438425 , n438424 );
buf ( n438426 , n438425 );
not ( n438427 , n438426 );
not ( n438428 , n438017 );
not ( n438429 , n438041 );
or ( n438430 , n438428 , n438429 );
and ( n438431 , n437600 , n438013 );
nor ( n438432 , n438431 , n438015 );
not ( n438433 , n438432 );
not ( n438434 , n438044 );
or ( n438435 , n438433 , n438434 );
nand ( n438436 , n438435 , n438111 );
nand ( n438437 , n438430 , n438436 );
buf ( n438438 , n438437 );
buf ( n438439 , n384644 );
not ( n438440 , n438439 );
buf ( n438441 , n36253 );
not ( n438442 , n438441 );
buf ( n438443 , n38823 );
not ( n438444 , n438443 );
or ( n438445 , n438442 , n438444 );
buf ( n438446 , n36068 );
buf ( n438447 , n36252 );
nand ( n438448 , n438446 , n438447 );
buf ( n438449 , n438448 );
buf ( n438450 , n438449 );
nand ( n438451 , n438445 , n438450 );
buf ( n438452 , n438451 );
buf ( n438453 , n438452 );
not ( n438454 , n438453 );
or ( n438455 , n438440 , n438454 );
buf ( n438456 , n437871 );
buf ( n438457 , n383897 );
nand ( n438458 , n438456 , n438457 );
buf ( n438459 , n438458 );
buf ( n438460 , n438459 );
nand ( n438461 , n438455 , n438460 );
buf ( n438462 , n438461 );
buf ( n438463 , n438462 );
buf ( n438464 , n438402 );
not ( n438465 , n438464 );
buf ( n438466 , n438110 );
not ( n438467 , n438466 );
or ( n438468 , n438465 , n438467 );
buf ( n438469 , n438110 );
buf ( n438470 , n438402 );
or ( n438471 , n438469 , n438470 );
buf ( n438472 , n438084 );
nand ( n438473 , n438471 , n438472 );
buf ( n438474 , n438473 );
buf ( n438475 , n438474 );
nand ( n438476 , n438468 , n438475 );
buf ( n438477 , n438476 );
buf ( n438478 , n438477 );
xor ( n438479 , n438463 , n438478 );
buf ( n438480 , n437963 );
not ( n438481 , n438480 );
buf ( n438482 , n386300 );
not ( n438483 , n438482 );
or ( n438484 , n438481 , n438483 );
buf ( n438485 , n386231 );
not ( n438486 , n438485 );
buf ( n438487 , n386310 );
nand ( n438488 , n438486 , n438487 );
buf ( n438489 , n438488 );
buf ( n438490 , n438489 );
nand ( n438491 , n438484 , n438490 );
buf ( n438492 , n438491 );
buf ( n438493 , n438492 );
buf ( n438494 , n383409 );
not ( n438495 , n438494 );
buf ( n438496 , n385729 );
not ( n438497 , n438496 );
buf ( n438498 , n384280 );
not ( n438499 , n438498 );
or ( n438500 , n438497 , n438499 );
buf ( n438501 , n384974 );
buf ( n438502 , n385633 );
nand ( n438503 , n438501 , n438502 );
buf ( n438504 , n438503 );
buf ( n438505 , n438504 );
nand ( n438506 , n438500 , n438505 );
buf ( n438507 , n438506 );
buf ( n438508 , n438507 );
not ( n438509 , n438508 );
or ( n438510 , n438495 , n438509 );
buf ( n438511 , n437981 );
not ( n438512 , n438511 );
buf ( n438513 , n385751 );
nand ( n438514 , n438512 , n438513 );
buf ( n438515 , n438514 );
buf ( n438516 , n438515 );
nand ( n438517 , n438510 , n438516 );
buf ( n438518 , n438517 );
buf ( n438519 , n438518 );
xor ( n438520 , n438493 , n438519 );
buf ( n438521 , n384557 );
not ( n438522 , n438521 );
buf ( n438523 , n384568 );
not ( n438524 , n438523 );
buf ( n438525 , n384211 );
not ( n438526 , n438525 );
or ( n438527 , n438524 , n438526 );
buf ( n438528 , n384189 );
buf ( n438529 , n384565 );
nand ( n438530 , n438528 , n438529 );
buf ( n438531 , n438530 );
buf ( n438532 , n438531 );
nand ( n438533 , n438527 , n438532 );
buf ( n438534 , n438533 );
buf ( n438535 , n438534 );
not ( n438536 , n438535 );
or ( n438537 , n438522 , n438536 );
buf ( n438538 , n384627 );
buf ( n438539 , n438077 );
nand ( n438540 , n438538 , n438539 );
buf ( n438541 , n438540 );
buf ( n438542 , n438541 );
nand ( n438543 , n438537 , n438542 );
buf ( n438544 , n438543 );
buf ( n438545 , n438544 );
xor ( n438546 , n438520 , n438545 );
buf ( n438547 , n438546 );
buf ( n438548 , n438547 );
xor ( n438549 , n438479 , n438548 );
buf ( n438550 , n438549 );
buf ( n438551 , n438550 );
xor ( n438552 , n438438 , n438551 );
buf ( n438553 , n438552 );
buf ( n438554 , n438553 );
not ( n438555 , n437799 );
buf ( n438556 , n437791 );
not ( n438557 , n438556 );
buf ( n438558 , n438557 );
not ( n438559 , n438558 );
or ( n438560 , n438555 , n438559 );
not ( n438561 , n437799 );
buf ( n438562 , n438561 );
not ( n438563 , n438562 );
buf ( n438564 , n437791 );
not ( n438565 , n438564 );
or ( n438566 , n438563 , n438565 );
buf ( n438567 , n437805 );
nand ( n438568 , n438566 , n438567 );
buf ( n438569 , n438568 );
nand ( n438570 , n438560 , n438569 );
buf ( n438571 , n438570 );
and ( n438572 , n438554 , n438571 );
not ( n438573 , n438554 );
buf ( n438574 , n438570 );
not ( n438575 , n438574 );
buf ( n438576 , n438575 );
buf ( n438577 , n438576 );
and ( n438578 , n438573 , n438577 );
nor ( n438579 , n438572 , n438578 );
buf ( n438580 , n438579 );
buf ( n438581 , n438580 );
buf ( n438582 , n438116 );
not ( n438583 , n438582 );
buf ( n438584 , n438132 );
not ( n438585 , n438584 );
or ( n438586 , n438583 , n438585 );
buf ( n438587 , n438146 );
nand ( n438588 , n438586 , n438587 );
buf ( n438589 , n438588 );
buf ( n438590 , n438589 );
not ( n438591 , n438116 );
nand ( n438592 , n438591 , n438127 );
buf ( n438593 , n438592 );
nand ( n438594 , n438590 , n438593 );
buf ( n438595 , n438594 );
buf ( n438596 , n438595 );
xor ( n438597 , n438581 , n438596 );
buf ( n438598 , n438597 );
buf ( n438599 , n437806 );
not ( n438600 , n438599 );
buf ( n438601 , n438001 );
not ( n438602 , n438601 );
or ( n438603 , n438600 , n438602 );
buf ( n438604 , n438001 );
buf ( n438605 , n437806 );
or ( n438606 , n438604 , n438605 );
buf ( n438607 , n437820 );
nand ( n438608 , n438606 , n438607 );
buf ( n438609 , n438608 );
buf ( n438610 , n438609 );
nand ( n438611 , n438603 , n438610 );
buf ( n438612 , n438611 );
and ( n438613 , n438598 , n438612 );
not ( n438614 , n438598 );
buf ( n438615 , n438612 );
not ( n438616 , n438615 );
buf ( n438617 , n438616 );
and ( n438618 , n438614 , n438617 );
nor ( n438619 , n438613 , n438618 );
not ( n438620 , n438619 );
buf ( n438621 , n438620 );
not ( n438622 , n438621 );
or ( n438623 , n438427 , n438622 );
nand ( n438624 , n438422 , n438619 );
buf ( n438625 , n438624 );
nand ( n438626 , n438623 , n438625 );
buf ( n438627 , n438626 );
buf ( n438628 , n438627 );
buf ( n438629 , n438011 );
not ( n438630 , n438629 );
buf ( n438631 , n438147 );
nand ( n438632 , n438630 , n438631 );
buf ( n438633 , n438632 );
buf ( n438634 , n438633 );
not ( n438635 , n438634 );
buf ( n438636 , n438159 );
not ( n438637 , n438636 );
buf ( n438638 , n438637 );
buf ( n438639 , n438638 );
not ( n438640 , n438639 );
or ( n438641 , n438635 , n438640 );
buf ( n438642 , n438147 );
not ( n438643 , n438642 );
buf ( n438644 , n438011 );
nand ( n438645 , n438643 , n438644 );
buf ( n438646 , n438645 );
buf ( n438647 , n438646 );
nand ( n438648 , n438641 , n438647 );
buf ( n438649 , n438648 );
buf ( n438650 , n438649 );
xnor ( n438651 , n438628 , n438650 );
buf ( n438652 , n438651 );
xor ( n438653 , n438003 , n438161 );
and ( n438654 , n438653 , n438181 );
and ( n438655 , n438003 , n438161 );
or ( n438656 , n438654 , n438655 );
buf ( n438657 , n438656 );
nand ( n438658 , n438652 , n438657 );
not ( n438659 , n438425 );
not ( n438660 , n438619 );
or ( n438661 , n438659 , n438660 );
buf ( n438662 , n438422 );
not ( n438663 , n438662 );
buf ( n438664 , n438620 );
not ( n438665 , n438664 );
or ( n438666 , n438663 , n438665 );
buf ( n438667 , n438649 );
nand ( n438668 , n438666 , n438667 );
buf ( n438669 , n438668 );
nand ( n438670 , n438661 , n438669 );
not ( n438671 , n438670 );
xor ( n438672 , n438344 , n438369 );
and ( n438673 , n438672 , n438404 );
and ( n438674 , n438344 , n438369 );
or ( n438675 , n438673 , n438674 );
buf ( n438676 , n438675 );
buf ( n438677 , n438676 );
buf ( n438678 , n438298 );
not ( n438679 , n438678 );
buf ( n438680 , n438283 );
not ( n438681 , n438680 );
buf ( n438682 , n438681 );
buf ( n438683 , n438682 );
not ( n438684 , n438683 );
or ( n438685 , n438679 , n438684 );
buf ( n438686 , n438310 );
nand ( n438687 , n438685 , n438686 );
buf ( n438688 , n438687 );
buf ( n438689 , n438688 );
buf ( n438690 , n438298 );
not ( n438691 , n438690 );
buf ( n438692 , n438283 );
nand ( n438693 , n438691 , n438692 );
buf ( n438694 , n438693 );
buf ( n438695 , n438694 );
nand ( n438696 , n438689 , n438695 );
buf ( n438697 , n438696 );
buf ( n438698 , n438697 );
xor ( n438699 , n438677 , n438698 );
buf ( n438700 , n438394 );
not ( n438701 , n438700 );
buf ( n438702 , n438381 );
not ( n438703 , n438702 );
or ( n438704 , n438701 , n438703 );
buf ( n438705 , n438389 );
not ( n438706 , n438705 );
buf ( n438707 , n438380 );
not ( n438708 , n438707 );
or ( n438709 , n438706 , n438708 );
buf ( n438710 , n438399 );
nand ( n438711 , n438709 , n438710 );
buf ( n438712 , n438711 );
buf ( n438713 , n438712 );
nand ( n438714 , n438704 , n438713 );
buf ( n438715 , n438714 );
buf ( n438716 , n438715 );
buf ( n438717 , n384369 );
not ( n438718 , n438717 );
buf ( n438719 , n438273 );
not ( n438720 , n438719 );
or ( n438721 , n438718 , n438720 );
buf ( n438722 , n386045 );
buf ( n438723 , n384416 );
nand ( n438724 , n438722 , n438723 );
buf ( n438725 , n438724 );
buf ( n438726 , n438725 );
nand ( n438727 , n438721 , n438726 );
buf ( n438728 , n438727 );
buf ( n438729 , n438728 );
xor ( n438730 , n438716 , n438729 );
buf ( n438731 , n386480 );
not ( n438732 , n438731 );
buf ( n438733 , n386516 );
not ( n438734 , n438733 );
or ( n438735 , n438732 , n438734 );
buf ( n438736 , n438358 );
buf ( n438737 , n386496 );
nand ( n438738 , n438736 , n438737 );
buf ( n438739 , n438738 );
buf ( n438740 , n438739 );
nand ( n438741 , n438735 , n438740 );
buf ( n438742 , n438741 );
buf ( n438743 , n438742 );
xor ( n438744 , n438730 , n438743 );
buf ( n438745 , n438744 );
buf ( n438746 , n438745 );
xor ( n438747 , n438699 , n438746 );
buf ( n438748 , n438747 );
buf ( n438749 , n438748 );
buf ( n438750 , n438316 );
not ( n438751 , n438750 );
buf ( n438752 , n438266 );
not ( n438753 , n438752 );
or ( n438754 , n438751 , n438753 );
buf ( n438755 , n438316 );
buf ( n438756 , n438266 );
or ( n438757 , n438755 , n438756 );
buf ( n438758 , n438406 );
nand ( n438759 , n438757 , n438758 );
buf ( n438760 , n438759 );
buf ( n438761 , n438760 );
nand ( n438762 , n438754 , n438761 );
buf ( n438763 , n438762 );
buf ( n438764 , n438763 );
xor ( n438765 , n438493 , n438519 );
and ( n438766 , n438765 , n438545 );
and ( n438767 , n438493 , n438519 );
or ( n438768 , n438766 , n438767 );
buf ( n438769 , n438768 );
buf ( n438770 , n438769 );
buf ( n438771 , n385269 );
not ( n438772 , n438771 );
buf ( n438773 , n438227 );
not ( n438774 , n438773 );
or ( n438775 , n438772 , n438774 );
buf ( n438776 , n39033 );
buf ( n438777 , n37695 );
nand ( n438778 , n438776 , n438777 );
buf ( n438779 , n438778 );
buf ( n438780 , n438779 );
nand ( n438781 , n438775 , n438780 );
buf ( n438782 , n438781 );
buf ( n438783 , n438782 );
xor ( n438784 , n438770 , n438783 );
buf ( n438785 , n384627 );
not ( n438786 , n438785 );
buf ( n438787 , n438534 );
not ( n438788 , n438787 );
or ( n438789 , n438786 , n438788 );
buf ( n438790 , n386122 );
buf ( n438791 , n384557 );
nand ( n438792 , n438790 , n438791 );
buf ( n438793 , n438792 );
buf ( n438794 , n438793 );
nand ( n438795 , n438789 , n438794 );
buf ( n438796 , n438795 );
buf ( n438797 , n438796 );
buf ( n438798 , n383482 );
not ( n438799 , n438798 );
buf ( n438800 , n438507 );
not ( n438801 , n438800 );
or ( n438802 , n438799 , n438801 );
buf ( n438803 , n386023 );
buf ( n438804 , n383409 );
nand ( n438805 , n438803 , n438804 );
buf ( n438806 , n438805 );
buf ( n438807 , n438806 );
nand ( n438808 , n438802 , n438807 );
buf ( n438809 , n438808 );
buf ( n438810 , n438809 );
xor ( n438811 , n438797 , n438810 );
buf ( n438812 , n384011 );
not ( n438813 , n438812 );
buf ( n438814 , n438333 );
not ( n438815 , n438814 );
or ( n438816 , n438813 , n438815 );
buf ( n438817 , n383943 );
not ( n438818 , n438817 );
buf ( n438819 , n386538 );
nand ( n438820 , n438818 , n438819 );
buf ( n438821 , n438820 );
buf ( n438822 , n438821 );
nand ( n438823 , n438816 , n438822 );
buf ( n438824 , n438823 );
buf ( n438825 , n438824 );
xor ( n438826 , n438811 , n438825 );
buf ( n438827 , n438826 );
buf ( n438828 , n438827 );
xor ( n438829 , n438784 , n438828 );
buf ( n438830 , n438829 );
buf ( n438831 , n438830 );
xor ( n438832 , n438764 , n438831 );
buf ( n438833 , n438832 );
buf ( n438834 , n438833 );
not ( n438835 , n438834 );
xor ( n438836 , n438749 , n438835 );
buf ( n438837 , n438836 );
buf ( n438838 , n438837 );
buf ( n438839 , n438580 );
buf ( n438840 , n438595 );
or ( n438841 , n438839 , n438840 );
buf ( n438842 , n438841 );
buf ( n438843 , n438842 );
buf ( n438844 , n438612 );
and ( n438845 , n438843 , n438844 );
and ( n438846 , n438581 , n438596 );
buf ( n438847 , n438846 );
buf ( n438848 , n438847 );
nor ( n438849 , n438845 , n438848 );
buf ( n438850 , n438849 );
buf ( n438851 , n438850 );
xor ( n438852 , n438838 , n438851 );
or ( n438853 , n438437 , n438550 );
buf ( n438854 , n438853 );
buf ( n438855 , n438570 );
and ( n438856 , n438854 , n438855 );
and ( n438857 , n438438 , n438551 );
buf ( n438858 , n438857 );
buf ( n438859 , n438858 );
nor ( n438860 , n438856 , n438859 );
buf ( n438861 , n438860 );
buf ( n438862 , n438861 );
xor ( n438863 , n438463 , n438478 );
and ( n438864 , n438863 , n438548 );
and ( n438865 , n438463 , n438478 );
or ( n438866 , n438864 , n438865 );
buf ( n438867 , n438866 );
xor ( n438868 , n386193 , n386217 );
xor ( n438869 , n438868 , n386250 );
buf ( n438870 , n438869 );
buf ( n438871 , n438870 );
buf ( n438872 , n383897 );
not ( n438873 , n438872 );
buf ( n438874 , n438452 );
not ( n438875 , n438874 );
or ( n438876 , n438873 , n438875 );
nand ( n438877 , n39055 , n384644 );
buf ( n438878 , n438877 );
nand ( n438879 , n438876 , n438878 );
buf ( n438880 , n438879 );
buf ( n438881 , n438880 );
xor ( n438882 , n438871 , n438881 );
buf ( n438883 , n385889 );
not ( n438884 , n438883 );
buf ( n438885 , n438205 );
not ( n438886 , n438885 );
buf ( n438887 , n438886 );
buf ( n438888 , n438887 );
not ( n438889 , n438888 );
or ( n438890 , n438884 , n438889 );
buf ( n438891 , n386086 );
buf ( n438892 , n38324 );
nand ( n438893 , n438891 , n438892 );
buf ( n438894 , n438893 );
buf ( n438895 , n438894 );
nand ( n438896 , n438890 , n438895 );
buf ( n438897 , n438896 );
buf ( n438898 , n438897 );
xor ( n438899 , n438882 , n438898 );
buf ( n438900 , n438899 );
buf ( n438901 , n438900 );
not ( n438902 , n438901 );
buf ( n438903 , n438902 );
and ( n438904 , n438867 , n438903 );
not ( n438905 , n438867 );
and ( n438906 , n438905 , n438900 );
nor ( n438907 , n438904 , n438906 );
buf ( n438908 , n438247 );
buf ( n438909 , n438213 );
buf ( n438910 , n438238 );
nand ( n438911 , n438909 , n438910 );
buf ( n438912 , n438911 );
buf ( n438913 , n438912 );
and ( n438914 , n438908 , n438913 );
buf ( n438915 , n438238 );
buf ( n438916 , n438213 );
nor ( n438917 , n438915 , n438916 );
buf ( n438918 , n438917 );
buf ( n438919 , n438918 );
nor ( n438920 , n438914 , n438919 );
buf ( n438921 , n438920 );
buf ( n438922 , n438921 );
not ( n438923 , n438922 );
buf ( n438924 , n438923 );
and ( n438925 , n438907 , n438924 );
not ( n438926 , n438907 );
and ( n438927 , n438926 , n438921 );
nor ( n438928 , n438925 , n438927 );
buf ( n438929 , n438928 );
xor ( n438930 , n438862 , n438929 );
buf ( n438931 , n438416 );
buf ( n438932 , n438250 );
nand ( n438933 , n438931 , n438932 );
buf ( n438934 , n438933 );
buf ( n438935 , n438934 );
buf ( n438936 , n438196 );
and ( n438937 , n438935 , n438936 );
buf ( n438938 , n438416 );
buf ( n438939 , n438250 );
nor ( n438940 , n438938 , n438939 );
buf ( n438941 , n438940 );
buf ( n438942 , n438941 );
nor ( n438943 , n438937 , n438942 );
buf ( n438944 , n438943 );
buf ( n438945 , n438944 );
xor ( n438946 , n438930 , n438945 );
buf ( n438947 , n438946 );
buf ( n438948 , n438947 );
xor ( n438949 , n438852 , n438948 );
buf ( n438950 , n438949 );
nand ( n438951 , n438671 , n438950 );
nand ( n438952 , n438191 , n438658 , n438951 );
buf ( n438953 , n438952 );
not ( n438954 , n438953 );
buf ( n438955 , n438954 );
buf ( n438956 , n386443 );
not ( n438957 , n438956 );
buf ( n438958 , n386372 );
not ( n438959 , n438958 );
or ( n438960 , n438957 , n438959 );
buf ( n438961 , n386372 );
buf ( n438962 , n386443 );
or ( n438963 , n438961 , n438962 );
nand ( n438964 , n438960 , n438963 );
buf ( n438965 , n438964 );
buf ( n438966 , n438965 );
buf ( n438967 , n386407 );
and ( n438968 , n438966 , n438967 );
not ( n438969 , n438966 );
buf ( n438970 , n386453 );
and ( n438971 , n438969 , n438970 );
nor ( n438972 , n438968 , n438971 );
buf ( n438973 , n438972 );
buf ( n438974 , n438973 );
buf ( n438975 , n386057 );
buf ( n438976 , n386062 );
xor ( n438977 , n438975 , n438976 );
buf ( n438978 , n386260 );
xnor ( n438979 , n438977 , n438978 );
buf ( n438980 , n438979 );
buf ( n438981 , n438980 );
xor ( n438982 , n438974 , n438981 );
xor ( n438983 , n438797 , n438810 );
and ( n438984 , n438983 , n438825 );
and ( n438985 , n438797 , n438810 );
or ( n438986 , n438984 , n438985 );
buf ( n438987 , n438986 );
buf ( n438988 , n438987 );
not ( n438989 , n438988 );
xor ( n438990 , n386093 , n386133 );
xor ( n438991 , n438990 , n386254 );
buf ( n438992 , n438991 );
nand ( n438993 , n438989 , n438992 );
buf ( n438994 , n438993 );
buf ( n438995 , n438994 );
xor ( n438996 , n438716 , n438729 );
and ( n438997 , n438996 , n438743 );
and ( n438998 , n438716 , n438729 );
or ( n438999 , n438997 , n438998 );
buf ( n439000 , n438999 );
buf ( n439001 , n439000 );
and ( n439002 , n438995 , n439001 );
buf ( n439003 , n438987 );
not ( n439004 , n439003 );
buf ( n439005 , n438991 );
nor ( n439006 , n439004 , n439005 );
buf ( n439007 , n439006 );
buf ( n439008 , n439007 );
nor ( n439009 , n439002 , n439008 );
buf ( n439010 , n439009 );
buf ( n439011 , n439010 );
and ( n439012 , n438982 , n439011 );
and ( n439013 , n438974 , n438981 );
or ( n439014 , n439012 , n439013 );
buf ( n439015 , n439014 );
not ( n439016 , n439015 );
buf ( n439017 , n386463 );
buf ( n439018 , n386615 );
and ( n439019 , n439017 , n439018 );
not ( n439020 , n439017 );
buf ( n439021 , n386618 );
and ( n439022 , n439020 , n439021 );
nor ( n439023 , n439019 , n439022 );
buf ( n439024 , n439023 );
buf ( n439025 , n439024 );
buf ( n439026 , n386274 );
and ( n439027 , n439025 , n439026 );
not ( n439028 , n439025 );
buf ( n439029 , n386274 );
not ( n439030 , n439029 );
buf ( n439031 , n439030 );
buf ( n439032 , n439031 );
and ( n439033 , n439028 , n439032 );
or ( n439034 , n439027 , n439033 );
buf ( n439035 , n439034 );
xor ( n439036 , n439016 , n439035 );
xor ( n439037 , n386551 , n386555 );
xor ( n439038 , n439037 , n386611 );
buf ( n439039 , n439038 );
buf ( n439040 , n439039 );
not ( n439041 , n439040 );
buf ( n439042 , n439041 );
buf ( n439043 , n439042 );
not ( n439044 , n439043 );
xor ( n439045 , n438987 , n439000 );
buf ( n439046 , n439045 );
buf ( n439047 , n438991 );
not ( n439048 , n439047 );
buf ( n439049 , n439048 );
buf ( n439050 , n439049 );
and ( n439051 , n439046 , n439050 );
not ( n439052 , n439046 );
buf ( n439053 , n438991 );
and ( n439054 , n439052 , n439053 );
nor ( n439055 , n439051 , n439054 );
buf ( n439056 , n439055 );
buf ( n439057 , n439056 );
not ( n439058 , n439057 );
buf ( n439059 , n386598 );
buf ( n439060 , n386575 );
and ( n439061 , n439059 , n439060 );
not ( n439062 , n439059 );
buf ( n439063 , n386578 );
and ( n439064 , n439062 , n439063 );
nor ( n439065 , n439061 , n439064 );
buf ( n439066 , n439065 );
buf ( n439067 , n439066 );
not ( n439068 , n439067 );
buf ( n439069 , n39060 );
buf ( n439070 , n439069 );
not ( n439071 , n439070 );
or ( n439072 , n439068 , n439071 );
buf ( n439073 , n439066 );
not ( n439074 , n439073 );
buf ( n439075 , n439074 );
buf ( n439076 , n439075 );
not ( n439077 , n439069 );
buf ( n439078 , n439077 );
nand ( n439079 , n439076 , n439078 );
buf ( n439080 , n439079 );
buf ( n439081 , n439080 );
nand ( n439082 , n439072 , n439081 );
buf ( n439083 , n439082 );
buf ( n439084 , n439083 );
not ( n439085 , n439084 );
or ( n439086 , n439058 , n439085 );
buf ( n439087 , n439056 );
buf ( n439088 , n439083 );
or ( n439089 , n439087 , n439088 );
xor ( n439090 , n438677 , n438698 );
and ( n439091 , n439090 , n438746 );
and ( n439092 , n438677 , n438698 );
or ( n439093 , n439091 , n439092 );
buf ( n439094 , n439093 );
buf ( n439095 , n439094 );
nand ( n439096 , n439089 , n439095 );
buf ( n439097 , n439096 );
buf ( n439098 , n439097 );
nand ( n439099 , n439086 , n439098 );
buf ( n439100 , n439099 );
buf ( n439101 , n439100 );
not ( n439102 , n439101 );
buf ( n439103 , n439102 );
buf ( n439104 , n439103 );
not ( n439105 , n439104 );
or ( n439106 , n439044 , n439105 );
xor ( n439107 , n386520 , n386524 );
xor ( n439108 , n439107 , n386546 );
buf ( n439109 , n439108 );
buf ( n439110 , n439109 );
xor ( n439111 , n438871 , n438881 );
and ( n439112 , n439111 , n438898 );
and ( n439113 , n438871 , n438881 );
or ( n439114 , n439112 , n439113 );
buf ( n439115 , n439114 );
buf ( n439116 , n439115 );
or ( n439117 , n439110 , n439116 );
xor ( n439118 , n438770 , n438783 );
and ( n439119 , n439118 , n438828 );
and ( n439120 , n438770 , n438783 );
or ( n439121 , n439119 , n439120 );
buf ( n439122 , n439121 );
buf ( n439123 , n439122 );
nand ( n439124 , n439117 , n439123 );
buf ( n439125 , n439124 );
buf ( n439126 , n439125 );
buf ( n439127 , n439115 );
buf ( n439128 , n439109 );
nand ( n439129 , n439127 , n439128 );
buf ( n439130 , n439129 );
buf ( n439131 , n439130 );
nand ( n439132 , n439126 , n439131 );
buf ( n439133 , n439132 );
buf ( n439134 , n439133 );
nand ( n439135 , n439106 , n439134 );
buf ( n439136 , n439135 );
buf ( n439137 , n439136 );
buf ( n439138 , n439100 );
buf ( n439139 , n439039 );
nand ( n439140 , n439138 , n439139 );
buf ( n439141 , n439140 );
buf ( n439142 , n439141 );
and ( n439143 , n439137 , n439142 );
buf ( n439144 , n439143 );
xnor ( n439145 , n439036 , n439144 );
xor ( n439146 , n438974 , n438981 );
xor ( n439147 , n439146 , n439011 );
buf ( n439148 , n439147 );
not ( n439149 , n438924 );
not ( n439150 , n438900 );
or ( n439151 , n439149 , n439150 );
not ( n439152 , n438921 );
not ( n439153 , n438903 );
or ( n439154 , n439152 , n439153 );
nand ( n439155 , n439154 , n438867 );
nand ( n439156 , n439151 , n439155 );
buf ( n439157 , n439156 );
not ( n439158 , n439157 );
buf ( n439159 , n439115 );
buf ( n439160 , n439109 );
xor ( n439161 , n439159 , n439160 );
buf ( n439162 , n439122 );
xnor ( n439163 , n439161 , n439162 );
buf ( n439164 , n439163 );
buf ( n439165 , n439164 );
not ( n439166 , n439165 );
buf ( n439167 , n439166 );
buf ( n439168 , n439167 );
not ( n439169 , n439168 );
or ( n439170 , n439158 , n439169 );
buf ( n439171 , n439156 );
not ( n439172 , n439171 );
buf ( n439173 , n439172 );
buf ( n439174 , n439173 );
not ( n439175 , n439174 );
buf ( n439176 , n439164 );
not ( n439177 , n439176 );
or ( n439178 , n439175 , n439177 );
buf ( n439179 , n438748 );
buf ( n439180 , n438830 );
or ( n439181 , n439179 , n439180 );
buf ( n439182 , n438763 );
nand ( n439183 , n439181 , n439182 );
buf ( n439184 , n439183 );
buf ( n439185 , n439184 );
buf ( n439186 , n438748 );
buf ( n439187 , n438830 );
nand ( n439188 , n439186 , n439187 );
buf ( n439189 , n439188 );
buf ( n439190 , n439189 );
nand ( n439191 , n439185 , n439190 );
buf ( n439192 , n439191 );
buf ( n439193 , n439192 );
nand ( n439194 , n439178 , n439193 );
buf ( n439195 , n439194 );
buf ( n439196 , n439195 );
nand ( n439197 , n439170 , n439196 );
buf ( n439198 , n439197 );
buf ( n439199 , n439198 );
not ( n439200 , n439199 );
buf ( n439201 , n439200 );
xor ( n439202 , n439148 , n439201 );
buf ( n439203 , n439039 );
buf ( n439204 , n439133 );
xor ( n439205 , n439203 , n439204 );
buf ( n439206 , n439205 );
buf ( n439207 , n439206 );
buf ( n439208 , n439103 );
and ( n439209 , n439207 , n439208 );
not ( n439210 , n439207 );
buf ( n439211 , n439100 );
and ( n439212 , n439210 , n439211 );
nor ( n439213 , n439209 , n439212 );
buf ( n439214 , n439213 );
and ( n439215 , n439202 , n439214 );
and ( n439216 , n439148 , n439201 );
or ( n439217 , n439215 , n439216 );
nand ( n439218 , n439145 , n439217 );
buf ( n439219 , n439083 );
buf ( n439220 , n439094 );
xor ( n439221 , n439219 , n439220 );
buf ( n439222 , n439056 );
xnor ( n439223 , n439221 , n439222 );
buf ( n439224 , n439223 );
buf ( n439225 , n439224 );
xor ( n439226 , n438862 , n438929 );
and ( n439227 , n439226 , n438945 );
and ( n439228 , n438862 , n438929 );
or ( n439229 , n439227 , n439228 );
buf ( n439230 , n439229 );
buf ( n439231 , n439230 );
xor ( n439232 , n439225 , n439231 );
buf ( n439233 , n439164 );
buf ( n439234 , n439173 );
and ( n439235 , n439233 , n439234 );
not ( n439236 , n439233 );
buf ( n439237 , n439156 );
and ( n439238 , n439236 , n439237 );
nor ( n439239 , n439235 , n439238 );
buf ( n439240 , n439239 );
buf ( n439241 , n439240 );
buf ( n439242 , n439192 );
not ( n439243 , n439242 );
buf ( n439244 , n439243 );
buf ( n439245 , n439244 );
and ( n439246 , n439241 , n439245 );
not ( n439247 , n439241 );
buf ( n439248 , n439192 );
and ( n439249 , n439247 , n439248 );
nor ( n439250 , n439246 , n439249 );
buf ( n439251 , n439250 );
buf ( n439252 , n439251 );
and ( n439253 , n439232 , n439252 );
and ( n439254 , n439225 , n439231 );
or ( n439255 , n439253 , n439254 );
buf ( n439256 , n439255 );
xor ( n439257 , n439148 , n439201 );
xor ( n439258 , n439257 , n439214 );
nand ( n439259 , n439256 , n439258 );
xor ( n439260 , n439225 , n439231 );
xor ( n439261 , n439260 , n439252 );
buf ( n439262 , n439261 );
xor ( n439263 , n438838 , n438851 );
and ( n439264 , n439263 , n438948 );
and ( n439265 , n438838 , n438851 );
or ( n439266 , n439264 , n439265 );
buf ( n439267 , n439266 );
nand ( n439268 , n439262 , n439267 );
nand ( n439269 , n439218 , n439259 , n439268 );
buf ( n439270 , n439269 );
buf ( n439271 , n439024 );
buf ( n439272 , n386274 );
and ( n439273 , n439271 , n439272 );
not ( n439274 , n439271 );
buf ( n439275 , n439031 );
and ( n439276 , n439274 , n439275 );
or ( n439277 , n439273 , n439276 );
buf ( n439278 , n439277 );
or ( n439279 , n439278 , n439015 );
and ( n439280 , n439279 , n439144 );
and ( n439281 , n439278 , n439015 );
nor ( n439282 , n439280 , n439281 );
not ( n439283 , n439282 );
not ( n439284 , n39124 );
not ( n439285 , n386631 );
not ( n439286 , n439285 );
or ( n439287 , n439284 , n439286 );
nand ( n439288 , n386631 , n386655 );
nand ( n439289 , n439287 , n439288 );
and ( n439290 , n439289 , n386649 );
not ( n439291 , n439289 );
and ( n439292 , n439291 , n39118 );
nor ( n439293 , n439290 , n439292 );
nand ( n439294 , n439283 , n439293 );
buf ( n439295 , n439294 );
not ( n439296 , n439295 );
buf ( n439297 , n439296 );
buf ( n439298 , n439297 );
nor ( n439299 , n439270 , n439298 );
buf ( n439300 , n439299 );
and ( n439301 , n435312 , n437326 , n438955 , n439300 );
nand ( n439302 , n433185 , n439301 );
buf ( n439303 , n437305 );
not ( n439304 , n439303 );
not ( n439305 , n437324 );
buf ( n439306 , n436343 );
buf ( n439307 , n436348 );
nand ( n439308 , n439306 , n439307 );
buf ( n439309 , n439308 );
or ( n439310 , n436337 , n439309 );
buf ( n439311 , n436309 );
buf ( n439312 , n436336 );
nand ( n439313 , n439311 , n439312 );
buf ( n439314 , n439313 );
nand ( n439315 , n439310 , n439314 );
not ( n439316 , n439315 );
or ( n439317 , n439305 , n439316 );
not ( n439318 , n437321 );
not ( n439319 , n437323 );
nand ( n439320 , n439318 , n439319 );
nand ( n439321 , n439317 , n439320 );
not ( n439322 , n439321 );
or ( n439323 , n439304 , n439322 );
nor ( n439324 , n439262 , n439267 );
not ( n439325 , n439324 );
not ( n439326 , n439259 );
or ( n439327 , n439325 , n439326 );
buf ( n439328 , n439258 );
not ( n439329 , n439328 );
buf ( n439330 , n439329 );
buf ( n439331 , n439256 );
not ( n439332 , n439331 );
buf ( n439333 , n439332 );
nand ( n439334 , n439330 , n439333 );
nand ( n439335 , n439327 , n439334 );
nand ( n439336 , n439335 , n439294 , n439218 );
nor ( n439337 , n439217 , n439145 );
and ( n439338 , n439337 , n439294 );
not ( n439339 , n439282 );
nor ( n439340 , n439339 , n439293 );
nor ( n439341 , n439338 , n439340 );
nand ( n439342 , n439336 , n439341 );
not ( n439343 , n437304 );
nand ( n439344 , n439343 , n437261 );
not ( n439345 , n439344 );
nor ( n439346 , n439342 , n439345 );
nand ( n439347 , n439323 , n439346 );
not ( n439348 , n438951 );
buf ( n439349 , n438658 );
not ( n439350 , n439349 );
not ( n439351 , n438189 );
not ( n439352 , n437331 );
nor ( n439353 , n439352 , n437772 );
not ( n439354 , n439353 );
or ( n439355 , n439351 , n439354 );
buf ( n439356 , n438183 );
not ( n439357 , n439356 );
buf ( n439358 , n439357 );
buf ( n439359 , n438188 );
not ( n439360 , n439359 );
buf ( n439361 , n439360 );
nand ( n439362 , n439358 , n439361 );
nand ( n439363 , n439355 , n439362 );
buf ( n439364 , n439363 );
not ( n439365 , n439364 );
or ( n439366 , n439350 , n439365 );
buf ( n439367 , n438652 );
buf ( n439368 , n438657 );
or ( n439369 , n439367 , n439368 );
buf ( n439370 , n439369 );
buf ( n439371 , n439370 );
nand ( n439372 , n439366 , n439371 );
buf ( n439373 , n439372 );
not ( n439374 , n439373 );
or ( n439375 , n439348 , n439374 );
not ( n439376 , n438950 );
nand ( n439377 , n439376 , n438670 );
nand ( n439378 , n439375 , n439377 );
nor ( n439379 , n439347 , n439378 );
not ( n439380 , n439379 );
not ( n439381 , n434262 );
buf ( n439382 , n434269 );
not ( n439383 , n439382 );
buf ( n439384 , n439383 );
nand ( n439385 , n439381 , n439384 );
nand ( n439386 , n433740 , n433199 );
nand ( n439387 , n439385 , n439386 );
not ( n439388 , n434270 );
nor ( n439389 , n434804 , n439388 );
not ( n439390 , n435309 );
nand ( n439391 , n439387 , n439389 , n439390 );
buf ( n439392 , n435301 );
buf ( n439393 , n435306 );
nand ( n439394 , n439392 , n439393 );
buf ( n439395 , n439394 );
not ( n439396 , n439395 );
nand ( n439397 , n434803 , n434281 );
not ( n439398 , n439397 );
or ( n439399 , n439396 , n439398 );
nand ( n439400 , n439399 , n439390 );
nand ( n439401 , n439391 , n439400 );
nand ( n439402 , n439401 , n437326 );
not ( n439403 , n439402 );
or ( n439404 , n439380 , n439403 );
not ( n439405 , n438951 );
not ( n439406 , n439373 );
or ( n439407 , n439405 , n439406 );
nand ( n439408 , n439407 , n439377 );
not ( n439409 , n439408 );
not ( n439410 , n439342 );
buf ( n439411 , n439410 );
buf ( n439412 , n438952 );
nand ( n439413 , n439411 , n439412 );
buf ( n439414 , n439413 );
not ( n439415 , n439414 );
and ( n439416 , n439409 , n439415 );
buf ( n439417 , n439300 );
buf ( n439418 , n439342 );
nor ( n439419 , n439417 , n439418 );
buf ( n439420 , n439419 );
nor ( n439421 , n439416 , n439420 );
nand ( n439422 , n439404 , n439421 );
not ( n439423 , n396187 );
nor ( n439424 , n52569 , n399870 );
nand ( n439425 , n51961 , n439424 );
not ( n439426 , n439425 );
not ( n439427 , n51960 );
not ( n439428 , n439427 );
not ( n439429 , n50675 );
not ( n439430 , n439429 );
or ( n439431 , n439428 , n439430 );
buf ( n439432 , n399921 );
not ( n439433 , n439432 );
buf ( n439434 , n439433 );
not ( n439435 , n52612 );
nand ( n439436 , n439434 , n439435 );
nand ( n439437 , n439431 , n439436 );
or ( n439438 , n439426 , n439437 );
nand ( n439439 , n399929 , n399934 );
and ( n439440 , n439439 , n52613 );
nand ( n439441 , n439438 , n439440 );
buf ( n439442 , n439441 );
or ( n439443 , n399929 , n399934 );
buf ( n439444 , n439443 );
nand ( n439445 , n439442 , n439444 );
buf ( n439446 , n439445 );
not ( n439447 , n439446 );
or ( n439448 , n439423 , n439447 );
buf ( n439449 , n393715 );
buf ( n439450 , n45580 );
nor ( n439451 , n439449 , n439450 );
buf ( n439452 , n439451 );
buf ( n439453 , n439452 );
buf ( n439454 , n47148 );
buf ( n439455 , n393722 );
nor ( n439456 , n439454 , n439455 );
buf ( n439457 , n439456 );
buf ( n439458 , n439457 );
nor ( n439459 , n439453 , n439458 );
buf ( n439460 , n439459 );
nor ( n439461 , n47154 , n395622 );
nand ( n439462 , n439461 , n394596 );
nand ( n439463 , n439460 , n439462 );
buf ( n439464 , n393718 );
buf ( n439465 , n396184 );
buf ( n439466 , n439465 );
buf ( n439467 , n439466 );
and ( n439468 , n439463 , n439464 , n439467 );
buf ( n439469 , n48191 );
not ( n439470 , n439469 );
buf ( n439471 , n396181 );
buf ( n439472 , n439471 );
nor ( n439473 , n439470 , n439472 );
buf ( n439474 , n439473 );
nor ( n439475 , n439468 , n439474 );
nand ( n439476 , n439448 , n439475 );
not ( n439477 , n439476 );
not ( n439478 , n439477 );
buf ( n439479 , n52572 );
buf ( n439480 , n52623 );
and ( n439481 , n439479 , n439480 );
buf ( n439482 , n439481 );
and ( n439483 , n439482 , n396187 );
nand ( n439484 , n410004 , n410013 );
not ( n439485 , n439484 );
nor ( n439486 , n58469 , n439485 );
not ( n439487 , n439486 );
buf ( n439488 , n60626 );
buf ( n439489 , n408538 );
nand ( n439490 , n439488 , n439489 );
buf ( n439491 , n439490 );
nand ( n439492 , n408546 , n62967 );
nand ( n439493 , n439491 , n439492 );
nand ( n439494 , n439493 , n62998 , n61500 );
buf ( n439495 , n63003 );
buf ( n439496 , n410010 );
nand ( n439497 , n439495 , n439496 );
buf ( n439498 , n439497 );
nand ( n439499 , n409985 , n62994 );
buf ( n439500 , n439499 );
nand ( n439501 , n439494 , n439498 , n439500 );
not ( n439502 , n439501 );
or ( n439503 , n439487 , n439502 );
buf ( n439504 , n54684 );
not ( n439505 , n439504 );
buf ( n439506 , n439505 );
nand ( n439507 , n56298 , n56302 );
buf ( n439508 , n403522 );
not ( n439509 , n439508 );
buf ( n439510 , n439509 );
nand ( n439511 , n439506 , n439507 , n439510 );
not ( n439512 , n56298 );
not ( n439513 , n56302 );
nand ( n439514 , n439512 , n439513 );
nand ( n439515 , n439511 , n439514 );
nor ( n439516 , n404445 , n58465 );
not ( n439517 , n439516 );
nand ( n439518 , n404440 , n404436 );
not ( n439519 , n439518 );
or ( n439520 , n439517 , n439519 );
buf ( n439521 , n404440 );
not ( n439522 , n439521 );
buf ( n439523 , n439522 );
buf ( n439524 , n404436 );
not ( n439525 , n439524 );
buf ( n439526 , n439525 );
nand ( n439527 , n439523 , n439526 );
nand ( n439528 , n439520 , n439527 );
nor ( n439529 , n439515 , n439528 );
nand ( n439530 , n439503 , n439529 );
not ( n439531 , n439514 );
buf ( n439532 , n56293 );
not ( n439533 , n439532 );
buf ( n439534 , n439533 );
not ( n439535 , n439534 );
or ( n439536 , n439531 , n439535 );
not ( n439537 , n56303 );
not ( n439538 , n439537 );
nand ( n439539 , n439536 , n439538 );
not ( n439540 , n439539 );
nand ( n439541 , n439483 , n439530 , n439540 );
not ( n439542 , n439541 );
or ( n439543 , n439478 , n439542 );
nand ( n439544 , n439543 , n439301 );
nand ( n439545 , n439302 , n439422 , n439544 );
not ( n439546 , n439545 );
or ( n439547 , n40563 , n439546 );
not ( n439548 , n40558 );
not ( n439549 , n387816 );
buf ( n439550 , n386989 );
not ( n439551 , n439550 );
buf ( n439552 , n385957 );
not ( n439553 , n439552 );
buf ( n439554 , n39146 );
buf ( n439555 , n39132 );
nand ( n439556 , n439554 , n439555 );
buf ( n439557 , n439556 );
or ( n439558 , n439557 , n39163 );
buf ( n439559 , n39152 );
buf ( n439560 , n386694 );
nand ( n439561 , n439559 , n439560 );
buf ( n439562 , n439561 );
nand ( n439563 , n439558 , n439562 );
buf ( n439564 , n439563 );
not ( n439565 , n439564 );
or ( n439566 , n439553 , n439565 );
buf ( n439567 , n385603 );
buf ( n439568 , n38410 );
or ( n439569 , n439567 , n439568 );
buf ( n439570 , n439569 );
buf ( n439571 , n439570 );
nand ( n439572 , n439566 , n439571 );
buf ( n439573 , n439572 );
buf ( n439574 , n439573 );
not ( n439575 , n439574 );
or ( n439576 , n439551 , n439575 );
buf ( n439577 , n386986 );
buf ( n439578 , n386980 );
or ( n439579 , n439577 , n439578 );
buf ( n439580 , n439579 );
buf ( n439581 , n439580 );
nand ( n439582 , n439576 , n439581 );
buf ( n439583 , n439582 );
not ( n439584 , n439583 );
or ( n439585 , n439549 , n439584 );
buf ( n439586 , n387753 );
not ( n439587 , n439586 );
not ( n439588 , n40040 );
buf ( n439589 , n387795 );
buf ( n439590 , n387811 );
buf ( n439591 , n40307 );
nand ( n439592 , n439590 , n439591 );
buf ( n439593 , n439592 );
buf ( n439594 , n439593 );
or ( n439595 , n439589 , n439594 );
buf ( n439596 , n40258 );
buf ( n439597 , n387792 );
nand ( n439598 , n439596 , n439597 );
buf ( n439599 , n439598 );
buf ( n439600 , n439599 );
nand ( n439601 , n439595 , n439600 );
buf ( n439602 , n439601 );
not ( n439603 , n439602 );
or ( n439604 , n439588 , n439603 );
buf ( n439605 , n387492 );
buf ( n439606 , n40039 );
or ( n439607 , n439605 , n439606 );
buf ( n439608 , n439607 );
nand ( n439609 , n439604 , n439608 );
buf ( n439610 , n439609 );
not ( n439611 , n439610 );
or ( n439612 , n439587 , n439611 );
buf ( n439613 , n387744 );
buf ( n439614 , n387750 );
or ( n439615 , n439613 , n439614 );
buf ( n439616 , n439615 );
buf ( n439617 , n439616 );
nand ( n439618 , n439612 , n439617 );
buf ( n439619 , n439618 );
buf ( n439620 , n439619 );
not ( n439621 , n439620 );
buf ( n439622 , n439621 );
nand ( n439623 , n439585 , n439622 );
not ( n439624 , n439623 );
or ( n439625 , n439548 , n439624 );
buf ( n439626 , n388038 );
not ( n439627 , n439626 );
nand ( n439628 , n387928 , n387835 );
or ( n439629 , n439628 , n387980 );
buf ( n439630 , n387971 );
buf ( n439631 , n387977 );
nand ( n439632 , n439630 , n439631 );
buf ( n439633 , n439632 );
nand ( n439634 , n439629 , n439633 );
buf ( n439635 , n439634 );
not ( n439636 , n439635 );
or ( n439637 , n439627 , n439636 );
buf ( n439638 , n388035 );
not ( n439639 , n439638 );
buf ( n439640 , n387991 );
nand ( n439641 , n439639 , n439640 );
buf ( n439642 , n439641 );
buf ( n439643 , n439642 );
nand ( n439644 , n439637 , n439643 );
buf ( n439645 , n439644 );
and ( n439646 , n439645 , n388052 );
buf ( n439647 , n388042 );
not ( n439648 , n439647 );
buf ( n439649 , n388049 );
nor ( n439650 , n439648 , n439649 );
buf ( n439651 , n439650 );
nor ( n439652 , n439646 , n439651 );
nand ( n439653 , n439625 , n439652 );
not ( n439654 , n439653 );
nand ( n439655 , n439547 , n439654 );
not ( n439656 , n439655 );
or ( n439657 , n36167 , n439656 );
not ( n439658 , n383736 );
and ( n439659 , n439658 , n383715 );
not ( n439660 , n439659 );
nand ( n439661 , n439657 , n439660 );
buf ( n439662 , n439661 );
and ( n439663 , n439662 , n383336 );
not ( n439664 , n439662 );
and ( n439665 , n439664 , n383332 );
nor ( n439666 , n439663 , n439665 );
buf ( n439667 , n439666 );
buf ( n439668 , n439651 );
not ( n439669 , n439668 );
buf ( n439670 , n388052 );
nand ( n439671 , n439669 , n439670 );
buf ( n439672 , n439671 );
buf ( n439673 , n439672 );
buf ( n439674 , n439672 );
not ( n439675 , n439674 );
buf ( n439676 , n439675 );
buf ( n439677 , n439676 );
buf ( n439678 , n388038 );
not ( n439679 , n439678 );
not ( n439680 , n387819 );
nor ( n439681 , n439680 , n387986 );
not ( n439682 , n439681 );
not ( n439683 , n439545 );
or ( n439684 , n439682 , n439683 );
not ( n439685 , n387986 );
nand ( n439686 , n439685 , n439623 );
nand ( n439687 , n439684 , n439686 );
buf ( n439688 , n439687 );
not ( n439689 , n439688 );
or ( n439690 , n439679 , n439689 );
buf ( n439691 , n439645 );
not ( n439692 , n439691 );
buf ( n439693 , n439692 );
buf ( n439694 , n439693 );
nand ( n439695 , n439690 , n439694 );
buf ( n439696 , n439695 );
buf ( n439697 , n439696 );
and ( n439698 , n439697 , n439677 );
not ( n439699 , n439697 );
and ( n439700 , n439699 , n439673 );
nor ( n439701 , n439698 , n439700 );
buf ( n439702 , n439701 );
buf ( n439703 , n439633 );
buf ( n439704 , n387983 );
nand ( n439705 , n439703 , n439704 );
buf ( n439706 , n439705 );
buf ( n439707 , n439706 );
buf ( n439708 , n439706 );
not ( n439709 , n439708 );
buf ( n439710 , n439709 );
buf ( n439711 , n439710 );
not ( n439712 , n387931 );
not ( n439713 , n387819 );
nand ( n439714 , n439302 , n439544 , n439422 );
not ( n439715 , n439714 );
or ( n439716 , n439713 , n439715 );
not ( n439717 , n439623 );
nand ( n439718 , n439716 , n439717 );
not ( n439719 , n439718 );
or ( n439720 , n439712 , n439719 );
buf ( n439721 , n439628 );
nand ( n439722 , n439720 , n439721 );
buf ( n439723 , n439722 );
and ( n439724 , n439723 , n439711 );
not ( n439725 , n439723 );
and ( n439726 , n439725 , n439707 );
nor ( n439727 , n439724 , n439726 );
buf ( n439728 , n439727 );
not ( n439729 , n387795 );
nand ( n439730 , n439729 , n439599 );
buf ( n439731 , n439730 );
buf ( n439732 , n439730 );
not ( n439733 , n439732 );
buf ( n439734 , n439733 );
buf ( n439735 , n439734 );
buf ( n439736 , n40311 );
not ( n439737 , n439736 );
not ( n439738 , n386992 );
not ( n439739 , n439714 );
or ( n439740 , n439738 , n439739 );
buf ( n439741 , n439583 );
not ( n439742 , n439741 );
buf ( n439743 , n439742 );
nand ( n439744 , n439740 , n439743 );
buf ( n439745 , n439744 );
not ( n439746 , n439745 );
or ( n439747 , n439737 , n439746 );
buf ( n439748 , n439593 );
buf ( n439749 , n439748 );
buf ( n439750 , n439749 );
buf ( n439751 , n439750 );
nand ( n439752 , n439747 , n439751 );
buf ( n439753 , n439752 );
buf ( n439754 , n439753 );
and ( n439755 , n439754 , n439735 );
not ( n439756 , n439754 );
and ( n439757 , n439756 , n439731 );
nor ( n439758 , n439755 , n439757 );
buf ( n439759 , n439758 );
buf ( n439760 , n388038 );
buf ( n439761 , n439642 );
nand ( n439762 , n439760 , n439761 );
buf ( n439763 , n439762 );
buf ( n439764 , n439763 );
not ( n439765 , n439764 );
buf ( n439766 , n439765 );
buf ( n439767 , n439766 );
buf ( n439768 , n439763 );
buf ( n439769 , n439687 );
buf ( n439770 , n439634 );
nor ( n439771 , n439769 , n439770 );
buf ( n439772 , n439771 );
buf ( n439773 , n439772 );
and ( n439774 , n439773 , n439768 );
not ( n439775 , n439773 );
and ( n439776 , n439775 , n439767 );
nor ( n439777 , n439774 , n439776 );
buf ( n439778 , n439777 );
buf ( n439779 , n40040 );
buf ( n439780 , n439608 );
nand ( n439781 , n439779 , n439780 );
buf ( n439782 , n439781 );
buf ( n439783 , n439782 );
not ( n439784 , n439783 );
buf ( n439785 , n439784 );
buf ( n439786 , n439785 );
buf ( n439787 , n439782 );
not ( n439788 , n386992 );
nor ( n439789 , n439788 , n40312 );
not ( n439790 , n439789 );
not ( n439791 , n439714 );
or ( n439792 , n439790 , n439791 );
not ( n439793 , n40312 );
nand ( n439794 , n439793 , n439583 );
nand ( n439795 , n439792 , n439794 );
buf ( n439796 , n439602 );
nor ( n439797 , n439795 , n439796 );
buf ( n439798 , n439797 );
and ( n439799 , n439798 , n439787 );
not ( n439800 , n439798 );
and ( n439801 , n439800 , n439786 );
nor ( n439802 , n439799 , n439801 );
buf ( n439803 , n439802 );
not ( n439804 , n439337 );
buf ( n439805 , n439218 );
nand ( n439806 , n439804 , n439805 );
buf ( n439807 , n439806 );
not ( n439808 , n439807 );
buf ( n439809 , n439808 );
buf ( n439810 , n439809 );
buf ( n439811 , n439806 );
nor ( n439812 , n436350 , n437325 , n437306 );
not ( n439813 , n439812 );
not ( n439814 , n438952 );
buf ( n439815 , n435312 );
buf ( n439816 , n439815 );
buf ( n439817 , n439816 );
nand ( n439818 , n439814 , n439817 );
nor ( n439819 , n439813 , n439818 );
not ( n439820 , n439819 );
nand ( n439821 , n439483 , n439530 , n439540 );
and ( n439822 , n433184 , n439477 , n439821 );
not ( n439823 , n439822 );
not ( n439824 , n439823 );
or ( n439825 , n439820 , n439824 );
and ( n439826 , n439321 , n439303 );
nor ( n439827 , n439826 , n439345 );
nand ( n439828 , n439827 , n439402 );
not ( n439829 , n438658 );
nor ( n439830 , n439829 , n438190 );
and ( n439831 , n439830 , n438951 );
and ( n439832 , n439828 , n439831 );
buf ( n439833 , n439408 );
nor ( n439834 , n439832 , n439833 );
nand ( n439835 , n439825 , n439834 );
and ( n439836 , n439268 , n439259 );
and ( n439837 , n439835 , n439836 );
buf ( n439838 , n439259 );
not ( n439839 , n439838 );
nor ( n439840 , n439262 , n439267 );
buf ( n439841 , n439840 );
not ( n439842 , n439841 );
or ( n439843 , n439839 , n439842 );
buf ( n439844 , n439334 );
nand ( n439845 , n439843 , n439844 );
buf ( n439846 , n439845 );
nor ( n439847 , n439837 , n439846 );
buf ( n439848 , n439847 );
and ( n439849 , n439848 , n439811 );
not ( n439850 , n439848 );
and ( n439851 , n439850 , n439810 );
nor ( n439852 , n439849 , n439851 );
buf ( n439853 , n439852 );
nand ( n439854 , n439562 , n39164 );
buf ( n439855 , n439854 );
buf ( n439856 , n439854 );
not ( n439857 , n439856 );
buf ( n439858 , n439857 );
buf ( n439859 , n439858 );
buf ( n439860 , n39148 );
not ( n439861 , n439860 );
buf ( n439862 , n439545 );
buf ( n439863 , n439862 );
not ( n439864 , n439863 );
or ( n439865 , n439861 , n439864 );
buf ( n439866 , n439557 );
buf ( n439867 , n439866 );
nand ( n439868 , n439865 , n439867 );
buf ( n439869 , n439868 );
buf ( n439870 , n439869 );
and ( n439871 , n439870 , n439859 );
not ( n439872 , n439870 );
and ( n439873 , n439872 , n439855 );
nor ( n439874 , n439871 , n439873 );
buf ( n439875 , n439874 );
nand ( n439876 , n387931 , n439721 );
buf ( n439877 , n439876 );
buf ( n439878 , n439876 );
not ( n439879 , n439878 );
buf ( n439880 , n439879 );
buf ( n439881 , n439880 );
buf ( n439882 , n439718 );
and ( n439883 , n439882 , n439881 );
not ( n439884 , n439882 );
and ( n439885 , n439884 , n439877 );
nor ( n439886 , n439883 , n439885 );
buf ( n439887 , n439886 );
buf ( n439888 , n439750 );
buf ( n439889 , n40311 );
nand ( n439890 , n439888 , n439889 );
buf ( n439891 , n439890 );
buf ( n439892 , n439891 );
buf ( n439893 , n439891 );
not ( n439894 , n439893 );
buf ( n439895 , n439894 );
buf ( n439896 , n439895 );
buf ( n439897 , n439744 );
and ( n439898 , n439897 , n439896 );
not ( n439899 , n439897 );
and ( n439900 , n439899 , n439892 );
nor ( n439901 , n439898 , n439900 );
buf ( n439902 , n439901 );
buf ( n439903 , n439580 );
buf ( n439904 , n386989 );
nand ( n439905 , n439903 , n439904 );
buf ( n439906 , n439905 );
buf ( n439907 , n439906 );
buf ( n439908 , n439906 );
not ( n439909 , n439908 );
buf ( n439910 , n439909 );
buf ( n439911 , n439910 );
buf ( n439912 , n386700 );
not ( n439913 , n439912 );
buf ( n439914 , n439862 );
not ( n439915 , n439914 );
or ( n439916 , n439913 , n439915 );
buf ( n439917 , n439573 );
not ( n439918 , n439917 );
buf ( n439919 , n439918 );
buf ( n439920 , n439919 );
nand ( n439921 , n439916 , n439920 );
buf ( n439922 , n439921 );
buf ( n439923 , n439922 );
and ( n439924 , n439923 , n439911 );
not ( n439925 , n439923 );
and ( n439926 , n439925 , n439907 );
nor ( n439927 , n439924 , n439926 );
buf ( n439928 , n439927 );
buf ( n439929 , n439570 );
buf ( n439930 , n385957 );
nand ( n439931 , n439929 , n439930 );
buf ( n439932 , n439931 );
buf ( n439933 , n439932 );
buf ( n439934 , n439932 );
not ( n439935 , n439934 );
buf ( n439936 , n439935 );
buf ( n439937 , n439936 );
buf ( n439938 , n39165 );
not ( n439939 , n439938 );
buf ( n439940 , n439939 );
buf ( n439941 , n439940 );
not ( n439942 , n439941 );
buf ( n439943 , n439862 );
not ( n439944 , n439943 );
or ( n439945 , n439942 , n439944 );
buf ( n439946 , n439563 );
buf ( n439947 , n439946 );
not ( n439948 , n439947 );
buf ( n439949 , n439948 );
buf ( n439950 , n439949 );
nand ( n439951 , n439945 , n439950 );
buf ( n439952 , n439951 );
buf ( n439953 , n439952 );
and ( n439954 , n439953 , n439937 );
not ( n439955 , n439953 );
and ( n439956 , n439955 , n439933 );
nor ( n439957 , n439954 , n439956 );
buf ( n439958 , n439957 );
not ( n439959 , n439340 );
nand ( n439960 , n439959 , n439294 );
buf ( n439961 , n439960 );
buf ( n439962 , n439960 );
not ( n439963 , n439962 );
buf ( n439964 , n439963 );
buf ( n439965 , n439964 );
buf ( n439966 , n439269 );
not ( n439967 , n439966 );
buf ( n439968 , n439967 );
buf ( n439969 , n439968 );
not ( n439970 , n439969 );
buf ( n439971 , n439835 );
not ( n439972 , n439971 );
or ( n439973 , n439970 , n439972 );
not ( n439974 , n439805 );
not ( n439975 , n439335 );
or ( n439976 , n439974 , n439975 );
nand ( n439977 , n439976 , n439804 );
buf ( n439978 , n439977 );
not ( n439979 , n439978 );
buf ( n439980 , n439979 );
buf ( n439981 , n439980 );
nand ( n439982 , n439973 , n439981 );
buf ( n439983 , n439982 );
buf ( n439984 , n439983 );
and ( n439985 , n439984 , n439965 );
not ( n439986 , n439984 );
and ( n439987 , n439986 , n439961 );
nor ( n439988 , n439985 , n439987 );
buf ( n439989 , n439988 );
buf ( n439990 , n439334 );
buf ( n439991 , n439259 );
nand ( n439992 , n439990 , n439991 );
buf ( n439993 , n439992 );
buf ( n439994 , n439993 );
buf ( n439995 , n439993 );
not ( n439996 , n439995 );
buf ( n439997 , n439996 );
buf ( n439998 , n439997 );
buf ( n439999 , n439268 );
not ( n440000 , n439999 );
buf ( n440001 , n439835 );
not ( n440002 , n440001 );
or ( n440003 , n440000 , n440002 );
buf ( n440004 , n439840 );
not ( n440005 , n440004 );
buf ( n440006 , n440005 );
buf ( n440007 , n440006 );
nand ( n440008 , n440003 , n440007 );
buf ( n440009 , n440008 );
buf ( n440010 , n440009 );
and ( n440011 , n440010 , n439998 );
not ( n440012 , n440010 );
and ( n440013 , n440012 , n439994 );
nor ( n440014 , n440011 , n440013 );
buf ( n440015 , n440014 );
buf ( n440016 , n440006 );
buf ( n440017 , n439268 );
nand ( n440018 , n440016 , n440017 );
buf ( n440019 , n440018 );
buf ( n440020 , n440019 );
buf ( n440021 , n440019 );
not ( n440022 , n440021 );
buf ( n440023 , n440022 );
buf ( n440024 , n440023 );
buf ( n440025 , n438955 );
not ( n440026 , n440025 );
and ( n440027 , n439812 , n439817 );
not ( n440028 , n440027 );
not ( n440029 , n439823 );
or ( n440030 , n440028 , n440029 );
not ( n440031 , n439828 );
nand ( n440032 , n440030 , n440031 );
buf ( n440033 , n440032 );
not ( n440034 , n440033 );
or ( n440035 , n440026 , n440034 );
not ( n440036 , n439833 );
buf ( n440037 , n440036 );
nand ( n440038 , n440035 , n440037 );
buf ( n440039 , n440038 );
buf ( n440040 , n440039 );
and ( n440041 , n440040 , n440024 );
not ( n440042 , n440040 );
and ( n440043 , n440042 , n440020 );
nor ( n440044 , n440041 , n440043 );
buf ( n440045 , n440044 );
buf ( n440046 , n439377 );
buf ( n440047 , n438951 );
nand ( n440048 , n440046 , n440047 );
buf ( n440049 , n440048 );
buf ( n440050 , n440049 );
buf ( n440051 , n440049 );
not ( n440052 , n440051 );
buf ( n440053 , n440052 );
buf ( n440054 , n440053 );
buf ( n440055 , n439830 );
not ( n440056 , n440055 );
buf ( n440057 , n440032 );
not ( n440058 , n440057 );
or ( n440059 , n440056 , n440058 );
buf ( n440060 , n439373 );
not ( n440061 , n440060 );
buf ( n440062 , n440061 );
buf ( n440063 , n440062 );
nand ( n440064 , n440059 , n440063 );
buf ( n440065 , n440064 );
buf ( n440066 , n440065 );
and ( n440067 , n440066 , n440054 );
not ( n440068 , n440066 );
and ( n440069 , n440068 , n440050 );
nor ( n440070 , n440067 , n440069 );
buf ( n440071 , n440070 );
nand ( n440072 , n439303 , n439344 );
buf ( n440073 , n440072 );
buf ( n440074 , n440072 );
not ( n440075 , n440074 );
buf ( n440076 , n440075 );
buf ( n440077 , n440076 );
nor ( n440078 , n436350 , n437325 );
not ( n440079 , n440078 );
not ( n440080 , n439817 );
not ( n440081 , n439823 );
or ( n440082 , n440080 , n440081 );
buf ( n440083 , n439401 );
buf ( n440084 , n440083 );
not ( n440085 , n440084 );
buf ( n440086 , n440085 );
nand ( n440087 , n440082 , n440086 );
not ( n440088 , n440087 );
or ( n440089 , n440079 , n440088 );
buf ( n440090 , n439321 );
not ( n440091 , n440090 );
buf ( n440092 , n440091 );
nand ( n440093 , n440089 , n440092 );
buf ( n440094 , n440093 );
and ( n440095 , n440094 , n440077 );
not ( n440096 , n440094 );
and ( n440097 , n440096 , n440073 );
nor ( n440098 , n440095 , n440097 );
buf ( n440099 , n440098 );
buf ( n440100 , n437324 );
buf ( n440101 , n439320 );
nand ( n440102 , n440100 , n440101 );
buf ( n440103 , n440102 );
buf ( n440104 , n440103 );
buf ( n440105 , n440103 );
not ( n440106 , n440105 );
buf ( n440107 , n440106 );
buf ( n440108 , n440107 );
not ( n440109 , n436350 );
not ( n440110 , n440109 );
not ( n440111 , n440087 );
or ( n440112 , n440110 , n440111 );
buf ( n440113 , n439315 );
not ( n440114 , n440113 );
nand ( n440115 , n440112 , n440114 );
buf ( n440116 , n440115 );
and ( n440117 , n440116 , n440108 );
not ( n440118 , n440116 );
and ( n440119 , n440118 , n440104 );
nor ( n440120 , n440117 , n440119 );
buf ( n440121 , n440120 );
buf ( n440122 , n439314 );
buf ( n440123 , n440122 );
buf ( n440124 , n436340 );
nand ( n440125 , n440123 , n440124 );
buf ( n440126 , n440125 );
buf ( n440127 , n440126 );
buf ( n440128 , n440126 );
not ( n440129 , n440128 );
buf ( n440130 , n440129 );
buf ( n440131 , n440130 );
buf ( n440132 , n436349 );
not ( n440133 , n440132 );
buf ( n440134 , n440087 );
not ( n440135 , n440134 );
or ( n440136 , n440133 , n440135 );
buf ( n440137 , n439309 );
buf ( n440138 , n440137 );
buf ( n440139 , n440138 );
buf ( n440140 , n440139 );
nand ( n440141 , n440136 , n440140 );
buf ( n440142 , n440141 );
buf ( n440143 , n440142 );
and ( n440144 , n440143 , n440131 );
not ( n440145 , n440143 );
and ( n440146 , n440145 , n440127 );
nor ( n440147 , n440144 , n440146 );
buf ( n440148 , n440147 );
buf ( n440149 , n439474 );
not ( n440150 , n440149 );
buf ( n440151 , n439467 );
nand ( n440152 , n440150 , n440151 );
buf ( n440153 , n440152 );
buf ( n440154 , n440153 );
buf ( n440155 , n440153 );
not ( n440156 , n440155 );
buf ( n440157 , n440156 );
buf ( n440158 , n440157 );
buf ( n440159 , n393718 );
buf ( n440160 , n394596 );
buf ( n440161 , n440160 );
buf ( n440162 , n48184 );
buf ( n440163 , n440162 );
and ( n440164 , n440159 , n440161 , n440163 );
buf ( n440165 , n440164 );
not ( n440166 , n440165 );
buf ( n440167 , n399939 );
buf ( n440168 , n440167 );
buf ( n440169 , n440168 );
buf ( n440170 , n440169 );
not ( n440171 , n440170 );
buf ( n440172 , n433183 );
buf ( n440173 , n63019 );
buf ( n440174 , n405627 );
nand ( n440175 , n440172 , n440173 , n440174 );
buf ( n440176 , n439528 );
buf ( n440177 , n440176 );
buf ( n440178 , n440177 );
buf ( n440179 , n403536 );
and ( n440180 , n440178 , n440179 );
buf ( n440181 , n439515 );
nor ( n440182 , n440180 , n440181 );
buf ( n440183 , n410016 );
not ( n440184 , n440183 );
nand ( n440185 , n439500 , n439494 );
buf ( n440186 , n440185 );
not ( n440187 , n440186 );
or ( n440188 , n440184 , n440187 );
buf ( n440189 , n439498 );
buf ( n440190 , n440189 );
nand ( n440191 , n440188 , n440190 );
buf ( n440192 , n440191 );
nand ( n440193 , n440174 , n440192 );
nand ( n440194 , n440175 , n440182 , n440193 );
buf ( n440195 , n440194 );
not ( n440196 , n440195 );
or ( n440197 , n440171 , n440196 );
buf ( n440198 , n439446 );
buf ( n440199 , n440198 );
buf ( n440200 , n440199 );
buf ( n440201 , n440200 );
not ( n440202 , n440201 );
buf ( n440203 , n440202 );
buf ( n440204 , n440203 );
nand ( n440205 , n440197 , n440204 );
buf ( n440206 , n440205 );
not ( n440207 , n440206 );
or ( n440208 , n440166 , n440207 );
nand ( n440209 , n439463 , n439464 );
nand ( n440210 , n440208 , n440209 );
buf ( n440211 , n440210 );
and ( n440212 , n440211 , n440158 );
not ( n440213 , n440211 );
and ( n440214 , n440213 , n440154 );
nor ( n440215 , n440212 , n440214 );
buf ( n440216 , n440215 );
buf ( n440217 , n439452 );
not ( n440218 , n440217 );
buf ( n440219 , n393718 );
buf ( n440220 , n440219 );
nand ( n440221 , n440218 , n440220 );
buf ( n440222 , n440221 );
buf ( n440223 , n440222 );
buf ( n440224 , n440222 );
not ( n440225 , n440224 );
buf ( n440226 , n440225 );
buf ( n440227 , n440226 );
not ( n440228 , n440160 );
buf ( n440229 , n440169 );
not ( n440230 , n440229 );
buf ( n440231 , n440162 );
not ( n440232 , n440231 );
buf ( n440233 , n440232 );
buf ( n440234 , n440233 );
nor ( n440235 , n440230 , n440234 );
buf ( n440236 , n440235 );
buf ( n440237 , n440236 );
not ( n440238 , n440237 );
nand ( n440239 , n440175 , n440193 );
buf ( n440240 , n440239 );
not ( n440241 , n440240 );
or ( n440242 , n440238 , n440241 );
buf ( n440243 , n440203 );
not ( n440244 , n440243 );
buf ( n440245 , n440233 );
not ( n440246 , n440245 );
and ( n440247 , n440244 , n440246 );
buf ( n440248 , n440182 );
not ( n440249 , n440248 );
buf ( n440250 , n440249 );
buf ( n440251 , n440250 );
buf ( n440252 , n440236 );
and ( n440253 , n440251 , n440252 );
nor ( n440254 , n440247 , n440253 );
buf ( n440255 , n440254 );
buf ( n440256 , n440255 );
nand ( n440257 , n440242 , n440256 );
buf ( n440258 , n440257 );
not ( n440259 , n440258 );
or ( n440260 , n440228 , n440259 );
not ( n440261 , n439462 );
buf ( n440262 , n439457 );
buf ( n440263 , n440262 );
nor ( n440264 , n440261 , n440263 );
nand ( n440265 , n440260 , n440264 );
buf ( n440266 , n440265 );
and ( n440267 , n440266 , n440227 );
not ( n440268 , n440266 );
and ( n440269 , n440268 , n440223 );
nor ( n440270 , n440267 , n440269 );
buf ( n440271 , n440270 );
buf ( n440272 , n440262 );
not ( n440273 , n440272 );
buf ( n440274 , n440160 );
nand ( n440275 , n440273 , n440274 );
buf ( n440276 , n440275 );
buf ( n440277 , n440276 );
not ( n440278 , n440277 );
buf ( n440279 , n440278 );
buf ( n440280 , n440279 );
buf ( n440281 , n440276 );
nor ( n440282 , n395622 , n47154 );
nor ( n440283 , n440258 , n440282 );
buf ( n440284 , n440283 );
and ( n440285 , n440284 , n440281 );
not ( n440286 , n440284 );
and ( n440287 , n440286 , n440280 );
nor ( n440288 , n440285 , n440287 );
buf ( n440289 , n440288 );
buf ( n440290 , n439385 );
not ( n440291 , n439388 );
buf ( n440292 , n440291 );
nand ( n440293 , n440290 , n440292 );
buf ( n440294 , n440293 );
buf ( n440295 , n440294 );
buf ( n440296 , n440294 );
not ( n440297 , n440296 );
buf ( n440298 , n440297 );
buf ( n440299 , n440298 );
buf ( n440300 , n433746 );
not ( n440301 , n440300 );
buf ( n440302 , n439823 );
not ( n440303 , n440302 );
or ( n440304 , n440301 , n440303 );
buf ( n440305 , n439386 );
buf ( n440306 , n440305 );
nand ( n440307 , n440304 , n440306 );
buf ( n440308 , n440307 );
buf ( n440309 , n440308 );
and ( n440310 , n440309 , n440299 );
not ( n440311 , n440309 );
and ( n440312 , n440311 , n440295 );
nor ( n440313 , n440310 , n440312 );
buf ( n440314 , n440313 );
buf ( n440315 , n439518 );
buf ( n440316 , n439527 );
nand ( n440317 , n440315 , n440316 );
buf ( n440318 , n440317 );
buf ( n440319 , n440317 );
not ( n440320 , n440319 );
buf ( n440321 , n440320 );
buf ( n440322 , n440321 );
nand ( n440323 , n414379 , n414384 );
not ( n440324 , n440323 );
nand ( n440325 , n409970 , n410016 , n409999 );
nor ( n440326 , n440324 , n440325 );
not ( n440327 , n440326 );
not ( n440328 , n67630 );
not ( n440329 , n67620 );
or ( n440330 , n440328 , n440329 );
nand ( n440331 , n433178 , n433171 );
nand ( n440332 , n440330 , n440331 );
not ( n440333 , n440332 );
or ( n440334 , n440327 , n440333 );
not ( n440335 , n433182 );
not ( n440336 , n440325 );
and ( n440337 , n440335 , n440336 );
nor ( n440338 , n440337 , n440192 );
nand ( n440339 , n440334 , n440338 );
buf ( n440340 , n440339 );
not ( n440341 , n440340 );
buf ( n440342 , n440341 );
buf ( n440343 , n440342 );
buf ( n440344 , n405619 );
not ( n440345 , n440344 );
buf ( n440346 , n440345 );
or ( n440347 , n440343 , n440346 );
buf ( n440348 , n439516 );
not ( n440349 , n440348 );
buf ( n440350 , n440349 );
buf ( n440351 , n440350 );
nand ( n440352 , n440347 , n440351 );
buf ( n440353 , n440352 );
buf ( n440354 , n440353 );
and ( n440355 , n440354 , n440322 );
not ( n440356 , n440354 );
and ( n440357 , n440356 , n440318 );
nor ( n440358 , n440355 , n440357 );
buf ( n440359 , n440358 );
buf ( n440360 , n56293 );
nand ( n440361 , n439506 , n439510 );
buf ( n440362 , n440361 );
nand ( n440363 , n440360 , n440362 );
buf ( n440364 , n440363 );
buf ( n440365 , n440364 );
buf ( n440366 , n440364 );
not ( n440367 , n440366 );
buf ( n440368 , n440367 );
buf ( n440369 , n440368 );
not ( n440370 , n58470 );
not ( n440371 , n440339 );
or ( n440372 , n440370 , n440371 );
buf ( n440373 , n440178 );
not ( n440374 , n440373 );
buf ( n440375 , n440374 );
nand ( n440376 , n440372 , n440375 );
buf ( n440377 , n440376 );
and ( n440378 , n440377 , n440369 );
not ( n440379 , n440377 );
and ( n440380 , n440379 , n440365 );
nor ( n440381 , n440378 , n440380 );
buf ( n440382 , n440381 );
nand ( n440383 , n439443 , n439439 );
buf ( n440384 , n440383 );
buf ( n440385 , n440383 );
not ( n440386 , n440385 );
buf ( n440387 , n440386 );
buf ( n440388 , n440387 );
buf ( n440389 , n52572 );
buf ( n440390 , n440389 );
buf ( n440391 , n440390 );
buf ( n440392 , n440391 );
buf ( n440393 , n52613 );
buf ( n440394 , n440393 );
and ( n440395 , n440392 , n440394 );
buf ( n440396 , n440395 );
buf ( n440397 , n440396 );
not ( n440398 , n440397 );
buf ( n440399 , n440239 );
not ( n440400 , n440399 );
or ( n440401 , n440398 , n440400 );
and ( n440402 , n440396 , n440250 );
not ( n440403 , n440393 );
buf ( n440404 , n439425 );
buf ( n440405 , n440404 );
nand ( n440406 , n439429 , n439427 );
buf ( n440407 , n440406 );
nand ( n440408 , n440405 , n440407 );
buf ( n440409 , n440408 );
not ( n440410 , n440409 );
or ( n440411 , n440403 , n440410 );
nand ( n440412 , n440411 , n439436 );
nor ( n440413 , n440402 , n440412 );
buf ( n440414 , n440413 );
nand ( n440415 , n440401 , n440414 );
buf ( n440416 , n440415 );
buf ( n440417 , n440416 );
and ( n440418 , n440417 , n440388 );
not ( n440419 , n440417 );
and ( n440420 , n440419 , n440384 );
nor ( n440421 , n440418 , n440420 );
buf ( n440422 , n440421 );
buf ( n440423 , n51961 );
nand ( n440424 , n440406 , n440423 );
buf ( n440425 , n440424 );
buf ( n440426 , n440424 );
not ( n440427 , n440426 );
buf ( n440428 , n440427 );
buf ( n440429 , n440428 );
buf ( n440430 , n52570 );
buf ( n440431 , n440430 );
buf ( n440432 , n440431 );
not ( n440433 , n440432 );
buf ( n440434 , n440194 );
not ( n440435 , n440434 );
or ( n440436 , n440433 , n440435 );
buf ( n440437 , n439424 );
buf ( n440438 , n440437 );
not ( n440439 , n440438 );
nand ( n440440 , n440436 , n440439 );
buf ( n440441 , n440440 );
and ( n440442 , n440441 , n440429 );
not ( n440443 , n440441 );
and ( n440444 , n440443 , n440425 );
nor ( n440445 , n440442 , n440444 );
buf ( n440446 , n440445 );
buf ( n440447 , n39148 );
buf ( n440448 , n439866 );
and ( n440449 , n440447 , n440448 );
buf ( n440450 , n440449 );
buf ( n440451 , n440450 );
buf ( n440452 , n439862 );
not ( n440453 , n440452 );
buf ( n440454 , n440453 );
buf ( n440455 , n440454 );
buf ( n440456 , n440450 );
buf ( n440457 , n440454 );
not ( n440458 , n440451 );
not ( n440459 , n440455 );
or ( n440460 , n440458 , n440459 );
or ( n440461 , n440456 , n440457 );
nand ( n440462 , n440460 , n440461 );
buf ( n440463 , n440462 );
buf ( n440464 , n437773 );
buf ( n440465 , n440464 );
not ( n440466 , n439353 );
buf ( n440467 , n440466 );
nand ( n440468 , n440465 , n440467 );
buf ( n440469 , n440468 );
buf ( n440470 , n440469 );
buf ( n440471 , n440032 );
buf ( n440472 , n440471 );
buf ( n440473 , n440469 );
buf ( n440474 , n440471 );
not ( n440475 , n440470 );
not ( n440476 , n440472 );
or ( n440477 , n440475 , n440476 );
or ( n440478 , n440473 , n440474 );
nand ( n440479 , n440477 , n440478 );
buf ( n440480 , n440479 );
buf ( n440481 , n440139 );
buf ( n440482 , n436349 );
nand ( n440483 , n440481 , n440482 );
buf ( n440484 , n440483 );
buf ( n440485 , n440484 );
buf ( n440486 , n440484 );
not ( n440487 , n440486 );
buf ( n440488 , n440487 );
buf ( n440489 , n440488 );
buf ( n440490 , n440087 );
and ( n440491 , n440490 , n440489 );
not ( n440492 , n440490 );
and ( n440493 , n440492 , n440485 );
nor ( n440494 , n440491 , n440493 );
buf ( n440495 , n440494 );
buf ( n440496 , n439436 );
buf ( n440497 , n440393 );
nand ( n440498 , n440496 , n440497 );
buf ( n440499 , n440498 );
buf ( n440500 , n440499 );
buf ( n440501 , n440499 );
not ( n440502 , n440501 );
buf ( n440503 , n440502 );
buf ( n440504 , n440503 );
buf ( n440505 , n440391 );
not ( n440506 , n440505 );
buf ( n440507 , n440434 );
not ( n440508 , n440507 );
or ( n440509 , n440506 , n440508 );
buf ( n440510 , n440409 );
not ( n440511 , n440510 );
buf ( n440512 , n440511 );
buf ( n440513 , n440512 );
nand ( n440514 , n440509 , n440513 );
buf ( n440515 , n440514 );
buf ( n440516 , n440515 );
and ( n440517 , n440516 , n440504 );
not ( n440518 , n440516 );
and ( n440519 , n440518 , n440500 );
nor ( n440520 , n440517 , n440519 );
buf ( n440521 , n440520 );
not ( n440522 , n440282 );
nand ( n440523 , n440522 , n440162 );
buf ( n440524 , n440523 );
buf ( n440525 , n440523 );
not ( n440526 , n440525 );
buf ( n440527 , n440526 );
buf ( n440528 , n440527 );
buf ( n440529 , n440206 );
and ( n440530 , n440529 , n440528 );
not ( n440531 , n440529 );
and ( n440532 , n440531 , n440524 );
nor ( n440533 , n440530 , n440532 );
buf ( n440534 , n440533 );
buf ( n440535 , n65799 );
buf ( n440536 , n414370 );
nand ( n440537 , n440535 , n440536 );
buf ( n440538 , n440537 );
buf ( n440539 , n440538 );
buf ( n440540 , n440538 );
not ( n440541 , n440540 );
buf ( n440542 , n440541 );
buf ( n440543 , n440542 );
buf ( n440544 , n67618 );
not ( n440545 , n433175 );
and ( n440546 , n440544 , n440545 );
buf ( n440547 , n67622 );
not ( n440548 , n417508 );
not ( n440549 , n433147 );
or ( n440550 , n440548 , n440549 );
nand ( n440551 , n440550 , n433170 );
nand ( n440552 , n440546 , n440547 , n440551 );
not ( n440553 , n67617 );
not ( n440554 , n440544 );
or ( n440555 , n440553 , n440554 );
buf ( n440556 , n412499 );
nand ( n440557 , n440556 , n412404 );
nand ( n440558 , n440555 , n440557 );
and ( n440559 , n440558 , n440547 );
nand ( n440560 , n65757 , n412587 );
not ( n440561 , n440560 );
nor ( n440562 , n440559 , n440561 );
nand ( n440563 , n440552 , n440562 );
buf ( n440564 , n440563 );
and ( n440565 , n440564 , n440543 );
not ( n440566 , n440564 );
and ( n440567 , n440566 , n440539 );
nor ( n440568 , n440565 , n440567 );
buf ( n440569 , n440568 );
buf ( n440570 , n440350 );
buf ( n440571 , n440344 );
nand ( n440572 , n440570 , n440571 );
buf ( n440573 , n440572 );
buf ( n440574 , n440573 );
not ( n440575 , n440574 );
buf ( n440576 , n440575 );
buf ( n440577 , n440576 );
buf ( n440578 , n440573 );
buf ( n440579 , n440342 );
and ( n440580 , n440579 , n440578 );
not ( n440581 , n440579 );
and ( n440582 , n440581 , n440577 );
nor ( n440583 , n440580 , n440582 );
buf ( n440584 , n440583 );
not ( n440585 , n440438 );
nand ( n440586 , n440585 , n440432 );
buf ( n440587 , n440586 );
buf ( n440588 , n440434 );
buf ( n440589 , n440586 );
buf ( n440590 , n440434 );
not ( n440591 , n440587 );
not ( n440592 , n440588 );
or ( n440593 , n440591 , n440592 );
or ( n440594 , n440589 , n440590 );
nand ( n440595 , n440593 , n440594 );
buf ( n440596 , n440595 );
buf ( n440597 , n409999 );
not ( n440598 , n440597 );
buf ( n440599 , n440598 );
not ( n440600 , n440599 );
nand ( n440601 , n440600 , n439500 );
buf ( n440602 , n440601 );
buf ( n440603 , n440601 );
not ( n440604 , n440603 );
buf ( n440605 , n440604 );
buf ( n440606 , n440605 );
buf ( n440607 , n409970 );
not ( n440608 , n440607 );
buf ( n440609 , n440172 );
not ( n440610 , n440609 );
or ( n440611 , n440608 , n440610 );
nand ( n440612 , n408541 , n60627 );
buf ( n440613 , n440612 );
buf ( n440614 , n439493 );
nand ( n440615 , n440613 , n440614 );
buf ( n440616 , n440615 );
nand ( n440617 , n440611 , n440616 );
buf ( n440618 , n440617 );
and ( n440619 , n440618 , n440606 );
not ( n440620 , n440618 );
and ( n440621 , n440620 , n440602 );
nor ( n440622 , n440619 , n440621 );
buf ( n440623 , n440622 );
buf ( n440624 , n440189 );
buf ( n440625 , n439484 );
nand ( n440626 , n440624 , n440625 );
buf ( n440627 , n440626 );
buf ( n440628 , n440627 );
buf ( n440629 , n440627 );
not ( n440630 , n440629 );
buf ( n440631 , n440630 );
buf ( n440632 , n440631 );
buf ( n440633 , n440607 );
not ( n440634 , n440633 );
buf ( n440635 , n440599 );
nor ( n440636 , n440634 , n440635 );
buf ( n440637 , n440636 );
not ( n440638 , n440637 );
not ( n440639 , n440609 );
or ( n440640 , n440638 , n440639 );
buf ( n440641 , n440185 );
not ( n440642 , n440641 );
buf ( n440643 , n440642 );
nand ( n440644 , n440640 , n440643 );
buf ( n440645 , n440644 );
and ( n440646 , n440645 , n440632 );
not ( n440647 , n440645 );
and ( n440648 , n440647 , n440628 );
nor ( n440649 , n440646 , n440648 );
buf ( n440650 , n440649 );
buf ( n440651 , n439823 );
buf ( n440652 , n440651 );
buf ( n440653 , n440652 );
buf ( n440654 , n433169 );
not ( n440655 , n440654 );
buf ( n440656 , n414401 );
buf ( n440657 , n440656 );
buf ( n440658 , n415763 );
nand ( n440659 , n440657 , n440658 );
buf ( n440660 , n440659 );
buf ( n440661 , n440660 );
nand ( n440662 , n440655 , n440661 );
buf ( n440663 , n440662 );
buf ( n440664 , n440663 );
buf ( n440665 , n440663 );
not ( n440666 , n440665 );
buf ( n440667 , n440666 );
buf ( n440668 , n440667 );
buf ( n440669 , n417505 );
buf ( n440670 , n432831 );
buf ( n440671 , n440670 );
buf ( n440672 , n432849 );
buf ( n440673 , n432854 );
nand ( n440674 , n440671 , n440672 , n440673 );
buf ( n440675 , n440674 );
buf ( n440676 , n440675 );
buf ( n440677 , n433015 );
buf ( n440678 , n433102 );
nand ( n440679 , n440676 , n440677 , n440678 );
buf ( n440680 , n440679 );
buf ( n440681 , n440680 );
buf ( n440682 , n433144 );
buf ( n440683 , n440682 );
buf ( n440684 , n440683 );
nand ( n440685 , n440681 , n440684 );
buf ( n440686 , n440685 );
buf ( n440687 , n440686 );
nand ( n440688 , n440669 , n440687 );
buf ( n440689 , n440688 );
buf ( n440690 , n415844 );
buf ( n440691 , n440690 );
buf ( n440692 , n440691 );
buf ( n440693 , n440692 );
not ( n440694 , n440693 );
buf ( n440695 , n440694 );
or ( n440696 , n440689 , n440695 );
not ( n440697 , n433167 );
nand ( n440698 , n440696 , n440697 );
buf ( n440699 , n440698 );
and ( n440700 , n440699 , n440668 );
not ( n440701 , n440699 );
and ( n440702 , n440701 , n440664 );
nor ( n440703 , n440700 , n440702 );
buf ( n440704 , n440703 );
buf ( n440705 , n433166 );
buf ( n440706 , n440692 );
nand ( n440707 , n440705 , n440706 );
buf ( n440708 , n440707 );
buf ( n440709 , n440708 );
buf ( n440710 , n440708 );
not ( n440711 , n440710 );
buf ( n440712 , n440711 );
buf ( n440713 , n440712 );
buf ( n440714 , n440689 );
buf ( n440715 , n433154 );
buf ( n440716 , n440715 );
not ( n440717 , n440716 );
buf ( n440718 , n440717 );
buf ( n440719 , n440718 );
nand ( n440720 , n440714 , n440719 );
buf ( n440721 , n440720 );
buf ( n440722 , n440721 );
and ( n440723 , n440722 , n440713 );
not ( n440724 , n440722 );
and ( n440725 , n440724 , n440709 );
nor ( n440726 , n440723 , n440725 );
buf ( n440727 , n440726 );
buf ( n440728 , n433143 );
buf ( n440729 , n433131 );
nand ( n440730 , n440728 , n440729 );
buf ( n440731 , n440730 );
buf ( n440732 , n440731 );
buf ( n440733 , n440731 );
not ( n440734 , n440733 );
buf ( n440735 , n440734 );
buf ( n440736 , n440735 );
buf ( n440737 , n432988 );
not ( n440738 , n440737 );
buf ( n440739 , n433125 );
not ( n440740 , n440739 );
buf ( n440741 , n433102 );
buf ( n440742 , n440670 );
buf ( n440743 , n432849 );
buf ( n440744 , n432854 );
nand ( n440745 , n440742 , n440743 , n440744 );
buf ( n440746 , n440745 );
buf ( n440747 , n440746 );
nand ( n440748 , n440741 , n440747 );
buf ( n440749 , n440748 );
buf ( n440750 , n440749 );
nand ( n440751 , n440740 , n440750 );
buf ( n440752 , n440751 );
buf ( n440753 , n440752 );
not ( n440754 , n440753 );
or ( n440755 , n440738 , n440754 );
buf ( n440756 , n432918 );
buf ( n440757 , n432982 );
nand ( n440758 , n440756 , n440757 );
buf ( n440759 , n440758 );
buf ( n440760 , n440759 );
nand ( n440761 , n440755 , n440760 );
buf ( n440762 , n440761 );
buf ( n440763 , n440762 );
and ( n440764 , n440763 , n440736 );
not ( n440765 , n440763 );
and ( n440766 , n440765 , n440732 );
nor ( n440767 , n440764 , n440766 );
buf ( n440768 , n440767 );
buf ( n440769 , n440759 );
buf ( n440770 , n432988 );
nand ( n440771 , n440769 , n440770 );
buf ( n440772 , n440771 );
buf ( n440773 , n440772 );
buf ( n440774 , n440772 );
not ( n440775 , n440774 );
buf ( n440776 , n440775 );
buf ( n440777 , n440776 );
buf ( n440778 , n440752 );
and ( n440779 , n440778 , n440777 );
not ( n440780 , n440778 );
and ( n440781 , n440780 , n440773 );
nor ( n440782 , n440779 , n440781 );
buf ( n440783 , n440782 );
buf ( n440784 , n433124 );
buf ( n440785 , n433099 );
nand ( n440786 , n440784 , n440785 );
buf ( n440787 , n440786 );
buf ( n440788 , n440787 );
buf ( n440789 , n440787 );
not ( n440790 , n440789 );
buf ( n440791 , n440790 );
buf ( n440792 , n440791 );
buf ( n440793 , n433075 );
not ( n440794 , n440793 );
buf ( n440795 , n440746 );
not ( n440796 , n440795 );
or ( n440797 , n440794 , n440796 );
buf ( n440798 , n433112 );
not ( n440799 , n440798 );
buf ( n440800 , n440799 );
buf ( n440801 , n440800 );
nand ( n440802 , n440797 , n440801 );
buf ( n440803 , n440802 );
buf ( n440804 , n440803 );
and ( n440805 , n440804 , n440792 );
not ( n440806 , n440804 );
and ( n440807 , n440806 , n440788 );
nor ( n440808 , n440805 , n440807 );
buf ( n440809 , n440808 );
buf ( n440810 , n432844 );
buf ( n440811 , n432806 );
nand ( n440812 , n440810 , n440811 );
buf ( n440813 , n440812 );
buf ( n440814 , n440813 );
buf ( n440815 , n440813 );
not ( n440816 , n440815 );
buf ( n440817 , n440816 );
buf ( n440818 , n440817 );
not ( n440819 , n432825 );
buf ( n440820 , n440819 );
not ( n440821 , n440820 );
not ( n440822 , n430929 );
not ( n440823 , n432167 );
or ( n440824 , n440822 , n440823 );
nand ( n440825 , n440824 , n432190 );
buf ( n440826 , n440825 );
not ( n440827 , n440826 );
or ( n440828 , n440821 , n440827 );
buf ( n440829 , n432837 );
not ( n440830 , n440829 );
buf ( n440831 , n440830 );
buf ( n440832 , n440831 );
nand ( n440833 , n440828 , n440832 );
buf ( n440834 , n440833 );
buf ( n440835 , n440834 );
and ( n440836 , n440835 , n440818 );
not ( n440837 , n440835 );
and ( n440838 , n440837 , n440814 );
nor ( n440839 , n440836 , n440838 );
buf ( n440840 , n440839 );
buf ( n440841 , n432178 );
buf ( n440842 , n431857 );
nand ( n440843 , n440841 , n440842 );
buf ( n440844 , n440843 );
buf ( n440845 , n440844 );
buf ( n440846 , n440844 );
not ( n440847 , n440846 );
buf ( n440848 , n440847 );
buf ( n440849 , n440848 );
buf ( n440850 , n431874 );
not ( n440851 , n440850 );
buf ( n440852 , n440851 );
not ( n440853 , n440852 );
buf ( n440854 , n430929 );
buf ( n440855 , n440854 );
buf ( n440856 , n440855 );
not ( n440857 , n440856 );
or ( n440858 , n440853 , n440857 );
not ( n440859 , n86947 );
nand ( n440860 , n440858 , n440859 );
buf ( n440861 , n440860 );
and ( n440862 , n440861 , n440849 );
not ( n440863 , n440861 );
and ( n440864 , n440863 , n440845 );
nor ( n440865 , n440862 , n440864 );
buf ( n440866 , n440865 );
buf ( n440867 , n440856 );
buf ( n440868 , n431857 );
buf ( n440869 , n440852 );
buf ( n440870 , n86954 );
and ( n440871 , n440867 , n440868 , n440869 );
nor ( n440872 , n440871 , n440870 );
buf ( n440873 , n440872 );
buf ( n440874 , n85470 );
buf ( n440875 , n80450 );
nand ( n440876 , n440874 , n440875 );
buf ( n440877 , n440876 );
buf ( n440878 , n440877 );
buf ( n440879 , n440877 );
not ( n440880 , n440879 );
buf ( n440881 , n440880 );
buf ( n440882 , n440881 );
buf ( n440883 , n425730 );
buf ( n440884 , n440883 );
buf ( n440885 , n440884 );
buf ( n440886 , n440885 );
not ( n440887 , n440886 );
buf ( n440888 , n426551 );
not ( n440889 , n440888 );
buf ( n440890 , n80454 );
not ( n440891 , n440890 );
buf ( n440892 , n440891 );
buf ( n440893 , n440892 );
not ( n440894 , n440893 );
buf ( n440895 , n85468 );
not ( n440896 , n440895 );
or ( n440897 , n440894 , n440896 );
buf ( n440898 , n80355 );
nand ( n440899 , n440897 , n440898 );
buf ( n440900 , n440899 );
buf ( n440901 , n440900 );
not ( n440902 , n440901 );
or ( n440903 , n440889 , n440902 );
buf ( n440904 , n425818 );
nand ( n440905 , n440903 , n440904 );
buf ( n440906 , n440905 );
buf ( n440907 , n440906 );
not ( n440908 , n440907 );
or ( n440909 , n440887 , n440908 );
buf ( n440910 , n426569 );
nand ( n440911 , n440909 , n440910 );
buf ( n440912 , n440911 );
buf ( n440913 , n440912 );
and ( n440914 , n440913 , n440882 );
not ( n440915 , n440913 );
and ( n440916 , n440915 , n440878 );
nor ( n440917 , n440914 , n440916 );
buf ( n440918 , n440917 );
buf ( n440919 , n426569 );
buf ( n440920 , n440885 );
nand ( n440921 , n440919 , n440920 );
buf ( n440922 , n440921 );
buf ( n440923 , n440922 );
buf ( n440924 , n440922 );
not ( n440925 , n440924 );
buf ( n440926 , n440925 );
buf ( n440927 , n440926 );
buf ( n440928 , n440906 );
and ( n440929 , n440928 , n440927 );
not ( n440930 , n440928 );
and ( n440931 , n440930 , n440923 );
nor ( n440932 , n440929 , n440931 );
buf ( n440933 , n440932 );
buf ( n440934 , n85520 );
buf ( n440935 , n85550 );
not ( n440936 , n440935 );
buf ( n440937 , n440936 );
buf ( n440938 , n440937 );
nand ( n440939 , n440934 , n440938 );
buf ( n440940 , n440939 );
buf ( n440941 , n425818 );
buf ( n440942 , n426551 );
nand ( n440943 , n440941 , n440942 );
buf ( n440944 , n440943 );
buf ( n440945 , n440944 );
buf ( n440946 , n440944 );
not ( n440947 , n440946 );
buf ( n440948 , n440947 );
buf ( n440949 , n440948 );
buf ( n440950 , n440900 );
and ( n440951 , n440950 , n440949 );
not ( n440952 , n440950 );
and ( n440953 , n440952 , n440945 );
nor ( n440954 , n440951 , n440953 );
buf ( n440955 , n440954 );
xor ( n440956 , n427610 , n427614 );
xor ( n440957 , n440956 , n430818 );
buf ( n440958 , n440957 );
buf ( n440959 , n432164 );
buf ( n440960 , n432186 );
nand ( n440961 , n440959 , n440960 );
buf ( n440962 , n440961 );
buf ( n440963 , n440831 );
buf ( n440964 , n440819 );
nand ( n440965 , n440963 , n440964 );
buf ( n440966 , n440965 );
buf ( n440967 , n440966 );
not ( n440968 , n440967 );
buf ( n440969 , n440968 );
xor ( n440970 , n427928 , n427932 );
xor ( n440971 , n440970 , n430813 );
buf ( n440972 , n440971 );
buf ( n440973 , n440800 );
buf ( n440974 , n433075 );
nand ( n440975 , n440973 , n440974 );
buf ( n440976 , n440975 );
buf ( n440977 , n440976 );
not ( n440978 , n440977 );
buf ( n440979 , n440978 );
buf ( n440980 , n440718 );
buf ( n440981 , n417505 );
nand ( n440982 , n440980 , n440981 );
buf ( n440983 , n440982 );
xor ( n440984 , n428051 , n428055 );
xor ( n440985 , n440984 , n430808 );
buf ( n440986 , n440985 );
buf ( n440987 , n440544 );
buf ( n440988 , n440557 );
nand ( n440989 , n440987 , n440988 );
buf ( n440990 , n440989 );
buf ( n440991 , n440990 );
not ( n440992 , n440991 );
buf ( n440993 , n440992 );
nand ( n440994 , n440560 , n440547 );
buf ( n440995 , n440994 );
not ( n440996 , n440995 );
buf ( n440997 , n440996 );
buf ( n440998 , n440892 );
buf ( n440999 , n80355 );
nand ( n441000 , n440998 , n440999 );
buf ( n441001 , n441000 );
xor ( n441002 , n428480 , n428484 );
xor ( n441003 , n441002 , n430803 );
buf ( n441004 , n441003 );
not ( n441005 , n440324 );
nand ( n441006 , n441005 , n433182 );
buf ( n441007 , n441006 );
not ( n441008 , n441007 );
buf ( n441009 , n441008 );
buf ( n441010 , n428928 );
buf ( n441011 , n430801 );
nand ( n441012 , n441010 , n441011 );
buf ( n441013 , n441012 );
buf ( n441014 , n430786 );
buf ( n441015 , n429088 );
not ( n441016 , n441014 );
nor ( n441017 , n441016 , n441015 );
buf ( n441018 , n441017 );
buf ( n441019 , n430754 );
buf ( n441020 , n430747 );
nand ( n441021 , n441019 , n441020 );
buf ( n441022 , n441021 );
buf ( n441023 , n441022 );
buf ( n441024 , n85328 );
buf ( n441025 , n85328 );
buf ( n441026 , n441022 );
not ( n441027 , n441023 );
not ( n441028 , n441024 );
or ( n441029 , n441027 , n441028 );
or ( n441030 , n441025 , n441026 );
nand ( n441031 , n441029 , n441030 );
buf ( n441032 , n441031 );
buf ( n441033 , n429674 );
buf ( n441034 , n430693 );
nand ( n441035 , n441033 , n441034 );
buf ( n441036 , n441035 );
buf ( n441037 , n430662 );
buf ( n441038 , n430665 );
buf ( n441039 , n430677 );
not ( n441040 , n441039 );
buf ( n441041 , n430683 );
nand ( n441042 , n441040 , n441041 );
buf ( n441043 , n441042 );
buf ( n441044 , n441043 );
and ( n441045 , n441044 , n441038 );
not ( n441046 , n441044 );
and ( n441047 , n441046 , n441037 );
nor ( n441048 , n441045 , n441047 );
buf ( n441049 , n441048 );
xor ( n441050 , n429969 , n430643 );
xor ( n441051 , n441050 , n430658 );
buf ( n441052 , n441051 );
buf ( n441053 , n430629 );
buf ( n441054 , n430641 );
nand ( n441055 , n441053 , n441054 );
buf ( n441056 , n441055 );
buf ( n441057 , n441056 );
buf ( n441058 , n430590 );
buf ( n441059 , n430590 );
buf ( n441060 , n441056 );
not ( n441061 , n441057 );
not ( n441062 , n441058 );
or ( n441063 , n441061 , n441062 );
or ( n441064 , n441059 , n441060 );
nand ( n441065 , n441063 , n441064 );
buf ( n441066 , n441065 );
buf ( n441067 , n440305 );
buf ( n441068 , n433746 );
and ( n441069 , n441067 , n441068 );
buf ( n441070 , n441069 );
buf ( n441071 , n430265 );
buf ( n441072 , n430542 );
nand ( n441073 , n441071 , n441072 );
buf ( n441074 , n441073 );
buf ( n441075 , n441074 );
buf ( n441076 , n85131 );
buf ( n441077 , n85131 );
buf ( n441078 , n441074 );
not ( n441079 , n441075 );
not ( n441080 , n441076 );
or ( n441081 , n441079 , n441080 );
or ( n441082 , n441077 , n441078 );
nand ( n441083 , n441081 , n441082 );
buf ( n441084 , n441083 );
buf ( n441085 , n435309 );
not ( n441086 , n441085 );
buf ( n441087 , n439395 );
nand ( n441088 , n441086 , n441087 );
buf ( n441089 , n441088 );
buf ( n441090 , n441089 );
not ( n441091 , n441090 );
buf ( n441092 , n441091 );
buf ( n441093 , n430536 );
buf ( n441094 , n430530 );
nand ( n441095 , n441093 , n441094 );
buf ( n441096 , n441095 );
buf ( n441097 , n441096 );
buf ( n441098 , n430509 );
buf ( n441099 , n430509 );
buf ( n441100 , n441096 );
not ( n441101 , n441097 );
not ( n441102 , n441098 );
or ( n441103 , n441101 , n441102 );
or ( n441104 , n441099 , n441100 );
nand ( n441105 , n441103 , n441104 );
buf ( n441106 , n441105 );
xor ( n441107 , n430454 , n430498 );
xor ( n441108 , n441107 , n430506 );
buf ( n441109 , n441108 );
xor ( n441110 , C0 , n430496 );
buf ( n441111 , n441110 );
xor ( n441112 , C0 , n430492 );
buf ( n441113 , n441112 );
buf ( n441114 , n430487 );
not ( n441115 , n441114 );
buf ( n441116 , n430488 );
nand ( n441117 , n441115 , n441116 );
buf ( n441118 , n441117 );
buf ( n441119 , n430479 );
buf ( n441120 , n441118 );
or ( n441121 , n441119 , n441120 );
nand ( n441122 , C1 , n441121 );
buf ( n441123 , n441122 );
xor ( n441124 , n430458 , n430476 );
xor ( n441125 , n441124 , n430478 );
buf ( n441126 , n441125 );
buf ( n441127 , n36166 );
buf ( n441128 , n439660 );
nand ( n441129 , n441127 , n441128 );
buf ( n441130 , n441129 );
buf ( n441131 , n441130 );
not ( n441132 , n441131 );
buf ( n441133 , n441132 );
xor ( n441134 , n430462 , n430472 );
xor ( n441135 , n441134 , n430474 );
buf ( n441136 , n441135 );
xor ( n441137 , n383207 , n383227 );
and ( n441138 , n441137 , n383285 );
and ( n441139 , n383207 , n383227 );
or ( n441140 , n441138 , n441139 );
buf ( n441141 , n441140 );
buf ( n441142 , n383206 );
not ( n441143 , n441142 );
buf ( n441144 , n383182 );
buf ( n441145 , n383200 );
nand ( n441146 , n441144 , n441145 );
buf ( n441147 , n441146 );
buf ( n441148 , n441147 );
not ( n441149 , n441148 );
buf ( n441150 , n383196 );
nor ( n441151 , n441149 , n441150 );
buf ( n441152 , n441151 );
buf ( n441153 , n382857 );
buf ( n441154 , n382538 );
and ( n441155 , n441153 , n441154 );
not ( n441156 , n441153 );
buf ( n441157 , n382551 );
and ( n441158 , n441156 , n441157 );
nor ( n441159 , n441155 , n441158 );
buf ( n441160 , n441159 );
buf ( n441161 , n441160 );
not ( n441162 , n441161 );
buf ( n441163 , n382950 );
nand ( n441164 , n441162 , n441163 );
buf ( n441165 , n441164 );
buf ( n441166 , n441165 );
nand ( n441167 , C1 , n441166 );
buf ( n441168 , n441167 );
buf ( n441169 , n441168 );
buf ( n441170 , n441152 );
or ( n441171 , n441169 , n441170 );
nand ( n441172 , C1 , n441171 );
buf ( n441173 , n441172 );
buf ( n441174 , n441173 );
not ( n441175 , n441174 );
or ( n441176 , n441143 , n441175 );
buf ( n441177 , n441173 );
buf ( n441178 , n383206 );
or ( n441179 , n441177 , n441178 );
nand ( n441180 , n441176 , n441179 );
buf ( n441181 , n441180 );
buf ( n441182 , C0 );
buf ( n441183 , C1 );
xor ( n441184 , n430464 , n430468 );
xor ( n441185 , n441184 , n430470 );
buf ( n441186 , n441185 );
buf ( n441187 , n430364 );
buf ( n441188 , n430376 );
xor ( n441189 , n441187 , n441188 );
buf ( n441190 , n441189 );
buf ( n441191 , n441141 );
buf ( n441192 , n441181 );
and ( n441193 , n441191 , n441192 );
buf ( n441194 , n441193 );
buf ( n441195 , n441070 );
buf ( n441196 , n440653 );
xor ( n441197 , n441195 , n441196 );
buf ( n441198 , n441197 );
buf ( n441199 , n440856 );
nand ( n441200 , n440852 , n440859 );
buf ( n441201 , n441200 );
xnor ( n441202 , n441199 , n441201 );
buf ( n441203 , n441202 );
buf ( n441204 , n440940 );
buf ( n441205 , n430909 );
buf ( n441206 , n85554 );
or ( n441207 , n441205 , n441206 );
buf ( n441208 , n441207 );
buf ( n441209 , n441208 );
xnor ( n441210 , n441204 , n441209 );
buf ( n441211 , n441210 );
buf ( n441212 , n440873 );
buf ( n441213 , n440962 );
xor ( n441214 , n441212 , n441213 );
buf ( n441215 , n441214 );
buf ( n441216 , n430882 );
buf ( n441217 , n440937 );
not ( n441218 , n441216 );
nand ( n441219 , n441218 , n441217 );
buf ( n441220 , n441219 );
buf ( n441221 , n428997 );
buf ( n441222 , n430793 );
not ( n441223 , n441221 );
nand ( n441224 , n441223 , n441222 );
buf ( n441225 , n441224 );
buf ( n441226 , n439492 );
buf ( n441227 , n441226 );
buf ( n441228 , n62969 );
nand ( n441229 , n441227 , n441228 );
buf ( n441230 , n441229 );
nand ( n441231 , n67616 , n440545 );
xnor ( n441232 , n440551 , n441231 );
buf ( n441233 , n440686 );
buf ( n441234 , n440983 );
xnor ( n441235 , n441233 , n441234 );
buf ( n441236 , n441235 );
buf ( n441237 , n85430 );
buf ( n441238 , n441013 );
xnor ( n441239 , n441237 , n441238 );
buf ( n441240 , n441239 );
buf ( n441241 , n439301 );
buf ( n441242 , n439823 );
buf ( n441243 , n439422 );
buf ( n441244 , n441243 );
not ( n441245 , n441241 );
not ( n441246 , n441242 );
or ( n441247 , n441245 , n441246 );
nand ( n441248 , n441247 , n441244 );
buf ( n441249 , n441248 );
buf ( n441250 , n430686 );
buf ( n441251 , n441036 );
buf ( n441252 , n430665 );
buf ( n441253 , n430677 );
or ( n441254 , n441252 , n441253 );
buf ( n441255 , n430683 );
nand ( n441256 , n441254 , n441255 );
buf ( n441257 , n441256 );
buf ( n441258 , n441257 );
buf ( n441259 , n441036 );
not ( n441260 , n441250 );
not ( n441261 , n441251 );
or ( n441262 , n441260 , n441261 );
or ( n441263 , n441258 , n441259 );
nand ( n441264 , n441262 , n441263 );
buf ( n441265 , n441264 );
nand ( n441266 , n439654 , n441133 );
or ( n441267 , n441249 , n441266 );
not ( n441268 , n388060 );
nor ( n441269 , n441268 , n441133 );
nand ( n441270 , n441269 , n441249 );
nor ( n441271 , n441266 , n388060 );
and ( n441272 , n439653 , n441130 );
nor ( n441273 , n441271 , n441272 );
nand ( n441274 , n441267 , n441270 , n441273 );
not ( n441275 , n434273 );
not ( n441276 , n439823 );
or ( n441277 , n441275 , n441276 );
nand ( n441278 , n439387 , n440291 );
nand ( n441279 , n441277 , n441278 );
not ( n441280 , n441279 );
not ( n441281 , n439397 );
nor ( n441282 , n441089 , n441281 );
nand ( n441283 , n441280 , n441282 );
not ( n441284 , n434804 );
not ( n441285 , n441284 );
nor ( n441286 , n441285 , n441092 );
nand ( n441287 , n441279 , n441286 );
not ( n441288 , n441092 );
not ( n441289 , n439397 );
and ( n441290 , n441288 , n441289 );
nor ( n441291 , n441089 , n441284 , n441281 );
nor ( n441292 , n441290 , n441291 );
nand ( n441293 , n441283 , n441287 , n441292 );
and ( n441294 , n440332 , n441009 );
not ( n441295 , n440332 );
and ( n441296 , n441295 , n441006 );
nor ( n441297 , n441294 , n441296 );
nand ( n441298 , n440612 , n439491 );
not ( n441299 , n441298 );
not ( n441300 , n62969 );
not ( n441301 , n440609 );
or ( n441302 , n441300 , n441301 );
nand ( n441303 , n441302 , n441226 );
not ( n441304 , n441303 );
or ( n441305 , n441299 , n441304 );
or ( n441306 , n441298 , n441303 );
nand ( n441307 , n441305 , n441306 );
nand ( n441308 , n439302 , n439544 , n439422 );
not ( n441309 , n35746 );
nand ( n441310 , n441309 , n36166 );
nor ( n441311 , n441310 , n441182 );
not ( n441312 , n441311 );
not ( n441313 , n441312 );
nand ( n441314 , n441313 , C1 );
nor ( n441315 , n40559 , n441314 );
nand ( n441316 , n441308 , n441315 );
not ( n441317 , n441309 );
not ( n441318 , n439659 );
or ( n441319 , n441317 , n441318 );
nand ( n441320 , n441319 , n383328 );
and ( n441321 , n441320 , n441183 );
nor ( n441322 , n441321 , n441194 );
and ( n441323 , n441322 , C1 );
not ( n441324 , n441323 );
not ( n441325 , n439654 );
or ( n441326 , n441324 , n441325 );
nand ( n441327 , n441326 , C1 );
nand ( n441328 , n441316 , n441327 );
and ( n441329 , n441328 , C1 );
not ( n441330 , n441328 );
and ( n441331 , n441330 , C0 );
nor ( n441332 , n441329 , n441331 );
not ( n441333 , n439609 );
nand ( n441334 , n439616 , n387753 );
not ( n441335 , n441334 );
nor ( n441336 , n40559 , n441312 );
not ( n441337 , n441336 );
not ( n441338 , n439862 );
or ( n441339 , n441337 , n441338 );
not ( n441340 , n441322 );
and ( n441341 , n439653 , n441311 );
nor ( n441342 , n441340 , n441341 );
nand ( n441343 , n441339 , n441342 );
and ( n441344 , n441343 , C1 );
not ( n441345 , n441343 );
and ( n441346 , n441345 , C0 );
nor ( n441347 , n441344 , n441346 );
not ( n441348 , n440464 );
not ( n441349 , n440032 );
or ( n441350 , n441348 , n441349 );
buf ( n441351 , n440466 );
nand ( n441352 , n441350 , n441351 );
buf ( n441353 , n438189 );
nand ( n441354 , n439362 , n441353 );
not ( n441355 , n441354 );
and ( n441356 , n441352 , n441355 );
not ( n441357 , n441352 );
and ( n441358 , n441357 , n441354 );
nor ( n441359 , n441356 , n441358 );
not ( n441360 , n438190 );
not ( n441361 , n441360 );
not ( n441362 , n440032 );
or ( n441363 , n441361 , n441362 );
not ( n441364 , n439363 );
nand ( n441365 , n441363 , n441364 );
buf ( n441366 , n439370 );
nand ( n441367 , n441366 , n438658 );
not ( n441368 , n441367 );
and ( n441369 , n441365 , n441368 );
not ( n441370 , n441365 );
and ( n441371 , n441370 , n441367 );
nor ( n441372 , n441369 , n441371 );
buf ( n441373 , n430827 );
or ( n441374 , n81036 , n81021 );
or ( n441375 , n441373 , n441374 );
nand ( n441376 , n81021 , n81036 );
or ( n441377 , n441376 , n441373 );
not ( n441378 , n85467 );
not ( n441379 , n81037 );
or ( n441380 , n441378 , n441379 );
nand ( n441381 , n441380 , n441373 );
nand ( n441382 , n441375 , n441377 , n441381 );
not ( n441383 , n56293 );
not ( n441384 , n440376 );
or ( n441385 , n441383 , n441384 );
nand ( n441386 , n441385 , n440361 );
not ( n441387 , n439537 );
nand ( n441388 , n441387 , n439514 );
not ( n441389 , n441388 );
and ( n441390 , n441386 , n441389 );
not ( n441391 , n441386 );
and ( n441392 , n441391 , n441388 );
nor ( n441393 , n441390 , n441392 );
nand ( n441394 , n441316 , n441327 , C1 );
nand ( n441395 , n441394 , C1 );
buf ( n441396 , n441395 );
and ( n441397 , n440551 , n440546 );
nor ( n441398 , n441397 , n440558 );
and ( n441399 , n441398 , n440994 );
not ( n441400 , n441398 );
and ( n441401 , n441400 , n440997 );
nor ( n441402 , n441399 , n441401 );
not ( n441403 , n440545 );
not ( n441404 , n440551 );
or ( n441405 , n441403 , n441404 );
nand ( n441406 , n441405 , n67616 );
and ( n441407 , n441406 , n440993 );
not ( n441408 , n441406 );
and ( n441409 , n441408 , n440990 );
nor ( n441410 , n441407 , n441409 );
not ( n441411 , n85414 );
and ( n441412 , n441225 , n85424 );
not ( n441413 , n441225 );
and ( n441414 , n441413 , n85423 );
nor ( n441415 , n441412 , n441414 );
not ( n441416 , n85417 );
not ( n441417 , n441018 );
or ( n441418 , n441416 , n441417 );
or ( n441419 , n441018 , n85417 );
nand ( n441420 , n441418 , n441419 );
not ( n441421 , n40040 );
nor ( n441422 , n441421 , n441335 );
not ( n441423 , n441333 );
nor ( n441424 , n441334 , n441423 , n40040 );
not ( n441425 , n441220 );
buf ( n441426 , n85471 );
not ( n441427 , n441426 );
or ( n441428 , n441425 , n441427 );
or ( n441429 , n441426 , n441220 );
nand ( n441430 , n441428 , n441429 );
not ( n441431 , n441230 );
not ( n441432 , n440609 );
or ( n441433 , n441431 , n441432 );
or ( n441434 , n441230 , n440609 );
nand ( n441435 , n441433 , n441434 );
buf ( n441436 , n440976 );
buf ( n441437 , n440979 );
buf ( n441438 , n440746 );
and ( n441439 , n441438 , n441437 );
not ( n441440 , n441438 );
and ( n441441 , n441440 , n441436 );
nor ( n441442 , n441439 , n441441 );
buf ( n441443 , n441442 );
xor ( n441444 , n422907 , n423399 );
xor ( n441445 , n441444 , n430925 );
buf ( n441446 , n441445 );
buf ( n441447 , n440966 );
buf ( n441448 , n440969 );
buf ( n441449 , n440825 );
and ( n441450 , n441449 , n441448 );
not ( n441451 , n441449 );
and ( n441452 , n441451 , n441447 );
nor ( n441453 , n441450 , n441452 );
buf ( n441454 , n441453 );
and ( n441455 , n430772 , n85413 );
not ( n441456 , n430772 );
and ( n441457 , n441456 , n430776 );
nor ( n441458 , n441455 , n441457 );
not ( n441459 , n441334 );
nand ( n441460 , n441459 , n441333 );
or ( n441461 , n441460 , n439795 );
nand ( n441462 , n439795 , n441422 );
not ( n441463 , n441335 );
not ( n441464 , n441333 );
and ( n441465 , n441463 , n441464 );
nor ( n441466 , n441465 , n441424 );
nand ( n441467 , n441461 , n441462 , n441466 );
buf ( n441468 , n432762 );
buf ( n441469 , n432854 );
nand ( n441470 , n441468 , n441469 );
buf ( n441471 , n441470 );
buf ( n441472 , n441471 );
buf ( n441473 , n441471 );
not ( n441474 , n441473 );
buf ( n441475 , n441474 );
buf ( n441476 , n441475 );
and ( n441477 , n440825 , n440819 , n432806 );
nor ( n441478 , n441477 , n432845 );
not ( n441479 , n441478 );
buf ( n441480 , n441479 );
and ( n441481 , n441480 , n441476 );
not ( n441482 , n441480 );
and ( n441483 , n441482 , n441472 );
nor ( n441484 , n441481 , n441483 );
buf ( n441485 , n441484 );
nand ( n441486 , n441284 , n439397 );
not ( n441487 , n441486 );
and ( n441488 , n441279 , n441487 );
not ( n441489 , n441279 );
and ( n441490 , n441489 , n441486 );
nor ( n441491 , n441488 , n441490 );
xor ( n441492 , n427447 , n427450 );
xor ( n441493 , n441492 , n430823 );
buf ( n441494 , n441493 );
buf ( n441495 , n85468 );
buf ( n441496 , n441001 );
xnor ( n441497 , n441495 , n441496 );
buf ( n441498 , n441497 );
nand ( n441499 , n430587 , n85192 );
not ( n441500 , n441499 );
nand ( n441501 , n430545 , n430265 );
not ( n441502 , n441501 );
or ( n441503 , n441500 , n441502 );
or ( n441504 , n441501 , n441499 );
nand ( n441505 , n441503 , n441504 );
not ( n441506 , n28556 );
xnor ( n441507 , n376032 , n372536 );
not ( n441508 , n441507 );
or ( n441509 , n441506 , n441508 );
or ( n441510 , n441507 , n28556 );
nand ( n441511 , n441509 , n441510 );
xor ( n441512 , n376064 , n376065 );
xor ( n441513 , n441512 , n376067 );
buf ( n441514 , n441513 );
not ( n441515 , n441411 );
not ( n441516 , n85391 );
or ( n441517 , n441515 , n441516 );
not ( n441518 , n85391 );
not ( n441519 , n441458 );
and ( n441520 , n441518 , n441519 );
and ( n441521 , n85391 , n85416 );
nor ( n441522 , n441520 , n441521 );
nand ( n441523 , n441517 , n441522 );
xor ( n441524 , n375860 , n376332 );
xor ( n441525 , n441524 , n376336 );
buf ( n441526 , n441525 );
xor ( n441527 , n375878 , n375882 );
xor ( n441528 , n441527 , n376327 );
buf ( n441529 , n441528 );
xor ( n441530 , n372360 , n24420 );
xor ( n441531 , n371212 , n371192 );
xor ( n441532 , n441531 , n24381 );
not ( n441533 , n441310 );
not ( n441534 , n441533 );
not ( n441535 , n439655 );
or ( n441536 , n441534 , n441535 );
not ( n441537 , n441320 );
nand ( n441538 , n441536 , n441537 );
nor ( n441539 , n441194 , n441182 );
and ( n441540 , n441538 , n441539 );
not ( n441541 , n441538 );
not ( n441542 , n441539 );
and ( n441543 , n441541 , n441542 );
nor ( n441544 , n441540 , n441543 );
xor ( n441545 , n372356 , n372021 );
xor ( n441546 , n371187 , n371164 );
not ( n441547 , n24377 );
xor ( n441548 , n441546 , n441547 );
not ( C0n , n0 );
and ( C0 , C0n , n0 );
not ( C1n , n0 );
or ( C1 , C1n , n0 );
endmodule
