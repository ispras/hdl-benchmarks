//
// Conformal-LEC Version 14.20-d237 ( 26-Mar-2015) ( 64 bit executable)
//
module top ( PI_clock , PI_reset , n0 , n1 , n2 , n3 , n4 , n5 , n6 , 
  n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , 
  n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , 
  n27 , n28 , n29 , n30 , n31 , DFF_state_reg_Q , n32 , n33 , n34 , n35 , 
  n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , 
  n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , 
  n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , 
  n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , 
  n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , 
  n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , 
  n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , 
  n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , 
  n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , 
  n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , 
  n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , 
  n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , 
  n156 , n157 , n158 , DFF_B_reg_Q , n159 , n160 , n161 , n162 , n163 , n164 , 
  n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , 
  n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , 
  n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , 
  n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , 
  n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , 
  n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , 
  n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , 
  n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , DFF_rd_reg_Q , DFF_wr_reg_Q , 
  n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , 
  n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , 
  n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , 
  n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , 
  n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , 
  n293 , n294 , PO_rd , PO_wr , DFF_state_reg_S , DFF_state_reg_R , DFF_state_reg_CK , DFF_state_reg_D , n295 , n296 , 
  n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , 
  n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , 
  n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , 
  n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , 
  n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , 
  n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , 
  n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , 
  n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , 
  n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , 
  n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , 
  n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , 
  n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , 
  n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , 
  n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , 
  n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , 
  n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , 
  n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , 
  n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , 
  n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , 
  n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , 
  n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , 
  n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , 
  n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , 
  n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , 
  n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , 
  n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , 
  n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , 
  n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , 
  n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , 
  n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , 
  n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , 
  n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , 
  n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , 
  n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , 
  n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , 
  n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , 
  n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , 
  n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , 
  n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , 
  n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , 
  n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , 
  n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , 
  n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , 
  n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , 
  n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , 
  n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , 
  n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , 
  n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , 
  n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , 
  n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , 
  n797 , n798 , n799 , n800 , n801 , n802 , DFF_B_reg_S , DFF_B_reg_R , DFF_B_reg_CK , DFF_B_reg_D , 
  n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , 
  n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , 
  n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , 
  n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , 
  n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , 
  n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , 
  n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , 
  n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , 
  n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , 
  n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , 
  n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , 
  n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , 
  n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , 
  n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , 
  n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , 
  n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , 
  n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , 
  n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , 
  n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , 
  n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , 
  n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , 
  n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , 
  n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , 
  n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , 
  n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , 
  n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , 
  n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , 
  n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , 
  n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , 
  n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , 
  n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , 
  n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , 
  n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , 
  n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , DFF_rd_reg_S , DFF_rd_reg_R , DFF_rd_reg_CK , DFF_rd_reg_D , 
  DFF_wr_reg_S , DFF_wr_reg_R , DFF_wr_reg_CK , DFF_wr_reg_D);
input PI_clock , PI_reset , n0 , n1 , n2 , n3 , n4 , n5 , n6 , 
  n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , 
  n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , 
  n27 , n28 , n29 , n30 , n31 , DFF_state_reg_Q , n32 , n33 , n34 , n35 , 
  n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , 
  n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , 
  n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , 
  n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , 
  n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , 
  n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , 
  n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , 
  n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , 
  n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , 
  n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , 
  n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , 
  n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , 
  n156 , n157 , n158 , DFF_B_reg_Q , n159 , n160 , n161 , n162 , n163 , n164 , 
  n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , 
  n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , 
  n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , 
  n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , 
  n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , 
  n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , 
  n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , 
  n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , DFF_rd_reg_Q , DFF_wr_reg_Q;
output n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , 
  n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , 
  n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , 
  n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , 
  n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , 
  n292 , n293 , n294 , PO_rd , PO_wr , DFF_state_reg_S , DFF_state_reg_R , DFF_state_reg_CK , DFF_state_reg_D , n295 , 
  n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , 
  n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , 
  n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , 
  n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , 
  n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , 
  n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , 
  n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , 
  n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , 
  n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , 
  n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , 
  n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , 
  n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , 
  n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , 
  n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , 
  n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , 
  n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , 
  n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , 
  n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , 
  n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , 
  n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , 
  n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , 
  n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , 
  n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , 
  n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , 
  n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , 
  n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , 
  n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , 
  n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , 
  n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , 
  n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , 
  n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , 
  n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , 
  n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , 
  n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , 
  n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , 
  n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , 
  n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , 
  n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , 
  n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , 
  n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , 
  n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , 
  n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , 
  n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , 
  n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , 
  n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , 
  n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , 
  n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , 
  n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , 
  n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , 
  n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , 
  n796 , n797 , n798 , n799 , n800 , n801 , n802 , DFF_B_reg_S , DFF_B_reg_R , DFF_B_reg_CK , 
  DFF_B_reg_D , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , 
  n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , 
  n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , 
  n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , 
  n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , 
  n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , 
  n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , 
  n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , 
  n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , 
  n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , 
  n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , 
  n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , 
  n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , 
  n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , 
  n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , 
  n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , 
  n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , 
  n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , 
  n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , 
  n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , 
  n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , 
  n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , 
  n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , 
  n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , 
  n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , 
  n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , 
  n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , 
  n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , 
  n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , 
  n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , 
  n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , 
  n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , 
  n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , 
  n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , DFF_rd_reg_S , DFF_rd_reg_R , DFF_rd_reg_CK , 
  DFF_rd_reg_D , DFF_wr_reg_S , DFF_wr_reg_R , DFF_wr_reg_CK , DFF_wr_reg_D;

wire n68421 , n68422 , n68423 , n68424 , n68425 , n68426 , n68427 , n68428 , n68429 , 
   n68430 , n68431 , n68432 , n68433 , n68434 , n68435 , n68436 , n68437 , n68438 , n68439 , 
   n68440 , n68441 , n68442 , n68443 , n68444 , n68445 , n68446 , n68447 , n68448 , n68449 , 
   n68450 , n68451 , n68452 , n68453 , n68454 , n68455 , n68456 , n68457 , n68458 , n68459 , 
   n68460 , n68461 , n68462 , n68463 , n68464 , n68465 , n68466 , n68467 , n68468 , n68469 , 
   n68470 , n68471 , n68472 , n68473 , n68474 , n68475 , n68476 , n68477 , n68478 , n68479 , 
   n68480 , n68481 , n68482 , n68483 , n68484 , n68485 , n68486 , n68487 , n68488 , n68489 , 
   n68490 , n68491 , n68492 , n68493 , n68494 , n68495 , n68496 , n68497 , n68498 , n68499 , 
   n68500 , n68501 , n68502 , n68503 , n68504 , n68505 , n68506 , n68507 , n68508 , n68509 , 
   n68510 , n68511 , n68512 , n68513 , n68514 , n68515 , n68516 , n68517 , n68518 , n68519 , 
   n68520 , n68521 , n68522 , n68523 , n68524 , n68525 , n68526 , n68527 , n68528 , n68529 , 
   n68530 , n68531 , n68532 , n68533 , n68534 , n68535 , n68536 , n68537 , n68538 , n68539 , 
   n68540 , n68541 , n68542 , n68543 , n68544 , n68545 , n68546 , n68547 , n68548 , n68549 , 
   n68550 , n68551 , n68552 , n68553 , n68554 , n68555 , n68556 , n68557 , n68558 , n68559 , 
   n68560 , n68561 , n68562 , n68563 , n68564 , n68565 , n68566 , n68567 , n68568 , n68569 , 
   n68570 , n68571 , n68572 , n68573 , n68574 , n68575 , n68576 , n68577 , n68578 , n68579 , 
   n68580 , n68581 , n68582 , n68583 , n68584 , n68585 , n68586 , n68587 , n68588 , n68589 , 
   n68590 , n68591 , n68592 , n68593 , n68594 , n68595 , n68596 , n68597 , n68598 , n68599 , 
   n68600 , n68601 , n68602 , n68603 , n68604 , n68605 , n68606 , n68607 , n68608 , n68609 , 
   n68610 , n68611 , n68612 , n68613 , n68614 , n68615 , n68616 , n68617 , n68618 , n68619 , 
   n68620 , n68621 , n68622 , n68623 , n68624 , n68625 , n68626 , n68627 , n68628 , n68629 , 
   n68630 , n68631 , n68632 , n68633 , n68634 , n68635 , n68636 , n68637 , n68638 , n68639 , 
   n68640 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n68648 , n68649 , 
   n68650 , n2508 , n2509 , n68653 , n68654 , n68655 , n2513 , n2514 , n2515 , n2516 , 
   n2517 , n2518 , n2519 , n68663 , n68664 , n68665 , n2523 , n2524 , n68668 , n68669 , 
   n68670 , n2528 , n2529 , n68673 , n68674 , n2532 , n2533 , n2534 , n68678 , n68679 , 
   n68680 , n2538 , n2539 , n68683 , n68684 , n68685 , n2543 , n2544 , n68688 , n68689 , 
   n2547 , n2548 , n2549 , n68693 , n68694 , n68695 , n2553 , n2554 , n68698 , n68699 , 
   n68700 , n2558 , n2559 , n68703 , n68704 , n2562 , n2563 , n2564 , n68708 , n68709 , 
   n68710 , n2568 , n2569 , n68713 , n68714 , n68715 , n2573 , n2574 , n68718 , n68719 , 
   n2577 , n2578 , n2579 , n68723 , n68724 , n68725 , n2583 , n2584 , n68728 , n68729 , 
   n68730 , n2588 , n2589 , n68733 , n68734 , n2592 , n2593 , n2594 , n68738 , n68739 , 
   n68740 , n2598 , n2599 , n68743 , n68744 , n68745 , n2603 , n2604 , n2605 , n2606 , 
   n68750 , n68751 , n2609 , n68753 , n68754 , n68755 , n2613 , n68757 , n68758 , n68759 , 
   n68760 , n2618 , n68762 , n68763 , n2621 , n2622 , n2623 , n2624 , n68768 , n68769 , 
   n68770 , n2628 , n2629 , n68773 , n68774 , n68775 , n2633 , n2634 , n2635 , n2636 , 
   n2637 , n2638 , n2639 , n68783 , n68784 , n68785 , n2643 , n2644 , n68788 , n68789 , 
   n68790 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n68798 , n68799 , 
   n68800 , n2658 , n2659 , n68803 , n68804 , n68805 , n2663 , n2664 , n2665 , n2666 , 
   n2667 , n2668 , n2669 , n68813 , n68814 , n68815 , n2673 , n2674 , n68818 , n68819 , 
   n68820 , n68821 , n68822 , n2680 , n2681 , n2682 , n68826 , n68827 , n68828 , n68829 , 
   n68830 , n2688 , n2689 , n68833 , n68834 , n68835 , n2693 , n2694 , n2695 , n2696 , 
   n2697 , n2698 , n68842 , n68843 , n68844 , n68845 , n2703 , n68847 , n68848 , n68849 , 
   n68850 , n68851 , n68852 , n2710 , n68854 , n68855 , n68856 , n68857 , n68858 , n68859 , 
   n68860 , n68861 , n68862 , n68863 , n68864 , n68865 , n68866 , n68867 , n68868 , n68869 , 
   n68870 , n2728 , n68872 , n68873 , n68874 , n68875 , n68876 , n2734 , n68878 , n68879 , 
   n68880 , n68881 , n68882 , n68883 , n68884 , n68885 , n68886 , n2744 , n68888 , n68889 , 
   n68890 , n68891 , n68892 , n68893 , n68894 , n68895 , n2753 , n68897 , n68898 , n68899 , 
   n68900 , n2758 , n68902 , n68903 , n68904 , n68905 , n68906 , n68907 , n68908 , n68909 , 
   n68910 , n68911 , n68912 , n68913 , n68914 , n68915 , n68916 , n2774 , n68918 , n68919 , 
   n68920 , n68921 , n68922 , n68923 , n68924 , n68925 , n68926 , n2784 , n68928 , n68929 , 
   n68930 , n68931 , n68932 , n68933 , n68934 , n68935 , n68936 , n68937 , n68938 , n68939 , 
   n68940 , n68941 , n68942 , n68943 , n68944 , n68945 , n68946 , n68947 , n68948 , n68949 , 
   n68950 , n68951 , n68952 , n68953 , n68954 , n68955 , n68956 , n68957 , n68958 , n68959 , 
   n68960 , n68961 , n68962 , n68963 , n68964 , n68965 , n68966 , n68967 , n68968 , n68969 , 
   n68970 , n68971 , n68972 , n68973 , n68974 , n68975 , n68976 , n68977 , n68978 , n68979 , 
   n68980 , n68981 , n68982 , n68983 , n68984 , n68985 , n68986 , n68987 , n68988 , n68989 , 
   n68990 , n68991 , n68992 , n68993 , n68994 , n68995 , n68996 , n68997 , n68998 , n68999 , 
   n69000 , n69001 , n69002 , n69003 , n69004 , n69005 , n69006 , n69007 , n69008 , n69009 , 
   n69010 , n69011 , n69012 , n69013 , n69014 , n69015 , n69016 , n69017 , n69018 , n69019 , 
   n69020 , n69021 , n69022 , n69023 , n69024 , n69025 , n69026 , n69027 , n69028 , n69029 , 
   n69030 , n69031 , n69032 , n69033 , n69034 , n69035 , n69036 , n69037 , n69038 , n69039 , 
   n69040 , n69041 , n69042 , n69043 , n69044 , n69045 , n69046 , n69047 , n69048 , n69049 , 
   n69050 , n69051 , n69052 , n69053 , n69054 , n69055 , n69056 , n69057 , n69058 , n69059 , 
   n69060 , n69061 , n69062 , n69063 , n69064 , n69065 , n69066 , n69067 , n69068 , n69069 , 
   n69070 , n69071 , n69072 , n69073 , n69074 , n69075 , n69076 , n69077 , n69078 , n69079 , 
   n69080 , n69081 , n69082 , n69083 , n69084 , n69085 , n69086 , n69087 , n69088 , n69089 , 
   n69090 , n69091 , n69092 , n69093 , n69094 , n69095 , n69096 , n69097 , n69098 , n69099 , 
   n69100 , n69101 , n69102 , n69103 , n69104 , n69105 , n69106 , n69107 , n69108 , n69109 , 
   n69110 , n69111 , n69112 , n69113 , n69114 , n69115 , n69116 , n69117 , n69118 , n69119 , 
   n69120 , n69121 , n69122 , n69123 , n69124 , n69125 , n69126 , n69127 , n69128 , n69129 , 
   n69130 , n69131 , n69132 , n69133 , n69134 , n69135 , n69136 , n69137 , n69138 , n69139 , 
   n69140 , n69141 , n69142 , n3000 , n69144 , n69145 , n69146 , n69147 , n69148 , n69149 , 
   n69150 , n69151 , n69152 , n69153 , n69154 , n69155 , n69156 , n69157 , n69158 , n69159 , 
   n69160 , n69161 , n69162 , n69163 , n69164 , n69165 , n69166 , n69167 , n69168 , n69169 , 
   n69170 , n69171 , n69172 , n69173 , n69174 , n69175 , n69176 , n69177 , n69178 , n69179 , 
   n69180 , n69181 , n69182 , n69183 , n69184 , n69185 , n69186 , n69187 , n69188 , n69189 , 
   n69190 , n69191 , n69192 , n69193 , n69194 , n69195 , n69196 , n69197 , n69198 , n69199 , 
   n69200 , n3058 , n3059 , n69203 , n69204 , n69205 , n69206 , n69207 , n69208 , n3066 , 
   n69210 , n69211 , n69212 , n69213 , n69214 , n69215 , n69216 , n69217 , n69218 , n69219 , 
   n69220 , n69221 , n69222 , n69223 , n69224 , n69225 , n69226 , n69227 , n69228 , n69229 , 
   n69230 , n69231 , n69232 , n69233 , n69234 , n69235 , n69236 , n69237 , n69238 , n69239 , 
   n69240 , n69241 , n69242 , n69243 , n69244 , n69245 , n69246 , n69247 , n69248 , n69249 , 
   n69250 , n69251 , n69252 , n69253 , n69254 , n69255 , n69256 , n69257 , n69258 , n69259 , 
   n69260 , n69261 , n69262 , n69263 , n69264 , n69265 , n69266 , n69267 , n69268 , n69269 , 
   n69270 , n69271 , n69272 , n69273 , n69274 , n69275 , n69276 , n69277 , n69278 , n69279 , 
   n69280 , n69281 , n69282 , n69283 , n69284 , n69285 , n69286 , n69287 , n69288 , n69289 , 
   n69290 , n69291 , n69292 , n69293 , n69294 , n69295 , n69296 , n69297 , n69298 , n69299 , 
   n69300 , n69301 , n69302 , n69303 , n69304 , n69305 , n69306 , n69307 , n69308 , n69309 , 
   n69310 , n69311 , n69312 , n69313 , n69314 , n69315 , n69316 , n69317 , n69318 , n69319 , 
   n69320 , n69321 , n69322 , n69323 , n69324 , n69325 , n69326 , n69327 , n69328 , n69329 , 
   n69330 , n69331 , n69332 , n69333 , n69334 , n69335 , n69336 , n69337 , n69338 , n69339 , 
   n69340 , n69341 , n69342 , n69343 , n69344 , n69345 , n69346 , n69347 , n69348 , n69349 , 
   n69350 , n69351 , n69352 , n69353 , n69354 , n69355 , n69356 , n69357 , n69358 , n69359 , 
   n69360 , n69361 , n69362 , n69363 , n69364 , n69365 , n69366 , n69367 , n69368 , n69369 , 
   n69370 , n69371 , n69372 , n69373 , n69374 , n69375 , n69376 , n69377 , n69378 , n69379 , 
   n69380 , n69381 , n69382 , n69383 , n69384 , n69385 , n69386 , n69387 , n69388 , n69389 , 
   n69390 , n69391 , n69392 , n69393 , n69394 , n69395 , n69396 , n69397 , n69398 , n69399 , 
   n69400 , n69401 , n69402 , n69403 , n69404 , n69405 , n69406 , n69407 , n69408 , n69409 , 
   n69410 , n69411 , n69412 , n69413 , n69414 , n69415 , n69416 , n69417 , n69418 , n3276 , 
   n69420 , n69421 , n69422 , n69423 , n69424 , n3282 , n69426 , n69427 , n69428 , n69429 , 
   n69430 , n3288 , n69432 , n69433 , n69434 , n3292 , n69436 , n69437 , n69438 , n69439 , 
   n69440 , n69441 , n69442 , n69443 , n3301 , n69445 , n69446 , n3304 , n69448 , n69449 , 
   n69450 , n69451 , n69452 , n69453 , n69454 , n69455 , n69456 , n69457 , n69458 , n3316 , 
   n69460 , n69461 , n69462 , n3320 , n69464 , n69465 , n69466 , n3324 , n69468 , n69469 , 
   n3327 , n69471 , n69472 , n69473 , n69474 , n69475 , n69476 , n69477 , n69478 , n3336 , 
   n69480 , n69481 , n69482 , n69483 , n69484 , n3342 , n69486 , n3344 , n69488 , n3346 , 
   n69490 , n69491 , n69492 , n3350 , n69494 , n69495 , n69496 , n69497 , n69498 , n3356 , 
   n69500 , n69501 , n3359 , n69503 , n69504 , n69505 , n69506 , n69507 , n69508 , n69509 , 
   n69510 , n69511 , n69512 , n69513 , n69514 , n69515 , n69516 , n69517 , n69518 , n69519 , 
   n69520 , n69521 , n69522 , n69523 , n69524 , n69525 , n69526 , n69527 , n69528 , n69529 , 
   n69530 , n69531 , n69532 , n69533 , n69534 , n69535 , n69536 , n69537 , n69538 , n69539 , 
   n69540 , n69541 , n69542 , n69543 , n69544 , n69545 , n69546 , n69547 , n3405 , n69549 , 
   n69550 , n69551 , n69552 , n69553 , n69554 , n3412 , n69556 , n69557 , n69558 , n69559 , 
   n69560 , n69561 , n69562 , n69563 , n69564 , n69565 , n69566 , n69567 , n69568 , n69569 , 
   n69570 , n69571 , n69572 , n69573 , n69574 , n69575 , n69576 , n69577 , n69578 , n69579 , 
   n69580 , n69581 , n69582 , n69583 , n69584 , n3442 , n69586 , n69587 , n69588 , n69589 , 
   n69590 , n69591 , n69592 , n3450 , n69594 , n69595 , n69596 , n3454 , n69598 , n69599 , 
   n69600 , n69601 , n69602 , n69603 , n69604 , n69605 , n69606 , n69607 , n69608 , n3466 , 
   n69610 , n69611 , n69612 , n3470 , n69614 , n69615 , n69616 , n69617 , n69618 , n69619 , 
   n69620 , n69621 , n69622 , n69623 , n69624 , n69625 , n69626 , n69627 , n69628 , n69629 , 
   n69630 , n69631 , n3489 , n69633 , n69634 , n69635 , n69636 , n69637 , n69638 , n69639 , 
   n69640 , n3498 , n69642 , n69643 , n69644 , n69645 , n69646 , n69647 , n69648 , n69649 , 
   n69650 , n69651 , n69652 , n3510 , n69654 , n69655 , n69656 , n3514 , n69658 , n69659 , 
   n69660 , n69661 , n69662 , n69663 , n69664 , n69665 , n69666 , n69667 , n69668 , n69669 , 
   n69670 , n69671 , n3529 , n69673 , n69674 , n69675 , n69676 , n69677 , n69678 , n69679 , 
   n69680 , n69681 , n69682 , n69683 , n69684 , n69685 , n69686 , n69687 , n69688 , n69689 , 
   n69690 , n69691 , n69692 , n69693 , n69694 , n3552 , n69696 , n69697 , n69698 , n69699 , 
   n69700 , n69701 , n69702 , n69703 , n3561 , n69705 , n69706 , n69707 , n69708 , n69709 , 
   n69710 , n69711 , n3569 , n69713 , n69714 , n69715 , n69716 , n69717 , n69718 , n69719 , 
   n69720 , n69721 , n69722 , n3580 , n69724 , n69725 , n69726 , n3584 , n69728 , n69729 , 
   n69730 , n69731 , n69732 , n69733 , n3591 , n69735 , n69736 , n69737 , n69738 , n69739 , 
   n69740 , n69741 , n69742 , n69743 , n69744 , n69745 , n69746 , n69747 , n69748 , n69749 , 
   n69750 , n69751 , n69752 , n69753 , n69754 , n69755 , n69756 , n69757 , n69758 , n69759 , 
   n69760 , n69761 , n69762 , n3620 , n69764 , n69765 , n69766 , n69767 , n69768 , n69769 , 
   n69770 , n69771 , n69772 , n69773 , n69774 , n69775 , n69776 , n69777 , n69778 , n3636 , 
   n69780 , n69781 , n69782 , n69783 , n69784 , n69785 , n69786 , n69787 , n69788 , n69789 , 
   n69790 , n69791 , n69792 , n69793 , n69794 , n69795 , n69796 , n69797 , n69798 , n69799 , 
   n69800 , n69801 , n69802 , n69803 , n69804 , n69805 , n69806 , n69807 , n69808 , n69809 , 
   n69810 , n69811 , n69812 , n69813 , n69814 , n69815 , n69816 , n69817 , n69818 , n69819 , 
   n69820 , n69821 , n69822 , n69823 , n69824 , n69825 , n69826 , n69827 , n69828 , n69829 , 
   n69830 , n69831 , n69832 , n69833 , n69834 , n69835 , n69836 , n69837 , n69838 , n69839 , 
   n69840 , n69841 , n69842 , n69843 , n69844 , n69845 , n69846 , n69847 , n69848 , n69849 , 
   n3707 , n69851 , n69852 , n69853 , n69854 , n69855 , n69856 , n69857 , n69858 , n69859 , 
   n69860 , n69861 , n69862 , n69863 , n3721 , n69865 , n69866 , n69867 , n69868 , n69869 , 
   n69870 , n69871 , n69872 , n69873 , n69874 , n69875 , n69876 , n69877 , n69878 , n69879 , 
   n69880 , n69881 , n69882 , n69883 , n69884 , n69885 , n69886 , n69887 , n69888 , n69889 , 
   n69890 , n69891 , n69892 , n69893 , n69894 , n69895 , n69896 , n69897 , n69898 , n69899 , 
   n69900 , n69901 , n69902 , n69903 , n69904 , n69905 , n69906 , n69907 , n69908 , n69909 , 
   n69910 , n69911 , n69912 , n69913 , n3771 , n69915 , n69916 , n69917 , n69918 , n69919 , 
   n69920 , n69921 , n69922 , n69923 , n69924 , n69925 , n69926 , n69927 , n69928 , n69929 , 
   n69930 , n69931 , n69932 , n69933 , n69934 , n69935 , n69936 , n69937 , n69938 , n69939 , 
   n69940 , n69941 , n3799 , n69943 , n69944 , n69945 , n69946 , n69947 , n69948 , n69949 , 
   n69950 , n69951 , n69952 , n69953 , n69954 , n69955 , n69956 , n69957 , n3815 , n69959 , 
   n69960 , n69961 , n69962 , n69963 , n69964 , n69965 , n69966 , n69967 , n69968 , n69969 , 
   n69970 , n69971 , n69972 , n69973 , n69974 , n69975 , n69976 , n69977 , n69978 , n69979 , 
   n69980 , n69981 , n69982 , n69983 , n69984 , n69985 , n69986 , n69987 , n69988 , n69989 , 
   n69990 , n69991 , n69992 , n69993 , n69994 , n69995 , n69996 , n69997 , n69998 , n69999 , 
   n70000 , n70001 , n70002 , n70003 , n70004 , n70005 , n70006 , n70007 , n70008 , n70009 , 
   n70010 , n70011 , n70012 , n70013 , n70014 , n70015 , n70016 , n70017 , n70018 , n70019 , 
   n70020 , n70021 , n70022 , n70023 , n70024 , n70025 , n70026 , n70027 , n70028 , n70029 , 
   n70030 , n70031 , n70032 , n70033 , n70034 , n70035 , n70036 , n70037 , n70038 , n70039 , 
   n70040 , n70041 , n70042 , n70043 , n70044 , n70045 , n70046 , n70047 , n70048 , n70049 , 
   n70050 , n70051 , n70052 , n70053 , n70054 , n70055 , n70056 , n70057 , n70058 , n70059 , 
   n70060 , n70061 , n70062 , n70063 , n70064 , n70065 , n70066 , n70067 , n70068 , n70069 , 
   n70070 , n70071 , n70072 , n70073 , n70074 , n70075 , n70076 , n70077 , n70078 , n70079 , 
   n70080 , n70081 , n70082 , n70083 , n70084 , n70085 , n70086 , n70087 , n70088 , n70089 , 
   n70090 , n70091 , n70092 , n70093 , n70094 , n70095 , n70096 , n70097 , n70098 , n70099 , 
   n70100 , n70101 , n70102 , n70103 , n70104 , n70105 , n70106 , n70107 , n70108 , n70109 , 
   n70110 , n70111 , n70112 , n70113 , n70114 , n70115 , n70116 , n70117 , n70118 , n70119 , 
   n70120 , n70121 , n70122 , n70123 , n70124 , n70125 , n70126 , n70127 , n70128 , n70129 , 
   n70130 , n70131 , n70132 , n70133 , n70134 , n70135 , n70136 , n70137 , n70138 , n70139 , 
   n70140 , n3998 , n70142 , n70143 , n70144 , n70145 , n70146 , n70147 , n70148 , n70149 , 
   n70150 , n70151 , n70152 , n70153 , n70154 , n4012 , n70156 , n70157 , n70158 , n70159 , 
   n70160 , n70161 , n70162 , n70163 , n70164 , n4022 , n70166 , n70167 , n70168 , n70169 , 
   n70170 , n70171 , n70172 , n4030 , n70174 , n70175 , n70176 , n70177 , n70178 , n70179 , 
   n70180 , n70181 , n70182 , n70183 , n70184 , n70185 , n70186 , n70187 , n70188 , n70189 , 
   n70190 , n70191 , n70192 , n70193 , n70194 , n70195 , n70196 , n70197 , n70198 , n70199 , 
   n70200 , n70201 , n70202 , n70203 , n70204 , n70205 , n70206 , n70207 , n70208 , n70209 , 
   n70210 , n70211 , n70212 , n70213 , n70214 , n70215 , n70216 , n70217 , n70218 , n70219 , 
   n70220 , n70221 , n70222 , n70223 , n70224 , n70225 , n70226 , n70227 , n70228 , n70229 , 
   n70230 , n70231 , n70232 , n70233 , n70234 , n70235 , n70236 , n70237 , n70238 , n70239 , 
   n70240 , n70241 , n70242 , n70243 , n70244 , n70245 , n70246 , n70247 , n70248 , n70249 , 
   n70250 , n70251 , n70252 , n70253 , n70254 , n70255 , n70256 , n70257 , n70258 , n70259 , 
   n70260 , n70261 , n70262 , n70263 , n70264 , n70265 , n70266 , n70267 , n70268 , n70269 , 
   n70270 , n70271 , n70272 , n70273 , n70274 , n70275 , n70276 , n70277 , n70278 , n70279 , 
   n70280 , n70281 , n70282 , n70283 , n70284 , n70285 , n70286 , n70287 , n70288 , n70289 , 
   n70290 , n70291 , n70292 , n70293 , n70294 , n70295 , n70296 , n70297 , n70298 , n70299 , 
   n70300 , n70301 , n70302 , n70303 , n70304 , n70305 , n70306 , n70307 , n70308 , n70309 , 
   n70310 , n70311 , n70312 , n70313 , n70314 , n70315 , n70316 , n70317 , n70318 , n70319 , 
   n70320 , n70321 , n70322 , n70323 , n70324 , n70325 , n70326 , n70327 , n70328 , n70329 , 
   n70330 , n70331 , n70332 , n70333 , n70334 , n70335 , n70336 , n70337 , n70338 , n70339 , 
   n70340 , n70341 , n70342 , n70343 , n70344 , n70345 , n70346 , n70347 , n70348 , n70349 , 
   n70350 , n70351 , n70352 , n70353 , n70354 , n70355 , n70356 , n70357 , n70358 , n70359 , 
   n70360 , n70361 , n70362 , n70363 , n70364 , n70365 , n70366 , n70367 , n70368 , n70369 , 
   n70370 , n70371 , n70372 , n70373 , n70374 , n70375 , n70376 , n70377 , n70378 , n70379 , 
   n70380 , n70381 , n70382 , n70383 , n70384 , n70385 , n70386 , n70387 , n70388 , n70389 , 
   n70390 , n70391 , n70392 , n70393 , n70394 , n70395 , n70396 , n70397 , n70398 , n70399 , 
   n70400 , n70401 , n70402 , n70403 , n70404 , n70405 , n70406 , n70407 , n70408 , n70409 , 
   n70410 , n70411 , n70412 , n70413 , n70414 , n70415 , n70416 , n70417 , n70418 , n70419 , 
   n70420 , n70421 , n70422 , n70423 , n70424 , n70425 , n70426 , n70427 , n70428 , n70429 , 
   n70430 , n70431 , n70432 , n70433 , n70434 , n70435 , n70436 , n70437 , n70438 , n70439 , 
   n70440 , n70441 , n70442 , n70443 , n70444 , n70445 , n70446 , n70447 , n70448 , n70449 , 
   n70450 , n70451 , n70452 , n70453 , n70454 , n70455 , n70456 , n70457 , n70458 , n70459 , 
   n70460 , n70461 , n70462 , n70463 , n70464 , n70465 , n70466 , n70467 , n70468 , n70469 , 
   n70470 , n70471 , n70472 , n70473 , n70474 , n70475 , n70476 , n70477 , n70478 , n70479 , 
   n70480 , n70481 , n70482 , n70483 , n70484 , n70485 , n70486 , n70487 , n70488 , n70489 , 
   n70490 , n70491 , n70492 , n70493 , n70494 , n70495 , n70496 , n70497 , n70498 , n70499 , 
   n70500 , n70501 , n70502 , n70503 , n70504 , n70505 , n70506 , n70507 , n70508 , n70509 , 
   n70510 , n70511 , n70512 , n70513 , n70514 , n70515 , n70516 , n70517 , n70518 , n70519 , 
   n70520 , n70521 , n70522 , n70523 , n70524 , n70525 , n70526 , n70527 , n70528 , n70529 , 
   n70530 , n70531 , n70532 , n70533 , n70534 , n70535 , n70536 , n70537 , n70538 , n70539 , 
   n70540 , n70541 , n70542 , n70543 , n70544 , n70545 , n70546 , n70547 , n70548 , n70549 , 
   n70550 , n70551 , n70552 , n70553 , n70554 , n70555 , n70556 , n70557 , n70558 , n70559 , 
   n70560 , n70561 , n70562 , n70563 , n70564 , n70565 , n70566 , n70567 , n70568 , n70569 , 
   n70570 , n70571 , n70572 , n70573 , n70574 , n70575 , n70576 , n70577 , n70578 , n70579 , 
   n70580 , n70581 , n70582 , n70583 , n70584 , n70585 , n70586 , n70587 , n70588 , n70589 , 
   n70590 , n70591 , n70592 , n70593 , n70594 , n70595 , n70596 , n70597 , n70598 , n70599 , 
   n70600 , n70601 , n70602 , n70603 , n70604 , n70605 , n70606 , n70607 , n70608 , n70609 , 
   n70610 , n70611 , n70612 , n70613 , n70614 , n70615 , n70616 , n70617 , n70618 , n70619 , 
   n70620 , n70621 , n70622 , n70623 , n70624 , n70625 , n70626 , n70627 , n70628 , n70629 , 
   n70630 , n70631 , n70632 , n70633 , n70634 , n70635 , n70636 , n70637 , n70638 , n70639 , 
   n70640 , n70641 , n70642 , n70643 , n70644 , n70645 , n70646 , n70647 , n70648 , n70649 , 
   n70650 , n70651 , n70652 , n70653 , n70654 , n70655 , n70656 , n70657 , n70658 , n70659 , 
   n70660 , n70661 , n70662 , n70663 , n70664 , n70665 , n70666 , n70667 , n70668 , n70669 , 
   n70670 , n70671 , n70672 , n70673 , n70674 , n70675 , n70676 , n70677 , n70678 , n70679 , 
   n70680 , n70681 , n70682 , n70683 , n70684 , n70685 , n70686 , n70687 , n70688 , n70689 , 
   n70690 , n70691 , n70692 , n70693 , n70694 , n70695 , n70696 , n70697 , n70698 , n70699 , 
   n70700 , n70701 , n70702 , n70703 , n70704 , n70705 , n70706 , n70707 , n70708 , n70709 , 
   n70710 , n70711 , n70712 , n70713 , n70714 , n70715 , n70716 , n70717 , n70718 , n70719 , 
   n70720 , n70721 , n70722 , n70723 , n70724 , n70725 , n70726 , n70727 , n70728 , n70729 , 
   n70730 , n70731 , n70732 , n70733 , n70734 , n70735 , n70736 , n70737 , n70738 , n70739 , 
   n70740 , n70741 , n70742 , n70743 , n70744 , n70745 , n70746 , n70747 , n70748 , n70749 , 
   n70750 , n70751 , n70752 , n70753 , n70754 , n70755 , n70756 , n70757 , n70758 , n70759 , 
   n70760 , n70761 , n70762 , n70763 , n70764 , n70765 , n70766 , n70767 , n70768 , n70769 , 
   n70770 , n70771 , n70772 , n70773 , n70774 , n70775 , n70776 , n70777 , n70778 , n70779 , 
   n70780 , n70781 , n70782 , n70783 , n70784 , n70785 , n70786 , n70787 , n70788 , n70789 , 
   n70790 , n70791 , n70792 , n70793 , n70794 , n70795 , n70796 , n70797 , n70798 , n70799 , 
   n70800 , n70801 , n70802 , n70803 , n70804 , n70805 , n70806 , n70807 , n70808 , n70809 , 
   n70810 , n70811 , n70812 , n70813 , n70814 , n70815 , n70816 , n70817 , n70818 , n70819 , 
   n70820 , n70821 , n70822 , n70823 , n70824 , n70825 , n70826 , n70827 , n70828 , n70829 , 
   n70830 , n70831 , n70832 , n70833 , n70834 , n70835 , n70836 , n70837 , n70838 , n70839 , 
   n70840 , n70841 , n70842 , n70843 , n70844 , n70845 , n70846 , n70847 , n70848 , n70849 , 
   n70850 , n70851 , n70852 , n70853 , n70854 , n70855 , n70856 , n70857 , n70858 , n70859 , 
   n70860 , n70861 , n70862 , n70863 , n70864 , n70865 , n70866 , n70867 , n70868 , n70869 , 
   n70870 , n70871 , n70872 , n70873 , n70874 , n70875 , n70876 , n70877 , n70878 , n70879 , 
   n70880 , n70881 , n70882 , n70883 , n70884 , n70885 , n70886 , n70887 , n70888 , n70889 , 
   n70890 , n70891 , n70892 , n70893 , n70894 , n70895 , n70896 , n70897 , n70898 , n70899 , 
   n70900 , n70901 , n70902 , n70903 , n70904 , n70905 , n70906 , n70907 , n70908 , n4766 , 
   n70910 , n70911 , n70912 , n4770 , n70914 , n70915 , n70916 , n70917 , n70918 , n70919 , 
   n70920 , n70921 , n70922 , n70923 , n70924 , n70925 , n70926 , n70927 , n70928 , n70929 , 
   n70930 , n70931 , n70932 , n70933 , n70934 , n70935 , n70936 , n70937 , n70938 , n70939 , 
   n70940 , n70941 , n70942 , n70943 , n70944 , n70945 , n70946 , n70947 , n70948 , n70949 , 
   n70950 , n70951 , n70952 , n70953 , n70954 , n70955 , n70956 , n70957 , n70958 , n70959 , 
   n70960 , n70961 , n70962 , n70963 , n70964 , n70965 , n70966 , n70967 , n70968 , n70969 , 
   n70970 , n70971 , n70972 , n70973 , n70974 , n70975 , n70976 , n70977 , n70978 , n70979 , 
   n70980 , n70981 , n70982 , n70983 , n70984 , n70985 , n70986 , n70987 , n70988 , n70989 , 
   n70990 , n70991 , n70992 , n70993 , n70994 , n70995 , n70996 , n70997 , n70998 , n70999 , 
   n71000 , n71001 , n71002 , n71003 , n71004 , n71005 , n71006 , n71007 , n71008 , n71009 , 
   n71010 , n71011 , n71012 , n71013 , n71014 , n71015 , n71016 , n71017 , n71018 , n71019 , 
   n71020 , n71021 , n71022 , n71023 , n4881 , n4882 , n71026 , n4884 , n4885 , n71029 , 
   n71030 , n71031 , n71032 , n71033 , n71034 , n71035 , n71036 , n71037 , n71038 , n71039 , 
   n71040 , n71041 , n71042 , n71043 , n71044 , n71045 , n71046 , n71047 , n71048 , n71049 , 
   n71050 , n71051 , n71052 , n71053 , n71054 , n71055 , n71056 , n71057 , n71058 , n71059 , 
   n71060 , n71061 , n71062 , n71063 , n71064 , n71065 , n71066 , n71067 , n71068 , n71069 , 
   n71070 , n71071 , n71072 , n71073 , n71074 , n71075 , n71076 , n71077 , n71078 , n71079 , 
   n71080 , n71081 , n71082 , n71083 , n71084 , n71085 , n71086 , n71087 , n71088 , n71089 , 
   n71090 , n71091 , n71092 , n71093 , n71094 , n71095 , n71096 , n71097 , n71098 , n71099 , 
   n71100 , n71101 , n71102 , n71103 , n71104 , n71105 , n71106 , n71107 , n71108 , n71109 , 
   n71110 , n71111 , n71112 , n71113 , n71114 , n71115 , n71116 , n71117 , n71118 , n71119 , 
   n71120 , n71121 , n71122 , n71123 , n71124 , n71125 , n71126 , n71127 , n71128 , n71129 , 
   n71130 , n71131 , n71132 , n71133 , n71134 , n71135 , n71136 , n71137 , n71138 , n71139 , 
   n71140 , n71141 , n71142 , n71143 , n71144 , n71145 , n71146 , n71147 , n71148 , n71149 , 
   n71150 , n71151 , n71152 , n71153 , n71154 , n71155 , n71156 , n71157 , n71158 , n71159 , 
   n71160 , n71161 , n71162 , n71163 , n71164 , n71165 , n71166 , n71167 , n71168 , n71169 , 
   n71170 , n71171 , n71172 , n71173 , n71174 , n71175 , n71176 , n71177 , n71178 , n71179 , 
   n71180 , n71181 , n71182 , n71183 , n71184 , n71185 , n71186 , n71187 , n71188 , n71189 , 
   n71190 , n71191 , n71192 , n71193 , n71194 , n71195 , n71196 , n71197 , n71198 , n71199 , 
   n71200 , n71201 , n71202 , n71203 , n71204 , n71205 , n71206 , n71207 , n71208 , n71209 , 
   n71210 , n71211 , n71212 , n71213 , n71214 , n5072 , n71216 , n71217 , n5075 , n71219 , 
   n71220 , n71221 , n71222 , n71223 , n71224 , n71225 , n71226 , n71227 , n71228 , n71229 , 
   n71230 , n71231 , n71232 , n71233 , n71234 , n71235 , n71236 , n71237 , n71238 , n71239 , 
   n71240 , n71241 , n71242 , n71243 , n71244 , n71245 , n71246 , n71247 , n71248 , n71249 , 
   n71250 , n71251 , n71252 , n71253 , n71254 , n71255 , n71256 , n71257 , n71258 , n71259 , 
   n71260 , n71261 , n71262 , n71263 , n71264 , n71265 , n71266 , n71267 , n71268 , n71269 , 
   n71270 , n5128 , n5129 , n71273 , n71274 , n71275 , n71276 , n71277 , n71278 , n71279 , 
   n71280 , n71281 , n71282 , n71283 , n71284 , n71285 , n71286 , n71287 , n71288 , n71289 , 
   n71290 , n71291 , n71292 , n71293 , n71294 , n71295 , n71296 , n71297 , n71298 , n71299 , 
   n71300 , n71301 , n71302 , n71303 , n71304 , n71305 , n71306 , n71307 , n71308 , n71309 , 
   n71310 , n71311 , n71312 , n71313 , n71314 , n71315 , n71316 , n71317 , n71318 , n71319 , 
   n71320 , n71321 , n71322 , n71323 , n71324 , n71325 , n71326 , n71327 , n71328 , n71329 , 
   n71330 , n71331 , n71332 , n71333 , n71334 , n71335 , n71336 , n71337 , n71338 , n71339 , 
   n71340 , n71341 , n71342 , n71343 , n71344 , n71345 , n71346 , n71347 , n71348 , n71349 , 
   n71350 , n71351 , n71352 , n71353 , n71354 , n71355 , n71356 , n71357 , n71358 , n71359 , 
   n71360 , n71361 , n71362 , n71363 , n71364 , n71365 , n71366 , n71367 , n71368 , n71369 , 
   n71370 , n71371 , n71372 , n71373 , n71374 , n71375 , n71376 , n71377 , n71378 , n71379 , 
   n71380 , n71381 , n71382 , n71383 , n71384 , n71385 , n71386 , n71387 , n71388 , n71389 , 
   n71390 , n71391 , n71392 , n71393 , n71394 , n71395 , n71396 , n71397 , n71398 , n71399 , 
   n71400 , n71401 , n71402 , n71403 , n71404 , n71405 , n71406 , n71407 , n71408 , n71409 , 
   n71410 , n71411 , n71412 , n71413 , n71414 , n71415 , n71416 , n71417 , n71418 , n71419 , 
   n71420 , n71421 , n71422 , n71423 , n71424 , n71425 , n71426 , n71427 , n71428 , n71429 , 
   n71430 , n71431 , n71432 , n71433 , n71434 , n71435 , n71436 , n71437 , n71438 , n71439 , 
   n71440 , n71441 , n71442 , n5300 , n5301 , n71445 , n71446 , n71447 , n71448 , n71449 , 
   n71450 , n71451 , n71452 , n71453 , n71454 , n71455 , n71456 , n71457 , n71458 , n71459 , 
   n71460 , n71461 , n71462 , n71463 , n71464 , n71465 , n71466 , n71467 , n71468 , n71469 , 
   n71470 , n71471 , n71472 , n71473 , n71474 , n71475 , n71476 , n71477 , n71478 , n71479 , 
   n71480 , n71481 , n71482 , n71483 , n71484 , n71485 , n71486 , n71487 , n71488 , n71489 , 
   n71490 , n71491 , n71492 , n71493 , n71494 , n71495 , n71496 , n71497 , n71498 , n71499 , 
   n71500 , n71501 , n71502 , n71503 , n71504 , n71505 , n71506 , n71507 , n71508 , n71509 , 
   n71510 , n71511 , n71512 , n71513 , n71514 , n71515 , n71516 , n71517 , n71518 , n5376 , 
   n71520 , n71521 , n71522 , n71523 , n71524 , n71525 , n71526 , n71527 , n71528 , n71529 , 
   n71530 , n71531 , n71532 , n71533 , n71534 , n71535 , n71536 , n71537 , n71538 , n71539 , 
   n71540 , n71541 , n71542 , n71543 , n71544 , n71545 , n71546 , n71547 , n71548 , n71549 , 
   n71550 , n71551 , n71552 , n71553 , n71554 , n71555 , n71556 , n71557 , n71558 , n71559 , 
   n71560 , n71561 , n71562 , n71563 , n71564 , n71565 , n71566 , n71567 , n71568 , n71569 , 
   n71570 , n71571 , n71572 , n71573 , n71574 , n71575 , n71576 , n71577 , n71578 , n71579 , 
   n71580 , n71581 , n71582 , n5440 , n71584 , n71585 , n71586 , n71587 , n71588 , n71589 , 
   n71590 , n71591 , n71592 , n71593 , n71594 , n71595 , n71596 , n71597 , n71598 , n71599 , 
   n71600 , n71601 , n71602 , n71603 , n71604 , n71605 , n71606 , n71607 , n71608 , n71609 , 
   n71610 , n71611 , n71612 , n71613 , n71614 , n71615 , n71616 , n71617 , n71618 , n71619 , 
   n71620 , n71621 , n71622 , n71623 , n71624 , n71625 , n71626 , n71627 , n71628 , n71629 , 
   n71630 , n71631 , n71632 , n71633 , n71634 , n71635 , n71636 , n71637 , n71638 , n71639 , 
   n71640 , n71641 , n71642 , n71643 , n71644 , n71645 , n71646 , n71647 , n71648 , n71649 , 
   n71650 , n71651 , n71652 , n71653 , n71654 , n71655 , n71656 , n71657 , n71658 , n71659 , 
   n71660 , n71661 , n71662 , n71663 , n71664 , n71665 , n71666 , n71667 , n71668 , n71669 , 
   n71670 , n71671 , n71672 , n71673 , n71674 , n71675 , n71676 , n71677 , n71678 , n71679 , 
   n71680 , n71681 , n71682 , n71683 , n71684 , n71685 , n71686 , n71687 , n71688 , n71689 , 
   n71690 , n71691 , n71692 , n71693 , n71694 , n71695 , n71696 , n71697 , n71698 , n71699 , 
   n71700 , n71701 , n71702 , n71703 , n71704 , n71705 , n71706 , n71707 , n71708 , n71709 , 
   n71710 , n71711 , n71712 , n71713 , n71714 , n71715 , n71716 , n71717 , n71718 , n71719 , 
   n71720 , n71721 , n71722 , n71723 , n71724 , n5582 , n5583 , n71727 , n71728 , n71729 , 
   n71730 , n71731 , n71732 , n71733 , n71734 , n5592 , n71736 , n71737 , n5595 , n71739 , 
   n71740 , n71741 , n71742 , n71743 , n71744 , n71745 , n5603 , n71747 , n71748 , n71749 , 
   n71750 , n71751 , n71752 , n71753 , n71754 , n71755 , n71756 , n71757 , n71758 , n71759 , 
   n71760 , n71761 , n71762 , n71763 , n71764 , n71765 , n71766 , n71767 , n71768 , n71769 , 
   n71770 , n71771 , n71772 , n71773 , n71774 , n71775 , n71776 , n71777 , n71778 , n71779 , 
   n71780 , n71781 , n71782 , n71783 , n71784 , n71785 , n71786 , n71787 , n5645 , n71789 , 
   n71790 , n71791 , n71792 , n71793 , n71794 , n71795 , n71796 , n71797 , n71798 , n71799 , 
   n71800 , n71801 , n71802 , n71803 , n71804 , n71805 , n5663 , n71807 , n71808 , n5666 , 
   n71810 , n71811 , n71812 , n71813 , n71814 , n71815 , n71816 , n71817 , n71818 , n71819 , 
   n71820 , n71821 , n71822 , n71823 , n71824 , n5682 , n71826 , n71827 , n71828 , n71829 , 
   n71830 , n71831 , n71832 , n71833 , n71834 , n71835 , n71836 , n71837 , n71838 , n71839 , 
   n71840 , n71841 , n71842 , n71843 , n71844 , n5702 , n71846 , n71847 , n71848 , n71849 , 
   n71850 , n71851 , n71852 , n71853 , n71854 , n71855 , n71856 , n71857 , n71858 , n5716 , 
   n71860 , n71861 , n71862 , n71863 , n71864 , n71865 , n71866 , n71867 , n71868 , n71869 , 
   n71870 , n71871 , n71872 , n71873 , n71874 , n71875 , n5733 , n71877 , n71878 , n5736 , 
   n71880 , n71881 , n71882 , n71883 , n71884 , n5742 , n5743 , n71887 , n5745 , n5746 , 
   n71890 , n71891 , n71892 , n71893 , n71894 , n5752 , n71896 , n71897 , n5755 , n71899 , 
   n71900 , n71901 , n71902 , n71903 , n71904 , n71905 , n71906 , n71907 , n71908 , n71909 , 
   n71910 , n71911 , n71912 , n71913 , n71914 , n71915 , n71916 , n71917 , n71918 , n71919 , 
   n71920 , n71921 , n71922 , n71923 , n71924 , n71925 , n71926 , n71927 , n71928 , n71929 , 
   n71930 , n71931 , n71932 , n71933 , n71934 , n71935 , n71936 , n71937 , n71938 , n71939 , 
   n71940 , n71941 , n71942 , n71943 , n71944 , n71945 , n71946 , n71947 , n71948 , n71949 , 
   n71950 , n71951 , n71952 , n71953 , n71954 , n71955 , n71956 , n71957 , n71958 , n71959 , 
   n71960 , n71961 , n71962 , n71963 , n71964 , n71965 , n71966 , n71967 , n71968 , n71969 , 
   n71970 , n71971 , n71972 , n71973 , n71974 , n71975 , n71976 , n71977 , n71978 , n71979 , 
   n71980 , n71981 , n71982 , n71983 , n71984 , n71985 , n71986 , n71987 , n71988 , n71989 , 
   n71990 , n71991 , n71992 , n71993 , n71994 , n71995 , n71996 , n71997 , n71998 , n71999 , 
   n72000 , n72001 , n72002 , n72003 , n72004 , n72005 , n72006 , n72007 , n72008 , n72009 , 
   n72010 , n72011 , n72012 , n72013 , n72014 , n72015 , n72016 , n72017 , n72018 , n72019 , 
   n72020 , n72021 , n72022 , n72023 , n72024 , n72025 , n72026 , n72027 , n72028 , n5886 , 
   n72030 , n72031 , n72032 , n5890 , n72034 , n72035 , n72036 , n72037 , n72038 , n72039 , 
   n72040 , n72041 , n72042 , n72043 , n72044 , n72045 , n72046 , n72047 , n72048 , n72049 , 
   n72050 , n72051 , n72052 , n72053 , n72054 , n72055 , n72056 , n72057 , n72058 , n72059 , 
   n72060 , n72061 , n72062 , n72063 , n72064 , n72065 , n72066 , n72067 , n72068 , n72069 , 
   n72070 , n72071 , n72072 , n72073 , n72074 , n72075 , n72076 , n72077 , n72078 , n72079 , 
   n72080 , n5938 , n72082 , n72083 , n5941 , n72085 , n72086 , n72087 , n72088 , n72089 , 
   n72090 , n72091 , n72092 , n72093 , n72094 , n72095 , n72096 , n72097 , n72098 , n72099 , 
   n72100 , n72101 , n72102 , n72103 , n72104 , n72105 , n72106 , n72107 , n72108 , n72109 , 
   n72110 , n72111 , n72112 , n72113 , n72114 , n72115 , n72116 , n72117 , n72118 , n72119 , 
   n72120 , n72121 , n72122 , n72123 , n72124 , n72125 , n72126 , n72127 , n72128 , n72129 , 
   n72130 , n72131 , n72132 , n72133 , n72134 , n72135 , n72136 , n72137 , n72138 , n72139 , 
   n72140 , n72141 , n72142 , n72143 , n72144 , n72145 , n72146 , n72147 , n72148 , n72149 , 
   n72150 , n72151 , n72152 , n72153 , n72154 , n72155 , n72156 , n72157 , n72158 , n72159 , 
   n6017 , n6018 , n72162 , n72163 , n72164 , n72165 , n72166 , n72167 , n72168 , n72169 , 
   n72170 , n72171 , n72172 , n72173 , n72174 , n72175 , n72176 , n72177 , n72178 , n72179 , 
   n72180 , n72181 , n72182 , n72183 , n72184 , n72185 , n72186 , n72187 , n72188 , n72189 , 
   n72190 , n72191 , n72192 , n72193 , n72194 , n72195 , n72196 , n72197 , n72198 , n72199 , 
   n72200 , n72201 , n72202 , n72203 , n72204 , n72205 , n72206 , n72207 , n72208 , n72209 , 
   n72210 , n72211 , n72212 , n72213 , n72214 , n72215 , n72216 , n72217 , n72218 , n72219 , 
   n6077 , n6078 , n72222 , n72223 , n72224 , n72225 , n72226 , n72227 , n72228 , n72229 , 
   n72230 , n72231 , n72232 , n72233 , n72234 , n72235 , n72236 , n72237 , n72238 , n72239 , 
   n72240 , n72241 , n72242 , n72243 , n72244 , n72245 , n72246 , n72247 , n72248 , n72249 , 
   n72250 , n72251 , n72252 , n72253 , n72254 , n72255 , n72256 , n72257 , n72258 , n72259 , 
   n72260 , n72261 , n72262 , n72263 , n72264 , n72265 , n72266 , n72267 , n72268 , n72269 , 
   n72270 , n72271 , n72272 , n72273 , n72274 , n72275 , n72276 , n72277 , n72278 , n72279 , 
   n6137 , n72281 , n72282 , n72283 , n72284 , n72285 , n72286 , n72287 , n72288 , n72289 , 
   n72290 , n72291 , n72292 , n72293 , n72294 , n72295 , n72296 , n72297 , n72298 , n72299 , 
   n72300 , n72301 , n72302 , n72303 , n72304 , n72305 , n72306 , n72307 , n72308 , n72309 , 
   n72310 , n72311 , n72312 , n72313 , n72314 , n72315 , n72316 , n72317 , n72318 , n72319 , 
   n72320 , n72321 , n72322 , n72323 , n72324 , n72325 , n72326 , n72327 , n6185 , n72329 , 
   n72330 , n72331 , n72332 , n72333 , n72334 , n72335 , n72336 , n72337 , n72338 , n72339 , 
   n72340 , n72341 , n72342 , n72343 , n72344 , n72345 , n72346 , n72347 , n72348 , n72349 , 
   n72350 , n72351 , n72352 , n72353 , n72354 , n72355 , n72356 , n72357 , n72358 , n72359 , 
   n72360 , n72361 , n72362 , n72363 , n72364 , n72365 , n72366 , n72367 , n72368 , n72369 , 
   n72370 , n72371 , n72372 , n72373 , n72374 , n72375 , n72376 , n72377 , n72378 , n72379 , 
   n72380 , n72381 , n72382 , n72383 , n72384 , n72385 , n72386 , n72387 , n72388 , n72389 , 
   n72390 , n72391 , n72392 , n72393 , n72394 , n72395 , n72396 , n72397 , n72398 , n72399 , 
   n72400 , n72401 , n72402 , n72403 , n72404 , n72405 , n72406 , n72407 , n72408 , n72409 , 
   n72410 , n72411 , n72412 , n72413 , n72414 , n72415 , n72416 , n72417 , n72418 , n72419 , 
   n72420 , n72421 , n72422 , n72423 , n72424 , n72425 , n72426 , n72427 , n72428 , n72429 , 
   n72430 , n72431 , n72432 , n72433 , n72434 , n72435 , n72436 , n72437 , n72438 , n72439 , 
   n72440 , n72441 , n72442 , n72443 , n72444 , n72445 , n72446 , n72447 , n72448 , n72449 , 
   n72450 , n72451 , n72452 , n72453 , n72454 , n72455 , n72456 , n72457 , n72458 , n72459 , 
   n72460 , n72461 , n72462 , n72463 , n72464 , n72465 , n72466 , n72467 , n72468 , n72469 , 
   n72470 , n72471 , n72472 , n72473 , n72474 , n72475 , n72476 , n72477 , n72478 , n72479 , 
   n72480 , n72481 , n72482 , n72483 , n72484 , n72485 , n72486 , n72487 , n72488 , n72489 , 
   n72490 , n72491 , n72492 , n72493 , n72494 , n72495 , n72496 , n72497 , n72498 , n72499 , 
   n72500 , n72501 , n72502 , n72503 , n72504 , n72505 , n72506 , n72507 , n72508 , n72509 , 
   n72510 , n72511 , n72512 , n72513 , n72514 , n72515 , n72516 , n72517 , n72518 , n72519 , 
   n72520 , n72521 , n72522 , n72523 , n72524 , n72525 , n72526 , n72527 , n72528 , n72529 , 
   n72530 , n72531 , n72532 , n72533 , n72534 , n72535 , n72536 , n72537 , n72538 , n72539 , 
   n72540 , n72541 , n72542 , n72543 , n72544 , n72545 , n72546 , n72547 , n72548 , n72549 , 
   n72550 , n72551 , n72552 , n72553 , n72554 , n72555 , n72556 , n72557 , n72558 , n72559 , 
   n72560 , n72561 , n72562 , n72563 , n72564 , n72565 , n72566 , n72567 , n72568 , n72569 , 
   n72570 , n72571 , n72572 , n72573 , n72574 , n72575 , n72576 , n72577 , n72578 , n72579 , 
   n72580 , n72581 , n72582 , n72583 , n72584 , n72585 , n72586 , n72587 , n72588 , n72589 , 
   n72590 , n72591 , n72592 , n72593 , n72594 , n72595 , n72596 , n72597 , n72598 , n72599 , 
   n72600 , n72601 , n72602 , n72603 , n72604 , n72605 , n72606 , n72607 , n72608 , n72609 , 
   n72610 , n72611 , n72612 , n72613 , n72614 , n72615 , n72616 , n72617 , n72618 , n72619 , 
   n72620 , n72621 , n72622 , n72623 , n72624 , n72625 , n72626 , n72627 , n72628 , n72629 , 
   n72630 , n72631 , n72632 , n72633 , n72634 , n72635 , n72636 , n72637 , n72638 , n72639 , 
   n72640 , n72641 , n72642 , n72643 , n72644 , n72645 , n72646 , n72647 , n72648 , n72649 , 
   n72650 , n72651 , n72652 , n72653 , n72654 , n72655 , n72656 , n72657 , n72658 , n72659 , 
   n72660 , n72661 , n72662 , n72663 , n72664 , n72665 , n72666 , n72667 , n72668 , n72669 , 
   n72670 , n72671 , n72672 , n72673 , n72674 , n72675 , n72676 , n72677 , n72678 , n72679 , 
   n72680 , n72681 , n72682 , n72683 , n72684 , n72685 , n72686 , n72687 , n72688 , n72689 , 
   n72690 , n72691 , n72692 , n72693 , n72694 , n72695 , n72696 , n72697 , n72698 , n72699 , 
   n72700 , n72701 , n72702 , n72703 , n72704 , n72705 , n72706 , n72707 , n72708 , n72709 , 
   n72710 , n72711 , n72712 , n72713 , n72714 , n72715 , n72716 , n72717 , n72718 , n72719 , 
   n72720 , n72721 , n72722 , n72723 , n72724 , n72725 , n72726 , n72727 , n72728 , n72729 , 
   n72730 , n72731 , n72732 , n72733 , n72734 , n72735 , n72736 , n72737 , n72738 , n72739 , 
   n72740 , n72741 , n72742 , n72743 , n72744 , n72745 , n72746 , n72747 , n72748 , n72749 , 
   n72750 , n72751 , n72752 , n72753 , n72754 , n72755 , n72756 , n72757 , n72758 , n72759 , 
   n72760 , n72761 , n72762 , n72763 , n72764 , n72765 , n72766 , n72767 , n72768 , n72769 , 
   n72770 , n72771 , n72772 , n72773 , n72774 , n72775 , n72776 , n72777 , n72778 , n72779 , 
   n72780 , n72781 , n72782 , n72783 , n72784 , n72785 , n72786 , n72787 , n72788 , n72789 , 
   n72790 , n72791 , n72792 , n72793 , n72794 , n72795 , n72796 , n72797 , n72798 , n72799 , 
   n72800 , n72801 , n72802 , n72803 , n72804 , n72805 , n72806 , n72807 , n72808 , n72809 , 
   n72810 , n72811 , n72812 , n72813 , n72814 , n72815 , n72816 , n72817 , n72818 , n72819 , 
   n72820 , n72821 , n72822 , n72823 , n72824 , n72825 , n72826 , n72827 , n72828 , n72829 , 
   n72830 , n72831 , n72832 , n72833 , n72834 , n72835 , n72836 , n72837 , n72838 , n6696 , 
   n6697 , n72841 , n72842 , n72843 , n72844 , n72845 , n72846 , n72847 , n72848 , n72849 , 
   n72850 , n72851 , n72852 , n72853 , n72854 , n72855 , n72856 , n72857 , n72858 , n72859 , 
   n72860 , n72861 , n72862 , n72863 , n72864 , n72865 , n72866 , n72867 , n72868 , n72869 , 
   n72870 , n72871 , n72872 , n72873 , n72874 , n72875 , n72876 , n72877 , n72878 , n72879 , 
   n72880 , n72881 , n72882 , n72883 , n72884 , n72885 , n72886 , n72887 , n72888 , n72889 , 
   n72890 , n72891 , n72892 , n72893 , n72894 , n72895 , n72896 , n72897 , n72898 , n72899 , 
   n72900 , n72901 , n72902 , n72903 , n72904 , n72905 , n72906 , n72907 , n72908 , n72909 , 
   n72910 , n72911 , n72912 , n72913 , n72914 , n72915 , n72916 , n72917 , n72918 , n72919 , 
   n6777 , n72921 , n72922 , n72923 , n72924 , n72925 , n72926 , n72927 , n72928 , n72929 , 
   n72930 , n72931 , n72932 , n72933 , n72934 , n72935 , n72936 , n72937 , n72938 , n72939 , 
   n72940 , n72941 , n72942 , n72943 , n72944 , n72945 , n72946 , n72947 , n72948 , n72949 , 
   n72950 , n72951 , n72952 , n72953 , n72954 , n72955 , n72956 , n72957 , n72958 , n72959 , 
   n72960 , n72961 , n72962 , n72963 , n72964 , n72965 , n72966 , n72967 , n72968 , n72969 , 
   n72970 , n72971 , n72972 , n72973 , n72974 , n72975 , n72976 , n72977 , n72978 , n72979 , 
   n72980 , n72981 , n72982 , n72983 , n72984 , n72985 , n72986 , n72987 , n72988 , n72989 , 
   n72990 , n72991 , n72992 , n72993 , n72994 , n6852 , n6853 , n72997 , n72998 , n72999 , 
   n73000 , n73001 , n73002 , n73003 , n73004 , n73005 , n73006 , n73007 , n73008 , n73009 , 
   n73010 , n73011 , n73012 , n73013 , n73014 , n73015 , n73016 , n73017 , n73018 , n73019 , 
   n73020 , n73021 , n73022 , n73023 , n73024 , n73025 , n73026 , n73027 , n73028 , n73029 , 
   n73030 , n73031 , n73032 , n73033 , n73034 , n73035 , n73036 , n73037 , n73038 , n73039 , 
   n73040 , n73041 , n73042 , n73043 , n73044 , n73045 , n73046 , n73047 , n73048 , n73049 , 
   n73050 , n73051 , n73052 , n73053 , n73054 , n73055 , n73056 , n73057 , n73058 , n73059 , 
   n73060 , n73061 , n73062 , n73063 , n73064 , n73065 , n73066 , n73067 , n73068 , n73069 , 
   n6927 , n73071 , n73072 , n73073 , n73074 , n73075 , n73076 , n73077 , n73078 , n73079 , 
   n73080 , n73081 , n73082 , n73083 , n73084 , n73085 , n73086 , n73087 , n73088 , n73089 , 
   n73090 , n73091 , n73092 , n73093 , n73094 , n73095 , n73096 , n73097 , n73098 , n73099 , 
   n73100 , n73101 , n73102 , n73103 , n73104 , n73105 , n73106 , n73107 , n73108 , n73109 , 
   n73110 , n73111 , n73112 , n73113 , n73114 , n73115 , n73116 , n73117 , n73118 , n73119 , 
   n73120 , n73121 , n73122 , n73123 , n73124 , n73125 , n73126 , n73127 , n73128 , n73129 , 
   n6987 , n6988 , n73132 , n73133 , n73134 , n73135 , n73136 , n73137 , n73138 , n73139 , 
   n73140 , n73141 , n73142 , n73143 , n73144 , n73145 , n73146 , n73147 , n73148 , n73149 , 
   n73150 , n73151 , n73152 , n73153 , n73154 , n73155 , n73156 , n73157 , n73158 , n73159 , 
   n73160 , n73161 , n73162 , n73163 , n73164 , n73165 , n73166 , n73167 , n73168 , n73169 , 
   n73170 , n73171 , n73172 , n73173 , n73174 , n73175 , n73176 , n73177 , n73178 , n73179 , 
   n73180 , n73181 , n73182 , n73183 , n73184 , n73185 , n73186 , n73187 , n73188 , n73189 , 
   n73190 , n73191 , n73192 , n73193 , n73194 , n73195 , n73196 , n73197 , n73198 , n73199 , 
   n73200 , n73201 , n73202 , n73203 , n73204 , n73205 , n73206 , n73207 , n73208 , n73209 , 
   n73210 , n73211 , n73212 , n73213 , n73214 , n73215 , n73216 , n73217 , n73218 , n73219 , 
   n73220 , n73221 , n73222 , n73223 , n73224 , n73225 , n73226 , n73227 , n73228 , n73229 , 
   n73230 , n73231 , n73232 , n73233 , n73234 , n73235 , n73236 , n73237 , n73238 , n73239 , 
   n73240 , n73241 , n73242 , n73243 , n73244 , n73245 , n73246 , n73247 , n73248 , n73249 , 
   n73250 , n73251 , n73252 , n73253 , n73254 , n73255 , n73256 , n73257 , n73258 , n73259 , 
   n73260 , n73261 , n73262 , n73263 , n73264 , n73265 , n73266 , n73267 , n73268 , n73269 , 
   n73270 , n73271 , n73272 , n73273 , n73274 , n73275 , n73276 , n73277 , n73278 , n73279 , 
   n73280 , n73281 , n7139 , n7140 , n73284 , n73285 , n73286 , n73287 , n73288 , n73289 , 
   n73290 , n73291 , n73292 , n73293 , n73294 , n73295 , n73296 , n73297 , n73298 , n73299 , 
   n73300 , n73301 , n73302 , n73303 , n73304 , n73305 , n73306 , n73307 , n73308 , n73309 , 
   n73310 , n73311 , n73312 , n73313 , n73314 , n73315 , n73316 , n73317 , n73318 , n73319 , 
   n73320 , n73321 , n73322 , n73323 , n73324 , n73325 , n73326 , n73327 , n73328 , n73329 , 
   n73330 , n73331 , n73332 , n73333 , n73334 , n73335 , n73336 , n73337 , n73338 , n73339 , 
   n73340 , n73341 , n73342 , n73343 , n73344 , n73345 , n73346 , n73347 , n73348 , n73349 , 
   n73350 , n7208 , n73352 , n73353 , n73354 , n73355 , n73356 , n73357 , n73358 , n73359 , 
   n73360 , n73361 , n73362 , n73363 , n73364 , n73365 , n73366 , n73367 , n73368 , n73369 , 
   n73370 , n73371 , n73372 , n73373 , n73374 , n73375 , n73376 , n73377 , n73378 , n73379 , 
   n73380 , n73381 , n73382 , n73383 , n73384 , n73385 , n73386 , n73387 , n73388 , n73389 , 
   n73390 , n73391 , n73392 , n73393 , n73394 , n73395 , n73396 , n73397 , n73398 , n73399 , 
   n73400 , n73401 , n73402 , n73403 , n73404 , n73405 , n73406 , n73407 , n73408 , n73409 , 
   n73410 , n73411 , n73412 , n73413 , n73414 , n73415 , n73416 , n73417 , n73418 , n73419 , 
   n73420 , n73421 , n73422 , n73423 , n73424 , n73425 , n73426 , n73427 , n73428 , n73429 , 
   n73430 , n73431 , n73432 , n73433 , n73434 , n73435 , n73436 , n73437 , n73438 , n73439 , 
   n73440 , n73441 , n73442 , n73443 , n73444 , n73445 , n73446 , n73447 , n73448 , n73449 , 
   n73450 , n73451 , n73452 , n73453 , n73454 , n73455 , n73456 , n73457 , n73458 , n73459 , 
   n73460 , n73461 , n73462 , n73463 , n73464 , n73465 , n73466 , n7324 , n73468 , n73469 , 
   n7327 , n7328 , n73472 , n73473 , n73474 , n73475 , n73476 , n73477 , n73478 , n73479 , 
   n73480 , n73481 , n73482 , n73483 , n73484 , n73485 , n73486 , n73487 , n73488 , n7346 , 
   n73490 , n73491 , n73492 , n7350 , n73494 , n73495 , n73496 , n73497 , n73498 , n73499 , 
   n73500 , n73501 , n73502 , n73503 , n73504 , n73505 , n73506 , n73507 , n73508 , n73509 , 
   n73510 , n73511 , n73512 , n73513 , n73514 , n73515 , n73516 , n73517 , n73518 , n73519 , 
   n73520 , n73521 , n73522 , n73523 , n73524 , n73525 , n73526 , n73527 , n73528 , n73529 , 
   n73530 , n7388 , n7389 , n73533 , n73534 , n7392 , n73536 , n73537 , n73538 , n73539 , 
   n73540 , n73541 , n73542 , n73543 , n73544 , n73545 , n73546 , n73547 , n73548 , n73549 , 
   n73550 , n73551 , n73552 , n73553 , n73554 , n73555 , n73556 , n73557 , n73558 , n73559 , 
   n73560 , n73561 , n73562 , n73563 , n73564 , n73565 , n73566 , n73567 , n73568 , n73569 , 
   n73570 , n73571 , n73572 , n73573 , n73574 , n73575 , n73576 , n73577 , n73578 , n73579 , 
   n73580 , n73581 , n73582 , n73583 , n73584 , n73585 , n73586 , n73587 , n73588 , n73589 , 
   n73590 , n73591 , n73592 , n73593 , n73594 , n73595 , n73596 , n73597 , n73598 , n73599 , 
   n73600 , n73601 , n73602 , n73603 , n73604 , n73605 , n73606 , n73607 , n73608 , n73609 , 
   n73610 , n73611 , n73612 , n73613 , n73614 , n73615 , n73616 , n73617 , n73618 , n73619 , 
   n73620 , n73621 , n73622 , n73623 , n73624 , n73625 , n73626 , n73627 , n73628 , n73629 , 
   n73630 , n73631 , n73632 , n73633 , n73634 , n73635 , n73636 , n73637 , n73638 , n73639 , 
   n73640 , n73641 , n73642 , n73643 , n73644 , n73645 , n73646 , n73647 , n73648 , n73649 , 
   n73650 , n73651 , n73652 , n73653 , n73654 , n73655 , n73656 , n73657 , n73658 , n73659 , 
   n73660 , n73661 , n73662 , n73663 , n73664 , n73665 , n73666 , n73667 , n73668 , n73669 , 
   n73670 , n73671 , n73672 , n73673 , n73674 , n73675 , n73676 , n73677 , n73678 , n7536 , 
   n7537 , n73681 , n73682 , n7540 , n73684 , n73685 , n73686 , n73687 , n73688 , n73689 , 
   n73690 , n73691 , n73692 , n73693 , n73694 , n73695 , n73696 , n73697 , n73698 , n73699 , 
   n73700 , n73701 , n73702 , n73703 , n73704 , n73705 , n73706 , n73707 , n73708 , n73709 , 
   n73710 , n73711 , n73712 , n73713 , n73714 , n73715 , n73716 , n73717 , n73718 , n73719 , 
   n73720 , n73721 , n73722 , n73723 , n73724 , n73725 , n73726 , n73727 , n73728 , n73729 , 
   n73730 , n73731 , n73732 , n73733 , n73734 , n73735 , n73736 , n73737 , n73738 , n73739 , 
   n73740 , n73741 , n73742 , n73743 , n73744 , n73745 , n73746 , n73747 , n73748 , n73749 , 
   n73750 , n73751 , n73752 , n73753 , n73754 , n73755 , n73756 , n73757 , n73758 , n73759 , 
   n73760 , n73761 , n7619 , n7620 , n73764 , n73765 , n7623 , n73767 , n73768 , n73769 , 
   n73770 , n73771 , n73772 , n73773 , n73774 , n73775 , n73776 , n73777 , n73778 , n73779 , 
   n73780 , n73781 , n73782 , n73783 , n7641 , n73785 , n73786 , n73787 , n73788 , n73789 , 
   n73790 , n73791 , n73792 , n73793 , n73794 , n73795 , n73796 , n73797 , n73798 , n73799 , 
   n73800 , n73801 , n73802 , n73803 , n73804 , n73805 , n73806 , n73807 , n73808 , n73809 , 
   n73810 , n73811 , n73812 , n73813 , n73814 , n73815 , n73816 , n73817 , n73818 , n7676 , 
   n7677 , n73821 , n73822 , n73823 , n73824 , n73825 , n73826 , n73827 , n73828 , n73829 , 
   n73830 , n73831 , n73832 , n73833 , n73834 , n73835 , n7693 , n73837 , n73838 , n73839 , 
   n73840 , n73841 , n73842 , n73843 , n73844 , n73845 , n73846 , n73847 , n73848 , n73849 , 
   n73850 , n73851 , n73852 , n73853 , n73854 , n73855 , n73856 , n73857 , n73858 , n73859 , 
   n73860 , n73861 , n73862 , n73863 , n73864 , n73865 , n73866 , n73867 , n73868 , n73869 , 
   n73870 , n73871 , n73872 , n73873 , n73874 , n73875 , n73876 , n73877 , n73878 , n73879 , 
   n73880 , n73881 , n73882 , n73883 , n73884 , n73885 , n73886 , n73887 , n73888 , n73889 , 
   n73890 , n73891 , n73892 , n7750 , n73894 , n7752 , n73896 , n73897 , n73898 , n73899 , 
   n73900 , n73901 , n73902 , n73903 , n73904 , n73905 , n73906 , n73907 , n73908 , n73909 , 
   n73910 , n73911 , n73912 , n73913 , n73914 , n73915 , n73916 , n73917 , n73918 , n73919 , 
   n73920 , n73921 , n73922 , n73923 , n73924 , n73925 , n73926 , n73927 , n73928 , n73929 , 
   n73930 , n73931 , n73932 , n73933 , n73934 , n73935 , n73936 , n73937 , n7795 , n73939 , 
   n73940 , n73941 , n73942 , n73943 , n73944 , n73945 , n73946 , n73947 , n73948 , n73949 , 
   n73950 , n73951 , n73952 , n73953 , n73954 , n73955 , n73956 , n73957 , n73958 , n73959 , 
   n73960 , n73961 , n73962 , n73963 , n73964 , n73965 , n73966 , n73967 , n73968 , n73969 , 
   n73970 , n73971 , n73972 , n7830 , n73974 , n7832 , n7833 , n73977 , n73978 , n73979 , 
   n73980 , n73981 , n73982 , n73983 , n73984 , n73985 , n73986 , n73987 , n73988 , n73989 , 
   n73990 , n73991 , n73992 , n73993 , n73994 , n73995 , n73996 , n73997 , n73998 , n73999 , 
   n74000 , n74001 , n74002 , n74003 , n74004 , n74005 , n74006 , n74007 , n74008 , n74009 , 
   n74010 , n74011 , n74012 , n74013 , n74014 , n74015 , n74016 , n74017 , n74018 , n74019 , 
   n74020 , n74021 , n74022 , n74023 , n74024 , n74025 , n74026 , n74027 , n74028 , n74029 , 
   n74030 , n74031 , n74032 , n74033 , n74034 , n74035 , n74036 , n74037 , n74038 , n74039 , 
   n74040 , n74041 , n74042 , n74043 , n74044 , n74045 , n74046 , n74047 , n74048 , n74049 , 
   n74050 , n74051 , n74052 , n74053 , n74054 , n74055 , n74056 , n74057 , n74058 , n74059 , 
   n74060 , n74061 , n74062 , n7920 , n7921 , n74065 , n74066 , n74067 , n74068 , n74069 , 
   n74070 , n74071 , n74072 , n74073 , n74074 , n74075 , n74076 , n74077 , n74078 , n74079 , 
   n7937 , n74081 , n74082 , n74083 , n74084 , n74085 , n74086 , n74087 , n74088 , n74089 , 
   n74090 , n74091 , n74092 , n74093 , n74094 , n74095 , n7953 , n7954 , n74098 , n74099 , 
   n74100 , n74101 , n74102 , n74103 , n74104 , n74105 , n74106 , n74107 , n74108 , n74109 , 
   n74110 , n74111 , n74112 , n74113 , n74114 , n7972 , n74116 , n7974 , n74118 , n74119 , 
   n74120 , n74121 , n74122 , n74123 , n74124 , n74125 , n74126 , n74127 , n74128 , n74129 , 
   n74130 , n74131 , n7989 , n74133 , n74134 , n74135 , n74136 , n74137 , n74138 , n74139 , 
   n74140 , n74141 , n74142 , n74143 , n74144 , n74145 , n74146 , n74147 , n74148 , n74149 , 
   n74150 , n74151 , n74152 , n74153 , n8011 , n74155 , n74156 , n74157 , n74158 , n74159 , 
   n74160 , n74161 , n74162 , n74163 , n74164 , n74165 , n74166 , n74167 , n74168 , n74169 , 
   n8027 , n74171 , n74172 , n74173 , n74174 , n74175 , n74176 , n74177 , n74178 , n74179 , 
   n74180 , n74181 , n74182 , n74183 , n74184 , n74185 , n74186 , n74187 , n74188 , n8046 , 
   n74190 , n8048 , n74192 , n74193 , n74194 , n74195 , n74196 , n74197 , n74198 , n74199 , 
   n74200 , n74201 , n74202 , n74203 , n74204 , n74205 , n74206 , n8064 , n74208 , n74209 , 
   n8067 , n8068 , n74212 , n74213 , n74214 , n74215 , n74216 , n74217 , n74218 , n74219 , 
   n74220 , n74221 , n74222 , n74223 , n74224 , n74225 , n74226 , n74227 , n74228 , n8086 , 
   n74230 , n74231 , n74232 , n74233 , n74234 , n74235 , n74236 , n74237 , n74238 , n74239 , 
   n74240 , n74241 , n74242 , n74243 , n74244 , n74245 , n74246 , n74247 , n74248 , n74249 , 
   n74250 , n74251 , n74252 , n74253 , n74254 , n74255 , n74256 , n74257 , n74258 , n74259 , 
   n74260 , n74261 , n74262 , n74263 , n74264 , n74265 , n74266 , n74267 , n74268 , n8126 , 
   n8127 , n74271 , n74272 , n74273 , n74274 , n74275 , n74276 , n74277 , n74278 , n74279 , 
   n74280 , n74281 , n74282 , n74283 , n74284 , n8142 , n8143 , n74287 , n74288 , n74289 , 
   n74290 , n74291 , n74292 , n74293 , n74294 , n74295 , n74296 , n74297 , n74298 , n74299 , 
   n74300 , n74301 , n74302 , n8160 , n74304 , n74305 , n74306 , n8164 , n74308 , n74309 , 
   n74310 , n74311 , n74312 , n74313 , n74314 , n74315 , n74316 , n74317 , n74318 , n74319 , 
   n74320 , n74321 , n74322 , n74323 , n74324 , n74325 , n74326 , n74327 , n74328 , n74329 , 
   n74330 , n74331 , n74332 , n74333 , n74334 , n74335 , n74336 , n74337 , n74338 , n74339 , 
   n74340 , n74341 , n74342 , n74343 , n8201 , n8202 , n74346 , n74347 , n74348 , n74349 , 
   n74350 , n74351 , n74352 , n74353 , n74354 , n74355 , n74356 , n74357 , n74358 , n74359 , 
   n8217 , n8218 , n74362 , n74363 , n74364 , n74365 , n74366 , n74367 , n74368 , n74369 , 
   n74370 , n74371 , n74372 , n74373 , n74374 , n74375 , n74376 , n74377 , n74378 , n74379 , 
   n74380 , n74381 , n8239 , n74383 , n74384 , n74385 , n74386 , n74387 , n74388 , n74389 , 
   n74390 , n74391 , n74392 , n74393 , n74394 , n74395 , n74396 , n74397 , n74398 , n74399 , 
   n74400 , n74401 , n74402 , n74403 , n74404 , n74405 , n74406 , n74407 , n74408 , n74409 , 
   n74410 , n74411 , n74412 , n74413 , n74414 , n74415 , n74416 , n8274 , n8275 , n74419 , 
   n8277 , n8278 , n74422 , n74423 , n74424 , n74425 , n74426 , n74427 , n74428 , n74429 , 
   n74430 , n74431 , n74432 , n74433 , n74434 , n8292 , n74436 , n74437 , n74438 , n8296 , 
   n74440 , n74441 , n74442 , n74443 , n74444 , n74445 , n74446 , n74447 , n74448 , n74449 , 
   n74450 , n74451 , n74452 , n74453 , n74454 , n74455 , n8313 , n74457 , n74458 , n74459 , 
   n74460 , n74461 , n74462 , n74463 , n74464 , n74465 , n74466 , n74467 , n74468 , n74469 , 
   n74470 , n74471 , n74472 , n74473 , n74474 , n74475 , n74476 , n74477 , n74478 , n74479 , 
   n74480 , n74481 , n74482 , n74483 , n74484 , n74485 , n74486 , n74487 , n74488 , n74489 , 
   n74490 , n74491 , n74492 , n74493 , n74494 , n8352 , n74496 , n74497 , n8355 , n74499 , 
   n74500 , n74501 , n74502 , n74503 , n74504 , n74505 , n74506 , n74507 , n74508 , n74509 , 
   n74510 , n74511 , n74512 , n74513 , n74514 , n74515 , n74516 , n74517 , n74518 , n74519 , 
   n74520 , n74521 , n74522 , n74523 , n74524 , n74525 , n74526 , n74527 , n74528 , n74529 , 
   n74530 , n74531 , n74532 , n74533 , n74534 , n74535 , n74536 , n74537 , n74538 , n74539 , 
   n8397 , n74541 , n74542 , n74543 , n74544 , n74545 , n74546 , n74547 , n74548 , n74549 , 
   n74550 , n74551 , n74552 , n74553 , n74554 , n74555 , n74556 , n74557 , n74558 , n74559 , 
   n8417 , n8418 , n74562 , n74563 , n74564 , n74565 , n74566 , n74567 , n74568 , n8426 , 
   n74570 , n74571 , n8429 , n74573 , n74574 , n74575 , n74576 , n74577 , n74578 , n74579 , 
   n74580 , n8438 , n8439 , n74583 , n74584 , n74585 , n74586 , n74587 , n74588 , n74589 , 
   n74590 , n74591 , n74592 , n74593 , n74594 , n74595 , n74596 , n74597 , n8455 , n8456 , 
   n74600 , n74601 , n74602 , n74603 , n74604 , n74605 , n74606 , n74607 , n74608 , n74609 , 
   n74610 , n74611 , n74612 , n74613 , n74614 , n74615 , n74616 , n74617 , n74618 , n74619 , 
   n74620 , n74621 , n74622 , n74623 , n74624 , n74625 , n74626 , n74627 , n74628 , n74629 , 
   n74630 , n74631 , n74632 , n74633 , n74634 , n74635 , n74636 , n74637 , n74638 , n74639 , 
   n74640 , n74641 , n8499 , n8500 , n74644 , n8502 , n8503 , n74647 , n74648 , n74649 , 
   n74650 , n74651 , n74652 , n74653 , n74654 , n74655 , n74656 , n74657 , n74658 , n74659 , 
   n74660 , n74661 , n8519 , n8520 , n74664 , n74665 , n74666 , n74667 , n74668 , n74669 , 
   n74670 , n74671 , n74672 , n74673 , n74674 , n74675 , n74676 , n74677 , n74678 , n74679 , 
   n74680 , n74681 , n74682 , n8540 , n74684 , n74685 , n74686 , n74687 , n74688 , n74689 , 
   n74690 , n74691 , n74692 , n74693 , n74694 , n74695 , n74696 , n74697 , n74698 , n74699 , 
   n74700 , n74701 , n74702 , n74703 , n74704 , n74705 , n74706 , n74707 , n74708 , n74709 , 
   n74710 , n74711 , n74712 , n74713 , n74714 , n74715 , n74716 , n74717 , n74718 , n74719 , 
   n74720 , n74721 , n74722 , n74723 , n74724 , n8582 , n74726 , n74727 , n74728 , n74729 , 
   n74730 , n74731 , n74732 , n74733 , n74734 , n74735 , n74736 , n74737 , n74738 , n74739 , 
   n74740 , n74741 , n74742 , n74743 , n74744 , n74745 , n8603 , n74747 , n74748 , n74749 , 
   n74750 , n74751 , n74752 , n74753 , n74754 , n74755 , n74756 , n74757 , n74758 , n74759 , 
   n74760 , n74761 , n8619 , n8620 , n74764 , n74765 , n74766 , n74767 , n74768 , n74769 , 
   n74770 , n74771 , n74772 , n74773 , n74774 , n74775 , n74776 , n74777 , n74778 , n74779 , 
   n74780 , n74781 , n8639 , n8640 , n74784 , n74785 , n74786 , n74787 , n74788 , n74789 , 
   n74790 , n74791 , n74792 , n74793 , n74794 , n74795 , n74796 , n74797 , n74798 , n74799 , 
   n74800 , n74801 , n74802 , n74803 , n8661 , n8662 , n74806 , n74807 , n74808 , n74809 , 
   n74810 , n74811 , n74812 , n74813 , n74814 , n74815 , n74816 , n74817 , n74818 , n74819 , 
   n74820 , n74821 , n74822 , n74823 , n74824 , n74825 , n8683 , n74827 , n74828 , n74829 , 
   n74830 , n74831 , n74832 , n74833 , n74834 , n74835 , n74836 , n74837 , n74838 , n74839 , 
   n74840 , n74841 , n74842 , n74843 , n74844 , n74845 , n74846 , n74847 , n74848 , n74849 , 
   n74850 , n74851 , n74852 , n74853 , n74854 , n74855 , n74856 , n74857 , n74858 , n74859 , 
   n74860 , n74861 , n74862 , n74863 , n8721 , n8722 , n74866 , n8724 , n8725 , n74869 , 
   n74870 , n74871 , n74872 , n74873 , n74874 , n74875 , n8733 , n74877 , n8735 , n8736 , 
   n74880 , n74881 , n74882 , n8740 , n8741 , n74885 , n8743 , n74887 , n74888 , n74889 , 
   n74890 , n74891 , n74892 , n74893 , n8751 , n8752 , n74896 , n74897 , n74898 , n8756 , 
   n8757 , n74901 , n74902 , n74903 , n74904 , n74905 , n74906 , n74907 , n74908 , n74909 , 
   n8767 , n8768 , n74912 , n74913 , n74914 , n74915 , n74916 , n74917 , n74918 , n74919 , 
   n74920 , n74921 , n74922 , n74923 , n74924 , n74925 , n74926 , n74927 , n74928 , n74929 , 
   n74930 , n74931 , n74932 , n74933 , n74934 , n74935 , n8793 , n8794 , n74938 , n74939 , 
   n74940 , n8798 , n8799 , n74943 , n74944 , n74945 , n74946 , n74947 , n74948 , n74949 , 
   n8807 , n74951 , n8809 , n8810 , n74954 , n74955 , n74956 , n8814 , n8815 , n74959 , 
   n8817 , n74961 , n74962 , n74963 , n74964 , n74965 , n74966 , n74967 , n8825 , n8826 , 
   n74970 , n74971 , n74972 , n74973 , n74974 , n74975 , n74976 , n74977 , n74978 , n8836 , 
   n74980 , n74981 , n74982 , n74983 , n8841 , n74985 , n74986 , n74987 , n74988 , n74989 , 
   n74990 , n74991 , n74992 , n74993 , n74994 , n74995 , n74996 , n74997 , n74998 , n74999 , 
   n75000 , n75001 , n75002 , n8860 , n75004 , n75005 , n75006 , n75007 , n75008 , n75009 , 
   n8867 , n8868 , n75012 , n75013 , n75014 , n8872 , n8873 , n75017 , n75018 , n75019 , 
   n75020 , n75021 , n75022 , n75023 , n8881 , n75025 , n8883 , n8884 , n75028 , n75029 , 
   n75030 , n8888 , n8889 , n75033 , n8891 , n75035 , n75036 , n75037 , n75038 , n75039 , 
   n75040 , n75041 , n8899 , n8900 , n75044 , n75045 , n75046 , n8904 , n8905 , n75049 , 
   n75050 , n75051 , n75052 , n75053 , n75054 , n75055 , n75056 , n75057 , n8915 , n8916 , 
   n75060 , n75061 , n75062 , n75063 , n75064 , n75065 , n75066 , n75067 , n75068 , n75069 , 
   n75070 , n75071 , n75072 , n75073 , n75074 , n75075 , n75076 , n75077 , n75078 , n8936 , 
   n75080 , n75081 , n75082 , n8940 , n75084 , n75085 , n75086 , n8944 , n75088 , n75089 , 
   n8947 , n75091 , n75092 , n75093 , n75094 , n8952 , n75096 , n75097 , n8955 , n8956 , 
   n75100 , n75101 , n75102 , n75103 , n75104 , n75105 , n8963 , n8964 , n75108 , n75109 , 
   n75110 , n75111 , n75112 , n75113 , n75114 , n75115 , n75116 , n75117 , n75118 , n75119 , 
   n75120 , n75121 , n8979 , n75123 , n75124 , n75125 , n75126 , n8984 , n8985 , n75129 , 
   n75130 , n75131 , n75132 , n75133 , n75134 , n75135 , n75136 , n75137 , n75138 , n75139 , 
   n75140 , n75141 , n75142 , n75143 , n75144 , n75145 , n75146 , n75147 , n75148 , n75149 , 
   n75150 , n75151 , n75152 , n75153 , n75154 , n75155 , n75156 , n9014 , n9015 , n75159 , 
   n75160 , n75161 , n75162 , n9020 , n9021 , n75165 , n75166 , n75167 , n75168 , n75169 , 
   n75170 , n75171 , n9029 , n9030 , n75174 , n9032 , n75176 , n75177 , n75178 , n75179 , 
   n75180 , n75181 , n75182 , n75183 , n75184 , n75185 , n75186 , n75187 , n75188 , n75189 , 
   n75190 , n75191 , n75192 , n75193 , n75194 , n9052 , n9053 , n75197 , n75198 , n75199 , 
   n75200 , n75201 , n75202 , n75203 , n75204 , n75205 , n75206 , n9064 , n75208 , n75209 , 
   n75210 , n75211 , n75212 , n75213 , n75214 , n75215 , n75216 , n75217 , n75218 , n75219 , 
   n75220 , n75221 , n75222 , n75223 , n75224 , n9082 , n9083 , n75227 , n75228 , n75229 , 
   n75230 , n75231 , n75232 , n75233 , n9091 , n9092 , n75236 , n75237 , n75238 , n75239 , 
   n75240 , n75241 , n75242 , n75243 , n75244 , n75245 , n75246 , n75247 , n75248 , n75249 , 
   n75250 , n75251 , n75252 , n75253 , n75254 , n75255 , n75256 , n75257 , n75258 , n75259 , 
   n75260 , n75261 , n75262 , n75263 , n75264 , n75265 , n75266 , n75267 , n9125 , n9126 , 
   n75270 , n75271 , n75272 , n75273 , n75274 , n75275 , n75276 , n75277 , n75278 , n75279 , 
   n75280 , n75281 , n75282 , n75283 , n75284 , n75285 , n75286 , n75287 , n75288 , n75289 , 
   n75290 , n75291 , n75292 , n75293 , n75294 , n75295 , n75296 , n75297 , n75298 , n75299 , 
   n75300 , n75301 , n75302 , n75303 , n75304 , n75305 , n75306 , n75307 , n75308 , n75309 , 
   n75310 , n75311 , n75312 , n75313 , n75314 , n75315 , n75316 , n75317 , n75318 , n75319 , 
   n75320 , n75321 , n75322 , n75323 , n75324 , n75325 , n75326 , n75327 , n75328 , n75329 , 
   n75330 , n75331 , n75332 , n75333 , n75334 , n75335 , n75336 , n75337 , n75338 , n75339 , 
   n75340 , n75341 , n75342 , n75343 , n75344 , n75345 , n75346 , n75347 , n75348 , n75349 , 
   n75350 , n75351 , n75352 , n75353 , n75354 , n75355 , n75356 , n75357 , n75358 , n75359 , 
   n75360 , n75361 , n75362 , n75363 , n75364 , n75365 , n75366 , n75367 , n75368 , n75369 , 
   n75370 , n75371 , n75372 , n75373 , n75374 , n75375 , n75376 , n75377 , n75378 , n75379 , 
   n75380 , n75381 , n75382 , n75383 , n75384 , n75385 , n75386 , n75387 , n75388 , n75389 , 
   n75390 , n75391 , n75392 , n75393 , n75394 , n75395 , n75396 , n75397 , n75398 , n75399 , 
   n75400 , n9258 , n9259 , n75403 , n75404 , n75405 , n75406 , n75407 , n75408 , n75409 , 
   n75410 , n75411 , n75412 , n75413 , n75414 , n75415 , n75416 , n75417 , n75418 , n75419 , 
   n75420 , n75421 , n75422 , n75423 , n75424 , n75425 , n75426 , n9284 , n75428 , n75429 , 
   n75430 , n75431 , n75432 , n75433 , n75434 , n75435 , n75436 , n75437 , n75438 , n75439 , 
   n75440 , n75441 , n75442 , n75443 , n75444 , n75445 , n75446 , n75447 , n75448 , n75449 , 
   n75450 , n75451 , n75452 , n75453 , n75454 , n75455 , n75456 , n75457 , n75458 , n75459 , 
   n9317 , n9318 , n75462 , n75463 , n75464 , n75465 , n75466 , n75467 , n75468 , n75469 , 
   n75470 , n75471 , n75472 , n75473 , n75474 , n75475 , n75476 , n75477 , n75478 , n75479 , 
   n75480 , n75481 , n75482 , n75483 , n75484 , n75485 , n75486 , n75487 , n75488 , n75489 , 
   n75490 , n75491 , n75492 , n75493 , n75494 , n75495 , n75496 , n75497 , n75498 , n75499 , 
   n75500 , n75501 , n75502 , n75503 , n75504 , n75505 , n75506 , n75507 , n75508 , n75509 , 
   n75510 , n75511 , n75512 , n75513 , n75514 , n75515 , n75516 , n75517 , n75518 , n75519 , 
   n75520 , n75521 , n75522 , n75523 , n75524 , n75525 , n75526 , n75527 , n75528 , n75529 , 
   n75530 , n75531 , n75532 , n75533 , n75534 , n75535 , n75536 , n75537 , n75538 , n75539 , 
   n75540 , n75541 , n75542 , n75543 , n75544 , n75545 , n75546 , n75547 , n75548 , n75549 , 
   n75550 , n75551 , n75552 , n75553 , n75554 , n75555 , n75556 , n75557 , n75558 , n75559 , 
   n75560 , n75561 , n75562 , n75563 , n75564 , n75565 , n75566 , n75567 , n75568 , n75569 , 
   n75570 , n75571 , n75572 , n75573 , n75574 , n75575 , n75576 , n75577 , n75578 , n75579 , 
   n75580 , n75581 , n75582 , n75583 , n75584 , n75585 , n75586 , n75587 , n75588 , n75589 , 
   n75590 , n75591 , n75592 , n75593 , n75594 , n75595 , n75596 , n75597 , n75598 , n75599 , 
   n75600 , n75601 , n75602 , n75603 , n75604 , n75605 , n75606 , n75607 , n75608 , n75609 , 
   n75610 , n75611 , n75612 , n75613 , n75614 , n75615 , n75616 , n75617 , n75618 , n75619 , 
   n75620 , n75621 , n75622 , n75623 , n75624 , n75625 , n75626 , n9484 , n75628 , n75629 , 
   n75630 , n9488 , n75632 , n75633 , n75634 , n75635 , n75636 , n75637 , n75638 , n75639 , 
   n75640 , n75641 , n75642 , n75643 , n75644 , n75645 , n75646 , n75647 , n75648 , n75649 , 
   n75650 , n75651 , n75652 , n75653 , n75654 , n75655 , n75656 , n75657 , n75658 , n75659 , 
   n75660 , n75661 , n75662 , n75663 , n75664 , n75665 , n75666 , n75667 , n75668 , n75669 , 
   n75670 , n75671 , n75672 , n75673 , n75674 , n75675 , n75676 , n75677 , n75678 , n75679 , 
   n75680 , n75681 , n75682 , n75683 , n75684 , n75685 , n75686 , n75687 , n75688 , n75689 , 
   n75690 , n75691 , n75692 , n75693 , n75694 , n75695 , n75696 , n75697 , n75698 , n75699 , 
   n75700 , n75701 , n75702 , n75703 , n75704 , n75705 , n75706 , n75707 , n75708 , n75709 , 
   n75710 , n75711 , n75712 , n75713 , n75714 , n75715 , n75716 , n75717 , n75718 , n75719 , 
   n75720 , n75721 , n75722 , n75723 , n75724 , n75725 , n75726 , n75727 , n75728 , n75729 , 
   n75730 , n75731 , n75732 , n75733 , n75734 , n75735 , n75736 , n75737 , n75738 , n75739 , 
   n75740 , n75741 , n75742 , n75743 , n75744 , n75745 , n75746 , n75747 , n75748 , n75749 , 
   n75750 , n75751 , n75752 , n75753 , n75754 , n75755 , n75756 , n75757 , n75758 , n75759 , 
   n75760 , n75761 , n75762 , n9620 , n75764 , n9622 , n9623 , n75767 , n75768 , n75769 , 
   n75770 , n75771 , n75772 , n75773 , n75774 , n75775 , n75776 , n75777 , n75778 , n75779 , 
   n75780 , n75781 , n75782 , n75783 , n75784 , n75785 , n75786 , n75787 , n75788 , n75789 , 
   n75790 , n75791 , n75792 , n75793 , n75794 , n75795 , n75796 , n75797 , n75798 , n9656 , 
   n9657 , n75801 , n75802 , n75803 , n75804 , n75805 , n75806 , n75807 , n75808 , n75809 , 
   n75810 , n75811 , n75812 , n75813 , n75814 , n75815 , n75816 , n75817 , n75818 , n75819 , 
   n75820 , n75821 , n75822 , n75823 , n75824 , n75825 , n75826 , n75827 , n75828 , n75829 , 
   n75830 , n75831 , n9689 , n9690 , n75834 , n75835 , n75836 , n75837 , n75838 , n75839 , 
   n75840 , n75841 , n75842 , n75843 , n75844 , n75845 , n75846 , n75847 , n75848 , n75849 , 
   n75850 , n75851 , n75852 , n75853 , n75854 , n75855 , n75856 , n75857 , n75858 , n75859 , 
   n75860 , n75861 , n75862 , n9720 , n9721 , n75865 , n9723 , n75867 , n75868 , n75869 , 
   n75870 , n75871 , n75872 , n75873 , n75874 , n75875 , n75876 , n75877 , n75878 , n75879 , 
   n75880 , n75881 , n75882 , n75883 , n75884 , n75885 , n75886 , n75887 , n75888 , n75889 , 
   n75890 , n75891 , n75892 , n75893 , n75894 , n75895 , n75896 , n75897 , n75898 , n75899 , 
   n75900 , n75901 , n75902 , n75903 , n75904 , n75905 , n75906 , n75907 , n75908 , n75909 , 
   n75910 , n75911 , n75912 , n75913 , n75914 , n75915 , n75916 , n75917 , n75918 , n75919 , 
   n75920 , n75921 , n75922 , n75923 , n75924 , n75925 , n75926 , n75927 , n75928 , n75929 , 
   n75930 , n75931 , n75932 , n75933 , n75934 , n75935 , n75936 , n75937 , n75938 , n75939 , 
   n75940 , n75941 , n75942 , n75943 , n75944 , n75945 , n75946 , n75947 , n75948 , n75949 , 
   n75950 , n75951 , n75952 , n75953 , n75954 , n75955 , n75956 , n75957 , n75958 , n75959 , 
   n75960 , n75961 , n75962 , n75963 , n75964 , n75965 , n75966 , n75967 , n75968 , n75969 , 
   n75970 , n75971 , n75972 , n75973 , n75974 , n75975 , n75976 , n75977 , n75978 , n75979 , 
   n75980 , n75981 , n75982 , n75983 , n75984 , n75985 , n75986 , n75987 , n75988 , n75989 , 
   n75990 , n75991 , n75992 , n75993 , n75994 , n75995 , n75996 , n75997 , n75998 , n75999 , 
   n76000 , n76001 , n76002 , n76003 , n76004 , n76005 , n76006 , n76007 , n76008 , n76009 , 
   n76010 , n76011 , n76012 , n76013 , n76014 , n76015 , n76016 , n76017 , n76018 , n76019 , 
   n76020 , n76021 , n76022 , n76023 , n76024 , n76025 , n76026 , n76027 , n76028 , n76029 , 
   n76030 , n76031 , n76032 , n76033 , n76034 , n76035 , n76036 , n76037 , n76038 , n76039 , 
   n76040 , n76041 , n76042 , n76043 , n76044 , n76045 , n76046 , n76047 , n76048 , n76049 , 
   n76050 , n76051 , n76052 , n76053 , n76054 , n76055 , n76056 , n76057 , n76058 , n76059 , 
   n76060 , n76061 , n76062 , n76063 , n76064 , n76065 , n76066 , n76067 , n76068 , n76069 , 
   n76070 , n76071 , n76072 , n76073 , n76074 , n76075 , n76076 , n76077 , n76078 , n76079 , 
   n76080 , n76081 , n76082 , n76083 , n76084 , n76085 , n76086 , n9944 , n76088 , n76089 , 
   n76090 , n76091 , n76092 , n9950 , n76094 , n9952 , n9953 , n76097 , n76098 , n76099 , 
   n76100 , n76101 , n76102 , n76103 , n76104 , n76105 , n76106 , n76107 , n76108 , n76109 , 
   n76110 , n76111 , n76112 , n76113 , n76114 , n76115 , n76116 , n76117 , n76118 , n76119 , 
   n76120 , n76121 , n9979 , n76123 , n76124 , n76125 , n9983 , n76127 , n76128 , n76129 , 
   n76130 , n76131 , n76132 , n76133 , n76134 , n76135 , n76136 , n76137 , n76138 , n76139 , 
   n76140 , n76141 , n76142 , n76143 , n76144 , n76145 , n76146 , n76147 , n76148 , n76149 , 
   n76150 , n76151 , n76152 , n10010 , n76154 , n10012 , n76156 , n76157 , n76158 , n76159 , 
   n76160 , n10018 , n10019 , n76163 , n76164 , n76165 , n76166 , n76167 , n76168 , n76169 , 
   n76170 , n76171 , n76172 , n76173 , n76174 , n76175 , n76176 , n76177 , n76178 , n76179 , 
   n76180 , n76181 , n76182 , n76183 , n76184 , n76185 , n76186 , n76187 , n76188 , n76189 , 
   n76190 , n76191 , n10049 , n10050 , n76194 , n76195 , n76196 , n76197 , n76198 , n76199 , 
   n76200 , n76201 , n10059 , n10060 , n76204 , n76205 , n76206 , n76207 , n76208 , n76209 , 
   n10067 , n76211 , n10069 , n10070 , n76214 , n76215 , n76216 , n76217 , n76218 , n10076 , 
   n76220 , n76221 , n76222 , n76223 , n76224 , n76225 , n76226 , n76227 , n76228 , n76229 , 
   n76230 , n76231 , n10089 , n10090 , n76234 , n76235 , n76236 , n76237 , n76238 , n10096 , 
   n76240 , n76241 , n76242 , n10100 , n76244 , n76245 , n76246 , n76247 , n76248 , n76249 , 
   n76250 , n76251 , n76252 , n76253 , n76254 , n76255 , n76256 , n76257 , n76258 , n76259 , 
   n76260 , n76261 , n10119 , n10120 , n76264 , n76265 , n76266 , n76267 , n76268 , n10126 , 
   n10127 , n76271 , n10129 , n10130 , n76274 , n76275 , n76276 , n76277 , n76278 , n76279 , 
   n10137 , n76281 , n10139 , n76283 , n76284 , n76285 , n76286 , n76287 , n76288 , n76289 , 
   n76290 , n76291 , n76292 , n76293 , n76294 , n76295 , n76296 , n76297 , n76298 , n10156 , 
   n10157 , n76301 , n76302 , n76303 , n76304 , n76305 , n76306 , n76307 , n76308 , n76309 , 
   n76310 , n76311 , n76312 , n76313 , n76314 , n76315 , n76316 , n76317 , n76318 , n76319 , 
   n76320 , n76321 , n76322 , n76323 , n76324 , n76325 , n76326 , n76327 , n76328 , n76329 , 
   n76330 , n76331 , n76332 , n10190 , n10191 , n76335 , n76336 , n76337 , n76338 , n10196 , 
   n10197 , n76341 , n10199 , n76343 , n76344 , n76345 , n76346 , n76347 , n76348 , n76349 , 
   n76350 , n76351 , n76352 , n76353 , n76354 , n76355 , n76356 , n76357 , n76358 , n76359 , 
   n76360 , n76361 , n76362 , n76363 , n76364 , n76365 , n76366 , n10224 , n76368 , n10226 , 
   n76370 , n76371 , n76372 , n76373 , n76374 , n10232 , n10233 , n76377 , n76378 , n76379 , 
   n76380 , n76381 , n76382 , n76383 , n76384 , n76385 , n76386 , n76387 , n76388 , n76389 , 
   n76390 , n76391 , n76392 , n76393 , n76394 , n76395 , n76396 , n76397 , n76398 , n76399 , 
   n76400 , n76401 , n76402 , n76403 , n76404 , n76405 , n76406 , n76407 , n76408 , n76409 , 
   n76410 , n76411 , n76412 , n76413 , n76414 , n76415 , n76416 , n76417 , n76418 , n76419 , 
   n76420 , n76421 , n76422 , n76423 , n76424 , n76425 , n76426 , n76427 , n76428 , n76429 , 
   n76430 , n76431 , n76432 , n76433 , n76434 , n76435 , n76436 , n76437 , n76438 , n76439 , 
   n76440 , n76441 , n76442 , n76443 , n76444 , n76445 , n76446 , n76447 , n76448 , n76449 , 
   n76450 , n76451 , n76452 , n76453 , n76454 , n76455 , n76456 , n76457 , n76458 , n76459 , 
   n76460 , n76461 , n76462 , n76463 , n76464 , n76465 , n76466 , n76467 , n76468 , n76469 , 
   n76470 , n76471 , n76472 , n76473 , n76474 , n76475 , n76476 , n76477 , n76478 , n76479 , 
   n76480 , n76481 , n76482 , n76483 , n76484 , n76485 , n76486 , n76487 , n76488 , n76489 , 
   n76490 , n76491 , n76492 , n76493 , n76494 , n76495 , n76496 , n76497 , n76498 , n76499 , 
   n76500 , n76501 , n76502 , n76503 , n76504 , n76505 , n76506 , n76507 , n76508 , n76509 , 
   n76510 , n76511 , n76512 , n76513 , n76514 , n76515 , n76516 , n76517 , n76518 , n76519 , 
   n76520 , n76521 , n76522 , n76523 , n76524 , n76525 , n76526 , n76527 , n76528 , n76529 , 
   n76530 , n76531 , n76532 , n76533 , n76534 , n76535 , n76536 , n76537 , n76538 , n76539 , 
   n76540 , n76541 , n76542 , n76543 , n76544 , n76545 , n76546 , n76547 , n76548 , n76549 , 
   n76550 , n76551 , n76552 , n76553 , n76554 , n76555 , n76556 , n76557 , n76558 , n76559 , 
   n76560 , n76561 , n76562 , n76563 , n76564 , n76565 , n76566 , n76567 , n76568 , n76569 , 
   n76570 , n76571 , n76572 , n76573 , n76574 , n76575 , n76576 , n76577 , n76578 , n76579 , 
   n76580 , n76581 , n76582 , n76583 , n76584 , n76585 , n76586 , n76587 , n76588 , n76589 , 
   n76590 , n76591 , n76592 , n76593 , n76594 , n76595 , n76596 , n76597 , n76598 , n76599 , 
   n76600 , n76601 , n76602 , n76603 , n76604 , n76605 , n76606 , n76607 , n76608 , n76609 , 
   n76610 , n76611 , n76612 , n76613 , n76614 , n76615 , n76616 , n76617 , n76618 , n76619 , 
   n76620 , n76621 , n76622 , n76623 , n76624 , n76625 , n76626 , n76627 , n76628 , n76629 , 
   n76630 , n76631 , n76632 , n76633 , n76634 , n76635 , n76636 , n76637 , n76638 , n76639 , 
   n76640 , n76641 , n76642 , n76643 , n76644 , n76645 , n76646 , n76647 , n76648 , n76649 , 
   n76650 , n76651 , n76652 , n76653 , n76654 , n76655 , n76656 , n76657 , n76658 , n76659 , 
   n76660 , n76661 , n76662 , n76663 , n76664 , n76665 , n76666 , n76667 , n76668 , n76669 , 
   n76670 , n76671 , n76672 , n76673 , n76674 , n76675 , n76676 , n76677 , n76678 , n76679 , 
   n76680 , n76681 , n76682 , n76683 , n76684 , n76685 , n76686 , n76687 , n76688 , n76689 , 
   n76690 , n76691 , n76692 , n76693 , n76694 , n76695 , n76696 , n76697 , n76698 , n76699 , 
   n76700 , n76701 , n76702 , n76703 , n76704 , n76705 , n76706 , n76707 , n76708 , n76709 , 
   n76710 , n76711 , n76712 , n76713 , n76714 , n76715 , n76716 , n76717 , n76718 , n76719 , 
   n76720 , n76721 , n76722 , n76723 , n76724 , n76725 , n76726 , n76727 , n76728 , n76729 , 
   n76730 , n76731 , n76732 , n76733 , n76734 , n76735 , n76736 , n76737 , n76738 , n76739 , 
   n76740 , n76741 , n76742 , n76743 , n76744 , n76745 , n76746 , n76747 , n76748 , n76749 , 
   n76750 , n76751 , n76752 , n76753 , n76754 , n76755 , n76756 , n76757 , n76758 , n76759 , 
   n76760 , n76761 , n76762 , n76763 , n76764 , n76765 , n76766 , n76767 , n76768 , n76769 , 
   n76770 , n76771 , n76772 , n76773 , n76774 , n76775 , n76776 , n76777 , n76778 , n76779 , 
   n76780 , n76781 , n76782 , n76783 , n76784 , n76785 , n76786 , n76787 , n76788 , n76789 , 
   n76790 , n76791 , n76792 , n76793 , n76794 , n76795 , n76796 , n76797 , n76798 , n76799 , 
   n76800 , n76801 , n76802 , n76803 , n76804 , n76805 , n76806 , n76807 , n76808 , n76809 , 
   n76810 , n76811 , n76812 , n76813 , n76814 , n76815 , n76816 , n76817 , n76818 , n76819 , 
   n76820 , n76821 , n76822 , n76823 , n76824 , n76825 , n76826 , n76827 , n76828 , n76829 , 
   n76830 , n76831 , n76832 , n76833 , n76834 , n76835 , n76836 , n76837 , n76838 , n76839 , 
   n76840 , n76841 , n76842 , n76843 , n76844 , n76845 , n76846 , n76847 , n76848 , n76849 , 
   n76850 , n76851 , n76852 , n76853 , n76854 , n76855 , n76856 , n76857 , n76858 , n76859 , 
   n76860 , n76861 , n76862 , n76863 , n76864 , n76865 , n76866 , n76867 , n76868 , n76869 , 
   n76870 , n76871 , n76872 , n76873 , n76874 , n76875 , n76876 , n76877 , n76878 , n76879 , 
   n76880 , n76881 , n76882 , n76883 , n76884 , n76885 , n76886 , n76887 , n76888 , n76889 , 
   n76890 , n76891 , n76892 , n76893 , n76894 , n76895 , n76896 , n76897 , n76898 , n76899 , 
   n76900 , n76901 , n76902 , n76903 , n76904 , n76905 , n76906 , n76907 , n76908 , n76909 , 
   n76910 , n76911 , n76912 , n76913 , n76914 , n76915 , n76916 , n76917 , n76918 , n76919 , 
   n76920 , n76921 , n76922 , n76923 , n76924 , n76925 , n76926 , n76927 , n76928 , n76929 , 
   n76930 , n76931 , n76932 , n76933 , n76934 , n76935 , n76936 , n76937 , n76938 , n76939 , 
   n76940 , n76941 , n76942 , n76943 , n76944 , n76945 , n76946 , n76947 , n76948 , n76949 , 
   n76950 , n76951 , n76952 , n76953 , n76954 , n76955 , n76956 , n76957 , n76958 , n76959 , 
   n76960 , n76961 , n76962 , n76963 , n76964 , n76965 , n76966 , n76967 , n76968 , n76969 , 
   n76970 , n76971 , n76972 , n76973 , n76974 , n76975 , n76976 , n76977 , n76978 , n76979 , 
   n76980 , n76981 , n76982 , n76983 , n76984 , n76985 , n76986 , n76987 , n76988 , n76989 , 
   n76990 , n76991 , n76992 , n76993 , n76994 , n76995 , n76996 , n76997 , n76998 , n76999 , 
   n77000 , n77001 , n77002 , n77003 , n77004 , n77005 , n77006 , n77007 , n77008 , n77009 , 
   n77010 , n77011 , n77012 , n77013 , n77014 , n77015 , n77016 , n77017 , n77018 , n77019 , 
   n77020 , n77021 , n77022 , n77023 , n77024 , n77025 , n77026 , n77027 , n77028 , n77029 , 
   n77030 , n77031 , n77032 , n77033 , n77034 , n77035 , n77036 , n77037 , n77038 , n77039 , 
   n77040 , n77041 , n77042 , n77043 , n77044 , n77045 , n77046 , n77047 , n77048 , n77049 , 
   n77050 , n77051 , n77052 , n77053 , n77054 , n77055 , n77056 , n77057 , n77058 , n77059 , 
   n77060 , n77061 , n77062 , n77063 , n77064 , n77065 , n77066 , n77067 , n77068 , n77069 , 
   n77070 , n77071 , n77072 , n77073 , n77074 , n77075 , n77076 , n77077 , n77078 , n77079 , 
   n77080 , n77081 , n77082 , n77083 , n77084 , n77085 , n77086 , n77087 , n77088 , n77089 , 
   n77090 , n77091 , n77092 , n77093 , n77094 , n77095 , n77096 , n77097 , n77098 , n77099 , 
   n77100 , n77101 , n77102 , n77103 , n77104 , n77105 , n77106 , n77107 , n77108 , n77109 , 
   n77110 , n77111 , n77112 , n77113 , n77114 , n77115 , n77116 , n77117 , n77118 , n77119 , 
   n77120 , n77121 , n77122 , n77123 , n77124 , n77125 , n77126 , n77127 , n77128 , n77129 , 
   n77130 , n77131 , n77132 , n77133 , n77134 , n77135 , n77136 , n77137 , n77138 , n77139 , 
   n77140 , n77141 , n77142 , n77143 , n77144 , n77145 , n77146 , n77147 , n77148 , n77149 , 
   n77150 , n77151 , n77152 , n77153 , n77154 , n77155 , n77156 , n77157 , n77158 , n77159 , 
   n77160 , n77161 , n77162 , n77163 , n77164 , n77165 , n77166 , n77167 , n77168 , n77169 , 
   n77170 , n77171 , n77172 , n77173 , n77174 , n77175 , n77176 , n77177 , n77178 , n77179 , 
   n77180 , n77181 , n77182 , n77183 , n77184 , n77185 , n77186 , n77187 , n77188 , n77189 , 
   n77190 , n77191 , n77192 , n77193 , n77194 , n77195 , n77196 , n77197 , n77198 , n77199 , 
   n77200 , n77201 , n77202 , n77203 , n77204 , n77205 , n77206 , n77207 , n77208 , n77209 , 
   n77210 , n77211 , n77212 , n77213 , n77214 , n77215 , n77216 , n77217 , n77218 , n77219 , 
   n77220 , n77221 , n77222 , n77223 , n77224 , n77225 , n77226 , n77227 , n77228 , n77229 , 
   n77230 , n77231 , n77232 , n77233 , n77234 , n77235 , n77236 , n77237 , n77238 , n77239 , 
   n77240 , n77241 , n77242 , n77243 , n77244 , n77245 , n77246 , n77247 , n77248 , n77249 , 
   n77250 , n77251 , n77252 , n77253 , n77254 , n77255 , n77256 , n77257 , n77258 , n77259 , 
   n77260 , n77261 , n77262 , n77263 , n77264 , n77265 , n77266 , n77267 , n77268 , n77269 , 
   n77270 , n77271 , n77272 , n77273 , n77274 , n77275 , n77276 , n77277 , n77278 , n77279 , 
   n77280 , n77281 , n77282 , n77283 , n77284 , n77285 , n77286 , n77287 , n77288 , n77289 , 
   n77290 , n77291 , n77292 , n77293 , n77294 , n77295 , n77296 , n77297 , n77298 , n77299 , 
   n77300 , n77301 , n77302 , n77303 , n77304 , n77305 , n77306 , n77307 , n77308 , n77309 , 
   n77310 , n77311 , n77312 , n77313 , n77314 , n77315 , n77316 , n77317 , n77318 , n77319 , 
   n77320 , n77321 , n77322 , n77323 , n77324 , n77325 , n77326 , n77327 , n77328 , n77329 , 
   n77330 , n77331 , n77332 , n77333 , n77334 , n77335 , n77336 , n77337 , n77338 , n77339 , 
   n77340 , n77341 , n77342 , n77343 , n77344 , n77345 , n77346 , n77347 , n77348 , n77349 , 
   n77350 , n77351 , n77352 , n77353 , n77354 , n77355 , n77356 , n77357 , n77358 , n77359 , 
   n77360 , n77361 , n77362 , n77363 , n77364 , n77365 , n77366 , n77367 , n77368 , n77369 , 
   n77370 , n77371 , n77372 , n77373 , n77374 , n77375 , n77376 , n77377 , n77378 , n77379 , 
   n77380 , n77381 , n77382 , n77383 , n77384 , n77385 , n77386 , n77387 , n77388 , n77389 , 
   n77390 , n77391 , n77392 , n77393 , n77394 , n77395 , n77396 , n77397 , n77398 , n77399 , 
   n77400 , n77401 , n77402 , n77403 , n77404 , n77405 , n77406 , n77407 , n77408 , n77409 , 
   n77410 , n77411 , n77412 , n77413 , n77414 , n77415 , n77416 , n77417 , n77418 , n77419 , 
   n77420 , n77421 , n77422 , n77423 , n77424 , n77425 , n77426 , n77427 , n77428 , n77429 , 
   n77430 , n77431 , n77432 , n77433 , n77434 , n77435 , n77436 , n77437 , n77438 , n77439 , 
   n77440 , n77441 , n77442 , n77443 , n77444 , n77445 , n77446 , n77447 , n77448 , n77449 , 
   n77450 , n77451 , n77452 , n77453 , n77454 , n77455 , n77456 , n77457 , n77458 , n77459 , 
   n77460 , n77461 , n77462 , n77463 , n77464 , n77465 , n77466 , n77467 , n77468 , n77469 , 
   n77470 , n77471 , n77472 , n77473 , n77474 , n77475 , n77476 , n77477 , n77478 , n77479 , 
   n77480 , n77481 , n77482 , n77483 , n77484 , n77485 , n77486 , n77487 , n77488 , n77489 , 
   n77490 , n77491 , n77492 , n77493 , n77494 , n77495 , n77496 , n77497 , n77498 , n77499 , 
   n77500 , n77501 , n77502 , n77503 , n77504 , n77505 , n77506 , n77507 , n77508 , n77509 , 
   n77510 , n77511 , n77512 , n77513 , n77514 , n77515 , n77516 , n77517 , n77518 , n77519 , 
   n77520 , n77521 , n77522 , n77523 , n77524 , n77525 , n77526 , n77527 , n77528 , n77529 , 
   n77530 , n77531 , n77532 , n77533 , n77534 , n77535 , n77536 , n77537 , n77538 , n77539 , 
   n77540 , n77541 , n77542 , n77543 , n77544 , n77545 , n77546 , n77547 , n77548 , n77549 , 
   n77550 , n77551 , n77552 , n77553 , n77554 , n77555 , n77556 , n77557 , n77558 , n77559 , 
   n77560 , n77561 , n77562 , n77563 , n77564 , n77565 , n77566 , n77567 , n77568 , n77569 , 
   n77570 , n77571 , n77572 , n77573 , n77574 , n77575 , n77576 , n77577 , n77578 , n77579 , 
   n77580 , n77581 , n77582 , n77583 , n77584 , n77585 , n77586 , n77587 , n77588 , n77589 , 
   n77590 , n77591 , n77592 , n77593 , n77594 , n77595 , n77596 , n77597 , n77598 , n77599 , 
   n77600 , n77601 , n77602 , n77603 , n77604 , n77605 , n77606 , n77607 , n77608 , n77609 , 
   n77610 , n77611 , n77612 , n77613 , n77614 , n77615 , n77616 , n77617 , n77618 , n77619 , 
   n77620 , n77621 , n77622 , n77623 , n77624 , n77625 , n77626 , n77627 , n77628 , n77629 , 
   n77630 , n77631 , n77632 , n77633 , n77634 , n77635 , n77636 , n77637 , n77638 , n77639 , 
   n77640 , n77641 , n77642 , n77643 , n77644 , n77645 , n77646 , n77647 , n77648 , n77649 , 
   n77650 , n77651 , n77652 , n77653 , n77654 , n77655 , n77656 , n77657 , n77658 , n77659 , 
   n77660 , n77661 , n77662 , n77663 , n77664 , n77665 , n77666 , n77667 , n77668 , n77669 , 
   n77670 , n77671 , n77672 , n77673 , n77674 , n77675 , n77676 , n77677 , n77678 , n77679 , 
   n77680 , n77681 , n77682 , n77683 , n77684 , n77685 , n77686 , n77687 , n77688 , n77689 , 
   n77690 , n77691 , n77692 , n77693 , n77694 , n77695 , n77696 , n77697 , n77698 , n77699 , 
   n77700 , n77701 , n77702 , n77703 , n77704 , n77705 , n77706 , n77707 , n77708 , n77709 , 
   n77710 , n77711 , n77712 , n77713 , n77714 , n77715 , n77716 , n77717 , n77718 , n77719 , 
   n77720 , n77721 , n77722 , n77723 , n77724 , n77725 , n77726 , n77727 , n77728 , n77729 , 
   n77730 , n77731 , n77732 , n77733 , n77734 , n77735 , n77736 , n77737 , n77738 , n77739 , 
   n77740 , n77741 , n77742 , n77743 , n77744 , n77745 , n77746 , n77747 , n77748 , n77749 , 
   n77750 , n77751 , n77752 , n77753 , n77754 , n77755 , n77756 , n77757 , n77758 , n77759 , 
   n77760 , n77761 , n77762 , n77763 , n77764 , n77765 , n77766 , n77767 , n77768 , n77769 , 
   n77770 , n77771 , n77772 , n77773 , n77774 , n77775 , n77776 , n77777 , n77778 , n77779 , 
   n77780 , n77781 , n77782 , n77783 , n77784 , n77785 , n77786 ;
buf ( n243 , n2533 );
buf ( n244 , n2538 );
buf ( n245 , n2543 );
buf ( n246 , n2548 );
buf ( n247 , n2553 );
buf ( n248 , n2558 );
buf ( n249 , n2563 );
buf ( n250 , n2568 );
buf ( n251 , n2573 );
buf ( n252 , n2578 );
buf ( n253 , n2583 );
buf ( n254 , n2588 );
buf ( n255 , n2593 );
buf ( n256 , n2598 );
buf ( n257 , n2603 );
buf ( n258 , n2605 );
buf ( n259 , n68753 );
buf ( n260 , n68755 );
buf ( n261 , n68760 );
buf ( n262 , n2622 );
buf ( n263 , n2624 );
buf ( n264 , n68769 );
buf ( n265 , n2628 );
buf ( n266 , n68773 );
buf ( n267 , n68775 );
buf ( n268 , n2634 );
buf ( n269 , n2636 );
buf ( n270 , n2638 );
buf ( n271 , n68783 );
buf ( n272 , n68785 );
buf ( n273 , n2644 );
buf ( n274 , n68789 );
buf ( n275 , n2648 );
buf ( n276 , n2650 );
buf ( n277 , n2652 );
buf ( n278 , n2654 );
buf ( n279 , n68799 );
buf ( n280 , n2658 );
buf ( n281 , n68803 );
buf ( n282 , n68805 );
buf ( n283 , n2664 );
buf ( n284 , n2666 );
buf ( n285 , n2668 );
buf ( n286 , n68813 );
buf ( n287 , n68815 );
buf ( n288 , n2674 );
buf ( n289 , n68819 );
buf ( n290 , n2681 );
buf ( n291 , n68829 );
buf ( n292 , n2688 );
buf ( n293 , n68833 );
buf ( n294 , n68835 );
buf ( PO_rd , n2694 );
buf ( PO_wr , n2696 );
buf ( DFF_state_reg_S , n71976 );
buf ( DFF_state_reg_R , n71978 );
buf ( DFF_state_reg_CK , n71979 );
buf ( DFF_state_reg_D , n71980 );
buf ( n295 , n76385 );
buf ( n296 , n76387 );
buf ( n297 , n76388 );
buf ( n298 , n76394 );
buf ( n299 , n10137 );
buf ( n300 , n10139 );
buf ( n301 , n76283 );
buf ( n302 , n76289 );
buf ( n303 , n76171 );
buf ( n304 , n76173 );
buf ( n305 , n76174 );
buf ( n306 , n76180 );
buf ( n307 , n76143 );
buf ( n308 , n76145 );
buf ( n309 , n76146 );
buf ( n310 , n76152 );
buf ( n311 , n76133 );
buf ( n312 , n76135 );
buf ( n313 , n76136 );
buf ( n314 , n76142 );
buf ( n315 , n76123 );
buf ( n316 , n76125 );
buf ( n317 , n9983 );
buf ( n318 , n76132 );
buf ( n319 , n76113 );
buf ( n320 , n76115 );
buf ( n321 , n76116 );
buf ( n322 , n9979 );
buf ( n323 , n76103 );
buf ( n324 , n76105 );
buf ( n325 , n76106 );
buf ( n326 , n76112 );
buf ( n327 , n9950 );
buf ( n328 , n9952 );
buf ( n329 , n9953 );
buf ( n330 , n76102 );
buf ( n331 , n76084 );
buf ( n332 , n76086 );
buf ( n333 , n9944 );
buf ( n334 , n76092 );
buf ( n335 , n10233 );
buf ( n336 , n76378 );
buf ( n337 , n76379 );
buf ( n338 , n76384 );
buf ( n339 , n10224 );
buf ( n340 , n10226 );
buf ( n341 , n76370 );
buf ( n342 , n10232 );
buf ( n343 , n76358 );
buf ( n344 , n76360 );
buf ( n345 , n76361 );
buf ( n346 , n76366 );
buf ( n347 , n76349 );
buf ( n348 , n76351 );
buf ( n349 , n76352 );
buf ( n350 , n76357 );
buf ( n351 , n10197 );
buf ( n352 , n10199 );
buf ( n353 , n76343 );
buf ( n354 , n76348 );
buf ( n355 , n76331 );
buf ( n356 , n10190 );
buf ( n357 , n10191 );
buf ( n358 , n10196 );
buf ( n359 , n76321 );
buf ( n360 , n76323 );
buf ( n361 , n76324 );
buf ( n362 , n76330 );
buf ( n363 , n76311 );
buf ( n364 , n76313 );
buf ( n365 , n76314 );
buf ( n366 , n76320 );
buf ( n367 , n10157 );
buf ( n368 , n76302 );
buf ( n369 , n76303 );
buf ( n370 , n76310 );
buf ( n371 , n76290 );
buf ( n372 , n76292 );
buf ( n373 , n76293 );
buf ( n374 , n10156 );
buf ( n375 , n10127 );
buf ( n376 , n10129 );
buf ( n377 , n10130 );
buf ( n378 , n76279 );
buf ( n379 , n76260 );
buf ( n380 , n10119 );
buf ( n381 , n10120 );
buf ( n382 , n10126 );
buf ( n383 , n76250 );
buf ( n384 , n76252 );
buf ( n385 , n76253 );
buf ( n386 , n76259 );
buf ( n387 , n76240 );
buf ( n388 , n76242 );
buf ( n389 , n10100 );
buf ( n390 , n76249 );
buf ( n391 , n76230 );
buf ( n392 , n10089 );
buf ( n393 , n10090 );
buf ( n394 , n10096 );
buf ( n395 , n76220 );
buf ( n396 , n76222 );
buf ( n397 , n76223 );
buf ( n398 , n76229 );
buf ( n399 , n10067 );
buf ( n400 , n10069 );
buf ( n401 , n10070 );
buf ( n402 , n10076 );
buf ( n403 , n76200 );
buf ( n404 , n10059 );
buf ( n405 , n10060 );
buf ( n406 , n76209 );
buf ( n407 , n76190 );
buf ( n408 , n10049 );
buf ( n409 , n10050 );
buf ( n410 , n76199 );
buf ( n411 , n76181 );
buf ( n412 , n76183 );
buf ( n413 , n76184 );
buf ( n414 , n76189 );
buf ( n415 , n10019 );
buf ( n416 , n76164 );
buf ( n417 , n76165 );
buf ( n418 , n76170 );
buf ( n419 , n10010 );
buf ( n420 , n10012 );
buf ( n421 , n76156 );
buf ( n422 , n10018 );
buf ( n423 , n75257 );
buf ( n424 , n75259 );
buf ( n425 , n75260 );
buf ( n426 , n75265 );
buf ( n427 , n75247 );
buf ( n428 , n75249 );
buf ( n429 , n75250 );
buf ( n430 , n75256 );
buf ( n431 , n73729 );
buf ( n432 , n73731 );
buf ( n433 , n73732 );
buf ( n434 , n7619 );
buf ( n435 , n73408 );
buf ( n436 , n73410 );
buf ( n437 , n73411 );
buf ( n438 , n73444 );
buf ( n439 , n72380 );
buf ( n440 , n72382 );
buf ( n441 , n72383 );
buf ( n442 , n72428 );
buf ( n443 , n6185 );
buf ( n444 , n72330 );
buf ( n445 , n72331 );
buf ( n446 , n72379 );
buf ( n447 , n6137 );
buf ( n448 , n72282 );
buf ( n449 , n72283 );
buf ( n450 , n72327 );
buf ( n451 , n72218 );
buf ( n452 , n6077 );
buf ( n453 , n6078 );
buf ( n454 , n72279 );
buf ( n455 , n6018 );
buf ( n456 , n72163 );
buf ( n457 , n72164 );
buf ( n458 , n72217 );
buf ( n459 , n72082 );
buf ( n460 , n5941 );
buf ( n461 , n72085 );
buf ( n462 , n6017 );
buf ( n463 , n72030 );
buf ( n464 , n72032 );
buf ( n465 , n5890 );
buf ( n466 , n5938 );
buf ( n467 , n71981 );
buf ( n468 , n71983 );
buf ( n469 , n71984 );
buf ( n470 , n5886 );
buf ( n471 , n73704 );
buf ( n472 , n73706 );
buf ( n473 , n73707 );
buf ( n474 , n73728 );
buf ( n475 , n7537 );
buf ( n476 , n73682 );
buf ( n477 , n7540 );
buf ( n478 , n73703 );
buf ( n479 , n73655 );
buf ( n480 , n73657 );
buf ( n481 , n73658 );
buf ( n482 , n7536 );
buf ( n483 , n73581 );
buf ( n484 , n73583 );
buf ( n485 , n73584 );
buf ( n486 , n73654 );
buf ( n487 , n73557 );
buf ( n488 , n73559 );
buf ( n489 , n73560 );
buf ( n490 , n73580 );
buf ( n491 , n7389 );
buf ( n492 , n73534 );
buf ( n493 , n7392 );
buf ( n494 , n73556 );
buf ( n495 , n73512 );
buf ( n496 , n73514 );
buf ( n497 , n73515 );
buf ( n498 , n7388 );
buf ( n499 , n73490 );
buf ( n500 , n73492 );
buf ( n501 , n7350 );
buf ( n502 , n73511 );
buf ( n503 , n73468 );
buf ( n504 , n7327 );
buf ( n505 , n7328 );
buf ( n506 , n7346 );
buf ( n507 , n73445 );
buf ( n508 , n73447 );
buf ( n509 , n73448 );
buf ( n510 , n7324 );
buf ( n511 , n7208 );
buf ( n512 , n73353 );
buf ( n513 , n73354 );
buf ( n514 , n73407 );
buf ( n515 , n73280 );
buf ( n516 , n7139 );
buf ( n517 , n7140 );
buf ( n518 , n73350 );
buf ( n519 , n73216 );
buf ( n520 , n73218 );
buf ( n521 , n73219 );
buf ( n522 , n73279 );
buf ( n523 , n6988 );
buf ( n524 , n73133 );
buf ( n525 , n73134 );
buf ( n526 , n73215 );
buf ( n527 , n6927 );
buf ( n528 , n73072 );
buf ( n529 , n73073 );
buf ( n530 , n6987 );
buf ( n531 , n6853 );
buf ( n532 , n72998 );
buf ( n533 , n72999 );
buf ( n534 , n73069 );
buf ( n535 , n6777 );
buf ( n536 , n72922 );
buf ( n537 , n72923 );
buf ( n538 , n6852 );
buf ( n539 , n72837 );
buf ( n540 , n6696 );
buf ( n541 , n6697 );
buf ( n542 , n72919 );
buf ( n543 , n72429 );
buf ( n544 , n72431 );
buf ( n545 , n72432 );
buf ( n546 , n72836 );
buf ( n547 , n74845 );
buf ( n548 , n74847 );
buf ( n549 , n74848 );
buf ( n550 , n8721 );
buf ( n551 , n8662 );
buf ( n552 , n74807 );
buf ( n553 , n74808 );
buf ( n554 , n74823 );
buf ( n555 , n74579 );
buf ( n556 , n8438 );
buf ( n557 , n8439 );
buf ( n558 , n8455 );
buf ( n559 , n8397 );
buf ( n560 , n74542 );
buf ( n561 , n74543 );
buf ( n562 , n8417 );
buf ( n563 , n74518 );
buf ( n564 , n74520 );
buf ( n565 , n74521 );
buf ( n566 , n74539 );
buf ( n567 , n74496 );
buf ( n568 , n8355 );
buf ( n569 , n74499 );
buf ( n570 , n74517 );
buf ( n571 , n74478 );
buf ( n572 , n74480 );
buf ( n573 , n74481 );
buf ( n574 , n8352 );
buf ( n575 , n74454 );
buf ( n576 , n8313 );
buf ( n577 , n74457 );
buf ( n578 , n74477 );
buf ( n579 , n74436 );
buf ( n580 , n74438 );
buf ( n581 , n8296 );
buf ( n582 , n74453 );
buf ( n583 , n70910 );
buf ( n584 , n70912 );
buf ( n585 , n4770 );
buf ( n586 , n4881 );
buf ( n587 , n71663 );
buf ( n588 , n71665 );
buf ( n589 , n71666 );
buf ( n590 , n71722 );
buf ( n591 , n5440 );
buf ( n592 , n71585 );
buf ( n593 , n71586 );
buf ( n594 , n71662 );
buf ( n595 , n71517 );
buf ( n596 , n5376 );
buf ( n597 , n71520 );
buf ( n598 , n71582 );
buf ( n599 , n74824 );
buf ( n600 , n8683 );
buf ( n601 , n74827 );
buf ( n602 , n74844 );
buf ( n603 , n5301 );
buf ( n604 , n71446 );
buf ( n605 , n71447 );
buf ( n606 , n71516 );
buf ( n607 , n71352 );
buf ( n608 , n71354 );
buf ( n609 , n71355 );
buf ( n610 , n5300 );
buf ( n611 , n71328 );
buf ( n612 , n71330 );
buf ( n613 , n71331 );
buf ( n614 , n71351 );
buf ( n615 , n5129 );
buf ( n616 , n71274 );
buf ( n617 , n71275 );
buf ( n618 , n71327 );
buf ( n619 , n5072 );
buf ( n620 , n71217 );
buf ( n621 , n5075 );
buf ( n622 , n5128 );
buf ( n623 , n4882 );
buf ( n624 , n4884 );
buf ( n625 , n4885 );
buf ( n626 , n71214 );
buf ( n627 , n8640 );
buf ( n628 , n74785 );
buf ( n629 , n74786 );
buf ( n630 , n8661 );
buf ( n631 , n8620 );
buf ( n632 , n74765 );
buf ( n633 , n74766 );
buf ( n634 , n8639 );
buf ( n635 , n74743 );
buf ( n636 , n74745 );
buf ( n637 , n8603 );
buf ( n638 , n8619 );
buf ( n639 , n74723 );
buf ( n640 , n8582 );
buf ( n641 , n74726 );
buf ( n642 , n74742 );
buf ( n643 , n74703 );
buf ( n644 , n74705 );
buf ( n645 , n74706 );
buf ( n646 , n74722 );
buf ( n647 , n8540 );
buf ( n648 , n74685 );
buf ( n649 , n74686 );
buf ( n650 , n74702 );
buf ( n651 , n8520 );
buf ( n652 , n74665 );
buf ( n653 , n74666 );
buf ( n654 , n74682 );
buf ( n655 , n8500 );
buf ( n656 , n8502 );
buf ( n657 , n8503 );
buf ( n658 , n8519 );
buf ( n659 , n74621 );
buf ( n660 , n74623 );
buf ( n661 , n74624 );
buf ( n662 , n8499 );
buf ( n663 , n8456 );
buf ( n664 , n74601 );
buf ( n665 , n74602 );
buf ( n666 , n74620 );
buf ( n667 , n74570 );
buf ( n668 , n8429 );
buf ( n669 , n74573 );
buf ( n670 , n74578 );
buf ( n671 , n8418 );
buf ( n672 , n74563 );
buf ( n673 , n74564 );
buf ( n674 , n8426 );
buf ( n675 , n75120 );
buf ( n676 , n8979 );
buf ( n677 , n75123 );
buf ( n678 , n8984 );
buf ( n679 , n8889 );
buf ( n680 , n8891 );
buf ( n681 , n75035 );
buf ( n682 , n75039 );
buf ( n683 , n8799 );
buf ( n684 , n74944 );
buf ( n685 , n74945 );
buf ( n686 , n74949 );
buf ( n687 , n74916 );
buf ( n688 , n74918 );
buf ( n689 , n74919 );
buf ( n690 , n74924 );
buf ( n691 , n74908 );
buf ( n692 , n8767 );
buf ( n693 , n8768 );
buf ( n694 , n74915 );
buf ( n695 , n8757 );
buf ( n696 , n74902 );
buf ( n697 , n74903 );
buf ( n698 , n74907 );
buf ( n699 , n74892 );
buf ( n700 , n8751 );
buf ( n701 , n8752 );
buf ( n702 , n8756 );
buf ( n703 , n8741 );
buf ( n704 , n8743 );
buf ( n705 , n74887 );
buf ( n706 , n74891 );
buf ( n707 , n8733 );
buf ( n708 , n8735 );
buf ( n709 , n8736 );
buf ( n710 , n8740 );
buf ( n711 , n8722 );
buf ( n712 , n8724 );
buf ( n713 , n8725 );
buf ( n714 , n74875 );
buf ( n715 , n75112 );
buf ( n716 , n75114 );
buf ( n717 , n75115 );
buf ( n718 , n75119 );
buf ( n719 , n75104 );
buf ( n720 , n8963 );
buf ( n721 , n8964 );
buf ( n722 , n75111 );
buf ( n723 , n75096 );
buf ( n724 , n8955 );
buf ( n725 , n8956 );
buf ( n726 , n75103 );
buf ( n727 , n75088 );
buf ( n728 , n8947 );
buf ( n729 , n75091 );
buf ( n730 , n8952 );
buf ( n731 , n75080 );
buf ( n732 , n75082 );
buf ( n733 , n8940 );
buf ( n734 , n8944 );
buf ( n735 , n75072 );
buf ( n736 , n75074 );
buf ( n737 , n75075 );
buf ( n738 , n8936 );
buf ( n739 , n75064 );
buf ( n740 , n75066 );
buf ( n741 , n75067 );
buf ( n742 , n75071 );
buf ( n743 , n75056 );
buf ( n744 , n8915 );
buf ( n745 , n8916 );
buf ( n746 , n75063 );
buf ( n747 , n8905 );
buf ( n748 , n75050 );
buf ( n749 , n75051 );
buf ( n750 , n75055 );
buf ( n751 , n75040 );
buf ( n752 , n8899 );
buf ( n753 , n8900 );
buf ( n754 , n8904 );
buf ( n755 , n8881 );
buf ( n756 , n8883 );
buf ( n757 , n8884 );
buf ( n758 , n8888 );
buf ( n759 , n8873 );
buf ( n760 , n75018 );
buf ( n761 , n75019 );
buf ( n762 , n75023 );
buf ( n763 , n75008 );
buf ( n764 , n8867 );
buf ( n765 , n8868 );
buf ( n766 , n8872 );
buf ( n767 , n75000 );
buf ( n768 , n75002 );
buf ( n769 , n8860 );
buf ( n770 , n75007 );
buf ( n771 , n74992 );
buf ( n772 , n74994 );
buf ( n773 , n74995 );
buf ( n774 , n74999 );
buf ( n775 , n8841 );
buf ( n776 , n74986 );
buf ( n777 , n74987 );
buf ( n778 , n74991 );
buf ( n779 , n74976 );
buf ( n780 , n74978 );
buf ( n781 , n8836 );
buf ( n782 , n74983 );
buf ( n783 , n74966 );
buf ( n784 , n8825 );
buf ( n785 , n8826 );
buf ( n786 , n74975 );
buf ( n787 , n8815 );
buf ( n788 , n8817 );
buf ( n789 , n74961 );
buf ( n790 , n74965 );
buf ( n791 , n8807 );
buf ( n792 , n8809 );
buf ( n793 , n8810 );
buf ( n794 , n8814 );
buf ( n795 , n74934 );
buf ( n796 , n8793 );
buf ( n797 , n8794 );
buf ( n798 , n8798 );
buf ( n799 , n74925 );
buf ( n800 , n74927 );
buf ( n801 , n74928 );
buf ( n802 , n74933 );
buf ( DFF_B_reg_S , n76395 );
buf ( DFF_B_reg_R , n76397 );
buf ( DFF_B_reg_CK , n76398 );
buf ( DFF_B_reg_D , n77769 );
buf ( n803 , n8275 );
buf ( n804 , n8277 );
buf ( n805 , n8278 );
buf ( n806 , n8292 );
buf ( n807 , n74227 );
buf ( n808 , n8086 );
buf ( n809 , n74230 );
buf ( n810 , n74247 );
buf ( n811 , n73956 );
buf ( n812 , n73958 );
buf ( n813 , n73959 );
buf ( n814 , n73972 );
buf ( n815 , n73877 );
buf ( n816 , n73879 );
buf ( n817 , n73880 );
buf ( n818 , n73892 );
buf ( n819 , n73854 );
buf ( n820 , n73856 );
buf ( n821 , n73857 );
buf ( n822 , n73876 );
buf ( n823 , n7693 );
buf ( n824 , n73838 );
buf ( n825 , n73839 );
buf ( n826 , n73853 );
buf ( n827 , n7677 );
buf ( n828 , n73822 );
buf ( n829 , n73823 );
buf ( n830 , n73835 );
buf ( n831 , n73804 );
buf ( n832 , n73806 );
buf ( n833 , n73807 );
buf ( n834 , n7676 );
buf ( n835 , n7641 );
buf ( n836 , n73786 );
buf ( n837 , n73787 );
buf ( n838 , n73803 );
buf ( n839 , n7620 );
buf ( n840 , n73765 );
buf ( n841 , n7623 );
buf ( n842 , n73783 );
buf ( n843 , n74399 );
buf ( n844 , n74401 );
buf ( n845 , n74402 );
buf ( n846 , n8274 );
buf ( n847 , n74380 );
buf ( n848 , n8239 );
buf ( n849 , n74383 );
buf ( n850 , n74398 );
buf ( n851 , n8218 );
buf ( n852 , n74363 );
buf ( n853 , n74364 );
buf ( n854 , n74379 );
buf ( n855 , n74342 );
buf ( n856 , n8201 );
buf ( n857 , n8202 );
buf ( n858 , n8217 );
buf ( n859 , n74323 );
buf ( n860 , n74325 );
buf ( n861 , n74326 );
buf ( n862 , n74341 );
buf ( n863 , n74304 );
buf ( n864 , n74306 );
buf ( n865 , n8164 );
buf ( n866 , n74322 );
buf ( n867 , n2698 );
buf ( n868 , n68844 );
buf ( n869 , n68845 );
buf ( n870 , n4766 );
buf ( n871 , n8143 );
buf ( n872 , n74288 );
buf ( n873 , n74289 );
buf ( n874 , n8160 );
buf ( n875 , n74267 );
buf ( n876 , n8126 );
buf ( n877 , n8127 );
buf ( n878 , n8142 );
buf ( n879 , n74248 );
buf ( n880 , n74250 );
buf ( n881 , n74251 );
buf ( n882 , n74266 );
buf ( n883 , n74208 );
buf ( n884 , n8067 );
buf ( n885 , n8068 );
buf ( n886 , n74226 );
buf ( n887 , n8046 );
buf ( n888 , n8048 );
buf ( n889 , n74192 );
buf ( n890 , n8064 );
buf ( n891 , n8027 );
buf ( n892 , n74172 );
buf ( n893 , n74173 );
buf ( n894 , n74188 );
buf ( n895 , n74151 );
buf ( n896 , n74153 );
buf ( n897 , n8011 );
buf ( n898 , n74169 );
buf ( n899 , n7989 );
buf ( n900 , n74134 );
buf ( n901 , n74135 );
buf ( n902 , n74150 );
buf ( n903 , n7972 );
buf ( n904 , n7974 );
buf ( n905 , n74118 );
buf ( n906 , n74131 );
buf ( n907 , n7954 );
buf ( n908 , n74099 );
buf ( n909 , n74100 );
buf ( n910 , n74114 );
buf ( n911 , n7937 );
buf ( n912 , n74082 );
buf ( n913 , n74083 );
buf ( n914 , n7953 );
buf ( n915 , n7921 );
buf ( n916 , n74066 );
buf ( n917 , n74067 );
buf ( n918 , n74079 );
buf ( n919 , n7830 );
buf ( n920 , n7832 );
buf ( n921 , n7833 );
buf ( n922 , n7920 );
buf ( n923 , n73936 );
buf ( n924 , n7795 );
buf ( n925 , n73939 );
buf ( n926 , n73955 );
buf ( n927 , n7750 );
buf ( n928 , n7752 );
buf ( n929 , n73896 );
buf ( n930 , n73935 );
buf ( n931 , n76070 );
buf ( n932 , n76072 );
buf ( n933 , n76073 );
buf ( n934 , n76083 );
buf ( n935 , n75612 );
buf ( n936 , n75614 );
buf ( n937 , n75615 );
buf ( n938 , n9484 );
buf ( n939 , n75582 );
buf ( n940 , n75584 );
buf ( n941 , n75585 );
buf ( n942 , n75611 );
buf ( n943 , n75555 );
buf ( n944 , n75557 );
buf ( n945 , n75558 );
buf ( n946 , n75581 );
buf ( n947 , n75519 );
buf ( n948 , n75521 );
buf ( n949 , n75522 );
buf ( n950 , n75554 );
buf ( n951 , n75488 );
buf ( n952 , n75490 );
buf ( n953 , n75491 );
buf ( n954 , n75518 );
buf ( n955 , n9318 );
buf ( n956 , n75463 );
buf ( n957 , n75464 );
buf ( n958 , n75487 );
buf ( n959 , n75424 );
buf ( n960 , n75426 );
buf ( n961 , n9284 );
buf ( n962 , n9317 );
buf ( n963 , n75399 );
buf ( n964 , n9258 );
buf ( n965 , n9259 );
buf ( n966 , n75423 );
buf ( n967 , n75266 );
buf ( n968 , n9125 );
buf ( n969 , n9126 );
buf ( n970 , n75398 );
buf ( n971 , n76042 );
buf ( n972 , n76044 );
buf ( n973 , n76045 );
buf ( n974 , n76069 );
buf ( n975 , n76004 );
buf ( n976 , n76006 );
buf ( n977 , n76007 );
buf ( n978 , n76041 );
buf ( n979 , n75978 );
buf ( n980 , n75980 );
buf ( n981 , n75981 );
buf ( n982 , n76003 );
buf ( n983 , n75944 );
buf ( n984 , n75946 );
buf ( n985 , n75947 );
buf ( n986 , n75977 );
buf ( n987 , n75914 );
buf ( n988 , n75916 );
buf ( n989 , n75917 );
buf ( n990 , n75943 );
buf ( n991 , n9721 );
buf ( n992 , n9723 );
buf ( n993 , n75867 );
buf ( n994 , n75913 );
buf ( n995 , n9690 );
buf ( n996 , n75835 );
buf ( n997 , n75836 );
buf ( n998 , n9720 );
buf ( n999 , n9657 );
buf ( n1000 , n75802 );
buf ( n1001 , n75803 );
buf ( n1002 , n9689 );
buf ( n1003 , n9620 );
buf ( n1004 , n9622 );
buf ( n1005 , n9623 );
buf ( n1006 , n9656 );
buf ( n1007 , n75628 );
buf ( n1008 , n75630 );
buf ( n1009 , n9488 );
buf ( n1010 , n75762 );
buf ( n1011 , n9092 );
buf ( n1012 , n75237 );
buf ( n1013 , n75238 );
buf ( n1014 , n75246 );
buf ( n1015 , n75223 );
buf ( n1016 , n9082 );
buf ( n1017 , n9083 );
buf ( n1018 , n9091 );
buf ( n1019 , n75193 );
buf ( n1020 , n9052 );
buf ( n1021 , n9053 );
buf ( n1022 , n75204 );
buf ( n1023 , n9030 );
buf ( n1024 , n9032 );
buf ( n1025 , n75176 );
buf ( n1026 , n75183 );
buf ( n1027 , n9021 );
buf ( n1028 , n75166 );
buf ( n1029 , n75167 );
buf ( n1030 , n9029 );
buf ( n1031 , n75155 );
buf ( n1032 , n9014 );
buf ( n1033 , n9015 );
buf ( n1034 , n9020 );
buf ( n1035 , n75146 );
buf ( n1036 , n75148 );
buf ( n1037 , n75149 );
buf ( n1038 , n75154 );
buf ( n1039 , n75137 );
buf ( n1040 , n75139 );
buf ( n1041 , n75140 );
buf ( n1042 , n75145 );
buf ( n1043 , n8985 );
buf ( n1044 , n75130 );
buf ( n1045 , n75131 );
buf ( n1046 , n75136 );
buf ( n1047 , n71723 );
buf ( n1048 , n5582 );
buf ( n1049 , n5583 );
buf ( n1050 , n71734 );
buf ( n1051 , n71967 );
buf ( n1052 , n71969 );
buf ( n1053 , n71970 );
buf ( n1054 , n71975 );
buf ( n1055 , n71958 );
buf ( n1056 , n71960 );
buf ( n1057 , n71961 );
buf ( n1058 , n71966 );
buf ( n1059 , n71949 );
buf ( n1060 , n71951 );
buf ( n1061 , n71952 );
buf ( n1062 , n71957 );
buf ( n1063 , n71940 );
buf ( n1064 , n71942 );
buf ( n1065 , n71943 );
buf ( n1066 , n71948 );
buf ( n1067 , n71931 );
buf ( n1068 , n71933 );
buf ( n1069 , n71934 );
buf ( n1070 , n71939 );
buf ( n1071 , n71922 );
buf ( n1072 , n71924 );
buf ( n1073 , n71925 );
buf ( n1074 , n71930 );
buf ( n1075 , n71913 );
buf ( n1076 , n71915 );
buf ( n1077 , n71916 );
buf ( n1078 , n71921 );
buf ( n1079 , n71904 );
buf ( n1080 , n71906 );
buf ( n1081 , n71907 );
buf ( n1082 , n71912 );
buf ( n1083 , n5752 );
buf ( n1084 , n71897 );
buf ( n1085 , n5755 );
buf ( n1086 , n71903 );
buf ( n1087 , n5743 );
buf ( n1088 , n5745 );
buf ( n1089 , n5746 );
buf ( n1090 , n71894 );
buf ( n1091 , n71877 );
buf ( n1092 , n5736 );
buf ( n1093 , n71880 );
buf ( n1094 , n5742 );
buf ( n1095 , n71860 );
buf ( n1096 , n71862 );
buf ( n1097 , n71863 );
buf ( n1098 , n5733 );
buf ( n1099 , n71842 );
buf ( n1100 , n71844 );
buf ( n1101 , n5702 );
buf ( n1102 , n5716 );
buf ( n1103 , n71822 );
buf ( n1104 , n71824 );
buf ( n1105 , n5682 );
buf ( n1106 , n71841 );
buf ( n1107 , n71807 );
buf ( n1108 , n5666 );
buf ( n1109 , n71810 );
buf ( n1110 , n71821 );
buf ( n1111 , n5645 );
buf ( n1112 , n71790 );
buf ( n1113 , n71791 );
buf ( n1114 , n5663 );
buf ( n1115 , n71771 );
buf ( n1116 , n71773 );
buf ( n1117 , n71774 );
buf ( n1118 , n71787 );
buf ( n1119 , n71744 );
buf ( n1120 , n5603 );
buf ( n1121 , n71747 );
buf ( n1122 , n71770 );
buf ( n1123 , n75214 );
buf ( n1124 , n75216 );
buf ( n1125 , n75217 );
buf ( n1126 , n75222 );
buf ( n1127 , n75205 );
buf ( n1128 , n9064 );
buf ( n1129 , n75208 );
buf ( n1130 , n75213 );
buf ( n1131 , n75184 );
buf ( n1132 , n75186 );
buf ( n1133 , n75187 );
buf ( n1134 , n75192 );
buf ( n1135 , n5592 );
buf ( n1136 , n71737 );
buf ( n1137 , n5595 );
buf ( n1138 , n71743 );
buf ( DFF_rd_reg_S , n77776 );
buf ( DFF_rd_reg_R , n77778 );
buf ( DFF_rd_reg_CK , n77779 );
buf ( DFF_rd_reg_D , n77786 );
buf ( DFF_wr_reg_S , n77770 );
buf ( DFF_wr_reg_R , n77773 );
buf ( DFF_wr_reg_CK , n77774 );
buf ( DFF_wr_reg_D , n77775 );
buf ( n68638 , PI_clock);
buf ( n68639 , PI_reset);
buf ( n68640 , n0 );
buf ( n2498 , n1 );
buf ( n2499 , n2 );
buf ( n2500 , n3 );
buf ( n2501 , n4 );
buf ( n2502 , n5 );
buf ( n2503 , n6 );
buf ( n2504 , n7 );
buf ( n68648 , n8 );
buf ( n68649 , n9 );
buf ( n68650 , n10 );
buf ( n2508 , n11 );
buf ( n2509 , n12 );
buf ( n68653 , n13 );
buf ( n68654 , n14 );
buf ( n68655 , n15 );
buf ( n2513 , n16 );
buf ( n2514 , n17 );
buf ( n2515 , n18 );
buf ( n2516 , n19 );
buf ( n2517 , n20 );
buf ( n2518 , n21 );
buf ( n2519 , n22 );
buf ( n68663 , n23 );
buf ( n68664 , n24 );
buf ( n68665 , n25 );
buf ( n2523 , n26 );
buf ( n2524 , n27 );
buf ( n68668 , n28 );
buf ( n68669 , n29 );
buf ( n68670 , n30 );
buf ( n2528 , n31 );
buf ( n2529 , n210 );
not ( n68673 , n2529 );
not ( n68674 , n68673 );
buf ( n2532 , n68674 );
buf ( n2533 , n2532 );
buf ( n2534 , n209 );
not ( n68678 , n2534 );
not ( n68679 , n68678 );
buf ( n68680 , n68679 );
buf ( n2538 , n68680 );
buf ( n2539 , n208 );
not ( n68683 , n2539 );
not ( n68684 , n68683 );
buf ( n68685 , n68684 );
buf ( n2543 , n68685 );
buf ( n2544 , n207 );
not ( n68688 , n2544 );
not ( n68689 , n68688 );
buf ( n2547 , n68689 );
buf ( n2548 , n2547 );
buf ( n2549 , n206 );
not ( n68693 , n2549 );
not ( n68694 , n68693 );
buf ( n68695 , n68694 );
buf ( n2553 , n68695 );
buf ( n2554 , n205 );
not ( n68698 , n2554 );
not ( n68699 , n68698 );
buf ( n68700 , n68699 );
buf ( n2558 , n68700 );
buf ( n2559 , n204 );
not ( n68703 , n2559 );
not ( n68704 , n68703 );
buf ( n2562 , n68704 );
buf ( n2563 , n2562 );
buf ( n2564 , n203 );
not ( n68708 , n2564 );
not ( n68709 , n68708 );
buf ( n68710 , n68709 );
buf ( n2568 , n68710 );
buf ( n2569 , n202 );
not ( n68713 , n2569 );
not ( n68714 , n68713 );
buf ( n68715 , n68714 );
buf ( n2573 , n68715 );
buf ( n2574 , n201 );
not ( n68718 , n2574 );
not ( n68719 , n68718 );
buf ( n2577 , n68719 );
buf ( n2578 , n2577 );
buf ( n2579 , n200 );
not ( n68723 , n2579 );
not ( n68724 , n68723 );
buf ( n68725 , n68724 );
buf ( n2583 , n68725 );
buf ( n2584 , n199 );
not ( n68728 , n2584 );
not ( n68729 , n68728 );
buf ( n68730 , n68729 );
buf ( n2588 , n68730 );
buf ( n2589 , n198 );
not ( n68733 , n2589 );
not ( n68734 , n68733 );
buf ( n2592 , n68734 );
buf ( n2593 , n2592 );
buf ( n2594 , n197 );
not ( n68738 , n2594 );
not ( n68739 , n68738 );
buf ( n68740 , n68739 );
buf ( n2598 , n68740 );
buf ( n2599 , n196 );
not ( n68743 , n2599 );
not ( n68744 , n68743 );
buf ( n68745 , n68744 );
buf ( n2603 , n68745 );
buf ( n2604 , n195 );
buf ( n2605 , n2604 );
buf ( n2606 , n194 );
not ( n68750 , n2606 );
not ( n68751 , n68750 );
buf ( n2609 , n68751 );
buf ( n68753 , n2609 );
buf ( n68754 , n193 );
buf ( n68755 , n68754 );
buf ( n2613 , n192 );
not ( n68757 , n2613 );
not ( n68758 , n68757 );
buf ( n68759 , n68758 );
buf ( n68760 , n68759 );
buf ( n2618 , n191 );
not ( n68762 , n2618 );
not ( n68763 , n68762 );
buf ( n2621 , n68763 );
buf ( n2622 , n2621 );
buf ( n2623 , n242 );
buf ( n2624 , n2623 );
buf ( n68768 , n241 );
buf ( n68769 , n68768 );
buf ( n68770 , n240 );
buf ( n2628 , n68770 );
buf ( n2629 , n239 );
buf ( n68773 , n2629 );
buf ( n68774 , n238 );
buf ( n68775 , n68774 );
buf ( n2633 , n237 );
buf ( n2634 , n2633 );
buf ( n2635 , n236 );
buf ( n2636 , n2635 );
buf ( n2637 , n235 );
buf ( n2638 , n2637 );
buf ( n2639 , n234 );
buf ( n68783 , n2639 );
buf ( n68784 , n233 );
buf ( n68785 , n68784 );
buf ( n2643 , n232 );
buf ( n2644 , n2643 );
buf ( n68788 , n231 );
buf ( n68789 , n68788 );
buf ( n68790 , n230 );
buf ( n2648 , n68790 );
buf ( n2649 , n229 );
buf ( n2650 , n2649 );
buf ( n2651 , n228 );
buf ( n2652 , n2651 );
buf ( n2653 , n227 );
buf ( n2654 , n2653 );
buf ( n68798 , n226 );
buf ( n68799 , n68798 );
buf ( n68800 , n225 );
buf ( n2658 , n68800 );
buf ( n2659 , n224 );
buf ( n68803 , n2659 );
buf ( n68804 , n223 );
buf ( n68805 , n68804 );
buf ( n2663 , n222 );
buf ( n2664 , n2663 );
buf ( n2665 , n221 );
buf ( n2666 , n2665 );
buf ( n2667 , n220 );
buf ( n2668 , n2667 );
buf ( n2669 , n219 );
buf ( n68813 , n2669 );
buf ( n68814 , n218 );
buf ( n68815 , n68814 );
buf ( n2673 , n217 );
buf ( n2674 , n2673 );
buf ( n68818 , n216 );
buf ( n68819 , n68818 );
buf ( n68820 , n215 );
not ( n68821 , n68820 );
not ( n68822 , n68821 );
buf ( n2680 , n68822 );
buf ( n2681 , n2680 );
buf ( n2682 , n214 );
not ( n68826 , n2682 );
not ( n68827 , n68826 );
buf ( n68828 , n68827 );
buf ( n68829 , n68828 );
buf ( n68830 , n213 );
buf ( n2688 , n68830 );
buf ( n2689 , n212 );
buf ( n68833 , n2689 );
buf ( n68834 , n211 );
buf ( n68835 , n68834 );
buf ( n2693 , DFF_rd_reg_Q);
buf ( n2694 , n2693 );
buf ( n2695 , DFF_wr_reg_Q);
buf ( n2696 , n2695 );
buf ( n2697 , n175 );
buf ( n2698 , 1'b0 );
not ( n68842 , n68639 );
not ( n68843 , n68842 );
buf ( n68844 , n68843 );
buf ( n68845 , n68638 );
buf ( n2703 , n63 );
not ( n68847 , n2703 );
not ( n68848 , n68847 );
not ( n68849 , n68848 );
buf ( n68850 , n36 );
not ( n68851 , n68850 );
not ( n68852 , n68851 );
buf ( n2710 , n37 );
not ( n68854 , n2710 );
not ( n68855 , n68854 );
not ( n68856 , n68855 );
not ( n68857 , n68856 );
nor ( n68858 , n68852 , n68857 );
buf ( n68859 , n39 );
not ( n68860 , n68859 );
not ( n68861 , n68860 );
not ( n68862 , n68861 );
not ( n68863 , n68862 );
buf ( n68864 , n38 );
not ( n68865 , n68864 );
not ( n68866 , n68865 );
not ( n68867 , n68866 );
not ( n68868 , n68867 );
nor ( n68869 , n68863 , n68868 );
nand ( n68870 , n68858 , n68869 );
buf ( n2728 , n32 );
not ( n68872 , n2728 );
buf ( n68873 , n33 );
not ( n68874 , n68873 );
nand ( n68875 , n68872 , n68874 );
not ( n68876 , n68875 );
buf ( n2734 , n34 );
not ( n68878 , n2734 );
not ( n68879 , n68878 );
buf ( n68880 , n35 );
not ( n68881 , n68880 );
not ( n68882 , n68881 );
nor ( n68883 , n68879 , n68882 );
nand ( n68884 , n68876 , n68883 );
or ( n68885 , n68870 , n68884 );
not ( n68886 , n68885 );
buf ( n2744 , n41 );
not ( n68888 , n2744 );
buf ( n68889 , n40 );
not ( n68890 , n68889 );
not ( n68891 , n68890 );
not ( n68892 , n68891 );
nand ( n68893 , n68888 , n68892 );
buf ( n68894 , n43 );
not ( n68895 , n68894 );
buf ( n2753 , n42 );
not ( n68897 , n2753 );
nand ( n68898 , n68895 , n68897 );
nor ( n68899 , n68893 , n68898 );
nand ( n68900 , n68886 , n68899 );
buf ( n2758 , n44 );
and ( n68902 , n68900 , n2758 );
not ( n68903 , n68900 );
not ( n68904 , n2758 );
and ( n68905 , n68903 , n68904 );
nor ( n68906 , n68902 , n68905 );
not ( n68907 , n68906 );
not ( n68908 , n68907 );
not ( n68909 , n68908 );
or ( n68910 , n68849 , n68909 );
nand ( n68911 , n68847 , n2758 );
nand ( n68912 , n68910 , n68911 );
not ( n68913 , n68912 );
not ( n68914 , n68913 );
not ( n68915 , n68847 );
not ( n68916 , n68915 );
buf ( n2774 , n47 );
not ( n68918 , n2774 );
not ( n68919 , n68918 );
not ( n68920 , n68884 );
not ( n68921 , n68870 );
nand ( n68922 , n68920 , n68921 );
not ( n68923 , n68922 );
buf ( n68924 , n45 );
not ( n68925 , n68924 );
nand ( n68926 , n68925 , n68904 );
buf ( n2784 , n46 );
nor ( n68928 , n68926 , n2784 );
and ( n68929 , n68899 , n68928 );
nand ( n68930 , n68923 , n68929 );
not ( n68931 , n68930 );
or ( n68932 , n68919 , n68931 );
or ( n68933 , n68930 , n68918 );
nand ( n68934 , n68932 , n68933 );
not ( n68935 , n68934 );
or ( n68936 , n68916 , n68935 );
nand ( n68937 , n68847 , n2774 );
nand ( n68938 , n68936 , n68937 );
nor ( n68939 , n68914 , n68938 );
not ( n68940 , n68848 );
not ( n68941 , n68899 );
nor ( n68942 , n68941 , n2758 );
nand ( n68943 , n68923 , n68942 );
and ( n68944 , n68943 , n68924 );
not ( n68945 , n68943 );
and ( n68946 , n68945 , n68925 );
nor ( n68947 , n68944 , n68946 );
not ( n68948 , n68947 );
or ( n68949 , n68940 , n68948 );
nand ( n68950 , n68847 , n68924 );
nand ( n68951 , n68949 , n68950 );
not ( n68952 , n68951 );
not ( n68953 , n68952 );
not ( n68954 , n68848 );
nor ( n68955 , n68941 , n68926 );
nand ( n68956 , n68923 , n68955 );
and ( n68957 , n68956 , n2784 );
not ( n68958 , n68956 );
not ( n68959 , n2784 );
and ( n68960 , n68958 , n68959 );
nor ( n68961 , n68957 , n68960 );
not ( n68962 , n68961 );
or ( n68963 , n68954 , n68962 );
nand ( n68964 , n68847 , n2784 );
nand ( n68965 , n68963 , n68964 );
nor ( n68966 , n68953 , n68965 );
not ( n68967 , n68848 );
not ( n68968 , n68897 );
nor ( n68969 , n68968 , n68893 );
nand ( n68970 , n68886 , n68969 );
not ( n68971 , n68895 );
and ( n68972 , n68970 , n68971 );
not ( n68973 , n68970 );
and ( n68974 , n68973 , n68895 );
nor ( n68975 , n68972 , n68974 );
not ( n68976 , n68975 );
not ( n68977 , n68976 );
not ( n68978 , n68977 );
or ( n68979 , n68967 , n68978 );
nand ( n68980 , n68847 , n68894 );
nand ( n68981 , n68979 , n68980 );
not ( n68982 , n68981 );
not ( n68983 , n68891 );
not ( n68984 , n68847 );
or ( n68985 , n68983 , n68984 );
not ( n68986 , n68891 );
not ( n68987 , n68886 );
or ( n68988 , n68986 , n68987 );
or ( n68989 , n68923 , n68891 );
nand ( n68990 , n68988 , n68989 );
nand ( n68991 , n68990 , n2703 );
nand ( n68992 , n68985 , n68991 );
and ( n68993 , n68847 , n68861 );
not ( n68994 , n68847 );
not ( n68995 , n68863 );
not ( n68996 , n68995 );
not ( n68997 , n68856 );
nor ( n68998 , n68997 , n68852 );
not ( n68999 , n68998 );
nor ( n69000 , n68999 , n68868 );
not ( n69001 , n68882 );
not ( n69002 , n68873 );
not ( n69003 , n2728 );
not ( n69004 , n68879 );
and ( n69005 , n69001 , n69002 , n69003 , n69004 );
nand ( n69006 , n69000 , n69005 );
not ( n69007 , n69006 );
or ( n69008 , n68996 , n69007 );
nand ( n69009 , n69005 , n69000 );
or ( n69010 , n69009 , n68995 );
nand ( n69011 , n69008 , n69010 );
and ( n69012 , n68994 , n69011 );
nor ( n69013 , n68993 , n69012 );
not ( n69014 , n69013 );
not ( n69015 , n69014 );
and ( n69016 , n68847 , n68855 );
not ( n69017 , n68847 );
not ( n69018 , n68997 );
not ( n69019 , n69018 );
not ( n69020 , n68852 );
nand ( n69021 , n69005 , n69020 );
not ( n69022 , n69021 );
or ( n69023 , n69019 , n69022 );
nand ( n69024 , n69005 , n69020 );
or ( n69025 , n69024 , n69018 );
nand ( n69026 , n69023 , n69025 );
and ( n69027 , n69017 , n69026 );
nor ( n69028 , n69016 , n69027 );
not ( n69029 , n69028 );
not ( n69030 , n69029 );
nand ( n69031 , n69015 , n69030 );
nor ( n69032 , n68992 , n69031 );
and ( n69033 , n68982 , n69032 );
nand ( n69034 , n68939 , n68966 , n69033 );
not ( n69035 , n69034 );
not ( n69036 , n68848 );
not ( n69037 , n68897 );
not ( n69038 , n68893 );
nand ( n69039 , n69038 , n68886 );
not ( n69040 , n69039 );
or ( n69041 , n69037 , n69040 );
or ( n69042 , n69039 , n68897 );
nand ( n69043 , n69041 , n69042 );
not ( n69044 , n69043 );
not ( n69045 , n69044 );
not ( n69046 , n69045 );
or ( n69047 , n69036 , n69046 );
nand ( n69048 , n68847 , n2753 );
nand ( n69049 , n69047 , n69048 );
not ( n69050 , n69049 );
and ( n69051 , n68847 , n68866 );
not ( n69052 , n68847 );
not ( n69053 , n68868 );
not ( n69054 , n69053 );
nand ( n69055 , n69005 , n68998 );
not ( n69056 , n69055 );
or ( n69057 , n69054 , n69056 );
nand ( n69058 , n69005 , n68998 );
or ( n69059 , n69058 , n69053 );
nand ( n69060 , n69057 , n69059 );
and ( n69061 , n69052 , n69060 );
nor ( n69062 , n69051 , n69061 );
not ( n69063 , n69062 );
not ( n69064 , n2703 );
and ( n69065 , n69064 , n68882 );
not ( n69066 , n69064 );
not ( n69067 , n69004 );
nor ( n69068 , n69067 , n68875 );
and ( n69069 , n69068 , n69001 );
not ( n69070 , n69068 );
not ( n69071 , n69001 );
and ( n69072 , n69070 , n69071 );
nor ( n69073 , n69069 , n69072 );
and ( n69074 , n69066 , n69073 );
nor ( n69075 , n69065 , n69074 );
not ( n69076 , n69075 );
not ( n69077 , n69076 );
not ( n69078 , n69020 );
not ( n69079 , n68884 );
or ( n69080 , n69078 , n69079 );
or ( n69081 , n69020 , n68884 );
nand ( n69082 , n69080 , n69081 );
and ( n69083 , n2703 , n69082 );
not ( n69084 , n2703 );
and ( n69085 , n69084 , n68852 );
nor ( n69086 , n69083 , n69085 );
not ( n69087 , n69086 );
not ( n69088 , n69087 );
not ( n69089 , n2703 );
not ( n69090 , n69004 );
not ( n69091 , n68875 );
or ( n69092 , n69090 , n69091 );
or ( n69093 , n68875 , n69004 );
nand ( n69094 , n69092 , n69093 );
not ( n69095 , n69094 );
or ( n69096 , n69089 , n69095 );
not ( n69097 , n2703 );
nand ( n69098 , n69097 , n68879 );
nand ( n69099 , n69096 , n69098 );
not ( n69100 , n2703 );
not ( n69101 , n69002 );
not ( n69102 , n69101 );
not ( n69103 , n69003 );
or ( n69104 , n69102 , n69103 );
or ( n69105 , n69101 , n69003 );
nand ( n69106 , n69104 , n69105 );
not ( n69107 , n69106 );
or ( n69108 , n69100 , n69107 );
nand ( n69109 , n69097 , n68873 );
nand ( n69110 , n69108 , n69109 );
not ( n69111 , n69110 );
not ( n69112 , n2728 );
nand ( n69113 , n69111 , n69112 );
nor ( n69114 , n69099 , n69113 );
nand ( n69115 , n69077 , n69088 , n69114 );
nor ( n69116 , n69063 , n69115 );
and ( n69117 , n69050 , n69116 );
not ( n69118 , n68848 );
nand ( n69119 , n68923 , n68892 );
and ( n69120 , n69119 , n2744 );
not ( n69121 , n69119 );
and ( n69122 , n69121 , n68888 );
nor ( n69123 , n69120 , n69122 );
not ( n69124 , n69123 );
or ( n69125 , n69118 , n69124 );
nand ( n69126 , n68847 , n2744 );
nand ( n69127 , n69125 , n69126 );
not ( n69128 , n69127 );
not ( n69129 , n68848 );
nand ( n69130 , n68897 , n68867 );
nand ( n69131 , n68895 , n68862 );
nor ( n69132 , n69130 , n69131 );
not ( n69133 , n68875 );
nor ( n69134 , n68891 , n68852 );
nand ( n69135 , n69132 , n69133 , n69134 );
nor ( n69136 , n68879 , n2758 );
nor ( n69137 , n68924 , n68882 );
nor ( n69138 , n2774 , n2784 );
nor ( n69139 , n2744 , n68855 );
nand ( n69140 , n69136 , n69137 , n69138 , n69139 );
nor ( n69141 , n69135 , n69140 );
buf ( n69142 , n49 );
buf ( n3000 , n48 );
not ( n69144 , n3000 );
not ( n69145 , n69144 );
nor ( n69146 , n69142 , n69145 );
not ( n69147 , n69146 );
not ( n69148 , n69147 );
nand ( n69149 , n69141 , n69148 );
buf ( n69150 , n50 );
not ( n69151 , n69150 );
not ( n69152 , n69151 );
and ( n69153 , n69149 , n69152 );
not ( n69154 , n69149 );
not ( n69155 , n69152 );
and ( n69156 , n69154 , n69155 );
nor ( n69157 , n69153 , n69156 );
not ( n69158 , n69157 );
or ( n69159 , n69129 , n69158 );
nand ( n69160 , n68847 , n69152 );
nand ( n69161 , n69159 , n69160 );
not ( n69162 , n69161 );
and ( n69163 , n69128 , n69162 );
not ( n69164 , n68848 );
not ( n69165 , n69141 );
nor ( n69166 , n69165 , n69145 );
or ( n69167 , n69166 , n69142 );
nand ( n69168 , n69137 , n69138 , n69134 , n69139 );
not ( n69169 , n69168 );
not ( n69170 , n69132 );
not ( n69171 , n69145 );
nand ( n69172 , n69171 , n69003 , n69002 , n69142 );
not ( n69173 , n69136 );
nor ( n69174 , n69170 , n69172 , n69173 );
nand ( n69175 , n69169 , n69174 );
nand ( n69176 , n69167 , n69175 );
not ( n69177 , n69176 );
or ( n69178 , n69164 , n69177 );
nand ( n69179 , n68847 , n69142 );
nand ( n69180 , n69178 , n69179 );
not ( n69181 , n69180 );
not ( n69182 , n69145 );
not ( n69183 , n68847 );
or ( n69184 , n69182 , n69183 );
not ( n69185 , n69145 );
not ( n69186 , n69141 );
or ( n69187 , n69185 , n69186 );
or ( n69188 , n69141 , n69145 );
nand ( n69189 , n69187 , n69188 );
nand ( n69190 , n69189 , n2703 );
nand ( n69191 , n69184 , n69190 );
not ( n69192 , n69191 );
and ( n69193 , n69181 , n69192 );
nand ( n69194 , n69117 , n69163 , n69193 );
not ( n69195 , n69194 );
and ( n69196 , n69035 , n69195 );
not ( n69197 , n69165 );
buf ( n69198 , n57 );
buf ( n69199 , n56 );
nor ( n69200 , n69198 , n69199 );
buf ( n3058 , n58 );
buf ( n3059 , n59 );
nor ( n69203 , n3058 , n3059 );
nand ( n69204 , n69200 , n69203 );
not ( n69205 , n69204 );
buf ( n69206 , n61 );
buf ( n69207 , n60 );
or ( n69208 , n69206 , n69207 );
buf ( n3066 , n62 );
nor ( n69210 , n69208 , n3066 );
nand ( n69211 , n69205 , n69210 );
buf ( n69212 , n53 );
not ( n69213 , n69212 );
not ( n69214 , n69213 );
buf ( n69215 , n51 );
nor ( n69216 , n69214 , n69215 );
buf ( n69217 , n54 );
nor ( n69218 , n69217 , n69145 );
buf ( n69219 , n55 );
nor ( n69220 , n69219 , n69142 );
buf ( n69221 , n52 );
not ( n69222 , n69221 );
not ( n69223 , n69222 );
nor ( n69224 , n69223 , n69152 );
nand ( n69225 , n69216 , n69218 , n69220 , n69224 );
nor ( n69226 , n69211 , n69225 );
nand ( n69227 , n69197 , n69226 );
and ( n69228 , n69227 , n2703 );
not ( n69229 , n69227 );
not ( n69230 , n2703 );
and ( n69231 , n69229 , n69230 );
nor ( n69232 , n69228 , n69231 );
nand ( n69233 , n69232 , n68848 );
not ( n69234 , n69233 );
not ( n69235 , n69234 );
nor ( n69236 , n69196 , n69235 );
not ( n69237 , n69215 );
not ( n69238 , n68847 );
or ( n69239 , n69237 , n69238 );
nor ( n69240 , n69147 , n69152 );
nand ( n69241 , n69141 , n69240 );
xor ( n69242 , n69241 , n69215 );
nand ( n69243 , n69242 , n68848 );
nand ( n69244 , n69239 , n69243 );
not ( n69245 , n69244 );
not ( n69246 , n68915 );
nor ( n69247 , n69152 , n69215 );
nand ( n69248 , n69146 , n69247 );
not ( n69249 , n69248 );
nand ( n69250 , n69249 , n69141 );
and ( n69251 , n69250 , n69223 );
not ( n69252 , n69250 );
not ( n69253 , n69223 );
and ( n69254 , n69252 , n69253 );
nor ( n69255 , n69251 , n69254 );
not ( n69256 , n69255 );
or ( n69257 , n69246 , n69256 );
not ( n69258 , n68848 );
nand ( n69259 , n69258 , n69223 );
nand ( n69260 , n69257 , n69259 );
not ( n69261 , n69260 );
not ( n69262 , n68915 );
nor ( n69263 , n69248 , n69223 );
nand ( n69264 , n69141 , n69263 );
xor ( n69265 , n69264 , n69214 );
not ( n69266 , n69265 );
or ( n69267 , n69262 , n69266 );
nand ( n69268 , n68847 , n69214 );
nand ( n69269 , n69267 , n69268 );
not ( n69270 , n69269 );
not ( n69271 , n68915 );
nor ( n69272 , n69214 , n69223 );
not ( n69273 , n69272 );
nor ( n69274 , n69273 , n69248 );
nand ( n69275 , n69141 , n69274 );
not ( n69276 , n69217 );
xnor ( n69277 , n69275 , n69276 );
not ( n69278 , n69277 );
or ( n69279 , n69271 , n69278 );
nand ( n69280 , n68847 , n69217 );
nand ( n69281 , n69279 , n69280 );
not ( n69282 , n69281 );
and ( n69283 , n69245 , n69261 , n69270 , n69282 );
not ( n69284 , n68848 );
nand ( n69285 , n69272 , n69276 );
nor ( n69286 , n69248 , n69285 );
nand ( n69287 , n69141 , n69286 );
not ( n69288 , n69219 );
xnor ( n69289 , n69287 , n69288 );
not ( n69290 , n69289 );
or ( n69291 , n69284 , n69290 );
nand ( n69292 , n69258 , n69219 );
nand ( n69293 , n69291 , n69292 );
not ( n69294 , n68915 );
nor ( n69295 , n69225 , n69199 );
nand ( n69296 , n69141 , n69295 );
not ( n69297 , n69198 );
xnor ( n69298 , n69296 , n69297 );
not ( n69299 , n69298 );
or ( n69300 , n69294 , n69299 );
nand ( n69301 , n68847 , n69198 );
nand ( n69302 , n69300 , n69301 );
not ( n69303 , n68915 );
not ( n69304 , n69199 );
not ( n69305 , n69304 );
not ( n69306 , n69225 );
nand ( n69307 , n69306 , n69141 );
not ( n69308 , n69307 );
or ( n69309 , n69305 , n69308 );
or ( n69310 , n69307 , n69304 );
nand ( n69311 , n69309 , n69310 );
not ( n69312 , n69311 );
or ( n69313 , n69303 , n69312 );
nand ( n69314 , n68847 , n69199 );
nand ( n69315 , n69313 , n69314 );
or ( n69316 , n69293 , n69302 , n69315 );
not ( n69317 , n68848 );
not ( n69318 , n69200 );
nor ( n69319 , n69318 , n69225 );
nand ( n69320 , n69141 , n69319 );
not ( n69321 , n3058 );
xnor ( n69322 , n69320 , n69321 );
not ( n69323 , n69322 );
not ( n69324 , n69323 );
not ( n69325 , n69324 );
or ( n69326 , n69317 , n69325 );
nand ( n69327 , n68847 , n3058 );
nand ( n69328 , n69326 , n69327 );
nor ( n69329 , n69316 , n69328 );
and ( n69330 , n69283 , n69329 );
nor ( n69331 , n69330 , n69235 );
nor ( n69332 , n69236 , n69331 );
not ( n69333 , n69332 );
not ( n69334 , n3059 );
not ( n69335 , n69258 );
or ( n69336 , n69334 , n69335 );
nand ( n69337 , n69200 , n69321 );
nor ( n69338 , n69225 , n69337 );
nand ( n69339 , n69141 , n69338 );
xor ( n69340 , n69339 , n3059 );
nand ( n69341 , n69340 , n68848 );
nand ( n69342 , n69336 , n69341 );
nand ( n69343 , n69333 , n69342 );
and ( n69344 , n68847 , n69207 );
not ( n69345 , n68847 );
nor ( n69346 , n69225 , n69204 );
nand ( n69347 , n69141 , n69346 );
not ( n69348 , n69207 );
not ( n69349 , n69348 );
and ( n69350 , n69347 , n69349 );
not ( n69351 , n69347 );
and ( n69352 , n69351 , n69348 );
nor ( n69353 , n69350 , n69352 );
and ( n69354 , n69345 , n69353 );
nor ( n69355 , n69344 , n69354 );
not ( n69356 , n69355 );
not ( n69357 , n69356 );
and ( n69358 , n69343 , n69357 );
not ( n69359 , n69343 );
and ( n69360 , n69359 , n69356 );
nor ( n69361 , n69358 , n69360 );
not ( n69362 , n69361 );
not ( n69363 , n69362 );
nand ( n69364 , n69190 , n69013 );
not ( n69365 , n69364 );
not ( n69366 , n68991 );
nand ( n69367 , n69062 , n69028 );
nor ( n69368 , n69366 , n69367 );
nor ( n69369 , n68934 , n69298 );
nand ( n69370 , n69365 , n69368 , n69369 );
nor ( n69371 , n69289 , n2728 );
nand ( n69372 , n69371 , n69323 , n69044 , n68907 );
nor ( n69373 , n69370 , n69372 );
nor ( n69374 , n69311 , n69265 );
nor ( n69375 , n69255 , n69157 );
nand ( n69376 , n69355 , n69341 , n69374 , n69375 );
not ( n69377 , n69376 );
not ( n69378 , n69123 );
nor ( n69379 , n69099 , n69110 );
and ( n69380 , n69086 , n69075 , n69379 );
nand ( n69381 , n69243 , n69378 , n68976 , n69380 );
nor ( n69382 , n68947 , n68961 );
nor ( n69383 , n69277 , n69176 );
nand ( n69384 , n69382 , n69383 );
nor ( n69385 , n69381 , n69384 );
nand ( n69386 , n69373 , n69377 , n69385 );
nand ( n69387 , n69205 , n69348 );
nor ( n69388 , n69387 , n69225 );
nand ( n69389 , n69197 , n69388 );
xor ( n69390 , n69389 , n69206 );
and ( n69391 , n69390 , n68915 );
and ( n69392 , n68847 , n69206 );
nor ( n69393 , n69391 , n69392 );
nor ( n69394 , n69393 , n69233 );
nand ( n69395 , n69386 , n69394 );
not ( n69396 , n69395 );
not ( n69397 , n69208 );
nand ( n69398 , n69397 , n69205 );
nor ( n69399 , n69398 , n69225 );
nand ( n69400 , n69197 , n69399 );
xor ( n69401 , n69400 , n3066 );
nand ( n69402 , n69401 , n68915 );
nand ( n69403 , n68847 , n3066 );
nand ( n69404 , n69402 , n69403 );
not ( n69405 , n69404 );
and ( n69406 , n69396 , n69405 );
and ( n69407 , n69395 , n69404 );
nor ( n69408 , n69406 , n69407 );
not ( n69409 , n69408 );
nand ( n69410 , n69386 , n69234 );
and ( n69411 , n69410 , n69393 );
not ( n69412 , n69410 );
not ( n69413 , n69393 );
and ( n69414 , n69412 , n69413 );
nor ( n69415 , n69411 , n69414 );
not ( n69416 , n69415 );
nand ( n69417 , n69409 , n69416 );
not ( n69418 , n69417 );
buf ( n3276 , n165 );
nand ( n69420 , n69418 , n3276 );
not ( n69421 , n69408 );
nor ( n69422 , n69416 , n69421 );
not ( n69423 , n69422 );
not ( n69424 , n69423 );
buf ( n3282 , n101 );
nand ( n69426 , n69424 , n3282 );
not ( n69427 , n69415 );
not ( n69428 , n69427 );
nand ( n69429 , n69409 , n69428 );
not ( n69430 , n69429 );
buf ( n3288 , n72 );
nand ( n69432 , n69430 , n3288 );
nand ( n69433 , n69408 , n69427 );
not ( n69434 , n69433 );
buf ( n3292 , n133 );
not ( n69436 , n3292 );
not ( n69437 , n69436 );
nand ( n69438 , n69434 , n69437 );
nand ( n69439 , n69420 , n69426 , n69432 , n69438 );
not ( n69440 , n69417 );
buf ( n69441 , n162 );
nand ( n69442 , n69440 , n69441 );
not ( n69443 , n69423 );
buf ( n3301 , n98 );
nand ( n69445 , n69443 , n3301 );
not ( n69446 , n69429 );
buf ( n3304 , n69 );
nand ( n69448 , n69446 , n3304 );
nand ( n69449 , n69408 , n69416 );
not ( n69450 , n69449 );
buf ( n69451 , n130 );
not ( n69452 , n69451 );
not ( n69453 , n69452 );
nand ( n69454 , n69450 , n69453 );
nand ( n69455 , n69442 , n69445 , n69448 , n69454 );
nand ( n69456 , n69439 , n69455 );
not ( n69457 , n69408 );
nor ( n69458 , n69457 , n69416 );
buf ( n3316 , n102 );
nand ( n69460 , n69458 , n3316 );
nand ( n69461 , n69421 , n69427 );
not ( n69462 , n69461 );
buf ( n3320 , n166 );
nand ( n69464 , n69462 , n3320 );
nand ( n69465 , n69428 , n69457 );
not ( n69466 , n69465 );
buf ( n3324 , n73 );
nand ( n69468 , n69466 , n3324 );
not ( n69469 , n69433 );
buf ( n3327 , n134 );
not ( n69471 , n3327 );
not ( n69472 , n69471 );
nand ( n69473 , n69469 , n69472 );
nand ( n69474 , n69460 , n69464 , n69468 , n69473 );
not ( n69475 , n69465 );
nand ( n69476 , n69474 , n69475 );
nor ( n69477 , n69456 , n69476 );
not ( n69478 , n69449 );
buf ( n3336 , n131 );
not ( n69480 , n3336 );
not ( n69481 , n69480 );
nand ( n69482 , n69478 , n69481 );
not ( n69483 , n69422 );
not ( n69484 , n69483 );
buf ( n3342 , n99 );
nand ( n69486 , n69484 , n3342 );
buf ( n3344 , n70 );
nand ( n69488 , n69430 , n3344 );
buf ( n3346 , n163 );
nand ( n69490 , n69418 , n3346 );
nand ( n69491 , n69482 , n69486 , n69488 , n69490 );
not ( n69492 , n69417 );
buf ( n3350 , n164 );
nand ( n69494 , n69492 , n3350 );
not ( n69495 , n69483 );
buf ( n69496 , n100 );
nand ( n69497 , n69495 , n69496 );
not ( n69498 , n69429 );
buf ( n3356 , n71 );
nand ( n69500 , n69498 , n3356 );
not ( n69501 , n69449 );
buf ( n3359 , n132 );
not ( n69503 , n3359 );
not ( n69504 , n69503 );
nand ( n69505 , n69501 , n69504 );
nand ( n69506 , n69494 , n69497 , n69500 , n69505 );
and ( n69507 , n69491 , n69506 );
nand ( n69508 , n69477 , n69507 );
not ( n69509 , n69508 );
not ( n69510 , n69461 );
buf ( n69511 , n170 );
nand ( n69512 , n69510 , n69511 );
buf ( n69513 , n106 );
nand ( n69514 , n69458 , n69513 );
not ( n69515 , n69465 );
buf ( n69516 , n77 );
nand ( n69517 , n69515 , n69516 );
not ( n69518 , n69433 );
buf ( n69519 , n138 );
not ( n69520 , n69519 );
not ( n69521 , n69520 );
nand ( n69522 , n69518 , n69521 );
nand ( n69523 , n69512 , n69514 , n69517 , n69522 );
buf ( n69524 , n76 );
nand ( n69525 , n69515 , n69524 );
buf ( n69526 , n169 );
nand ( n69527 , n69510 , n69526 );
buf ( n69528 , n105 );
nand ( n69529 , n69458 , n69528 );
not ( n69530 , n69433 );
buf ( n69531 , n137 );
not ( n69532 , n69531 );
not ( n69533 , n69532 );
nand ( n69534 , n69530 , n69533 );
nand ( n69535 , n69525 , n69527 , n69529 , n69534 );
nand ( n69536 , n69523 , n69535 );
buf ( n69537 , n168 );
nand ( n69538 , n69462 , n69537 );
buf ( n69539 , n104 );
nand ( n69540 , n69458 , n69539 );
buf ( n69541 , n75 );
nand ( n69542 , n69466 , n69541 );
buf ( n69543 , n136 );
not ( n69544 , n69543 );
not ( n69545 , n69544 );
nand ( n69546 , n69434 , n69545 );
nand ( n69547 , n69538 , n69540 , n69542 , n69546 );
buf ( n3405 , n167 );
nand ( n69549 , n69462 , n3405 );
buf ( n69550 , n103 );
nand ( n69551 , n69458 , n69550 );
not ( n69552 , n69465 );
buf ( n69553 , n74 );
nand ( n69554 , n69552 , n69553 );
buf ( n3412 , n135 );
nand ( n69556 , n69434 , n3412 );
nand ( n69557 , n69549 , n69551 , n69554 , n69556 );
nand ( n69558 , n69547 , n69557 );
nor ( n69559 , n69536 , n69558 );
not ( n69560 , n69461 );
not ( n69561 , n69560 );
buf ( n69562 , n172 );
not ( n69563 , n69562 );
nor ( n69564 , n69561 , n69563 );
not ( n69565 , n69458 );
buf ( n69566 , n108 );
not ( n69567 , n69566 );
nor ( n69568 , n69565 , n69567 );
nor ( n69569 , n69564 , n69568 );
not ( n69570 , n69465 );
buf ( n69571 , n79 );
and ( n69572 , n69570 , n69571 );
not ( n69573 , n69434 );
buf ( n69574 , n140 );
not ( n69575 , n69574 );
not ( n69576 , n69575 );
not ( n69577 , n69576 );
nor ( n69578 , n69573 , n69577 );
nor ( n69579 , n69572 , n69578 );
nand ( n69580 , n69569 , n69579 );
buf ( n69581 , n171 );
nand ( n69582 , n69510 , n69581 );
buf ( n69583 , n107 );
nand ( n69584 , n69458 , n69583 );
buf ( n3442 , n78 );
nand ( n69586 , n69515 , n3442 );
buf ( n69587 , n139 );
not ( n69588 , n69587 );
not ( n69589 , n69588 );
nand ( n69590 , n69530 , n69589 );
nand ( n69591 , n69582 , n69584 , n69586 , n69590 );
nand ( n69592 , n69580 , n69591 );
buf ( n3450 , n173 );
nand ( n69594 , n69560 , n3450 );
buf ( n69595 , n109 );
nand ( n69596 , n69458 , n69595 );
buf ( n3454 , n80 );
nand ( n69598 , n69430 , n3454 );
buf ( n69599 , n141 );
not ( n69600 , n69599 );
not ( n69601 , n69600 );
nand ( n69602 , n69478 , n69601 );
nand ( n69603 , n69594 , n69596 , n69598 , n69602 );
not ( n69604 , n69603 );
nor ( n69605 , n69592 , n69604 );
nand ( n69606 , n69509 , n69559 , n69605 );
buf ( n69607 , n81 );
nand ( n69608 , n69475 , n69607 );
buf ( n3466 , n174 );
nand ( n69610 , n69418 , n3466 );
buf ( n69611 , n110 );
nand ( n69612 , n69424 , n69611 );
buf ( n3470 , n142 );
not ( n69614 , n3470 );
not ( n69615 , n69614 );
nand ( n69616 , n69478 , n69615 );
nand ( n69617 , n69608 , n69610 , n69612 , n69616 );
not ( n69618 , n69617 );
and ( n69619 , n69606 , n69618 );
not ( n69620 , n69606 );
and ( n69621 , n69620 , n69617 );
nor ( n69622 , n69619 , n69621 );
not ( n69623 , n69622 );
not ( n69624 , n69623 );
and ( n69625 , n69363 , n69624 );
not ( n69626 , n69363 );
nand ( n69627 , n69506 , n69557 , n69491 , n69547 );
nor ( n69628 , n69627 , n69592 );
nand ( n69629 , n69617 , n69603 );
nor ( n69630 , n69536 , n69629 );
and ( n69631 , n69628 , n69630 , n69477 );
buf ( n3489 , n143 );
not ( n69633 , n3489 );
not ( n69634 , n69633 );
nand ( n69635 , n69530 , n69634 );
not ( n69636 , n69462 );
not ( n69637 , n69636 );
nand ( n69638 , n69637 , n2697 );
not ( n69639 , n69458 );
not ( n69640 , n69639 );
buf ( n3498 , n111 );
nand ( n69642 , n69640 , n3498 );
buf ( n69643 , n82 );
nand ( n69644 , n69475 , n69643 );
nand ( n69645 , n69635 , n69638 , n69642 , n69644 );
nand ( n69646 , n69631 , n69645 );
buf ( n69647 , n144 );
not ( n69648 , n69647 );
not ( n69649 , n69648 );
nand ( n69650 , n69530 , n69649 );
not ( n69651 , n69458 );
not ( n69652 , n69651 );
buf ( n3510 , n112 );
nand ( n69654 , n69652 , n3510 );
buf ( n69655 , n176 );
nand ( n69656 , n69637 , n69655 );
buf ( n3514 , n83 );
nand ( n69658 , n69475 , n3514 );
nand ( n69659 , n69650 , n69654 , n69656 , n69658 );
not ( n69660 , n69659 );
and ( n69661 , n69646 , n69660 );
not ( n69662 , n69646 );
and ( n69663 , n69662 , n69659 );
nor ( n69664 , n69661 , n69663 );
not ( n69665 , n69664 );
not ( n69666 , n69565 );
buf ( n69667 , n121 );
not ( n69668 , n69667 );
not ( n69669 , n69668 );
and ( n69670 , n69666 , n69669 );
not ( n69671 , n69510 );
buf ( n3529 , n185 );
not ( n69673 , n3529 );
not ( n69674 , n69673 );
not ( n69675 , n69674 );
nor ( n69676 , n69671 , n69675 );
nor ( n69677 , n69670 , n69676 );
buf ( n69678 , n92 );
not ( n69679 , n69678 );
not ( n69680 , n69679 );
and ( n69681 , n69570 , n69680 );
not ( n69682 , n69434 );
buf ( n69683 , n153 );
not ( n69684 , n69683 );
not ( n69685 , n69684 );
not ( n69686 , n69685 );
nor ( n69687 , n69682 , n69686 );
nor ( n69688 , n69681 , n69687 );
nand ( n69689 , n69677 , n69688 );
buf ( n69690 , n186 );
not ( n69691 , n69690 );
not ( n69692 , n69691 );
not ( n69693 , n69692 );
nor ( n69694 , n69461 , n69693 );
buf ( n3552 , n122 );
not ( n69696 , n3552 );
not ( n69697 , n69696 );
not ( n69698 , n69697 );
nor ( n69699 , n69565 , n69698 );
nor ( n69700 , n69694 , n69699 );
buf ( n69701 , n154 );
not ( n69702 , n69701 );
nor ( n69703 , n69573 , n69702 );
buf ( n3561 , n93 );
not ( n69705 , n3561 );
not ( n69706 , n69705 );
not ( n69707 , n69706 );
nor ( n69708 , n69465 , n69707 );
nor ( n69709 , n69703 , n69708 );
nand ( n69710 , n69700 , n69709 );
nand ( n69711 , n69689 , n69710 );
buf ( n3569 , n187 );
not ( n69713 , n3569 );
not ( n69714 , n69713 );
not ( n69715 , n69714 );
nor ( n69716 , n69461 , n69715 );
buf ( n69717 , n123 );
not ( n69718 , n69717 );
not ( n69719 , n69718 );
not ( n69720 , n69719 );
nor ( n69721 , n69565 , n69720 );
nor ( n69722 , n69716 , n69721 );
buf ( n3580 , n94 );
not ( n69724 , n3580 );
not ( n69725 , n69724 );
and ( n69726 , n69570 , n69725 );
buf ( n3584 , n155 );
not ( n69728 , n3584 );
not ( n69729 , n69728 );
not ( n69730 , n69729 );
nor ( n69731 , n69682 , n69730 );
nor ( n69732 , n69726 , n69731 );
nand ( n69733 , n69722 , n69732 );
buf ( n3591 , n156 );
not ( n69735 , n3591 );
not ( n69736 , n69735 );
nand ( n69737 , n69530 , n69736 );
not ( n69738 , n69565 );
buf ( n69739 , n124 );
not ( n69740 , n69739 );
not ( n69741 , n69740 );
nand ( n69742 , n69738 , n69741 );
buf ( n69743 , n188 );
not ( n69744 , n69743 );
not ( n69745 , n69744 );
nand ( n69746 , n69510 , n69745 );
nand ( n69747 , n69737 , n69742 , n69746 );
nand ( n69748 , n69733 , n69747 );
nor ( n69749 , n69711 , n69748 );
not ( n69750 , n69561 );
buf ( n69751 , n182 );
not ( n69752 , n69751 );
not ( n69753 , n69752 );
not ( n69754 , n69753 );
not ( n69755 , n69754 );
and ( n69756 , n69750 , n69755 );
buf ( n69757 , n118 );
not ( n69758 , n69757 );
not ( n69759 , n69758 );
and ( n69760 , n69640 , n69759 );
nor ( n69761 , n69756 , n69760 );
not ( n69762 , n69433 );
buf ( n3620 , n150 );
not ( n69764 , n3620 );
not ( n69765 , n69764 );
not ( n69766 , n69765 );
not ( n69767 , n69766 );
and ( n69768 , n69762 , n69767 );
not ( n69769 , n69465 );
buf ( n69770 , n89 );
and ( n69771 , n69769 , n69770 );
nor ( n69772 , n69768 , n69771 );
nand ( n69773 , n69761 , n69772 );
buf ( n69774 , n88 );
not ( n69775 , n69774 );
not ( n69776 , n69775 );
not ( n69777 , n69776 );
nor ( n69778 , n69465 , n69777 );
buf ( n3636 , n117 );
not ( n69780 , n3636 );
not ( n69781 , n69780 );
not ( n69782 , n69781 );
nor ( n69783 , n69651 , n69782 );
nor ( n69784 , n69778 , n69783 );
buf ( n69785 , n181 );
not ( n69786 , n69785 );
not ( n69787 , n69786 );
not ( n69788 , n69787 );
nor ( n69789 , n69461 , n69788 );
buf ( n69790 , n149 );
not ( n69791 , n69790 );
not ( n69792 , n69791 );
not ( n69793 , n69792 );
nor ( n69794 , n69433 , n69793 );
nor ( n69795 , n69789 , n69794 );
nand ( n69796 , n69784 , n69795 );
nand ( n69797 , n69773 , n69796 );
buf ( n69798 , n146 );
not ( n69799 , n69798 );
not ( n69800 , n69799 );
nand ( n69801 , n69434 , n69800 );
buf ( n69802 , n178 );
nand ( n69803 , n69560 , n69802 );
buf ( n69804 , n114 );
nand ( n69805 , n69640 , n69804 );
buf ( n69806 , n85 );
nand ( n69807 , n69570 , n69806 );
nand ( n69808 , n69801 , n69803 , n69805 , n69807 );
not ( n69809 , n69636 );
buf ( n69810 , n177 );
not ( n69811 , n69810 );
not ( n69812 , n69811 );
and ( n69813 , n69809 , n69812 );
buf ( n69814 , n113 );
and ( n69815 , n69652 , n69814 );
nor ( n69816 , n69813 , n69815 );
buf ( n69817 , n145 );
not ( n69818 , n69817 );
not ( n69819 , n69818 );
not ( n69820 , n69819 );
nor ( n69821 , n69433 , n69820 );
buf ( n69822 , n84 );
not ( n69823 , n69822 );
nor ( n69824 , n69465 , n69823 );
nor ( n69825 , n69821 , n69824 );
nand ( n69826 , n69816 , n69825 );
nand ( n69827 , n69808 , n69826 );
nor ( n69828 , n69797 , n69827 );
nand ( n69829 , n69749 , n69828 );
nand ( n69830 , n69659 , n69645 );
not ( n69831 , n69830 );
not ( n69832 , n69461 );
buf ( n69833 , n184 );
not ( n69834 , n69833 );
not ( n69835 , n69834 );
not ( n69836 , n69835 );
not ( n69837 , n69836 );
and ( n69838 , n69832 , n69837 );
buf ( n69839 , n120 );
not ( n69840 , n69839 );
not ( n69841 , n69840 );
and ( n69842 , n69666 , n69841 );
nor ( n69843 , n69838 , n69842 );
buf ( n69844 , n152 );
not ( n69845 , n69844 );
not ( n69846 , n69845 );
not ( n69847 , n69846 );
nor ( n69848 , n69573 , n69847 );
not ( n69849 , n69570 );
buf ( n3707 , n91 );
not ( n69851 , n3707 );
nor ( n69852 , n69849 , n69851 );
nor ( n69853 , n69848 , n69852 );
nand ( n69854 , n69843 , n69853 );
buf ( n69855 , n86 );
not ( n69856 , n69855 );
nor ( n69857 , n69465 , n69856 );
buf ( n69858 , n115 );
not ( n69859 , n69858 );
not ( n69860 , n69859 );
not ( n69861 , n69860 );
nor ( n69862 , n69639 , n69861 );
nor ( n69863 , n69857 , n69862 );
buf ( n3721 , n179 );
not ( n69865 , n3721 );
not ( n69866 , n69865 );
not ( n69867 , n69866 );
nor ( n69868 , n69461 , n69867 );
buf ( n69869 , n147 );
not ( n69870 , n69869 );
not ( n69871 , n69870 );
not ( n69872 , n69871 );
nor ( n69873 , n69433 , n69872 );
nor ( n69874 , n69868 , n69873 );
nand ( n69875 , n69863 , n69874 );
and ( n69876 , n69854 , n69875 );
not ( n69877 , n69461 );
buf ( n69878 , n180 );
not ( n69879 , n69878 );
not ( n69880 , n69879 );
not ( n69881 , n69880 );
not ( n69882 , n69881 );
and ( n69883 , n69877 , n69882 );
buf ( n69884 , n116 );
not ( n69885 , n69884 );
not ( n69886 , n69885 );
and ( n69887 , n69640 , n69886 );
nor ( n69888 , n69883 , n69887 );
buf ( n69889 , n87 );
not ( n69890 , n69889 );
not ( n69891 , n69890 );
not ( n69892 , n69891 );
nor ( n69893 , n69465 , n69892 );
buf ( n69894 , n148 );
not ( n69895 , n69894 );
not ( n69896 , n69895 );
not ( n69897 , n69896 );
nor ( n69898 , n69433 , n69897 );
nor ( n69899 , n69893 , n69898 );
nand ( n69900 , n69888 , n69899 );
buf ( n69901 , n125 );
not ( n69902 , n69901 );
not ( n69903 , n69902 );
nand ( n69904 , n69666 , n69903 );
not ( n69905 , n69461 );
buf ( n69906 , n189 );
nand ( n69907 , n69905 , n69906 );
buf ( n69908 , n157 );
not ( n69909 , n69908 );
not ( n69910 , n69909 );
nand ( n69911 , n69530 , n69910 );
nand ( n69912 , n69904 , n69907 , n69911 );
and ( n69913 , n69900 , n69912 );
buf ( n3771 , n119 );
not ( n69915 , n3771 );
not ( n69916 , n69915 );
and ( n69917 , n69738 , n69916 );
buf ( n69918 , n183 );
not ( n69919 , n69918 );
not ( n69920 , n69919 );
not ( n69921 , n69920 );
nor ( n69922 , n69671 , n69921 );
nor ( n69923 , n69917 , n69922 );
not ( n69924 , n69530 );
buf ( n69925 , n151 );
not ( n69926 , n69925 );
not ( n69927 , n69926 );
not ( n69928 , n69927 );
nor ( n69929 , n69924 , n69928 );
buf ( n69930 , n90 );
not ( n69931 , n69930 );
not ( n69932 , n69931 );
not ( n69933 , n69932 );
nor ( n69934 , n69465 , n69933 );
nor ( n69935 , n69929 , n69934 );
nand ( n69936 , n69923 , n69935 );
nand ( n69937 , n69831 , n69876 , n69913 , n69936 );
nor ( n69938 , n69829 , n69937 );
nand ( n69939 , n69631 , n69938 );
buf ( n69940 , n126 );
nand ( n69941 , n69738 , n69940 );
buf ( n3799 , n158 );
nand ( n69943 , n69530 , n3799 );
buf ( n69944 , n190 );
nand ( n69945 , n69510 , n69944 );
nand ( n69946 , n69941 , n69943 , n69945 );
not ( n69947 , n69946 );
and ( n69948 , n69939 , n69947 );
not ( n69949 , n69939 );
and ( n69950 , n69949 , n69946 );
nor ( n69951 , n69948 , n69950 );
buf ( n69952 , n66 );
not ( n69953 , n69952 );
not ( n69954 , n69953 );
not ( n69955 , n69954 );
not ( n69956 , n69475 );
or ( n69957 , n69955 , n69956 );
buf ( n3815 , n159 );
nand ( n69959 , n69905 , n3815 );
nand ( n69960 , n69957 , n69959 );
buf ( n69961 , n95 );
not ( n69962 , n69961 );
not ( n69963 , n69640 );
or ( n69964 , n69962 , n69963 );
buf ( n69965 , n127 );
not ( n69966 , n69965 );
not ( n69967 , n69966 );
nand ( n69968 , n69434 , n69967 );
nand ( n69969 , n69964 , n69968 );
nor ( n69970 , n69960 , n69969 );
not ( n69971 , n69970 );
nand ( n69972 , n69951 , n69971 );
not ( n69973 , n69972 );
not ( n69974 , n69973 );
not ( n69975 , n69974 );
not ( n69976 , n69645 );
not ( n69977 , n69631 );
not ( n69978 , n69977 );
or ( n69979 , n69976 , n69978 );
or ( n69980 , n69977 , n69645 );
nand ( n69981 , n69979 , n69980 );
not ( n69982 , n69981 );
not ( n69983 , n69592 );
nand ( n69984 , n69983 , n69509 , n69559 );
xor ( n69985 , n69984 , n69604 );
nand ( n69986 , n69622 , n69985 );
nor ( n69987 , n69982 , n69986 );
not ( n69988 , n69987 );
nand ( n69989 , n69509 , n69559 );
not ( n69990 , n69591 );
and ( n69991 , n69989 , n69990 );
not ( n69992 , n69989 );
and ( n69993 , n69992 , n69591 );
nor ( n69994 , n69991 , n69993 );
not ( n69995 , n69558 );
not ( n69996 , n69995 );
not ( n69997 , n69535 );
nor ( n69998 , n69996 , n69997 );
nand ( n69999 , n69509 , n69998 );
not ( n70000 , n69523 );
and ( n70001 , n69999 , n70000 );
not ( n70002 , n69999 );
and ( n70003 , n70002 , n69523 );
nor ( n70004 , n70001 , n70003 );
nand ( n70005 , n69994 , n70004 );
nand ( n70006 , n69509 , n69557 );
not ( n70007 , n69547 );
and ( n70008 , n70006 , n70007 );
not ( n70009 , n70006 );
and ( n70010 , n70009 , n69547 );
nor ( n70011 , n70008 , n70010 );
nand ( n70012 , n69509 , n69995 );
not ( n70013 , n69535 );
and ( n70014 , n70012 , n70013 );
not ( n70015 , n70012 );
and ( n70016 , n70015 , n69535 );
nor ( n70017 , n70014 , n70016 );
and ( n70018 , n70011 , n70017 );
not ( n70019 , n70018 );
nor ( n70020 , n70005 , n70019 );
nand ( n70021 , n69455 , n69475 );
not ( n70022 , n69491 );
or ( n70023 , n70021 , n70022 );
not ( n70024 , n69506 );
and ( n70025 , n70023 , n70024 );
not ( n70026 , n70023 );
and ( n70027 , n70026 , n69506 );
nor ( n70028 , n70025 , n70027 );
not ( n70029 , n69507 );
or ( n70030 , n70021 , n70029 );
not ( n70031 , n69439 );
and ( n70032 , n70030 , n70031 );
not ( n70033 , n70030 );
and ( n70034 , n70033 , n69439 );
nor ( n70035 , n70032 , n70034 );
nand ( n70036 , n70028 , n70035 );
not ( n70037 , n69491 );
nand ( n70038 , n69455 , n69475 );
not ( n70039 , n70038 );
or ( n70040 , n70037 , n70039 );
or ( n70041 , n70038 , n69491 );
nand ( n70042 , n70040 , n70041 );
or ( n70043 , n69455 , n69475 );
and ( n70044 , n70038 , n70043 );
buf ( n70045 , n67 );
nand ( n70046 , n69475 , n70045 );
buf ( n70047 , n128 );
not ( n70048 , n70047 );
not ( n70049 , n70048 );
nand ( n70050 , n69434 , n70049 );
buf ( n70051 , n96 );
not ( n70052 , n70051 );
not ( n70053 , n70052 );
nand ( n70054 , n69640 , n70053 );
buf ( n70055 , n160 );
nand ( n70056 , n69905 , n70055 );
nand ( n70057 , n70046 , n70050 , n70054 , n70056 );
buf ( n70058 , n68 );
not ( n70059 , n70058 );
not ( n70060 , n69475 );
or ( n70061 , n70059 , n70060 );
buf ( n70062 , n161 );
nand ( n70063 , n69905 , n70062 );
nand ( n70064 , n70061 , n70063 );
buf ( n70065 , n129 );
not ( n70066 , n70065 );
not ( n70067 , n70066 );
not ( n70068 , n70067 );
not ( n70069 , n69434 );
or ( n70070 , n70068 , n70069 );
buf ( n70071 , n97 );
not ( n70072 , n70071 );
not ( n70073 , n70072 );
nand ( n70074 , n69640 , n70073 );
nand ( n70075 , n70070 , n70074 );
nor ( n70076 , n70064 , n70075 );
not ( n70077 , n70076 );
and ( n70078 , n70057 , n70077 );
nand ( n70079 , n70042 , n70044 , n70078 );
nor ( n70080 , n70036 , n70079 );
not ( n70081 , n69557 );
not ( n70082 , n69509 );
not ( n70083 , n70082 );
or ( n70084 , n70081 , n70083 );
or ( n70085 , n70082 , n69557 );
nand ( n70086 , n70084 , n70085 );
not ( n70087 , n69474 );
not ( n70088 , n70038 );
nor ( n70089 , n70029 , n70031 );
nand ( n70090 , n70088 , n70089 );
not ( n70091 , n70090 );
or ( n70092 , n70087 , n70091 );
or ( n70093 , n70090 , n69474 );
nand ( n70094 , n70092 , n70093 );
nand ( n70095 , n70080 , n70086 , n70094 );
not ( n70096 , n70095 );
nand ( n70097 , n69509 , n69559 , n69591 );
not ( n70098 , n69580 );
and ( n70099 , n70097 , n70098 );
not ( n70100 , n70097 );
and ( n70101 , n70100 , n69580 );
nor ( n70102 , n70099 , n70101 );
nand ( n70103 , n70020 , n70096 , n70102 );
not ( n70104 , n70103 );
not ( n70105 , n70104 );
nor ( n70106 , n69988 , n70105 );
nand ( n70107 , n69975 , n70106 );
not ( n70108 , n70107 );
or ( n70109 , n69665 , n70108 );
or ( n70110 , n70107 , n69664 );
nand ( n70111 , n70109 , n70110 );
and ( n70112 , n69626 , n70111 );
nor ( n70113 , n69625 , n70112 );
not ( n70114 , n69302 );
not ( n70115 , n69293 );
not ( n70116 , n69234 );
or ( n70117 , n70115 , n70116 );
not ( n70118 , n69034 );
not ( n70119 , n69194 );
and ( n70120 , n70118 , n70119 );
nor ( n70121 , n70120 , n69235 );
nor ( n70122 , n69283 , n69235 );
nor ( n70123 , n70121 , n70122 );
nand ( n70124 , n70117 , n70123 );
nand ( n70125 , n70124 , n69315 );
nor ( n70126 , n70114 , n70125 );
xor ( n70127 , n70126 , n69328 );
not ( n70128 , n70125 );
not ( n70129 , n69302 );
and ( n70130 , n70128 , n70129 );
and ( n70131 , n70125 , n69302 );
nor ( n70132 , n70130 , n70131 );
and ( n70133 , n70124 , n69315 );
not ( n70134 , n70124 );
not ( n70135 , n69315 );
and ( n70136 , n70134 , n70135 );
nor ( n70137 , n70133 , n70136 );
not ( n70138 , n70137 );
nor ( n70139 , n70132 , n70138 );
nand ( n70140 , n70127 , n70139 );
buf ( n3998 , DFF_state_reg_Q);
not ( n70142 , n3998 );
not ( n70143 , n70142 );
and ( n70144 , n70140 , n70143 );
not ( n70145 , n70144 );
not ( n70146 , n70123 );
not ( n70147 , n69293 );
and ( n70148 , n70146 , n70147 );
and ( n70149 , n70123 , n69293 );
nor ( n70150 , n70148 , n70149 );
not ( n70151 , n70150 );
nor ( n70152 , n70145 , n70151 );
not ( n70153 , n70132 );
not ( n70154 , n70153 );
buf ( n4012 , DFF_B_reg_Q);
not ( n70156 , n4012 );
nand ( n70157 , n70154 , n70156 );
not ( n70158 , n70157 );
not ( n70159 , n70127 );
or ( n70160 , n70158 , n70159 );
nand ( n70161 , n70160 , n70137 );
not ( n70162 , n70137 );
nand ( n70163 , n70162 , n4012 );
nor ( n70164 , n70153 , n70163 );
buf ( n4022 , n64 );
or ( n70166 , n70164 , n4022 );
nand ( n70167 , n70166 , n70127 );
nand ( n70168 , n70161 , n70167 );
not ( n70169 , n70153 );
not ( n70170 , n70127 );
not ( n70171 , n70170 );
or ( n70172 , n70169 , n70171 );
buf ( n4030 , n65 );
not ( n70174 , n4030 );
not ( n70175 , n70174 );
nand ( n70176 , n70137 , n70156 );
not ( n70177 , n70176 );
not ( n70178 , n70163 );
or ( n70179 , n70177 , n70178 );
nand ( n70180 , n70179 , n70154 );
not ( n70181 , n70180 );
or ( n70182 , n70175 , n70181 );
nand ( n70183 , n70182 , n70127 );
nand ( n70184 , n70172 , n70183 );
not ( n70185 , n70184 );
nor ( n70186 , n70168 , n70185 );
nand ( n70187 , n70152 , n70186 );
not ( n70188 , n69245 );
nand ( n70189 , n70121 , n70188 );
nor ( n70190 , n70189 , n69261 );
nand ( n70191 , n70190 , n69269 );
xor ( n70192 , n70191 , n69282 );
not ( n70193 , n69269 );
nor ( n70194 , n70193 , n70190 );
not ( n70195 , n70194 );
not ( n70196 , n69269 );
nand ( n70197 , n70196 , n70190 );
nand ( n70198 , n70195 , n70197 );
nand ( n70199 , n70192 , n70198 );
not ( n70200 , n70199 );
not ( n70201 , n69261 );
not ( n70202 , n70201 );
not ( n70203 , n70189 );
or ( n70204 , n70202 , n70203 );
or ( n70205 , n70189 , n70201 );
nand ( n70206 , n70204 , n70205 );
and ( n70207 , n70121 , n70188 );
not ( n70208 , n70121 );
and ( n70209 , n70208 , n69245 );
nor ( n70210 , n70207 , n70209 );
nor ( n70211 , n70206 , n70210 );
nand ( n70212 , n70200 , n70211 );
nor ( n70213 , n70187 , n70212 );
not ( n70214 , n70213 );
or ( n70215 , n70113 , n70214 );
not ( n70216 , n69645 );
not ( n70217 , n69332 );
not ( n70218 , n69342 );
and ( n70219 , n70217 , n70218 );
and ( n70220 , n69332 , n69342 );
nor ( n70221 , n70219 , n70220 );
and ( n70222 , n69342 , n69357 );
not ( n70223 , n69342 );
and ( n70224 , n70223 , n69356 );
nor ( n70225 , n70222 , n70224 );
nand ( n70226 , n70221 , n70225 );
or ( n70227 , n70226 , n69192 );
nand ( n70228 , n70226 , n68655 );
nand ( n70229 , n70227 , n70228 );
not ( n70230 , n70229 );
or ( n70231 , n70216 , n70230 );
not ( n70232 , n69645 );
not ( n70233 , n70229 );
nand ( n70234 , n70232 , n70233 );
nand ( n70235 , n70231 , n70234 );
not ( n70236 , n70226 );
not ( n70237 , n68938 );
not ( n70238 , n70237 );
and ( n70239 , n70236 , n70238 );
and ( n70240 , n70226 , n2513 );
nor ( n70241 , n70239 , n70240 );
not ( n70242 , n70241 );
not ( n70243 , n70242 );
and ( n70244 , n70243 , n69617 );
nor ( n70245 , n70235 , n70244 );
not ( n70246 , n70245 );
nand ( n70247 , n70235 , n70244 );
nand ( n70248 , n70246 , n70247 );
not ( n70249 , n70248 );
not ( n70250 , n69535 );
not ( n70251 , n70226 );
not ( n70252 , n69049 );
not ( n70253 , n70252 );
and ( n70254 , n70251 , n70253 );
and ( n70255 , n70226 , n2518 );
nor ( n70256 , n70254 , n70255 );
not ( n70257 , n70256 );
not ( n70258 , n70257 );
or ( n70259 , n70250 , n70258 );
not ( n70260 , n70257 );
not ( n70261 , n69535 );
nand ( n70262 , n70260 , n70261 );
nand ( n70263 , n70259 , n70262 );
nor ( n70264 , n70226 , n69128 );
not ( n70265 , n70264 );
nand ( n70266 , n70226 , n2519 );
nand ( n70267 , n70265 , n70266 );
not ( n70268 , n70267 );
and ( n70269 , n69547 , n70268 );
and ( n70270 , n70263 , n70269 );
not ( n70271 , n70270 );
not ( n70272 , n70226 );
not ( n70273 , n68982 );
and ( n70274 , n70272 , n70273 );
and ( n70275 , n70226 , n2517 );
nor ( n70276 , n70274 , n70275 );
not ( n70277 , n70276 );
not ( n70278 , n70277 );
not ( n70279 , n69523 );
or ( n70280 , n70278 , n70279 );
not ( n70281 , n70277 );
not ( n70282 , n69523 );
nand ( n70283 , n70281 , n70282 );
nand ( n70284 , n70280 , n70283 );
nor ( n70285 , n70257 , n70261 );
nor ( n70286 , n70284 , n70285 );
not ( n70287 , n70286 );
not ( n70288 , n70287 );
or ( n70289 , n70271 , n70288 );
nand ( n70290 , n70284 , n70285 );
nand ( n70291 , n70289 , n70290 );
not ( n70292 , n70291 );
not ( n70293 , n69580 );
not ( n70294 , n70293 );
not ( n70295 , n70226 );
not ( n70296 , n68952 );
and ( n70297 , n70295 , n70296 );
and ( n70298 , n70226 , n2515 );
nor ( n70299 , n70297 , n70298 );
not ( n70300 , n70299 );
not ( n70301 , n70300 );
not ( n70302 , n70301 );
or ( n70303 , n70294 , n70302 );
nand ( n70304 , n69580 , n70300 );
nand ( n70305 , n70303 , n70304 );
not ( n70306 , n69591 );
not ( n70307 , n70226 );
not ( n70308 , n68913 );
and ( n70309 , n70307 , n70308 );
and ( n70310 , n70226 , n2516 );
nor ( n70311 , n70309 , n70310 );
not ( n70312 , n70311 );
nor ( n70313 , n70306 , n70312 );
nor ( n70314 , n70305 , n70313 );
not ( n70315 , n69591 );
not ( n70316 , n70312 );
or ( n70317 , n70315 , n70316 );
not ( n70318 , n70312 );
not ( n70319 , n69591 );
nand ( n70320 , n70318 , n70319 );
nand ( n70321 , n70317 , n70320 );
nand ( n70322 , n69523 , n70281 );
not ( n70323 , n70322 );
nor ( n70324 , n70321 , n70323 );
nor ( n70325 , n70314 , n70324 );
not ( n70326 , n69603 );
not ( n70327 , n68965 );
nor ( n70328 , n70226 , n70327 );
not ( n70329 , n70328 );
nand ( n70330 , n70226 , n2514 );
nand ( n70331 , n70329 , n70330 );
not ( n70332 , n70331 );
or ( n70333 , n70326 , n70332 );
not ( n70334 , n69603 );
not ( n70335 , n70331 );
nand ( n70336 , n70334 , n70335 );
nand ( n70337 , n70333 , n70336 );
not ( n70338 , n69580 );
nor ( n70339 , n70338 , n70300 );
nor ( n70340 , n70337 , n70339 );
not ( n70341 , n69617 );
not ( n70342 , n70242 );
or ( n70343 , n70341 , n70342 );
not ( n70344 , n69617 );
nand ( n70345 , n70344 , n70243 );
nand ( n70346 , n70343 , n70345 );
nand ( n70347 , n70335 , n69603 );
not ( n70348 , n70347 );
nor ( n70349 , n70346 , n70348 );
nor ( n70350 , n70340 , n70349 );
and ( n70351 , n70325 , n70350 );
not ( n70352 , n70351 );
or ( n70353 , n70292 , n70352 );
not ( n70354 , n70350 );
nand ( n70355 , n70321 , n70323 );
not ( n70356 , n70355 );
not ( n70357 , n70356 );
not ( n70358 , n70314 );
not ( n70359 , n70358 );
or ( n70360 , n70357 , n70359 );
nand ( n70361 , n70305 , n70313 );
nand ( n70362 , n70360 , n70361 );
not ( n70363 , n70362 );
or ( n70364 , n70354 , n70363 );
not ( n70365 , n70349 );
nand ( n70366 , n70337 , n70339 );
not ( n70367 , n70366 );
and ( n70368 , n70365 , n70367 );
nand ( n70369 , n70346 , n70348 );
not ( n70370 , n70369 );
nor ( n70371 , n70368 , n70370 );
nand ( n70372 , n70364 , n70371 );
not ( n70373 , n70372 );
nand ( n70374 , n70353 , n70373 );
not ( n70375 , n70374 );
nor ( n70376 , n70263 , n70269 );
nor ( n70377 , n70376 , n70286 );
not ( n70378 , n69557 );
not ( n70379 , n68992 );
or ( n70380 , n70226 , n70379 );
nand ( n70381 , n70226 , n68663 );
nand ( n70382 , n70380 , n70381 );
not ( n70383 , n70382 );
or ( n70384 , n70378 , n70383 );
not ( n70385 , n70382 );
not ( n70386 , n69557 );
nand ( n70387 , n70385 , n70386 );
nand ( n70388 , n70384 , n70387 );
not ( n70389 , n70388 );
or ( n70390 , n70226 , n69015 );
nand ( n70391 , n70226 , n68664 );
nand ( n70392 , n70390 , n70391 );
not ( n70393 , n69474 );
nor ( n70394 , n70392 , n70393 );
not ( n70395 , n70394 );
nand ( n70396 , n70389 , n70395 );
xor ( n70397 , n69547 , n70268 );
not ( n70398 , n70397 );
nor ( n70399 , n70382 , n70386 );
not ( n70400 , n70399 );
nand ( n70401 , n70398 , n70400 );
and ( n70402 , n70396 , n70401 );
not ( n70403 , n69491 );
not ( n70404 , n70226 );
not ( n70405 , n69088 );
and ( n70406 , n70404 , n70405 );
and ( n70407 , n70226 , n2524 );
nor ( n70408 , n70406 , n70407 );
not ( n70409 , n70408 );
not ( n70410 , n70409 );
or ( n70411 , n70403 , n70410 );
or ( n70412 , n70409 , n69491 );
nand ( n70413 , n70411 , n70412 );
not ( n70414 , n69475 );
not ( n70415 , n70414 );
not ( n70416 , n69455 );
not ( n70417 , n70416 );
or ( n70418 , n70415 , n70417 );
not ( n70419 , n69076 );
not ( n70420 , n70226 );
not ( n70421 , n70420 );
or ( n70422 , n70419 , n70421 );
nand ( n70423 , n70226 , n68668 );
nand ( n70424 , n70422 , n70423 );
not ( n70425 , n70424 );
nand ( n70426 , n70418 , n70425 );
not ( n70427 , n70416 );
nand ( n70428 , n70427 , n69475 );
nand ( n70429 , n70426 , n70428 );
nor ( n70430 , n70413 , n70429 );
not ( n70431 , n69506 );
not ( n70432 , n69029 );
not ( n70433 , n70420 );
or ( n70434 , n70432 , n70433 );
nand ( n70435 , n70226 , n2523 );
nand ( n70436 , n70434 , n70435 );
not ( n70437 , n70436 );
or ( n70438 , n70431 , n70437 );
not ( n70439 , n70436 );
not ( n70440 , n69506 );
nand ( n70441 , n70439 , n70440 );
nand ( n70442 , n70438 , n70441 );
not ( n70443 , n69491 );
nor ( n70444 , n70443 , n70409 );
nor ( n70445 , n70442 , n70444 );
nor ( n70446 , n70430 , n70445 );
not ( n70447 , n69475 );
not ( n70448 , n69455 );
not ( n70449 , n70448 );
or ( n70450 , n70447 , n70449 );
nand ( n70451 , n69455 , n70414 );
nand ( n70452 , n70450 , n70451 );
and ( n70453 , n70452 , n70425 );
not ( n70454 , n70452 );
and ( n70455 , n70454 , n70424 );
nor ( n70456 , n70453 , n70455 );
not ( n70457 , n70226 );
not ( n70458 , n69099 );
not ( n70459 , n70458 );
and ( n70460 , n70457 , n70459 );
and ( n70461 , n70226 , n68669 );
nor ( n70462 , n70460 , n70461 );
not ( n70463 , n70462 );
not ( n70464 , n70463 );
and ( n70465 , n70077 , n70464 );
nor ( n70466 , n70456 , n70465 );
not ( n70467 , n70466 );
and ( n70468 , n70377 , n70402 , n70446 , n70467 );
not ( n70469 , n70393 );
not ( n70470 , n70392 );
not ( n70471 , n70470 );
or ( n70472 , n70469 , n70471 );
nand ( n70473 , n70392 , n69474 );
nand ( n70474 , n70472 , n70473 );
not ( n70475 , n70226 );
not ( n70476 , n69063 );
not ( n70477 , n70476 );
and ( n70478 , n70475 , n70477 );
and ( n70479 , n70226 , n68665 );
nor ( n70480 , n70478 , n70479 );
not ( n70481 , n70480 );
not ( n70482 , n69439 );
nor ( n70483 , n70481 , n70482 );
nor ( n70484 , n70474 , n70483 );
not ( n70485 , n69439 );
not ( n70486 , n70481 );
or ( n70487 , n70485 , n70486 );
not ( n70488 , n70481 );
nand ( n70489 , n70488 , n70482 );
nand ( n70490 , n70487 , n70489 );
nor ( n70491 , n70436 , n70440 );
nand ( n70492 , n70490 , n70491 );
nor ( n70493 , n70484 , n70492 );
and ( n70494 , n70474 , n70483 );
nor ( n70495 , n70493 , n70494 );
or ( n70496 , n70474 , n70483 );
not ( n70497 , n70490 );
not ( n70498 , n70491 );
nand ( n70499 , n70497 , n70498 );
nand ( n70500 , n70496 , n70499 );
nand ( n70501 , n70495 , n70500 );
not ( n70502 , n70226 );
not ( n70503 , n69111 );
and ( n70504 , n70502 , n70503 );
and ( n70505 , n70226 , n68670 );
nor ( n70506 , n70504 , n70505 );
not ( n70507 , n70506 );
or ( n70508 , n70507 , n70057 );
nand ( n70509 , n70057 , n70507 );
nand ( n70510 , n70508 , n70509 );
nor ( n70511 , n70510 , n69971 );
not ( n70512 , n70464 );
not ( n70513 , n70077 );
not ( n70514 , n70513 );
or ( n70515 , n70512 , n70514 );
nand ( n70516 , n70077 , n70463 );
nand ( n70517 , n70515 , n70516 );
not ( n70518 , n70057 );
nor ( n70519 , n70518 , n70507 );
nor ( n70520 , n70517 , n70519 );
nor ( n70521 , n70511 , n70520 );
nand ( n70522 , n70510 , n69971 );
not ( n70523 , n69971 );
or ( n70524 , n70226 , n69112 );
nand ( n70525 , n70226 , n2528 );
nand ( n70526 , n70524 , n70525 );
not ( n70527 , n70526 );
nand ( n70528 , n70523 , n70527 );
nand ( n70529 , n70522 , n70528 );
nand ( n70530 , n70521 , n70529 );
nand ( n70531 , n70456 , n70465 );
nand ( n70532 , n70517 , n70519 );
and ( n70533 , n70531 , n70532 );
nand ( n70534 , n70530 , n70533 );
nand ( n70535 , n70468 , n70501 , n70351 , n70534 );
not ( n70536 , n70376 );
and ( n70537 , n70536 , n70287 , n70396 , n70401 );
not ( n70538 , n70493 );
nand ( n70539 , n70429 , n70413 );
not ( n70540 , n70539 );
not ( n70541 , n70442 );
not ( n70542 , n70444 );
nand ( n70543 , n70541 , n70542 );
nand ( n70544 , n70540 , n70543 );
not ( n70545 , n70494 );
nand ( n70546 , n70442 , n70444 );
nand ( n70547 , n70538 , n70544 , n70545 , n70546 );
nand ( n70548 , n70351 , n70501 , n70537 , n70547 );
and ( n70549 , n70388 , n70394 );
not ( n70550 , n70549 );
not ( n70551 , n70401 );
or ( n70552 , n70550 , n70551 );
or ( n70553 , n70398 , n70400 );
nand ( n70554 , n70552 , n70553 );
and ( n70555 , n70554 , n70377 );
nand ( n70556 , n70351 , n70555 );
nand ( n70557 , n70375 , n70535 , n70548 , n70556 );
not ( n70558 , n70557 );
or ( n70559 , n70249 , n70558 );
or ( n70560 , n70557 , n70248 );
nand ( n70561 , n70559 , n70560 );
not ( n70562 , n70192 );
not ( n70563 , n70198 );
nand ( n70564 , n70562 , n70563 );
nand ( n70565 , n70564 , n70199 );
and ( n70566 , n70192 , n70210 );
not ( n70567 , n70192 );
and ( n70568 , n70567 , n70206 );
nor ( n70569 , n70566 , n70568 );
nor ( n70570 , n70565 , n70569 );
not ( n70571 , n70570 );
nor ( n70572 , n70571 , n70187 );
and ( n70573 , n70561 , n70572 );
not ( n70574 , n70569 );
nor ( n70575 , n70574 , n70565 );
not ( n70576 , n70575 );
nor ( n70577 , n70576 , n70187 );
not ( n70578 , n70577 );
not ( n70579 , n70229 );
not ( n70580 , n69645 );
not ( n70581 , n70580 );
or ( n70582 , n70579 , n70581 );
not ( n70583 , n70229 );
nand ( n70584 , n70583 , n69645 );
nand ( n70585 , n70582 , n70584 );
not ( n70586 , n70585 );
and ( n70587 , n69617 , n70242 );
not ( n70588 , n70587 );
nand ( n70589 , n70586 , n70588 );
nand ( n70590 , n70585 , n70587 );
and ( n70591 , n70589 , n70590 );
not ( n70592 , n70591 );
not ( n70593 , n69439 );
not ( n70594 , n70481 );
not ( n70595 , n70594 );
or ( n70596 , n70593 , n70595 );
not ( n70597 , n69439 );
nand ( n70598 , n70597 , n70481 );
nand ( n70599 , n70596 , n70598 );
and ( n70600 , n70436 , n69506 );
nand ( n70601 , n70599 , n70600 );
not ( n70602 , n70601 );
not ( n70603 , n69474 );
not ( n70604 , n70392 );
not ( n70605 , n70604 );
or ( n70606 , n70603 , n70605 );
not ( n70607 , n69474 );
nand ( n70608 , n70607 , n70392 );
nand ( n70609 , n70606 , n70608 );
nand ( n70610 , n70481 , n69439 );
not ( n70611 , n70610 );
nor ( n70612 , n70609 , n70611 );
not ( n70613 , n70612 );
and ( n70614 , n70602 , n70613 );
nand ( n70615 , n70609 , n70611 );
not ( n70616 , n70615 );
nor ( n70617 , n70614 , n70616 );
not ( n70618 , n70599 );
not ( n70619 , n70600 );
nand ( n70620 , n70618 , n70619 );
not ( n70621 , n70612 );
nand ( n70622 , n70620 , n70621 );
nand ( n70623 , n70617 , n70622 );
not ( n70624 , n69547 );
not ( n70625 , n70624 );
not ( n70626 , n70267 );
or ( n70627 , n70625 , n70626 );
not ( n70628 , n70267 );
nand ( n70629 , n70628 , n69547 );
nand ( n70630 , n70627 , n70629 );
not ( n70631 , n70630 );
and ( n70632 , n70382 , n69557 );
not ( n70633 , n70632 );
nand ( n70634 , n70631 , n70633 );
not ( n70635 , n69557 );
not ( n70636 , n70382 );
not ( n70637 , n70636 );
or ( n70638 , n70635 , n70637 );
not ( n70639 , n69557 );
nand ( n70640 , n70382 , n70639 );
nand ( n70641 , n70638 , n70640 );
not ( n70642 , n70641 );
and ( n70643 , n70392 , n69474 );
not ( n70644 , n70643 );
nand ( n70645 , n70642 , n70644 );
nand ( n70646 , n70634 , n70645 );
not ( n70647 , n70277 );
not ( n70648 , n69523 );
not ( n70649 , n70648 );
or ( n70650 , n70647 , n70649 );
not ( n70651 , n70277 );
nand ( n70652 , n69523 , n70651 );
nand ( n70653 , n70650 , n70652 );
not ( n70654 , n70653 );
and ( n70655 , n70257 , n69535 );
not ( n70656 , n70655 );
nand ( n70657 , n70654 , n70656 );
xor ( n70658 , n69535 , n70257 );
not ( n70659 , n70658 );
and ( n70660 , n69547 , n70267 );
not ( n70661 , n70660 );
nand ( n70662 , n70659 , n70661 );
nand ( n70663 , n70657 , n70662 );
nor ( n70664 , n70646 , n70663 );
not ( n70665 , n69580 );
not ( n70666 , n70300 );
not ( n70667 , n70666 );
or ( n70668 , n70665 , n70667 );
not ( n70669 , n69580 );
nand ( n70670 , n70669 , n70300 );
nand ( n70671 , n70668 , n70670 );
nand ( n70672 , n70312 , n69591 );
not ( n70673 , n70672 );
nor ( n70674 , n70671 , n70673 );
not ( n70675 , n70312 );
not ( n70676 , n69591 );
not ( n70677 , n70676 );
or ( n70678 , n70675 , n70677 );
not ( n70679 , n70312 );
nand ( n70680 , n70679 , n69591 );
nand ( n70681 , n70678 , n70680 );
and ( n70682 , n70277 , n69523 );
nor ( n70683 , n70681 , n70682 );
nor ( n70684 , n70674 , n70683 );
not ( n70685 , n70242 );
not ( n70686 , n70685 );
not ( n70687 , n69617 );
or ( n70688 , n70686 , n70687 );
not ( n70689 , n69617 );
nand ( n70690 , n70689 , n70242 );
nand ( n70691 , n70688 , n70690 );
nand ( n70692 , n69603 , n70331 );
not ( n70693 , n70692 );
nor ( n70694 , n70691 , n70693 );
not ( n70695 , n69603 );
not ( n70696 , n70695 );
not ( n70697 , n70331 );
or ( n70698 , n70696 , n70697 );
not ( n70699 , n70331 );
nand ( n70700 , n70699 , n69603 );
nand ( n70701 , n70698 , n70700 );
and ( n70702 , n69580 , n70300 );
nor ( n70703 , n70701 , n70702 );
nor ( n70704 , n70694 , n70703 );
nand ( n70705 , n70623 , n70664 , n70684 , n70704 );
not ( n70706 , n70705 );
not ( n70707 , n70706 );
not ( n70708 , n70463 );
not ( n70709 , n70077 );
not ( n70710 , n70709 );
or ( n70711 , n70708 , n70710 );
not ( n70712 , n70463 );
nand ( n70713 , n70712 , n70077 );
nand ( n70714 , n70711 , n70713 );
not ( n70715 , n70714 );
not ( n70716 , n70057 );
not ( n70717 , n70507 );
nor ( n70718 , n70716 , n70717 );
not ( n70719 , n70718 );
nand ( n70720 , n70715 , n70719 );
not ( n70721 , n70507 );
not ( n70722 , n70057 );
not ( n70723 , n70722 );
or ( n70724 , n70721 , n70723 );
nand ( n70725 , n70057 , n70717 );
nand ( n70726 , n70724 , n70725 );
not ( n70727 , n69971 );
not ( n70728 , n70526 );
nor ( n70729 , n70727 , n70728 );
nand ( n70730 , n70726 , n70729 );
not ( n70731 , n70730 );
nand ( n70732 , n70720 , n70731 );
xor ( n70733 , n69475 , n69455 );
xor ( n70734 , n70733 , n70424 );
and ( n70735 , n70077 , n70463 );
nand ( n70736 , n70734 , n70735 );
nand ( n70737 , n70714 , n70718 );
nand ( n70738 , n70732 , n70736 , n70737 );
not ( n70739 , n69506 );
not ( n70740 , n70436 );
not ( n70741 , n70740 );
or ( n70742 , n70739 , n70741 );
not ( n70743 , n69506 );
nand ( n70744 , n70436 , n70743 );
nand ( n70745 , n70742 , n70744 );
not ( n70746 , n70745 );
and ( n70747 , n70409 , n69491 );
not ( n70748 , n70747 );
nand ( n70749 , n70746 , n70748 );
xor ( n70750 , n69475 , n69455 );
and ( n70751 , n70750 , n70424 );
and ( n70752 , n69475 , n69455 );
or ( n70753 , n70751 , n70752 );
not ( n70754 , n70753 );
not ( n70755 , n69491 );
not ( n70756 , n70409 );
not ( n70757 , n70756 );
or ( n70758 , n70755 , n70757 );
not ( n70759 , n69491 );
nand ( n70760 , n70759 , n70409 );
nand ( n70761 , n70758 , n70760 );
not ( n70762 , n70761 );
nand ( n70763 , n70754 , n70762 );
and ( n70764 , n70749 , n70763 );
or ( n70765 , n70734 , n70735 );
nand ( n70766 , n70738 , n70764 , n70765 );
and ( n70767 , n70753 , n70761 );
not ( n70768 , n70767 );
not ( n70769 , n70749 );
or ( n70770 , n70768 , n70769 );
not ( n70771 , n70748 );
nand ( n70772 , n70771 , n70745 );
nand ( n70773 , n70770 , n70772 );
not ( n70774 , n70617 );
nor ( n70775 , n70773 , n70774 );
nand ( n70776 , n70766 , n70775 );
not ( n70777 , n70776 );
or ( n70778 , n70707 , n70777 );
not ( n70779 , n70701 );
not ( n70780 , n70702 );
nor ( n70781 , n70779 , n70780 );
not ( n70782 , n70781 );
not ( n70783 , n70694 );
not ( n70784 , n70783 );
or ( n70785 , n70782 , n70784 );
nand ( n70786 , n70691 , n70693 );
nand ( n70787 , n70785 , n70786 );
nand ( n70788 , n70681 , n70682 );
or ( n70789 , n70674 , n70788 );
nand ( n70790 , n70671 , n70673 );
nand ( n70791 , n70789 , n70790 );
nor ( n70792 , n70787 , n70791 );
not ( n70793 , n70792 );
nand ( n70794 , n70653 , n70655 );
nand ( n70795 , n70663 , n70794 );
nand ( n70796 , n70658 , n70660 );
nand ( n70797 , n70630 , n70632 );
nand ( n70798 , n70796 , n70794 , n70797 );
not ( n70799 , n70798 );
and ( n70800 , n70641 , n70643 );
nand ( n70801 , n70634 , n70800 );
nand ( n70802 , n70799 , n70801 );
nand ( n70803 , n70795 , n70802 , n70684 );
not ( n70804 , n70803 );
or ( n70805 , n70793 , n70804 );
or ( n70806 , n70787 , n70704 );
nand ( n70807 , n70805 , n70806 );
nand ( n70808 , n70778 , n70807 );
not ( n70809 , n70808 );
not ( n70810 , n70809 );
or ( n70811 , n70592 , n70810 );
nand ( n70812 , n70706 , n70776 );
nand ( n70813 , n70807 , n70812 );
not ( n70814 , n70813 );
or ( n70815 , n70814 , n70591 );
nand ( n70816 , n70811 , n70815 );
not ( n70817 , n70816 );
or ( n70818 , n70578 , n70817 );
not ( n70819 , n70229 );
nor ( n70820 , n70392 , n70436 );
not ( n70821 , n70409 );
not ( n70822 , n70821 );
nor ( n70823 , n70481 , n70822 );
nor ( n70824 , n70331 , n70242 );
nor ( n70825 , n70424 , n70463 );
nand ( n70826 , n70820 , n70823 , n70824 , n70825 );
not ( n70827 , n70826 );
nor ( n70828 , n70267 , n70382 );
not ( n70829 , n70257 );
not ( n70830 , n70277 );
and ( n70831 , n70828 , n70829 , n70830 );
nor ( n70832 , n70300 , n70312 );
not ( n70833 , n70507 );
not ( n70834 , n70833 );
nor ( n70835 , n70834 , n70526 );
nand ( n70836 , n70827 , n70831 , n70832 , n70835 );
not ( n70837 , n70836 );
not ( n70838 , n70837 );
or ( n70839 , n70819 , n70838 );
or ( n70840 , n70837 , n70229 );
nand ( n70841 , n70839 , n70840 );
nor ( n70842 , n70192 , n70198 );
nand ( n70843 , n70842 , n70211 );
nor ( n70844 , n70187 , n70843 );
nand ( n70845 , n70841 , n70844 );
not ( n70846 , n70187 );
not ( n70847 , n70198 );
not ( n70848 , n70206 );
nor ( n70849 , n70848 , n70192 );
nand ( n70850 , n70847 , n70849 );
not ( n70851 , n70850 );
nand ( n70852 , n70846 , n70851 );
not ( n70853 , n70852 );
nand ( n70854 , n70853 , n70229 );
not ( n70855 , n70849 );
nor ( n70856 , n70206 , n70210 );
not ( n70857 , n70856 );
nand ( n70858 , n70565 , n70855 , n70857 );
not ( n70859 , n70858 );
not ( n70860 , n70168 );
or ( n70861 , n70859 , n70860 );
or ( n70862 , n70199 , n70211 );
not ( n70863 , n70143 );
not ( n70864 , n70863 );
nand ( n70865 , n70140 , n70864 );
not ( n70866 , n70865 );
not ( n70867 , n70151 );
nand ( n70868 , n70862 , n70866 , n70867 );
not ( n70869 , n70210 );
nor ( n70870 , n70206 , n70869 );
and ( n70871 , n70842 , n70870 );
nor ( n70872 , n70871 , n70184 );
nor ( n70873 , n70868 , n70872 );
nand ( n70874 , n70861 , n70873 );
and ( n70875 , n70874 , n2697 );
not ( n70876 , n70564 );
nand ( n70877 , n70870 , n70143 );
not ( n70878 , n70877 );
nand ( n70879 , n70140 , n70876 , n70878 , n70867 );
not ( n70880 , n70879 );
not ( n70881 , n3356 );
nand ( n70882 , n3304 , n3344 );
nor ( n70883 , n70881 , n70882 );
nand ( n70884 , n70883 , n3288 );
not ( n70885 , n3324 );
nor ( n70886 , n70884 , n70885 );
nand ( n70887 , n70886 , n69553 );
not ( n70888 , n69541 );
nor ( n70889 , n70887 , n70888 );
nand ( n70890 , n70889 , n69524 );
not ( n70891 , n69516 );
nor ( n70892 , n70890 , n70891 );
and ( n70893 , n70892 , n3442 );
nand ( n70894 , n70893 , n69571 );
not ( n70895 , n3454 );
nor ( n70896 , n70894 , n70895 );
nand ( n70897 , n70896 , n69607 );
not ( n70898 , n69643 );
and ( n70899 , n70897 , n70898 );
not ( n70900 , n70897 );
and ( n70901 , n70900 , n69643 );
nor ( n70902 , n70899 , n70901 );
and ( n70903 , n70880 , n70902 );
nor ( n70904 , n70875 , n70903 );
and ( n70905 , n70845 , n70854 , n70904 );
nand ( n70906 , n70818 , n70905 );
nor ( n70907 , n70573 , n70906 );
nand ( n70908 , n70215 , n70907 );
buf ( n4766 , n70908 );
buf ( n70910 , 1'b0 );
not ( n70911 , n68842 );
buf ( n70912 , n70911 );
buf ( n4770 , n68638 );
not ( n70914 , n69362 );
not ( n70915 , n70017 );
nand ( n70916 , n69973 , n70096 );
not ( n70917 , n70916 );
nand ( n70918 , n70917 , n70011 );
not ( n70919 , n70918 );
or ( n70920 , n70915 , n70919 );
or ( n70921 , n70918 , n70017 );
nand ( n70922 , n70920 , n70921 );
not ( n70923 , n70922 );
or ( n70924 , n70914 , n70923 );
nand ( n70925 , n70086 , n69363 );
nand ( n70926 , n70924 , n70925 );
not ( n70927 , n70199 );
and ( n70928 , n70926 , n70927 );
not ( n70929 , n70210 );
not ( n70930 , n70192 );
or ( n70931 , n70929 , n70930 );
or ( n70932 , n70876 , n70855 );
nand ( n70933 , n70931 , n70932 );
not ( n70934 , n70933 );
not ( n70935 , n70934 );
not ( n70936 , n70935 );
nand ( n70937 , n70401 , n70553 );
not ( n70938 , n70937 );
not ( n70939 , n70396 );
not ( n70940 , n70446 );
nor ( n70941 , n70500 , n70940 );
not ( n70942 , n70941 );
not ( n70943 , n70467 );
not ( n70944 , n70530 );
not ( n70945 , n70944 );
or ( n70946 , n70943 , n70945 );
not ( n70947 , n70532 );
and ( n70948 , n70467 , n70947 );
not ( n70949 , n70531 );
nor ( n70950 , n70948 , n70949 );
nand ( n70951 , n70946 , n70950 );
not ( n70952 , n70951 );
or ( n70953 , n70942 , n70952 );
nand ( n70954 , n70544 , n70546 );
not ( n70955 , n70954 );
not ( n70956 , n70500 );
not ( n70957 , n70956 );
or ( n70958 , n70955 , n70957 );
nand ( n70959 , n70958 , n70495 );
not ( n70960 , n70959 );
nand ( n70961 , n70953 , n70960 );
not ( n70962 , n70961 );
or ( n70963 , n70939 , n70962 );
not ( n70964 , n70549 );
nand ( n70965 , n70963 , n70964 );
not ( n70966 , n70965 );
or ( n70967 , n70938 , n70966 );
or ( n70968 , n70965 , n70937 );
nand ( n70969 , n70967 , n70968 );
not ( n70970 , n70969 );
or ( n70971 , n70936 , n70970 );
nand ( n70972 , n70634 , n70797 );
not ( n70973 , n70972 );
not ( n70974 , n70645 );
not ( n70975 , n70764 );
nor ( n70976 , n70975 , n70622 );
not ( n70977 , n70976 );
not ( n70978 , n70732 );
nand ( n70979 , n70978 , n70765 );
not ( n70980 , n70737 );
nand ( n70981 , n70765 , n70980 );
nand ( n70982 , n70979 , n70981 , n70736 );
not ( n70983 , n70982 );
or ( n70984 , n70977 , n70983 );
not ( n70985 , n70622 );
and ( n70986 , n70773 , n70985 );
nor ( n70987 , n70986 , n70774 );
nand ( n70988 , n70984 , n70987 );
not ( n70989 , n70988 );
or ( n70990 , n70974 , n70989 );
not ( n70991 , n70800 );
nand ( n70992 , n70990 , n70991 );
not ( n70993 , n70992 );
or ( n70994 , n70973 , n70993 );
or ( n70995 , n70992 , n70972 );
nand ( n70996 , n70994 , n70995 );
and ( n70997 , n70996 , n70575 );
not ( n70998 , n70856 );
nor ( n70999 , n70998 , n70564 );
not ( n71000 , n70999 );
not ( n71001 , n70267 );
not ( n71002 , n71001 );
not ( n71003 , n70382 );
and ( n71004 , n70835 , n70825 );
and ( n71005 , n70823 , n70820 );
nand ( n71006 , n71004 , n71005 );
not ( n71007 , n71006 );
nand ( n71008 , n71003 , n71007 );
not ( n71009 , n71008 );
or ( n71010 , n71002 , n71009 );
or ( n71011 , n71008 , n71001 );
nand ( n71012 , n71010 , n71011 );
not ( n71013 , n71012 );
or ( n71014 , n71000 , n71013 );
nand ( n71015 , n70851 , n70267 );
nand ( n71016 , n71014 , n71015 );
nor ( n71017 , n70997 , n71016 );
nand ( n71018 , n70971 , n71017 );
nor ( n71019 , n70928 , n71018 );
nand ( n71020 , n70152 , n70168 , n70185 , n70858 );
or ( n71021 , n71019 , n71020 );
nand ( n71022 , n71020 , n69539 );
nand ( n71023 , n71021 , n71022 );
buf ( n4881 , n71023 );
buf ( n4882 , 1'b0 );
not ( n71026 , n68842 );
buf ( n4884 , n71026 );
buf ( n4885 , n68638 );
not ( n71029 , n71020 );
not ( n71030 , n69804 );
or ( n71031 , n71029 , n71030 );
not ( n71032 , n69362 );
nor ( n71033 , n69827 , n69830 );
not ( n71034 , n71033 );
not ( n71035 , n71034 );
nand ( n71036 , n71035 , n69631 );
not ( n71037 , n69875 );
and ( n71038 , n71036 , n71037 );
not ( n71039 , n71036 );
and ( n71040 , n71039 , n69875 );
nor ( n71041 , n71038 , n71040 );
not ( n71042 , n71041 );
nand ( n71043 , n69987 , n69664 );
nor ( n71044 , n70103 , n71043 );
nand ( n71045 , n69975 , n71044 );
nand ( n71046 , n69631 , n69831 );
not ( n71047 , n69826 );
and ( n71048 , n71046 , n71047 );
not ( n71049 , n71046 );
and ( n71050 , n71049 , n69826 );
nor ( n71051 , n71048 , n71050 );
not ( n71052 , n71051 );
nor ( n71053 , n71045 , n71052 );
not ( n71054 , n69808 );
not ( n71055 , n69831 );
nor ( n71056 , n71055 , n71047 );
nand ( n71057 , n69631 , n71056 );
not ( n71058 , n71057 );
or ( n71059 , n71054 , n71058 );
nand ( n71060 , n69631 , n71056 );
or ( n71061 , n71060 , n69808 );
nand ( n71062 , n71059 , n71061 );
nand ( n71063 , n71053 , n71062 );
not ( n71064 , n71063 );
or ( n71065 , n71042 , n71064 );
or ( n71066 , n71063 , n71041 );
nand ( n71067 , n71065 , n71066 );
not ( n71068 , n71067 );
or ( n71069 , n71032 , n71068 );
nand ( n71070 , n71051 , n69363 );
nand ( n71071 , n71069 , n71070 );
and ( n71072 , n71071 , n70927 );
not ( n71073 , n69180 );
not ( n71074 , n70226 );
not ( n71075 , n71074 );
or ( n71076 , n71073 , n71075 );
nand ( n71077 , n70226 , n68654 );
nand ( n71078 , n71076 , n71077 );
not ( n71079 , n71078 );
not ( n71080 , n71079 );
not ( n71081 , n69659 );
not ( n71082 , n71081 );
or ( n71083 , n71080 , n71082 );
nand ( n71084 , n69659 , n71078 );
nand ( n71085 , n71083 , n71084 );
nand ( n71086 , n70233 , n69645 );
not ( n71087 , n71086 );
nor ( n71088 , n71085 , n71087 );
nor ( n71089 , n71088 , n70245 );
not ( n71090 , n71089 );
not ( n71091 , n69826 );
not ( n71092 , n69161 );
not ( n71093 , n71074 );
or ( n71094 , n71092 , n71093 );
nand ( n71095 , n70226 , n68653 );
nand ( n71096 , n71094 , n71095 );
not ( n71097 , n71096 );
or ( n71098 , n71091 , n71097 );
not ( n71099 , n71096 );
not ( n71100 , n69826 );
nand ( n71101 , n71099 , n71100 );
nand ( n71102 , n71098 , n71101 );
and ( n71103 , n71079 , n69659 );
nor ( n71104 , n71102 , n71103 );
nor ( n71105 , n71090 , n71104 );
not ( n71106 , n71105 );
not ( n71107 , n70557 );
or ( n71108 , n71106 , n71107 );
not ( n71109 , n71104 );
not ( n71110 , n71109 );
or ( n71111 , n70247 , n71088 );
nand ( n71112 , n71085 , n71087 );
nand ( n71113 , n71111 , n71112 );
not ( n71114 , n71113 );
or ( n71115 , n71110 , n71114 );
nand ( n71116 , n71102 , n71103 );
nand ( n71117 , n71115 , n71116 );
not ( n71118 , n71117 );
nand ( n71119 , n71108 , n71118 );
not ( n71120 , n69808 );
not ( n71121 , n70226 );
not ( n71122 , n69245 );
and ( n71123 , n71121 , n71122 );
and ( n71124 , n70226 , n2509 );
nor ( n71125 , n71123 , n71124 );
not ( n71126 , n71125 );
not ( n71127 , n71126 );
or ( n71128 , n71120 , n71127 );
not ( n71129 , n71126 );
not ( n71130 , n69808 );
nand ( n71131 , n71129 , n71130 );
nand ( n71132 , n71128 , n71131 );
not ( n71133 , n69826 );
nor ( n71134 , n71133 , n71096 );
nor ( n71135 , n71132 , n71134 );
and ( n71136 , n71132 , n71134 );
or ( n71137 , n71135 , n71136 );
xnor ( n71138 , n71119 , n71137 );
nand ( n71139 , n71138 , n70933 );
not ( n71140 , n71126 );
not ( n71141 , n71140 );
not ( n71142 , n69808 );
or ( n71143 , n71141 , n71142 );
not ( n71144 , n69808 );
nand ( n71145 , n71144 , n71126 );
nand ( n71146 , n71143 , n71145 );
nand ( n71147 , n71096 , n69826 );
not ( n71148 , n71147 );
and ( n71149 , n71146 , n71148 );
nor ( n71150 , n71146 , n71148 );
or ( n71151 , n71149 , n71150 );
not ( n71152 , n71151 );
not ( n71153 , n69659 );
not ( n71154 , n71078 );
not ( n71155 , n71154 );
or ( n71156 , n71153 , n71155 );
not ( n71157 , n69659 );
nand ( n71158 , n71157 , n71078 );
nand ( n71159 , n71156 , n71158 );
nand ( n71160 , n69645 , n70229 );
not ( n71161 , n71160 );
nor ( n71162 , n71159 , n71161 );
not ( n71163 , n71162 );
nand ( n71164 , n71163 , n70589 );
not ( n71165 , n69826 );
not ( n71166 , n71096 );
not ( n71167 , n71166 );
or ( n71168 , n71165 , n71167 );
not ( n71169 , n69826 );
nand ( n71170 , n71096 , n71169 );
nand ( n71171 , n71168 , n71170 );
and ( n71172 , n69659 , n71078 );
nor ( n71173 , n71171 , n71172 );
nor ( n71174 , n71164 , n71173 );
not ( n71175 , n71174 );
not ( n71176 , n70808 );
or ( n71177 , n71175 , n71176 );
not ( n71178 , n71173 );
not ( n71179 , n71178 );
or ( n71180 , n71162 , n70590 );
nand ( n71181 , n71159 , n71161 );
nand ( n71182 , n71180 , n71181 );
not ( n71183 , n71182 );
or ( n71184 , n71179 , n71183 );
nand ( n71185 , n71171 , n71172 );
nand ( n71186 , n71184 , n71185 );
not ( n71187 , n71186 );
nand ( n71188 , n71177 , n71187 );
not ( n71189 , n71188 );
or ( n71190 , n71152 , n71189 );
or ( n71191 , n71188 , n71151 );
nand ( n71192 , n71190 , n71191 );
and ( n71193 , n71192 , n70575 );
not ( n71194 , n70999 );
not ( n71195 , n71126 );
not ( n71196 , n70229 );
not ( n71197 , n71078 );
nand ( n71198 , n71196 , n71197 );
or ( n71199 , n71198 , n71096 );
nor ( n71200 , n70836 , n71199 );
not ( n71201 , n71200 );
or ( n71202 , n71195 , n71201 );
or ( n71203 , n71200 , n71126 );
nand ( n71204 , n71202 , n71203 );
not ( n71205 , n71204 );
or ( n71206 , n71194 , n71205 );
nand ( n71207 , n70851 , n71126 );
nand ( n71208 , n71206 , n71207 );
nor ( n71209 , n71193 , n71208 );
nand ( n71210 , n71139 , n71209 );
nor ( n71211 , n71072 , n71210 );
or ( n71212 , n71211 , n71020 );
nand ( n71213 , n71031 , n71212 );
buf ( n71214 , n71213 );
buf ( n5072 , 1'b0 );
not ( n71216 , n68842 );
buf ( n71217 , n71216 );
buf ( n5075 , n68638 );
not ( n71219 , n69362 );
not ( n71220 , n71062 );
not ( n71221 , n71220 );
not ( n71222 , n71053 );
or ( n71223 , n71221 , n71222 );
or ( n71224 , n71053 , n71220 );
nand ( n71225 , n71223 , n71224 );
not ( n71226 , n71225 );
or ( n71227 , n71219 , n71226 );
nand ( n71228 , n69664 , n69363 );
nand ( n71229 , n71227 , n71228 );
and ( n71230 , n71229 , n70927 );
not ( n71231 , n71089 );
not ( n71232 , n70557 );
or ( n71233 , n71231 , n71232 );
not ( n71234 , n71113 );
nand ( n71235 , n71233 , n71234 );
nand ( n71236 , n71109 , n71116 );
xnor ( n71237 , n71235 , n71236 );
not ( n71238 , n71237 );
not ( n71239 , n70933 );
or ( n71240 , n71238 , n71239 );
nand ( n71241 , n71178 , n71185 );
not ( n71242 , n71241 );
not ( n71243 , n71164 );
not ( n71244 , n71243 );
not ( n71245 , n70808 );
or ( n71246 , n71244 , n71245 );
not ( n71247 , n71182 );
nand ( n71248 , n71246 , n71247 );
not ( n71249 , n71248 );
or ( n71250 , n71242 , n71249 );
or ( n71251 , n71248 , n71241 );
nand ( n71252 , n71250 , n71251 );
and ( n71253 , n71252 , n70575 );
not ( n71254 , n70999 );
not ( n71255 , n71096 );
nor ( n71256 , n70836 , n71198 );
not ( n71257 , n71256 );
or ( n71258 , n71255 , n71257 );
or ( n71259 , n71256 , n71096 );
nand ( n71260 , n71258 , n71259 );
not ( n71261 , n71260 );
or ( n71262 , n71254 , n71261 );
nand ( n71263 , n70851 , n71096 );
nand ( n71264 , n71262 , n71263 );
nor ( n71265 , n71253 , n71264 );
nand ( n71266 , n71240 , n71265 );
nor ( n71267 , n71230 , n71266 );
or ( n71268 , n71267 , n71020 );
nand ( n71269 , n71020 , n69814 );
nand ( n71270 , n71268 , n71269 );
buf ( n5128 , n71270 );
buf ( n5129 , 1'b0 );
not ( n71273 , n68842 );
buf ( n71274 , n71273 );
buf ( n71275 , n68638 );
not ( n71276 , n69362 );
and ( n71277 , n71276 , n69981 );
not ( n71278 , n71276 );
not ( n71279 , n71051 );
not ( n71280 , n71045 );
or ( n71281 , n71279 , n71280 );
or ( n71282 , n71045 , n71051 );
nand ( n71283 , n71281 , n71282 );
and ( n71284 , n71278 , n71283 );
nor ( n71285 , n71277 , n71284 );
not ( n71286 , n71285 );
and ( n71287 , n71286 , n70927 );
not ( n71288 , n70933 );
not ( n71289 , n70246 );
not ( n71290 , n70557 );
or ( n71291 , n71289 , n71290 );
nand ( n71292 , n71291 , n70247 );
not ( n71293 , n71088 );
nand ( n71294 , n71293 , n71112 );
xnor ( n71295 , n71292 , n71294 );
not ( n71296 , n71295 );
or ( n71297 , n71288 , n71296 );
not ( n71298 , n71162 );
nand ( n71299 , n71298 , n71181 );
not ( n71300 , n71299 );
not ( n71301 , n70589 );
not ( n71302 , n70808 );
or ( n71303 , n71301 , n71302 );
nand ( n71304 , n71303 , n70590 );
not ( n71305 , n71304 );
or ( n71306 , n71300 , n71305 );
or ( n71307 , n71304 , n71299 );
nand ( n71308 , n71306 , n71307 );
and ( n71309 , n71308 , n70575 );
not ( n71310 , n70999 );
not ( n71311 , n71078 );
nor ( n71312 , n70836 , n70229 );
not ( n71313 , n71312 );
or ( n71314 , n71311 , n71313 );
or ( n71315 , n71312 , n71078 );
nand ( n71316 , n71314 , n71315 );
not ( n71317 , n71316 );
or ( n71318 , n71310 , n71317 );
nand ( n71319 , n70851 , n71078 );
nand ( n71320 , n71318 , n71319 );
nor ( n71321 , n71309 , n71320 );
nand ( n71322 , n71297 , n71321 );
nor ( n71323 , n71287 , n71322 );
or ( n71324 , n71323 , n71020 );
nand ( n71325 , n71020 , n3510 );
nand ( n71326 , n71324 , n71325 );
buf ( n71327 , n71326 );
buf ( n71328 , 1'b0 );
not ( n71329 , n68842 );
buf ( n71330 , n71329 );
buf ( n71331 , n68638 );
not ( n71332 , n70113 );
and ( n71333 , n71332 , n70200 );
not ( n71334 , n70935 );
not ( n71335 , n70561 );
or ( n71336 , n71334 , n71335 );
and ( n71337 , n70816 , n70575 );
not ( n71338 , n70999 );
not ( n71339 , n70841 );
or ( n71340 , n71338 , n71339 );
nand ( n71341 , n70229 , n70851 );
nand ( n71342 , n71340 , n71341 );
nor ( n71343 , n71337 , n71342 );
nand ( n71344 , n71336 , n71343 );
nor ( n71345 , n71333 , n71344 );
or ( n71346 , n71345 , n71020 );
not ( n71347 , n71020 );
not ( n71348 , n71347 );
nand ( n71349 , n71348 , n3498 );
nand ( n71350 , n71346 , n71349 );
buf ( n71351 , n71350 );
buf ( n71352 , 1'b0 );
not ( n71353 , n68842 );
buf ( n71354 , n71353 );
buf ( n71355 , n68638 );
not ( n71356 , n69362 );
not ( n71357 , n69982 );
not ( n71358 , n71357 );
nor ( n71359 , n70105 , n69986 );
nand ( n71360 , n69973 , n71359 );
not ( n71361 , n71360 );
or ( n71362 , n71358 , n71361 );
or ( n71363 , n71360 , n71357 );
nand ( n71364 , n71362 , n71363 );
not ( n71365 , n71364 );
or ( n71366 , n71356 , n71365 );
nand ( n71367 , n69985 , n71276 );
nand ( n71368 , n71366 , n71367 );
and ( n71369 , n71368 , n70200 );
not ( n71370 , n70935 );
not ( n71371 , n70349 );
nand ( n71372 , n71371 , n70369 );
not ( n71373 , n71372 );
not ( n71374 , n70340 );
nand ( n71375 , n70325 , n71374 );
not ( n71376 , n70537 );
nor ( n71377 , n71375 , n71376 );
not ( n71378 , n71377 );
not ( n71379 , n70961 );
or ( n71380 , n71378 , n71379 );
nor ( n71381 , n70291 , n70555 );
not ( n71382 , n71381 );
not ( n71383 , n71375 );
and ( n71384 , n71382 , n71383 );
not ( n71385 , n71374 );
not ( n71386 , n70362 );
or ( n71387 , n71385 , n71386 );
nand ( n71388 , n71387 , n70366 );
nor ( n71389 , n71384 , n71388 );
nand ( n71390 , n71380 , n71389 );
not ( n71391 , n71390 );
or ( n71392 , n71373 , n71391 );
or ( n71393 , n71390 , n71372 );
nand ( n71394 , n71392 , n71393 );
not ( n71395 , n71394 );
or ( n71396 , n71370 , n71395 );
nand ( n71397 , n70783 , n70786 );
not ( n71398 , n71397 );
not ( n71399 , n70703 );
nand ( n71400 , n70684 , n71399 );
not ( n71401 , n70664 );
nor ( n71402 , n71400 , n71401 );
not ( n71403 , n71402 );
not ( n71404 , n70988 );
or ( n71405 , n71403 , n71404 );
nand ( n71406 , n70802 , n70795 );
not ( n71407 , n71406 );
not ( n71408 , n71400 );
and ( n71409 , n71407 , n71408 );
not ( n71410 , n71399 );
not ( n71411 , n70791 );
or ( n71412 , n71410 , n71411 );
not ( n71413 , n70781 );
nand ( n71414 , n71412 , n71413 );
nor ( n71415 , n71409 , n71414 );
nand ( n71416 , n71405 , n71415 );
not ( n71417 , n71416 );
or ( n71418 , n71398 , n71417 );
or ( n71419 , n71416 , n71397 );
nand ( n71420 , n71418 , n71419 );
and ( n71421 , n71420 , n70575 );
not ( n71422 , n70999 );
not ( n71423 , n70242 );
not ( n71424 , n71423 );
not ( n71425 , n70331 );
nand ( n71426 , n70831 , n70832 , n71425 );
not ( n71427 , n71426 );
nand ( n71428 , n71427 , n71007 );
not ( n71429 , n71428 );
or ( n71430 , n71424 , n71429 );
or ( n71431 , n71428 , n71423 );
nand ( n71432 , n71430 , n71431 );
not ( n71433 , n71432 );
or ( n71434 , n71422 , n71433 );
nand ( n71435 , n70242 , n70851 );
nand ( n71436 , n71434 , n71435 );
nor ( n71437 , n71421 , n71436 );
nand ( n71438 , n71396 , n71437 );
nor ( n71439 , n71369 , n71438 );
or ( n71440 , n71439 , n71020 );
nand ( n71441 , n71020 , n69611 );
nand ( n71442 , n71440 , n71441 );
buf ( n5300 , n71442 );
buf ( n5301 , 1'b0 );
not ( n71445 , n68842 );
buf ( n71446 , n71445 );
buf ( n71447 , n68638 );
not ( n71448 , n69362 );
not ( n71449 , n69622 );
not ( n71450 , n71449 );
nand ( n71451 , n69973 , n70104 );
not ( n71452 , n69985 );
nor ( n71453 , n71451 , n71452 );
not ( n71454 , n71453 );
or ( n71455 , n71450 , n71454 );
or ( n71456 , n71453 , n71449 );
nand ( n71457 , n71455 , n71456 );
not ( n71458 , n71457 );
or ( n71459 , n71448 , n71458 );
nand ( n71460 , n70102 , n69363 );
nand ( n71461 , n71459 , n71460 );
and ( n71462 , n71461 , n70927 );
not ( n71463 , n70933 );
nand ( n71464 , n71374 , n70366 );
not ( n71465 , n71464 );
not ( n71466 , n70325 );
nor ( n71467 , n71376 , n71466 );
not ( n71468 , n71467 );
not ( n71469 , n70961 );
or ( n71470 , n71468 , n71469 );
or ( n71471 , n71381 , n71466 );
not ( n71472 , n70362 );
nand ( n71473 , n71471 , n71472 );
not ( n71474 , n71473 );
nand ( n71475 , n71470 , n71474 );
not ( n71476 , n71475 );
or ( n71477 , n71465 , n71476 );
or ( n71478 , n71475 , n71464 );
nand ( n71479 , n71477 , n71478 );
not ( n71480 , n71479 );
or ( n71481 , n71463 , n71480 );
nand ( n71482 , n71399 , n71413 );
not ( n71483 , n71482 );
not ( n71484 , n70684 );
nor ( n71485 , n71484 , n71401 );
not ( n71486 , n71485 );
not ( n71487 , n70988 );
or ( n71488 , n71486 , n71487 );
not ( n71489 , n70803 );
nor ( n71490 , n71489 , n70791 );
nand ( n71491 , n71488 , n71490 );
not ( n71492 , n71491 );
or ( n71493 , n71483 , n71492 );
or ( n71494 , n71491 , n71482 );
nand ( n71495 , n71493 , n71494 );
and ( n71496 , n71495 , n70575 );
not ( n71497 , n70999 );
not ( n71498 , n71425 );
nand ( n71499 , n70831 , n70832 );
not ( n71500 , n71499 );
nand ( n71501 , n71500 , n71007 );
not ( n71502 , n71501 );
or ( n71503 , n71498 , n71502 );
or ( n71504 , n71501 , n71425 );
nand ( n71505 , n71503 , n71504 );
not ( n71506 , n71505 );
or ( n71507 , n71497 , n71506 );
nand ( n71508 , n70331 , n70851 );
nand ( n71509 , n71507 , n71508 );
nor ( n71510 , n71496 , n71509 );
nand ( n71511 , n71481 , n71510 );
nor ( n71512 , n71462 , n71511 );
or ( n71513 , n71512 , n71020 );
nand ( n71514 , n71020 , n69595 );
nand ( n71515 , n71513 , n71514 );
buf ( n71516 , n71515 );
buf ( n71517 , 1'b0 );
not ( n71518 , n68842 );
buf ( n5376 , n71518 );
buf ( n71520 , n68638 );
not ( n71521 , n69362 );
not ( n71522 , n70102 );
not ( n71523 , n70019 );
not ( n71524 , n70005 );
and ( n71525 , n70096 , n71523 , n71524 );
nand ( n71526 , n69975 , n71525 );
not ( n71527 , n71526 );
or ( n71528 , n71522 , n71527 );
or ( n71529 , n71526 , n70102 );
nand ( n71530 , n71528 , n71529 );
not ( n71531 , n71530 );
or ( n71532 , n71521 , n71531 );
not ( n71533 , n70004 );
not ( n71534 , n71533 );
nand ( n71535 , n71534 , n69363 );
nand ( n71536 , n71532 , n71535 );
and ( n71537 , n71536 , n70927 );
not ( n71538 , n70935 );
not ( n71539 , n70324 );
nand ( n71540 , n71539 , n70355 );
not ( n71541 , n71540 );
not ( n71542 , n70537 );
not ( n71543 , n70961 );
or ( n71544 , n71542 , n71543 );
nand ( n71545 , n71544 , n71381 );
not ( n71546 , n71545 );
or ( n71547 , n71541 , n71546 );
or ( n71548 , n71545 , n71540 );
nand ( n71549 , n71547 , n71548 );
not ( n71550 , n71549 );
or ( n71551 , n71538 , n71550 );
not ( n71552 , n70683 );
nand ( n71553 , n71552 , n70788 );
not ( n71554 , n71553 );
not ( n71555 , n70664 );
not ( n71556 , n70988 );
or ( n71557 , n71555 , n71556 );
nand ( n71558 , n71557 , n71406 );
not ( n71559 , n71558 );
or ( n71560 , n71554 , n71559 );
or ( n71561 , n71558 , n71553 );
nand ( n71562 , n71560 , n71561 );
and ( n71563 , n71562 , n70575 );
not ( n71564 , n70999 );
not ( n71565 , n70312 );
not ( n71566 , n71565 );
nand ( n71567 , n71007 , n70831 );
not ( n71568 , n71567 );
or ( n71569 , n71566 , n71568 );
or ( n71570 , n71567 , n71565 );
nand ( n71571 , n71569 , n71570 );
not ( n71572 , n71571 );
or ( n71573 , n71564 , n71572 );
nand ( n71574 , n70312 , n70851 );
nand ( n71575 , n71573 , n71574 );
nor ( n71576 , n71563 , n71575 );
nand ( n71577 , n71551 , n71576 );
nor ( n71578 , n71537 , n71577 );
or ( n71579 , n71578 , n71020 );
nand ( n71580 , n71020 , n69583 );
nand ( n71581 , n71579 , n71580 );
buf ( n71582 , n71581 );
buf ( n5440 , 1'b0 );
not ( n71584 , n68842 );
buf ( n71585 , n71584 );
buf ( n71586 , n68638 );
not ( n71587 , n69362 );
not ( n71588 , n69994 );
not ( n71589 , n71588 );
not ( n71590 , n70095 );
and ( n71591 , n71590 , n70018 );
nand ( n71592 , n69973 , n71591 );
not ( n71593 , n70004 );
nor ( n71594 , n71592 , n71593 );
not ( n71595 , n71594 );
or ( n71596 , n71589 , n71595 );
or ( n71597 , n71594 , n71588 );
nand ( n71598 , n71596 , n71597 );
not ( n71599 , n71598 );
or ( n71600 , n71587 , n71599 );
nand ( n71601 , n70017 , n69363 );
nand ( n71602 , n71600 , n71601 );
and ( n71603 , n71602 , n70200 );
not ( n71604 , n70935 );
nand ( n71605 , n70287 , n70290 );
not ( n71606 , n71605 );
not ( n71607 , n70402 );
nor ( n71608 , n71607 , n70376 );
not ( n71609 , n71608 );
not ( n71610 , n70961 );
or ( n71611 , n71609 , n71610 );
not ( n71612 , n70536 );
not ( n71613 , n70554 );
or ( n71614 , n71612 , n71613 );
not ( n71615 , n70270 );
nand ( n71616 , n71614 , n71615 );
not ( n71617 , n71616 );
nand ( n71618 , n71611 , n71617 );
not ( n71619 , n71618 );
or ( n71620 , n71606 , n71619 );
or ( n71621 , n71618 , n71605 );
nand ( n71622 , n71620 , n71621 );
not ( n71623 , n71622 );
or ( n71624 , n71604 , n71623 );
nand ( n71625 , n70657 , n70794 );
not ( n71626 , n71625 );
not ( n71627 , n70662 );
nor ( n71628 , n71627 , n70646 );
not ( n71629 , n71628 );
not ( n71630 , n70988 );
or ( n71631 , n71629 , n71630 );
not ( n71632 , n70662 );
nand ( n71633 , n70801 , n70797 );
not ( n71634 , n71633 );
or ( n71635 , n71632 , n71634 );
nand ( n71636 , n71635 , n70796 );
not ( n71637 , n71636 );
nand ( n71638 , n71631 , n71637 );
not ( n71639 , n71638 );
or ( n71640 , n71626 , n71639 );
or ( n71641 , n71638 , n71625 );
nand ( n71642 , n71640 , n71641 );
and ( n71643 , n71642 , n70575 );
not ( n71644 , n70999 );
not ( n71645 , n70830 );
and ( n71646 , n70828 , n70829 );
nand ( n71647 , n71007 , n71646 );
not ( n71648 , n71647 );
or ( n71649 , n71645 , n71648 );
or ( n71650 , n71647 , n70830 );
nand ( n71651 , n71649 , n71650 );
not ( n71652 , n71651 );
or ( n71653 , n71644 , n71652 );
nand ( n71654 , n70277 , n70851 );
nand ( n71655 , n71653 , n71654 );
nor ( n71656 , n71643 , n71655 );
nand ( n71657 , n71624 , n71656 );
nor ( n71658 , n71603 , n71657 );
or ( n71659 , n71658 , n71020 );
nand ( n71660 , n71020 , n69513 );
nand ( n71661 , n71659 , n71660 );
buf ( n71662 , n71661 );
buf ( n71663 , 1'b0 );
not ( n71664 , n68842 );
buf ( n71665 , n71664 );
buf ( n71666 , n68638 );
not ( n71667 , n69362 );
not ( n71668 , n70004 );
not ( n71669 , n71592 );
or ( n71670 , n71668 , n71669 );
or ( n71671 , n71592 , n70004 );
nand ( n71672 , n71670 , n71671 );
not ( n71673 , n71672 );
or ( n71674 , n71667 , n71673 );
nand ( n71675 , n70011 , n69363 );
nand ( n71676 , n71674 , n71675 );
and ( n71677 , n71676 , n70200 );
not ( n71678 , n70933 );
nand ( n71679 , n70536 , n71615 );
not ( n71680 , n71679 );
not ( n71681 , n70402 );
not ( n71682 , n70961 );
or ( n71683 , n71681 , n71682 );
not ( n71684 , n70554 );
nand ( n71685 , n71683 , n71684 );
not ( n71686 , n71685 );
or ( n71687 , n71680 , n71686 );
or ( n71688 , n71685 , n71679 );
nand ( n71689 , n71687 , n71688 );
not ( n71690 , n71689 );
or ( n71691 , n71678 , n71690 );
nand ( n71692 , n70662 , n70796 );
not ( n71693 , n71692 );
not ( n71694 , n70646 );
not ( n71695 , n71694 );
not ( n71696 , n70988 );
or ( n71697 , n71695 , n71696 );
not ( n71698 , n71633 );
nand ( n71699 , n71697 , n71698 );
not ( n71700 , n71699 );
or ( n71701 , n71693 , n71700 );
or ( n71702 , n71699 , n71692 );
nand ( n71703 , n71701 , n71702 );
and ( n71704 , n71703 , n70575 );
not ( n71705 , n70999 );
not ( n71706 , n70829 );
nand ( n71707 , n71007 , n70828 );
not ( n71708 , n71707 );
or ( n71709 , n71706 , n71708 );
or ( n71710 , n71707 , n70829 );
nand ( n71711 , n71709 , n71710 );
not ( n71712 , n71711 );
or ( n71713 , n71705 , n71712 );
nand ( n71714 , n70257 , n70851 );
nand ( n71715 , n71713 , n71714 );
nor ( n71716 , n71704 , n71715 );
nand ( n71717 , n71691 , n71716 );
nor ( n71718 , n71677 , n71717 );
or ( n71719 , n71718 , n71020 );
nand ( n71720 , n71020 , n69528 );
nand ( n71721 , n71719 , n71720 );
buf ( n71722 , n71721 );
buf ( n71723 , 1'b0 );
not ( n71724 , n68842 );
buf ( n5582 , n71724 );
buf ( n5583 , n68638 );
nand ( n71727 , n70150 , n70864 );
nor ( n71728 , n70140 , n71727 );
not ( n71729 , n71728 );
and ( n71730 , n71729 , n2667 );
not ( n71731 , n71729 );
and ( n71732 , n71731 , n70011 );
or ( n71733 , n71730 , n71732 );
buf ( n71734 , n71733 );
buf ( n5592 , 1'b0 );
not ( n71736 , n68842 );
buf ( n71737 , n71736 );
buf ( n5595 , n68638 );
and ( n71739 , n71729 , n2623 );
not ( n71740 , n71729 );
and ( n71741 , n71740 , n69951 );
or ( n71742 , n71739 , n71741 );
buf ( n71743 , n71742 );
buf ( n71744 , 1'b0 );
not ( n71745 , n68842 );
buf ( n5603 , n71745 );
buf ( n71747 , n68638 );
and ( n71748 , n71729 , n68774 );
not ( n71749 , n71729 );
not ( n71750 , n69631 );
not ( n71751 , n71750 );
nand ( n71752 , n69900 , n69875 );
nor ( n71753 , n71752 , n69797 );
nand ( n71754 , n71033 , n71753 );
not ( n71755 , n71754 );
not ( n71756 , n69936 );
not ( n71757 , n69854 );
nor ( n71758 , n71756 , n71757 );
not ( n71759 , n71758 );
not ( n71760 , n69689 );
nor ( n71761 , n71759 , n71760 );
nand ( n71762 , n71751 , n71755 , n71761 );
not ( n71763 , n69710 );
and ( n71764 , n71762 , n71763 );
not ( n71765 , n71762 );
and ( n71766 , n71765 , n69710 );
nor ( n71767 , n71764 , n71766 );
and ( n71768 , n71749 , n71767 );
or ( n71769 , n71748 , n71768 );
buf ( n71770 , n71769 );
buf ( n71771 , 1'b0 );
not ( n71772 , n68842 );
buf ( n71773 , n71772 );
buf ( n71774 , n68638 );
and ( n71775 , n71729 , n2633 );
not ( n71776 , n71729 );
not ( n71777 , n71759 );
nand ( n71778 , n71777 , n71755 , n69631 );
and ( n71779 , n71778 , n71760 );
not ( n71780 , n71778 );
and ( n71781 , n71780 , n69689 );
nor ( n71782 , n71779 , n71781 );
not ( n71783 , n71782 );
not ( n71784 , n71783 );
and ( n71785 , n71776 , n71784 );
or ( n71786 , n71775 , n71785 );
buf ( n71787 , n71786 );
buf ( n5645 , 1'b0 );
not ( n71789 , n68842 );
buf ( n71790 , n71789 );
buf ( n71791 , n68638 );
and ( n71792 , n71729 , n2635 );
not ( n71793 , n71729 );
not ( n71794 , n69631 );
not ( n71795 , n71794 );
nand ( n71796 , n71795 , n71755 , n69936 );
and ( n71797 , n71796 , n71757 );
not ( n71798 , n71796 );
not ( n71799 , n71757 );
and ( n71800 , n71798 , n71799 );
nor ( n71801 , n71797 , n71800 );
not ( n71802 , n71801 );
not ( n71803 , n71802 );
and ( n71804 , n71793 , n71803 );
or ( n71805 , n71792 , n71804 );
buf ( n5663 , n71805 );
buf ( n71807 , 1'b0 );
not ( n71808 , n68842 );
buf ( n5666 , n71808 );
buf ( n71810 , n68638 );
and ( n71811 , n71729 , n2637 );
not ( n71812 , n71729 );
nand ( n71813 , n71755 , n69631 );
not ( n71814 , n69936 );
and ( n71815 , n71813 , n71814 );
not ( n71816 , n71813 );
and ( n71817 , n71816 , n69936 );
nor ( n71818 , n71815 , n71817 );
and ( n71819 , n71812 , n71818 );
or ( n71820 , n71811 , n71819 );
buf ( n71821 , n71820 );
buf ( n71822 , 1'b0 );
not ( n71823 , n68842 );
buf ( n71824 , n71823 );
buf ( n5682 , n68638 );
and ( n71826 , n71729 , n2639 );
not ( n71827 , n71729 );
not ( n71828 , n71752 );
nand ( n71829 , n71828 , n69796 );
nor ( n71830 , n71034 , n71829 );
nand ( n71831 , n69631 , n71830 );
not ( n71832 , n69773 );
and ( n71833 , n71831 , n71832 );
not ( n71834 , n71831 );
and ( n71835 , n71834 , n69773 );
nor ( n71836 , n71833 , n71835 );
not ( n71837 , n71836 );
not ( n71838 , n71837 );
and ( n71839 , n71827 , n71838 );
or ( n71840 , n71826 , n71839 );
buf ( n71841 , n71840 );
buf ( n71842 , 1'b0 );
not ( n71843 , n68842 );
buf ( n71844 , n71843 );
buf ( n5702 , n68638 );
not ( n71846 , n71729 );
not ( n71847 , n71846 );
and ( n71848 , n71847 , n68784 );
not ( n71849 , n71847 );
nor ( n71850 , n71034 , n71752 );
nand ( n71851 , n69631 , n71850 );
not ( n71852 , n69796 );
and ( n71853 , n71851 , n71852 );
not ( n71854 , n71851 );
and ( n71855 , n71854 , n69796 );
nor ( n71856 , n71853 , n71855 );
and ( n71857 , n71849 , n71856 );
or ( n71858 , n71848 , n71857 );
buf ( n5716 , n71858 );
buf ( n71860 , 1'b0 );
not ( n71861 , n68842 );
buf ( n71862 , n71861 );
buf ( n71863 , n68638 );
and ( n71864 , n71729 , n2643 );
not ( n71865 , n71729 );
not ( n71866 , n69900 );
and ( n71867 , n71033 , n69875 );
nand ( n71868 , n71867 , n69631 );
not ( n71869 , n71868 );
or ( n71870 , n71866 , n71869 );
nand ( n71871 , n69631 , n71867 );
or ( n71872 , n71871 , n69900 );
nand ( n71873 , n71870 , n71872 );
and ( n71874 , n71865 , n71873 );
or ( n71875 , n71864 , n71874 );
buf ( n5733 , n71875 );
buf ( n71877 , 1'b0 );
not ( n71878 , n68842 );
buf ( n5736 , n71878 );
buf ( n71880 , n68638 );
and ( n71881 , n71847 , n68788 );
not ( n71882 , n71847 );
and ( n71883 , n71882 , n71041 );
or ( n71884 , n71881 , n71883 );
buf ( n5742 , n71884 );
buf ( n5743 , 1'b0 );
not ( n71887 , n68842 );
buf ( n5745 , n71887 );
buf ( n5746 , n68638 );
and ( n71890 , n71847 , n68790 );
not ( n71891 , n71847 );
and ( n71892 , n71891 , n71062 );
or ( n71893 , n71890 , n71892 );
buf ( n71894 , n71893 );
buf ( n5752 , 1'b0 );
not ( n71896 , n68842 );
buf ( n71897 , n71896 );
buf ( n5755 , n68638 );
and ( n71899 , n71847 , n2649 );
not ( n71900 , n71847 );
and ( n71901 , n71900 , n71051 );
or ( n71902 , n71899 , n71901 );
buf ( n71903 , n71902 );
buf ( n71904 , 1'b0 );
not ( n71905 , n68842 );
buf ( n71906 , n71905 );
buf ( n71907 , n68638 );
and ( n71908 , n71847 , n2651 );
not ( n71909 , n71847 );
and ( n71910 , n71909 , n69664 );
or ( n71911 , n71908 , n71910 );
buf ( n71912 , n71911 );
buf ( n71913 , 1'b0 );
not ( n71914 , n68842 );
buf ( n71915 , n71914 );
buf ( n71916 , n68638 );
and ( n71917 , n71847 , n2653 );
not ( n71918 , n71847 );
and ( n71919 , n71918 , n69981 );
or ( n71920 , n71917 , n71919 );
buf ( n71921 , n71920 );
buf ( n71922 , 1'b0 );
not ( n71923 , n68842 );
buf ( n71924 , n71923 );
buf ( n71925 , n68638 );
and ( n71926 , n71729 , n68798 );
not ( n71927 , n71729 );
and ( n71928 , n71927 , n69624 );
or ( n71929 , n71926 , n71928 );
buf ( n71930 , n71929 );
buf ( n71931 , 1'b0 );
not ( n71932 , n68842 );
buf ( n71933 , n71932 );
buf ( n71934 , n68638 );
and ( n71935 , n71729 , n68800 );
not ( n71936 , n71729 );
and ( n71937 , n71936 , n69985 );
or ( n71938 , n71935 , n71937 );
buf ( n71939 , n71938 );
buf ( n71940 , 1'b0 );
not ( n71941 , n68842 );
buf ( n71942 , n71941 );
buf ( n71943 , n68638 );
and ( n71944 , n71729 , n2659 );
not ( n71945 , n71729 );
and ( n71946 , n71945 , n70102 );
or ( n71947 , n71944 , n71946 );
buf ( n71948 , n71947 );
buf ( n71949 , 1'b0 );
not ( n71950 , n68842 );
buf ( n71951 , n71950 );
buf ( n71952 , n68638 );
and ( n71953 , n71729 , n68804 );
not ( n71954 , n71729 );
and ( n71955 , n71954 , n69994 );
or ( n71956 , n71953 , n71955 );
buf ( n71957 , n71956 );
buf ( n71958 , 1'b0 );
not ( n71959 , n68842 );
buf ( n71960 , n71959 );
buf ( n71961 , n68638 );
and ( n71962 , n71729 , n2663 );
not ( n71963 , n71729 );
and ( n71964 , n71963 , n71534 );
or ( n71965 , n71962 , n71964 );
buf ( n71966 , n71965 );
buf ( n71967 , 1'b0 );
not ( n71968 , n68842 );
buf ( n71969 , n71968 );
buf ( n71970 , n68638 );
and ( n71971 , n71729 , n2665 );
not ( n71972 , n71729 );
and ( n71973 , n71972 , n70017 );
or ( n71974 , n71971 , n71973 );
buf ( n71975 , n71974 );
buf ( n71976 , 1'b0 );
not ( n71977 , n68842 );
buf ( n71978 , n71977 );
buf ( n71979 , n68638 );
buf ( n71980 , n70863 );
buf ( n71981 , 1'b0 );
not ( n71982 , n68842 );
buf ( n71983 , n71982 );
buf ( n71984 , n68638 );
not ( n71985 , n70926 );
nand ( n71986 , n70168 , n70184 , n70867 );
and ( n71987 , n70211 , n70143 );
nand ( n71988 , n70140 , n70200 , n71987 );
nor ( n71989 , n71986 , n71988 );
not ( n71990 , n71989 );
or ( n71991 , n71985 , n71990 );
not ( n71992 , n70866 );
nor ( n71993 , n71992 , n71986 );
nand ( n71994 , n71993 , n70575 );
nand ( n71995 , n71993 , n70570 );
not ( n71996 , n70143 );
nor ( n71997 , n71989 , n71996 );
nand ( n71998 , n71994 , n71995 , n71997 );
not ( n71999 , n71998 );
not ( n72000 , n70851 );
not ( n72001 , n71993 );
or ( n72002 , n72000 , n72001 );
nand ( n72003 , n72002 , n70879 );
nand ( n72004 , n70140 , n70876 , n71987 );
nor ( n72005 , n71986 , n72004 );
nor ( n72006 , n72003 , n72005 );
nand ( n72007 , n71999 , n72006 );
not ( n72008 , n72007 );
and ( n72009 , n70887 , n69541 );
not ( n72010 , n70887 );
and ( n72011 , n72010 , n70888 );
nor ( n72012 , n72009 , n72011 );
not ( n72013 , n72012 );
and ( n72014 , n72008 , n72013 );
not ( n72015 , n71995 );
and ( n72016 , n70969 , n72015 );
nor ( n72017 , n72014 , n72016 );
not ( n72018 , n71994 );
and ( n72019 , n70996 , n72018 );
not ( n72020 , n72005 );
not ( n72021 , n72020 );
nand ( n72022 , n71012 , n72021 );
nand ( n72023 , n72003 , n70267 );
nand ( n72024 , n69541 , n70863 );
nand ( n72025 , n72022 , n72023 , n72024 );
nor ( n72026 , n72019 , n72025 );
and ( n72027 , n72017 , n72026 );
nand ( n72028 , n71991 , n72027 );
buf ( n5886 , n72028 );
buf ( n72030 , 1'b0 );
not ( n72031 , n68842 );
buf ( n72032 , n72031 );
buf ( n5890 , n68638 );
not ( n72034 , n69362 );
not ( n72035 , n70011 );
nand ( n72036 , n69975 , n70096 );
not ( n72037 , n72036 );
or ( n72038 , n72035 , n72037 );
or ( n72039 , n72036 , n70011 );
nand ( n72040 , n72038 , n72039 );
not ( n72041 , n72040 );
or ( n72042 , n72034 , n72041 );
nand ( n72043 , n70094 , n71276 );
nand ( n72044 , n72042 , n72043 );
not ( n72045 , n72044 );
or ( n72046 , n72045 , n71990 );
nand ( n72047 , n70645 , n70991 );
not ( n72048 , n72047 );
not ( n72049 , n70988 );
or ( n72050 , n72048 , n72049 );
or ( n72051 , n70988 , n72047 );
nand ( n72052 , n72050 , n72051 );
nand ( n72053 , n72052 , n72018 );
nand ( n72054 , n70396 , n70964 );
not ( n72055 , n72054 );
not ( n72056 , n70961 );
or ( n72057 , n72055 , n72056 );
or ( n72058 , n70961 , n72054 );
nand ( n72059 , n72057 , n72058 );
nand ( n72060 , n72059 , n72015 );
not ( n72061 , n72007 );
and ( n72062 , n70886 , n69553 );
not ( n72063 , n70886 );
not ( n72064 , n69553 );
and ( n72065 , n72063 , n72064 );
nor ( n72066 , n72062 , n72065 );
nand ( n72067 , n72061 , n72066 );
nand ( n72068 , n72003 , n70382 );
not ( n72069 , n70382 );
not ( n72070 , n71007 );
or ( n72071 , n72069 , n72070 );
or ( n72072 , n71007 , n70382 );
nand ( n72073 , n72071 , n72072 );
nand ( n72074 , n72073 , n72021 );
not ( n72075 , n70863 );
nor ( n72076 , n72064 , n72075 );
not ( n72077 , n72076 );
and ( n72078 , n72068 , n72074 , n72077 );
and ( n72079 , n72053 , n72060 , n72067 , n72078 );
nand ( n72080 , n72046 , n72079 );
buf ( n5938 , n72080 );
buf ( n72082 , 1'b0 );
not ( n72083 , n68842 );
buf ( n5941 , n72083 );
buf ( n72085 , n68638 );
and ( n72086 , n71276 , n70035 );
not ( n72087 , n71276 );
not ( n72088 , n70086 );
not ( n72089 , n72088 );
nand ( n72090 , n69975 , n70080 );
not ( n72091 , n70094 );
nor ( n72092 , n72090 , n72091 );
not ( n72093 , n72092 );
or ( n72094 , n72089 , n72093 );
or ( n72095 , n72092 , n72088 );
nand ( n72096 , n72094 , n72095 );
and ( n72097 , n72087 , n72096 );
nor ( n72098 , n72086 , n72097 );
or ( n72099 , n72098 , n71990 );
not ( n72100 , n70484 );
nand ( n72101 , n72100 , n70545 );
not ( n72102 , n72101 );
not ( n72103 , n70499 );
nor ( n72104 , n70940 , n72103 );
not ( n72105 , n72104 );
not ( n72106 , n70951 );
or ( n72107 , n72105 , n72106 );
not ( n72108 , n70954 );
or ( n72109 , n72108 , n72103 );
nand ( n72110 , n72109 , n70492 );
not ( n72111 , n72110 );
nand ( n72112 , n72107 , n72111 );
not ( n72113 , n72112 );
or ( n72114 , n72102 , n72113 );
or ( n72115 , n72112 , n72101 );
nand ( n72116 , n72114 , n72115 );
nand ( n72117 , n72116 , n72015 );
nand ( n72118 , n70621 , n70615 );
not ( n72119 , n72118 );
not ( n72120 , n70620 );
nor ( n72121 , n72120 , n70975 );
not ( n72122 , n72121 );
not ( n72123 , n70982 );
or ( n72124 , n72122 , n72123 );
not ( n72125 , n70620 );
not ( n72126 , n70773 );
or ( n72127 , n72125 , n72126 );
nand ( n72128 , n72127 , n70601 );
not ( n72129 , n72128 );
nand ( n72130 , n72124 , n72129 );
not ( n72131 , n72130 );
or ( n72132 , n72119 , n72131 );
or ( n72133 , n72130 , n72118 );
nand ( n72134 , n72132 , n72133 );
nand ( n72135 , n72134 , n72018 );
and ( n72136 , n70884 , n70885 );
not ( n72137 , n70884 );
and ( n72138 , n72137 , n3324 );
nor ( n72139 , n72136 , n72138 );
nand ( n72140 , n72061 , n72139 );
and ( n72141 , n72003 , n70392 );
nor ( n72142 , n70885 , n72075 );
not ( n72143 , n72142 );
not ( n72144 , n70392 );
not ( n72145 , n71004 );
not ( n72146 , n70436 );
not ( n72147 , n70822 );
nand ( n72148 , n72146 , n72147 );
or ( n72149 , n72148 , n70481 );
nor ( n72150 , n72145 , n72149 );
not ( n72151 , n72150 );
or ( n72152 , n72144 , n72151 );
or ( n72153 , n72150 , n70392 );
nand ( n72154 , n72152 , n72153 );
nand ( n72155 , n72154 , n72021 );
nand ( n72156 , n72143 , n72155 );
nor ( n72157 , n72141 , n72156 );
and ( n72158 , n72117 , n72135 , n72140 , n72157 );
nand ( n72159 , n72099 , n72158 );
buf ( n6017 , n72159 );
buf ( n6018 , 1'b0 );
not ( n72162 , n68842 );
buf ( n72163 , n72162 );
buf ( n72164 , n68638 );
and ( n72165 , n69363 , n70028 );
not ( n72166 , n69363 );
not ( n72167 , n70094 );
not ( n72168 , n72090 );
or ( n72169 , n72167 , n72168 );
or ( n72170 , n72090 , n70094 );
nand ( n72171 , n72169 , n72170 );
and ( n72172 , n72166 , n72171 );
nor ( n72173 , n72165 , n72172 );
or ( n72174 , n72173 , n71990 );
nand ( n72175 , n70620 , n70601 );
not ( n72176 , n72175 );
not ( n72177 , n70773 );
nand ( n72178 , n72177 , n70766 );
not ( n72179 , n72178 );
or ( n72180 , n72176 , n72179 );
or ( n72181 , n72178 , n72175 );
nand ( n72182 , n72180 , n72181 );
nand ( n72183 , n72182 , n72018 );
not ( n72184 , n72103 );
nand ( n72185 , n72184 , n70492 );
not ( n72186 , n72185 );
nor ( n72187 , n70940 , n70466 );
not ( n72188 , n72187 );
not ( n72189 , n70534 );
or ( n72190 , n72188 , n72189 );
nand ( n72191 , n72190 , n72108 );
not ( n72192 , n72191 );
or ( n72193 , n72186 , n72192 );
or ( n72194 , n72191 , n72185 );
nand ( n72195 , n72193 , n72194 );
nand ( n72196 , n72195 , n72015 );
and ( n72197 , n70883 , n3288 );
not ( n72198 , n70883 );
not ( n72199 , n3288 );
and ( n72200 , n72198 , n72199 );
nor ( n72201 , n72197 , n72200 );
nand ( n72202 , n72061 , n72201 );
and ( n72203 , n72003 , n70481 );
nor ( n72204 , n72199 , n72075 );
not ( n72205 , n72204 );
not ( n72206 , n70481 );
nor ( n72207 , n72145 , n72148 );
not ( n72208 , n72207 );
or ( n72209 , n72206 , n72208 );
or ( n72210 , n72207 , n70481 );
nand ( n72211 , n72209 , n72210 );
nand ( n72212 , n72211 , n72021 );
nand ( n72213 , n72205 , n72212 );
nor ( n72214 , n72203 , n72213 );
and ( n72215 , n72183 , n72196 , n72202 , n72214 );
nand ( n72216 , n72174 , n72215 );
buf ( n72217 , n72216 );
buf ( n72218 , 1'b0 );
not ( n72219 , n68842 );
buf ( n6077 , n72219 );
buf ( n6078 , n68638 );
and ( n72222 , n71276 , n70042 );
not ( n72223 , n71276 );
not ( n72224 , n70035 );
not ( n72225 , n70079 );
nand ( n72226 , n72225 , n69975 );
not ( n72227 , n72226 );
nand ( n72228 , n72227 , n70028 );
not ( n72229 , n72228 );
or ( n72230 , n72224 , n72229 );
or ( n72231 , n72228 , n70035 );
nand ( n72232 , n72230 , n72231 );
and ( n72233 , n72223 , n72232 );
nor ( n72234 , n72222 , n72233 );
or ( n72235 , n72234 , n71990 );
nand ( n72236 , n70543 , n70546 );
not ( n72237 , n72236 );
not ( n72238 , n70430 );
not ( n72239 , n72238 );
not ( n72240 , n70951 );
or ( n72241 , n72239 , n72240 );
nand ( n72242 , n72241 , n70539 );
not ( n72243 , n72242 );
or ( n72244 , n72237 , n72243 );
or ( n72245 , n72242 , n72236 );
nand ( n72246 , n72244 , n72245 );
nand ( n72247 , n72246 , n72015 );
nand ( n72248 , n70749 , n70772 );
not ( n72249 , n72248 );
not ( n72250 , n70763 );
not ( n72251 , n70982 );
or ( n72252 , n72250 , n72251 );
not ( n72253 , n70767 );
nand ( n72254 , n72252 , n72253 );
not ( n72255 , n72254 );
or ( n72256 , n72249 , n72255 );
or ( n72257 , n72254 , n72248 );
nand ( n72258 , n72256 , n72257 );
nand ( n72259 , n72258 , n72018 );
and ( n72260 , n70882 , n70881 );
not ( n72261 , n70882 );
and ( n72262 , n72261 , n3356 );
nor ( n72263 , n72260 , n72262 );
nand ( n72264 , n72061 , n72263 );
and ( n72265 , n72003 , n70436 );
nor ( n72266 , n70881 , n72075 );
not ( n72267 , n72266 );
not ( n72268 , n70436 );
nor ( n72269 , n72145 , n70822 );
not ( n72270 , n72269 );
or ( n72271 , n72268 , n72270 );
or ( n72272 , n72269 , n70436 );
nand ( n72273 , n72271 , n72272 );
nand ( n72274 , n72273 , n72021 );
nand ( n72275 , n72267 , n72274 );
nor ( n72276 , n72265 , n72275 );
and ( n72277 , n72247 , n72259 , n72264 , n72276 );
nand ( n72278 , n72235 , n72277 );
buf ( n72279 , n72278 );
buf ( n6137 , 1'b0 );
not ( n72281 , n68842 );
buf ( n72282 , n72281 );
buf ( n72283 , n68638 );
not ( n72284 , n69362 );
not ( n72285 , n70028 );
not ( n72286 , n72226 );
or ( n72287 , n72285 , n72286 );
or ( n72288 , n72226 , n70028 );
nand ( n72289 , n72287 , n72288 );
not ( n72290 , n72289 );
or ( n72291 , n72284 , n72290 );
nand ( n72292 , n70044 , n71276 );
nand ( n72293 , n72291 , n72292 );
not ( n72294 , n72293 );
or ( n72295 , n72294 , n71990 );
nand ( n72296 , n72238 , n70539 );
xnor ( n72297 , n70951 , n72296 );
nand ( n72298 , n72297 , n72015 );
nand ( n72299 , n70763 , n72253 );
not ( n72300 , n72299 );
not ( n72301 , n70982 );
or ( n72302 , n72300 , n72301 );
or ( n72303 , n70982 , n72299 );
nand ( n72304 , n72302 , n72303 );
nand ( n72305 , n72304 , n72018 );
not ( n72306 , n70821 );
and ( n72307 , n72003 , n72306 );
and ( n72308 , n71004 , n72147 );
not ( n72309 , n71004 );
and ( n72310 , n72309 , n70822 );
nor ( n72311 , n72308 , n72310 );
not ( n72312 , n72311 );
not ( n72313 , n72021 );
or ( n72314 , n72312 , n72313 );
nand ( n72315 , n3344 , n70863 );
nand ( n72316 , n72314 , n72315 );
nor ( n72317 , n72307 , n72316 );
nand ( n72318 , n72298 , n72305 , n72317 );
not ( n72319 , n3344 );
and ( n72320 , n72319 , n3304 );
not ( n72321 , n3304 );
and ( n72322 , n72321 , n3344 );
nor ( n72323 , n72320 , n72322 );
nor ( n72324 , n72007 , n72323 );
nor ( n72325 , n72318 , n72324 );
nand ( n72326 , n72295 , n72325 );
buf ( n72327 , n72326 );
buf ( n6185 , 1'b0 );
not ( n72329 , n68842 );
buf ( n72330 , n72329 );
buf ( n72331 , n68638 );
and ( n72332 , n69363 , n70077 );
not ( n72333 , n69363 );
not ( n72334 , n70077 );
nand ( n72335 , n69973 , n70057 );
nor ( n72336 , n72334 , n72335 );
nand ( n72337 , n72336 , n70044 );
not ( n72338 , n70042 );
and ( n72339 , n72337 , n72338 );
not ( n72340 , n72337 );
and ( n72341 , n72340 , n70042 );
nor ( n72342 , n72339 , n72341 );
and ( n72343 , n72333 , n72342 );
nor ( n72344 , n72332 , n72343 );
or ( n72345 , n72344 , n71990 );
not ( n72346 , n70944 );
nand ( n72347 , n72346 , n70532 );
nand ( n72348 , n70467 , n70531 );
xnor ( n72349 , n72347 , n72348 );
and ( n72350 , n72349 , n72015 );
and ( n72351 , n72003 , n70424 );
nor ( n72352 , n72350 , n72351 );
not ( n72353 , n70978 );
nand ( n72354 , n72353 , n70737 );
not ( n72355 , n72354 );
nand ( n72356 , n70765 , n70736 );
not ( n72357 , n72356 );
or ( n72358 , n72355 , n72357 );
or ( n72359 , n72356 , n72354 );
nand ( n72360 , n72358 , n72359 );
and ( n72361 , n72360 , n72018 );
not ( n72362 , n72021 );
not ( n72363 , n70424 );
not ( n72364 , n70835 );
nor ( n72365 , n72364 , n70463 );
not ( n72366 , n72365 );
or ( n72367 , n72363 , n72366 );
or ( n72368 , n72365 , n70424 );
nand ( n72369 , n72367 , n72368 );
not ( n72370 , n72369 );
or ( n72371 , n72362 , n72370 );
nor ( n72372 , n72321 , n72075 );
not ( n72373 , n72372 );
nand ( n72374 , n72371 , n72373 );
nor ( n72375 , n72361 , n72374 );
nand ( n72376 , n72061 , n72321 );
and ( n72377 , n72352 , n72375 , n72376 );
nand ( n72378 , n72345 , n72377 );
buf ( n72379 , n72378 );
buf ( n72380 , 1'b0 );
not ( n72381 , n68842 );
buf ( n72382 , n72381 );
buf ( n72383 , n68638 );
and ( n72384 , n71276 , n70057 );
not ( n72385 , n71276 );
xor ( n72386 , n70044 , n72336 );
and ( n72387 , n72385 , n72386 );
nor ( n72388 , n72384 , n72387 );
or ( n72389 , n72388 , n71990 );
nand ( n72390 , n72007 , n72075 );
and ( n72391 , n72390 , n70058 );
not ( n72392 , n72020 );
not ( n72393 , n70463 );
not ( n72394 , n70835 );
or ( n72395 , n72393 , n72394 );
or ( n72396 , n70835 , n70463 );
nand ( n72397 , n72395 , n72396 );
not ( n72398 , n72397 );
not ( n72399 , n72398 );
and ( n72400 , n72392 , n72399 );
not ( n72401 , n70520 );
nand ( n72402 , n72401 , n70532 );
not ( n72403 , n72402 );
or ( n72404 , n70511 , n70528 );
nand ( n72405 , n72404 , n70522 );
not ( n72406 , n72405 );
or ( n72407 , n72403 , n72406 );
or ( n72408 , n72402 , n72405 );
nand ( n72409 , n72407 , n72408 );
and ( n72410 , n72409 , n72015 );
nor ( n72411 , n72400 , n72410 );
not ( n72412 , n72003 );
not ( n72413 , n72412 );
not ( n72414 , n70463 );
not ( n72415 , n72414 );
and ( n72416 , n72413 , n72415 );
not ( n72417 , n70731 );
nand ( n72418 , n70720 , n70737 );
not ( n72419 , n72418 );
or ( n72420 , n72417 , n72419 );
or ( n72421 , n72418 , n70731 );
nand ( n72422 , n72420 , n72421 );
and ( n72423 , n72422 , n72018 );
nor ( n72424 , n72416 , n72423 );
nand ( n72425 , n72411 , n72424 );
nor ( n72426 , n72391 , n72425 );
nand ( n72427 , n72389 , n72426 );
buf ( n72428 , n72427 );
buf ( n72429 , 1'b0 );
not ( n72430 , n68842 );
buf ( n72431 , n72430 );
buf ( n72432 , n68638 );
and ( n72433 , n71276 , n71767 );
not ( n72434 , n71276 );
not ( n72435 , n71818 );
nand ( n72436 , n71856 , n71836 );
nor ( n72437 , n72435 , n72436 );
and ( n72438 , n71591 , n72437 , n71524 );
nand ( n72439 , n71041 , n71873 );
not ( n72440 , n72439 );
nand ( n72441 , n69664 , n71062 );
not ( n72442 , n72441 );
nand ( n72443 , n69981 , n70102 );
nor ( n72444 , n69986 , n72443 );
nand ( n72445 , n72440 , n72442 , n72444 , n71051 );
nor ( n72446 , n69974 , n72445 );
not ( n72447 , n71767 );
nand ( n72448 , n71801 , n71782 );
nor ( n72449 , n72447 , n72448 );
nand ( n72450 , n72438 , n72446 , n72449 );
not ( n72451 , n71750 );
not ( n72452 , n69711 );
nand ( n72453 , n72452 , n71758 );
not ( n72454 , n72453 );
nand ( n72455 , n72451 , n71755 , n72454 );
xnor ( n72456 , n72455 , n69733 );
not ( n72457 , n72456 );
nor ( n72458 , n72450 , n72457 );
not ( n72459 , n72458 );
not ( n72460 , n69747 );
not ( n72461 , n69733 );
nor ( n72462 , n72461 , n72453 );
nand ( n72463 , n72451 , n71755 , n72462 );
not ( n72464 , n72463 );
or ( n72465 , n72460 , n72464 );
or ( n72466 , n72463 , n69747 );
nand ( n72467 , n72465 , n72466 );
not ( n72468 , n72467 );
and ( n72469 , n72459 , n72468 );
not ( n72470 , n72459 );
and ( n72471 , n72470 , n72467 );
nor ( n72472 , n72469 , n72471 );
and ( n72473 , n72434 , n72472 );
nor ( n72474 , n72433 , n72473 );
or ( n72475 , n72474 , n71990 );
nor ( n72476 , n71135 , n71104 );
and ( n72477 , n72476 , n71089 );
nand ( n72478 , n70226 , n68650 );
not ( n72479 , n72478 );
not ( n72480 , n72479 );
not ( n72481 , n72480 );
not ( n72482 , n69900 );
not ( n72483 , n72482 );
or ( n72484 , n72481 , n72483 );
nand ( n72485 , n69900 , n72479 );
nand ( n72486 , n72484 , n72485 );
not ( n72487 , n69875 );
nand ( n72488 , n70226 , n2508 );
not ( n72489 , n72488 );
nor ( n72490 , n72487 , n72489 );
nor ( n72491 , n72486 , n72490 );
not ( n72492 , n72489 );
not ( n72493 , n69875 );
or ( n72494 , n72492 , n72493 );
not ( n72495 , n72489 );
not ( n72496 , n69875 );
nand ( n72497 , n72495 , n72496 );
nand ( n72498 , n72494 , n72497 );
nor ( n72499 , n71130 , n71126 );
nor ( n72500 , n72498 , n72499 );
nor ( n72501 , n72491 , n72500 );
nand ( n72502 , n70226 , n68649 );
not ( n72503 , n72502 );
not ( n72504 , n72503 );
not ( n72505 , n69796 );
or ( n72506 , n72504 , n72505 );
not ( n72507 , n72503 );
not ( n72508 , n69796 );
nand ( n72509 , n72507 , n72508 );
nand ( n72510 , n72506 , n72509 );
and ( n72511 , n69900 , n72480 );
nor ( n72512 , n72510 , n72511 );
nand ( n72513 , n70226 , n68648 );
not ( n72514 , n72513 );
not ( n72515 , n72514 );
not ( n72516 , n69773 );
or ( n72517 , n72515 , n72516 );
not ( n72518 , n69773 );
not ( n72519 , n72514 );
nand ( n72520 , n72518 , n72519 );
nand ( n72521 , n72517 , n72520 );
nor ( n72522 , n72508 , n72503 );
nor ( n72523 , n72521 , n72522 );
nor ( n72524 , n72512 , n72523 );
and ( n72525 , n72501 , n72524 );
nand ( n72526 , n72477 , n72525 );
and ( n72527 , n70226 , n2501 );
not ( n72528 , n72527 );
not ( n72529 , n69710 );
or ( n72530 , n72528 , n72529 );
not ( n72531 , n72527 );
not ( n72532 , n69710 );
nand ( n72533 , n72531 , n72532 );
nand ( n72534 , n72530 , n72533 );
not ( n72535 , n69689 );
not ( n72536 , n71074 );
nand ( n72537 , n72536 , n2502 );
not ( n72538 , n72537 );
nor ( n72539 , n72535 , n72538 );
nor ( n72540 , n72534 , n72539 );
not ( n72541 , n72538 );
not ( n72542 , n69689 );
or ( n72543 , n72541 , n72542 );
not ( n72544 , n72538 );
not ( n72545 , n69689 );
nand ( n72546 , n72544 , n72545 );
nand ( n72547 , n72543 , n72546 );
and ( n72548 , n70226 , n2503 );
not ( n72549 , n72548 );
and ( n72550 , n69854 , n72549 );
nor ( n72551 , n72547 , n72550 );
nor ( n72552 , n72540 , n72551 );
not ( n72553 , n72548 );
not ( n72554 , n69854 );
or ( n72555 , n72553 , n72554 );
not ( n72556 , n69854 );
nand ( n72557 , n72556 , n72549 );
nand ( n72558 , n72555 , n72557 );
not ( n72559 , n69936 );
nand ( n72560 , n72536 , n2504 );
not ( n72561 , n72560 );
nor ( n72562 , n72559 , n72561 );
nor ( n72563 , n72558 , n72562 );
not ( n72564 , n72561 );
not ( n72565 , n69936 );
or ( n72566 , n72564 , n72565 );
not ( n72567 , n72561 );
not ( n72568 , n69936 );
nand ( n72569 , n72567 , n72568 );
nand ( n72570 , n72566 , n72569 );
and ( n72571 , n69773 , n72519 );
nor ( n72572 , n72570 , n72571 );
nor ( n72573 , n72563 , n72572 );
nand ( n72574 , n72552 , n72573 );
nor ( n72575 , n72526 , n72574 );
not ( n72576 , n72575 );
not ( n72577 , n70557 );
or ( n72578 , n72576 , n72577 );
not ( n72579 , n72574 );
not ( n72580 , n72579 );
not ( n72581 , n72525 );
not ( n72582 , n71113 );
not ( n72583 , n72476 );
or ( n72584 , n72582 , n72583 );
not ( n72585 , n71135 );
not ( n72586 , n71116 );
and ( n72587 , n72585 , n72586 );
nor ( n72588 , n72587 , n71136 );
nand ( n72589 , n72584 , n72588 );
not ( n72590 , n72589 );
or ( n72591 , n72581 , n72590 );
not ( n72592 , n72524 );
and ( n72593 , n72498 , n72499 );
not ( n72594 , n72593 );
not ( n72595 , n72491 );
not ( n72596 , n72595 );
or ( n72597 , n72594 , n72596 );
nand ( n72598 , n72486 , n72490 );
nand ( n72599 , n72597 , n72598 );
not ( n72600 , n72599 );
or ( n72601 , n72592 , n72600 );
nand ( n72602 , n72510 , n72511 );
nor ( n72603 , n72523 , n72602 );
and ( n72604 , n72521 , n72522 );
nor ( n72605 , n72603 , n72604 );
nand ( n72606 , n72601 , n72605 );
not ( n72607 , n72606 );
nand ( n72608 , n72591 , n72607 );
not ( n72609 , n72608 );
or ( n72610 , n72580 , n72609 );
not ( n72611 , n72552 );
nand ( n72612 , n72570 , n72571 );
or ( n72613 , n72563 , n72612 );
nand ( n72614 , n72558 , n72562 );
nand ( n72615 , n72613 , n72614 );
not ( n72616 , n72615 );
or ( n72617 , n72611 , n72616 );
not ( n72618 , n72540 );
nand ( n72619 , n72547 , n72550 );
not ( n72620 , n72619 );
and ( n72621 , n72618 , n72620 );
and ( n72622 , n72534 , n72539 );
nor ( n72623 , n72621 , n72622 );
nand ( n72624 , n72617 , n72623 );
not ( n72625 , n72624 );
nand ( n72626 , n72610 , n72625 );
not ( n72627 , n72626 );
nand ( n72628 , n72578 , n72627 );
nand ( n72629 , n70226 , n2500 );
not ( n72630 , n72629 );
not ( n72631 , n72630 );
not ( n72632 , n69733 );
not ( n72633 , n72632 );
not ( n72634 , n72633 );
or ( n72635 , n72631 , n72634 );
not ( n72636 , n72630 );
not ( n72637 , n72633 );
nand ( n72638 , n72636 , n72637 );
nand ( n72639 , n72635 , n72638 );
not ( n72640 , n69710 );
nor ( n72641 , n72640 , n72527 );
nor ( n72642 , n72639 , n72641 );
not ( n72643 , n72642 );
nand ( n72644 , n72639 , n72641 );
nand ( n72645 , n72643 , n72644 );
not ( n72646 , n72645 );
and ( n72647 , n72628 , n72646 );
not ( n72648 , n72628 );
and ( n72649 , n72648 , n72645 );
nor ( n72650 , n72647 , n72649 );
nand ( n72651 , n72650 , n72015 );
xor ( n72652 , n72527 , n69710 );
and ( n72653 , n69689 , n72538 );
nor ( n72654 , n72652 , n72653 );
not ( n72655 , n69689 );
not ( n72656 , n72538 );
not ( n72657 , n72656 );
or ( n72658 , n72655 , n72657 );
not ( n72659 , n69689 );
nand ( n72660 , n72659 , n72538 );
nand ( n72661 , n72658 , n72660 );
and ( n72662 , n72548 , n69854 );
nor ( n72663 , n72661 , n72662 );
nor ( n72664 , n72654 , n72663 );
xor ( n72665 , n72548 , n69854 );
and ( n72666 , n69936 , n72561 );
nor ( n72667 , n72665 , n72666 );
not ( n72668 , n72561 );
not ( n72669 , n72668 );
not ( n72670 , n69936 );
or ( n72671 , n72669 , n72670 );
not ( n72672 , n69936 );
nand ( n72673 , n72672 , n72561 );
nand ( n72674 , n72671 , n72673 );
and ( n72675 , n69773 , n72514 );
nor ( n72676 , n72674 , n72675 );
nor ( n72677 , n72667 , n72676 );
and ( n72678 , n72664 , n72677 );
not ( n72679 , n72678 );
not ( n72680 , n72479 );
not ( n72681 , n69900 );
not ( n72682 , n72681 );
or ( n72683 , n72680 , n72682 );
not ( n72684 , n72479 );
nand ( n72685 , n72684 , n69900 );
nand ( n72686 , n72683 , n72685 );
and ( n72687 , n69875 , n72489 );
nor ( n72688 , n72686 , n72687 );
not ( n72689 , n72688 );
not ( n72690 , n72489 );
not ( n72691 , n69875 );
not ( n72692 , n72691 );
or ( n72693 , n72690 , n72692 );
not ( n72694 , n72489 );
nand ( n72695 , n72694 , n69875 );
nand ( n72696 , n72693 , n72695 );
not ( n72697 , n72696 );
and ( n72698 , n69808 , n71126 );
not ( n72699 , n72698 );
nand ( n72700 , n72697 , n72699 );
nand ( n72701 , n72689 , n72700 );
not ( n72702 , n72701 );
not ( n72703 , n72503 );
not ( n72704 , n69796 );
not ( n72705 , n72704 );
or ( n72706 , n72703 , n72705 );
not ( n72707 , n72503 );
nand ( n72708 , n69796 , n72707 );
nand ( n72709 , n72706 , n72708 );
and ( n72710 , n69900 , n72479 );
nor ( n72711 , n72709 , n72710 );
not ( n72712 , n72514 );
not ( n72713 , n72712 );
not ( n72714 , n69773 );
or ( n72715 , n72713 , n72714 );
not ( n72716 , n69773 );
nand ( n72717 , n72716 , n72514 );
nand ( n72718 , n72715 , n72717 );
nand ( n72719 , n69796 , n72503 );
not ( n72720 , n72719 );
nor ( n72721 , n72718 , n72720 );
nor ( n72722 , n72711 , n72721 );
nand ( n72723 , n72702 , n72722 );
not ( n72724 , n72723 );
nor ( n72725 , n71173 , n71150 );
not ( n72726 , n72725 );
nor ( n72727 , n72726 , n71164 );
nand ( n72728 , n72724 , n72727 );
nor ( n72729 , n72679 , n72728 );
not ( n72730 , n72729 );
not ( n72731 , n70813 );
or ( n72732 , n72730 , n72731 );
nand ( n72733 , n72709 , n72710 );
or ( n72734 , n72721 , n72733 );
nand ( n72735 , n72718 , n72720 );
nand ( n72736 , n72734 , n72735 );
not ( n72737 , n72736 );
not ( n72738 , n72722 );
and ( n72739 , n72737 , n72738 );
nand ( n72740 , n72696 , n72698 );
or ( n72741 , n72688 , n72740 );
nand ( n72742 , n72686 , n72687 );
nand ( n72743 , n72741 , n72742 );
nor ( n72744 , n72736 , n72743 );
and ( n72745 , n72744 , n72701 );
nor ( n72746 , n72739 , n72745 );
nand ( n72747 , n71182 , n72725 );
not ( n72748 , n71150 );
not ( n72749 , n71185 );
and ( n72750 , n72748 , n72749 );
nor ( n72751 , n72750 , n71149 );
nand ( n72752 , n72744 , n72747 , n72751 );
nand ( n72753 , n72746 , n72752 );
not ( n72754 , n72753 );
and ( n72755 , n72754 , n72678 );
not ( n72756 , n72664 );
nand ( n72757 , n72674 , n72675 );
or ( n72758 , n72667 , n72757 );
nand ( n72759 , n72665 , n72666 );
nand ( n72760 , n72758 , n72759 );
not ( n72761 , n72760 );
or ( n72762 , n72756 , n72761 );
not ( n72763 , n72654 );
nand ( n72764 , n72661 , n72662 );
not ( n72765 , n72764 );
and ( n72766 , n72763 , n72765 );
nand ( n72767 , n72652 , n72653 );
not ( n72768 , n72767 );
nor ( n72769 , n72766 , n72768 );
nand ( n72770 , n72762 , n72769 );
nor ( n72771 , n72755 , n72770 );
nand ( n72772 , n72732 , n72771 );
xor ( n72773 , n72630 , n69733 );
and ( n72774 , n72527 , n69710 );
or ( n72775 , n72773 , n72774 );
nand ( n72776 , n72773 , n72774 );
nand ( n72777 , n72775 , n72776 );
not ( n72778 , n72777 );
and ( n72779 , n72772 , n72778 );
not ( n72780 , n72772 );
and ( n72781 , n72780 , n72777 );
nor ( n72782 , n72779 , n72781 );
and ( n72783 , n72782 , n72018 );
not ( n72784 , n69724 );
not ( n72785 , n69706 );
nor ( n72786 , n70897 , n70898 );
nand ( n72787 , n72786 , n3514 );
not ( n72788 , n69822 );
nor ( n72789 , n72787 , n72788 );
nand ( n72790 , n72789 , n69806 );
not ( n72791 , n69855 );
nor ( n72792 , n72790 , n72791 );
and ( n72793 , n72792 , n69891 );
nand ( n72794 , n72793 , n69776 );
not ( n72795 , n69770 );
nor ( n72796 , n72794 , n72795 );
nand ( n72797 , n72796 , n69932 );
not ( n72798 , n3707 );
nor ( n72799 , n72797 , n72798 );
nand ( n72800 , n72799 , n69680 );
nor ( n72801 , n72785 , n72800 );
not ( n72802 , n72801 );
or ( n72803 , n72784 , n72802 );
or ( n72804 , n72801 , n69724 );
nand ( n72805 , n72803 , n72804 );
not ( n72806 , n72805 );
or ( n72807 , n72806 , n72007 );
not ( n72808 , n72630 );
not ( n72809 , n71096 );
not ( n72810 , n71126 );
nand ( n72811 , n72809 , n72810 );
nor ( n72812 , n72811 , n71198 );
nor ( n72813 , n72503 , n72514 );
nor ( n72814 , n72489 , n72479 );
and ( n72815 , n72813 , n72814 );
and ( n72816 , n72812 , n72815 );
nor ( n72817 , n72561 , n72548 );
not ( n72818 , n72527 );
not ( n72819 , n72818 );
nor ( n72820 , n72819 , n72538 );
and ( n72821 , n72817 , n72820 );
nand ( n72822 , n72816 , n72821 );
nor ( n72823 , n70836 , n72822 );
not ( n72824 , n72823 );
or ( n72825 , n72808 , n72824 );
or ( n72826 , n72823 , n72630 );
nand ( n72827 , n72825 , n72826 );
nand ( n72828 , n72827 , n72021 );
nand ( n72829 , n72003 , n72630 );
nand ( n72830 , n69725 , n70863 );
and ( n72831 , n72828 , n72829 , n72830 );
nand ( n72832 , n72807 , n72831 );
nor ( n72833 , n72783 , n72832 );
and ( n72834 , n72651 , n72833 );
nand ( n72835 , n72475 , n72834 );
buf ( n72836 , n72835 );
buf ( n72837 , 1'b0 );
not ( n72838 , n68842 );
buf ( n6696 , n72838 );
buf ( n6697 , n68638 );
and ( n72841 , n69363 , n71784 );
not ( n72842 , n69363 );
and ( n72843 , n72450 , n72457 );
not ( n72844 , n72450 );
not ( n72845 , n72457 );
and ( n72846 , n72844 , n72845 );
nor ( n72847 , n72843 , n72846 );
and ( n72848 , n72842 , n72847 );
nor ( n72849 , n72841 , n72848 );
or ( n72850 , n72849 , n71990 );
not ( n72851 , n72551 );
and ( n72852 , n72573 , n72851 );
not ( n72853 , n72852 );
nor ( n72854 , n72526 , n72853 );
not ( n72855 , n72854 );
not ( n72856 , n70557 );
or ( n72857 , n72855 , n72856 );
not ( n72858 , n72852 );
not ( n72859 , n72608 );
or ( n72860 , n72858 , n72859 );
not ( n72861 , n72851 );
not ( n72862 , n72615 );
or ( n72863 , n72861 , n72862 );
nand ( n72864 , n72863 , n72619 );
not ( n72865 , n72864 );
nand ( n72866 , n72860 , n72865 );
not ( n72867 , n72866 );
nand ( n72868 , n72857 , n72867 );
or ( n72869 , n72540 , n72622 );
xnor ( n72870 , n72868 , n72869 );
nand ( n72871 , n72870 , n72015 );
not ( n72872 , n72654 );
nand ( n72873 , n72872 , n72767 );
not ( n72874 , n72873 );
not ( n72875 , n72663 );
nand ( n72876 , n72677 , n72875 );
nor ( n72877 , n72728 , n72876 );
not ( n72878 , n72877 );
not ( n72879 , n70808 );
or ( n72880 , n72878 , n72879 );
not ( n72881 , n72753 );
not ( n72882 , n72876 );
and ( n72883 , n72881 , n72882 );
not ( n72884 , n72875 );
not ( n72885 , n72760 );
or ( n72886 , n72884 , n72885 );
nand ( n72887 , n72886 , n72764 );
nor ( n72888 , n72883 , n72887 );
nand ( n72889 , n72880 , n72888 );
not ( n72890 , n72889 );
or ( n72891 , n72874 , n72890 );
or ( n72892 , n72889 , n72873 );
nand ( n72893 , n72891 , n72892 );
and ( n72894 , n72893 , n72018 );
and ( n72895 , n72800 , n69706 );
not ( n72896 , n72800 );
and ( n72897 , n72896 , n69705 );
nor ( n72898 , n72895 , n72897 );
or ( n72899 , n72007 , n72898 );
not ( n72900 , n72819 );
not ( n72901 , n72561 );
nor ( n72902 , n72811 , n70229 );
nor ( n72903 , n72548 , n72538 );
and ( n72904 , n72813 , n72903 , n71197 );
nand ( n72905 , n72901 , n72902 , n72904 , n72814 );
nor ( n72906 , n70836 , n72905 );
not ( n72907 , n72906 );
or ( n72908 , n72900 , n72907 );
or ( n72909 , n72906 , n72819 );
nand ( n72910 , n72908 , n72909 );
and ( n72911 , n72910 , n72021 );
nor ( n72912 , n69705 , n72075 );
nor ( n72913 , n72911 , n72912 );
nand ( n72914 , n72003 , n72819 );
nand ( n72915 , n72899 , n72913 , n72914 );
nor ( n72916 , n72894 , n72915 );
and ( n72917 , n72871 , n72916 );
nand ( n72918 , n72850 , n72917 );
buf ( n72919 , n72918 );
buf ( n6777 , 1'b0 );
not ( n72921 , n68842 );
buf ( n72922 , n72921 );
buf ( n72923 , n68638 );
and ( n72924 , n71276 , n71803 );
not ( n72925 , n71276 );
not ( n72926 , n72445 );
nand ( n72927 , n72926 , n72438 );
not ( n72928 , n72927 );
not ( n72929 , n72448 );
nand ( n72930 , n72928 , n69973 , n72929 );
not ( n72931 , n71767 );
and ( n72932 , n72930 , n72931 );
not ( n72933 , n72930 );
and ( n72934 , n72933 , n71767 );
nor ( n72935 , n72932 , n72934 );
and ( n72936 , n72925 , n72935 );
nor ( n72937 , n72924 , n72936 );
or ( n72938 , n72937 , n71990 );
not ( n72939 , n72573 );
nor ( n72940 , n72939 , n72526 );
not ( n72941 , n72940 );
not ( n72942 , n70557 );
or ( n72943 , n72941 , n72942 );
not ( n72944 , n72573 );
not ( n72945 , n72608 );
or ( n72946 , n72944 , n72945 );
not ( n72947 , n72615 );
nand ( n72948 , n72946 , n72947 );
not ( n72949 , n72948 );
nand ( n72950 , n72943 , n72949 );
nand ( n72951 , n72851 , n72619 );
not ( n72952 , n72951 );
and ( n72953 , n72950 , n72952 );
not ( n72954 , n72950 );
and ( n72955 , n72954 , n72951 );
nor ( n72956 , n72953 , n72955 );
nand ( n72957 , n72956 , n72015 );
not ( n72958 , n72677 );
nor ( n72959 , n72728 , n72958 );
not ( n72960 , n72959 );
not ( n72961 , n70808 );
or ( n72962 , n72960 , n72961 );
and ( n72963 , n72754 , n72677 );
nor ( n72964 , n72963 , n72760 );
nand ( n72965 , n72962 , n72964 );
nand ( n72966 , n72875 , n72764 );
not ( n72967 , n72966 );
and ( n72968 , n72965 , n72967 );
not ( n72969 , n72965 );
and ( n72970 , n72969 , n72966 );
nor ( n72971 , n72968 , n72970 );
and ( n72972 , n72971 , n72018 );
and ( n72973 , n72799 , n69679 );
not ( n72974 , n72799 );
and ( n72975 , n72974 , n69680 );
nor ( n72976 , n72973 , n72975 );
or ( n72977 , n72007 , n72976 );
not ( n72978 , n72538 );
not ( n72979 , n72811 );
not ( n72980 , n71198 );
nand ( n72981 , n72979 , n72980 , n72815 , n72817 );
nor ( n72982 , n70836 , n72981 );
not ( n72983 , n72982 );
or ( n72984 , n72978 , n72983 );
or ( n72985 , n72982 , n72538 );
nand ( n72986 , n72984 , n72985 );
and ( n72987 , n72986 , n72021 );
nor ( n72988 , n69679 , n72075 );
nor ( n72989 , n72987 , n72988 );
nand ( n72990 , n72003 , n72538 );
nand ( n72991 , n72977 , n72989 , n72990 );
nor ( n72992 , n72972 , n72991 );
and ( n72993 , n72957 , n72992 );
nand ( n72994 , n72938 , n72993 );
buf ( n6852 , n72994 );
buf ( n6853 , 1'b0 );
not ( n72997 , n68842 );
buf ( n72998 , n72997 );
buf ( n72999 , n68638 );
and ( n73000 , n69363 , n71818 );
not ( n73001 , n69363 );
not ( n73002 , n69973 );
nor ( n73003 , n72927 , n73002 );
nand ( n73004 , n73003 , n71801 );
not ( n73005 , n71782 );
and ( n73006 , n73004 , n73005 );
not ( n73007 , n73004 );
and ( n73008 , n73007 , n71782 );
nor ( n73009 , n73006 , n73008 );
and ( n73010 , n73001 , n73009 );
nor ( n73011 , n73000 , n73010 );
or ( n73012 , n73011 , n71990 );
nor ( n73013 , n72526 , n72572 );
not ( n73014 , n73013 );
not ( n73015 , n70557 );
or ( n73016 , n73014 , n73015 );
not ( n73017 , n72572 );
not ( n73018 , n73017 );
not ( n73019 , n72608 );
or ( n73020 , n73018 , n73019 );
nand ( n73021 , n73020 , n72612 );
not ( n73022 , n73021 );
nand ( n73023 , n73016 , n73022 );
not ( n73024 , n72563 );
nand ( n73025 , n73024 , n72614 );
xnor ( n73026 , n73023 , n73025 );
nand ( n73027 , n73026 , n72015 );
not ( n73028 , n72667 );
nand ( n73029 , n73028 , n72759 );
not ( n73030 , n73029 );
nor ( n73031 , n72728 , n72676 );
not ( n73032 , n73031 );
not ( n73033 , n70808 );
or ( n73034 , n73032 , n73033 );
not ( n73035 , n72753 );
not ( n73036 , n72676 );
and ( n73037 , n73035 , n73036 );
not ( n73038 , n72757 );
nor ( n73039 , n73037 , n73038 );
nand ( n73040 , n73034 , n73039 );
not ( n73041 , n73040 );
or ( n73042 , n73030 , n73041 );
or ( n73043 , n73040 , n73029 );
nand ( n73044 , n73042 , n73043 );
and ( n73045 , n73044 , n72018 );
and ( n73046 , n72797 , n3707 );
not ( n73047 , n72797 );
and ( n73048 , n73047 , n72798 );
nor ( n73049 , n73046 , n73048 );
or ( n73050 , n72007 , n73049 );
not ( n73051 , n72548 );
not ( n73052 , n72503 );
and ( n73053 , n72814 , n73052 );
nor ( n73054 , n71078 , n72561 , n72514 );
nand ( n73055 , n72902 , n73053 , n73054 );
nor ( n73056 , n70836 , n73055 );
not ( n73057 , n73056 );
or ( n73058 , n73051 , n73057 );
or ( n73059 , n73056 , n72548 );
nand ( n73060 , n73058 , n73059 );
and ( n73061 , n73060 , n72021 );
nor ( n73062 , n72798 , n72075 );
nor ( n73063 , n73061 , n73062 );
nand ( n73064 , n72003 , n72548 );
nand ( n73065 , n73050 , n73063 , n73064 );
nor ( n73066 , n73045 , n73065 );
and ( n73067 , n73027 , n73066 );
nand ( n73068 , n73012 , n73067 );
buf ( n73069 , n73068 );
buf ( n6927 , 1'b0 );
not ( n73071 , n68842 );
buf ( n73072 , n73071 );
buf ( n73073 , n68638 );
and ( n73074 , n71276 , n71838 );
not ( n73075 , n71276 );
not ( n73076 , n73003 );
not ( n73077 , n71801 );
and ( n73078 , n73076 , n73077 );
not ( n73079 , n73076 );
and ( n73080 , n73079 , n71801 );
nor ( n73081 , n73078 , n73080 );
and ( n73082 , n73075 , n73081 );
nor ( n73083 , n73074 , n73082 );
or ( n73084 , n73083 , n71990 );
not ( n73085 , n72526 );
not ( n73086 , n73085 );
not ( n73087 , n70557 );
or ( n73088 , n73086 , n73087 );
not ( n73089 , n72608 );
nand ( n73090 , n73088 , n73089 );
nand ( n73091 , n73017 , n72612 );
not ( n73092 , n73091 );
and ( n73093 , n73090 , n73092 );
not ( n73094 , n73090 );
and ( n73095 , n73094 , n73091 );
nor ( n73096 , n73093 , n73095 );
nand ( n73097 , n73096 , n72015 );
not ( n73098 , n72728 );
not ( n73099 , n73098 );
not ( n73100 , n70813 );
or ( n73101 , n73099 , n73100 );
nand ( n73102 , n73101 , n72753 );
nor ( n73103 , n73038 , n72676 );
and ( n73104 , n73102 , n73103 );
not ( n73105 , n73102 );
not ( n73106 , n73103 );
and ( n73107 , n73105 , n73106 );
nor ( n73108 , n73104 , n73107 );
and ( n73109 , n73108 , n72018 );
and ( n73110 , n72796 , n69931 );
not ( n73111 , n72796 );
and ( n73112 , n73111 , n69932 );
nor ( n73113 , n73110 , n73112 );
or ( n73114 , n72007 , n73113 );
not ( n73115 , n72561 );
not ( n73116 , n72816 );
nor ( n73117 , n73116 , n70836 );
not ( n73118 , n73117 );
or ( n73119 , n73115 , n73118 );
or ( n73120 , n73117 , n72561 );
nand ( n73121 , n73119 , n73120 );
and ( n73122 , n73121 , n72021 );
nor ( n73123 , n69931 , n72075 );
nor ( n73124 , n73122 , n73123 );
nand ( n73125 , n72003 , n72561 );
nand ( n73126 , n73114 , n73124 , n73125 );
nor ( n73127 , n73109 , n73126 );
and ( n73128 , n73097 , n73127 );
nand ( n73129 , n73084 , n73128 );
buf ( n6987 , n73129 );
buf ( n6988 , 1'b0 );
not ( n73132 , n68842 );
buf ( n73133 , n73132 );
buf ( n73134 , n68638 );
and ( n73135 , n69363 , n71856 );
not ( n73136 , n69363 );
nor ( n73137 , n72445 , n71526 );
nand ( n73138 , n73137 , n71856 );
not ( n73139 , n73138 );
nand ( n73140 , n73139 , n71836 );
not ( n73141 , n71818 );
and ( n73142 , n73140 , n73141 );
not ( n73143 , n73140 );
and ( n73144 , n73143 , n71818 );
nor ( n73145 , n73142 , n73144 );
and ( n73146 , n73136 , n73145 );
nor ( n73147 , n73135 , n73146 );
or ( n73148 , n73147 , n71990 );
not ( n73149 , n72477 );
not ( n73150 , n72512 );
and ( n73151 , n72501 , n73150 );
not ( n73152 , n73151 );
nor ( n73153 , n73149 , n73152 );
not ( n73154 , n73153 );
not ( n73155 , n70557 );
or ( n73156 , n73154 , n73155 );
and ( n73157 , n73151 , n72589 );
not ( n73158 , n73150 );
not ( n73159 , n72599 );
or ( n73160 , n73158 , n73159 );
nand ( n73161 , n73160 , n72602 );
nor ( n73162 , n73157 , n73161 );
nand ( n73163 , n73156 , n73162 );
or ( n73164 , n72604 , n72523 );
xnor ( n73165 , n73163 , n73164 );
nand ( n73166 , n73165 , n72015 );
not ( n73167 , n72721 );
nand ( n73168 , n73167 , n72735 );
not ( n73169 , n73168 );
nor ( n73170 , n72701 , n72711 );
not ( n73171 , n73170 );
not ( n73172 , n72727 );
nor ( n73173 , n73171 , n73172 );
not ( n73174 , n73173 );
not ( n73175 , n70813 );
or ( n73176 , n73174 , n73175 );
not ( n73177 , n73170 );
nand ( n73178 , n72747 , n72751 );
not ( n73179 , n73178 );
or ( n73180 , n73177 , n73179 );
not ( n73181 , n72711 );
not ( n73182 , n73181 );
not ( n73183 , n72743 );
or ( n73184 , n73182 , n73183 );
nand ( n73185 , n73184 , n72733 );
not ( n73186 , n73185 );
nand ( n73187 , n73180 , n73186 );
not ( n73188 , n73187 );
nand ( n73189 , n73176 , n73188 );
not ( n73190 , n73189 );
or ( n73191 , n73169 , n73190 );
or ( n73192 , n73189 , n73168 );
nand ( n73193 , n73191 , n73192 );
and ( n73194 , n73193 , n72018 );
and ( n73195 , n72794 , n69770 );
not ( n73196 , n72794 );
and ( n73197 , n73196 , n72795 );
nor ( n73198 , n73195 , n73197 );
or ( n73199 , n72007 , n73198 );
not ( n73200 , n72514 );
nand ( n73201 , n72812 , n73053 );
nor ( n73202 , n70836 , n73201 );
not ( n73203 , n73202 );
or ( n73204 , n73200 , n73203 );
or ( n73205 , n73202 , n72514 );
nand ( n73206 , n73204 , n73205 );
and ( n73207 , n73206 , n72021 );
nor ( n73208 , n72795 , n72075 );
nor ( n73209 , n73207 , n73208 );
nand ( n73210 , n72003 , n72514 );
nand ( n73211 , n73199 , n73209 , n73210 );
nor ( n73212 , n73194 , n73211 );
and ( n73213 , n73166 , n73212 );
nand ( n73214 , n73148 , n73213 );
buf ( n73215 , n73214 );
buf ( n73216 , 1'b0 );
not ( n73217 , n68842 );
buf ( n73218 , n73217 );
buf ( n73219 , n68638 );
and ( n73220 , n71276 , n71873 );
not ( n73221 , n71276 );
not ( n73222 , n71836 );
and ( n73223 , n73138 , n73222 );
not ( n73224 , n73138 );
and ( n73225 , n73224 , n71836 );
nor ( n73226 , n73223 , n73225 );
and ( n73227 , n73221 , n73226 );
nor ( n73228 , n73220 , n73227 );
or ( n73229 , n73228 , n71990 );
not ( n73230 , n72501 );
nor ( n73231 , n73149 , n73230 );
not ( n73232 , n73231 );
not ( n73233 , n70557 );
or ( n73234 , n73232 , n73233 );
and ( n73235 , n72501 , n72589 );
nor ( n73236 , n73235 , n72599 );
nand ( n73237 , n73234 , n73236 );
nand ( n73238 , n73150 , n72602 );
not ( n73239 , n73238 );
and ( n73240 , n73237 , n73239 );
not ( n73241 , n73237 );
and ( n73242 , n73241 , n73238 );
nor ( n73243 , n73240 , n73242 );
nand ( n73244 , n73243 , n72015 );
nor ( n73245 , n73172 , n72701 );
not ( n73246 , n73245 );
not ( n73247 , n70813 );
or ( n73248 , n73246 , n73247 );
and ( n73249 , n72702 , n73178 );
nor ( n73250 , n73249 , n72743 );
nand ( n73251 , n73248 , n73250 );
nand ( n73252 , n73181 , n72733 );
not ( n73253 , n73252 );
and ( n73254 , n73251 , n73253 );
not ( n73255 , n73251 );
and ( n73256 , n73255 , n73252 );
nor ( n73257 , n73254 , n73256 );
and ( n73258 , n73257 , n72018 );
and ( n73259 , n72793 , n69775 );
not ( n73260 , n72793 );
and ( n73261 , n73260 , n69776 );
nor ( n73262 , n73259 , n73261 );
or ( n73263 , n72007 , n73262 );
not ( n73264 , n72503 );
nand ( n73265 , n72812 , n72814 );
nor ( n73266 , n70836 , n73265 );
not ( n73267 , n73266 );
or ( n73268 , n73264 , n73267 );
or ( n73269 , n73266 , n72503 );
nand ( n73270 , n73268 , n73269 );
and ( n73271 , n73270 , n72021 );
nor ( n73272 , n69775 , n72075 );
nor ( n73273 , n73271 , n73272 );
nand ( n73274 , n72003 , n72503 );
nand ( n73275 , n73263 , n73273 , n73274 );
nor ( n73276 , n73258 , n73275 );
and ( n73277 , n73244 , n73276 );
nand ( n73278 , n73229 , n73277 );
buf ( n73279 , n73278 );
buf ( n73280 , 1'b0 );
not ( n73281 , n68842 );
buf ( n7139 , n73281 );
buf ( n7140 , n68638 );
and ( n73284 , n69363 , n71041 );
not ( n73285 , n69363 );
not ( n73286 , n71856 );
not ( n73287 , n73137 );
not ( n73288 , n73287 );
or ( n73289 , n73286 , n73288 );
or ( n73290 , n71856 , n73287 );
nand ( n73291 , n73289 , n73290 );
and ( n73292 , n73285 , n73291 );
nor ( n73293 , n73284 , n73292 );
or ( n73294 , n73293 , n71990 );
nor ( n73295 , n73149 , n72500 );
not ( n73296 , n73295 );
not ( n73297 , n70557 );
or ( n73298 , n73296 , n73297 );
not ( n73299 , n72500 );
not ( n73300 , n73299 );
not ( n73301 , n72589 );
or ( n73302 , n73300 , n73301 );
not ( n73303 , n72593 );
nand ( n73304 , n73302 , n73303 );
not ( n73305 , n73304 );
nand ( n73306 , n73298 , n73305 );
nand ( n73307 , n72595 , n72598 );
xnor ( n73308 , n73306 , n73307 );
nand ( n73309 , n73308 , n72015 );
not ( n73310 , n72688 );
nand ( n73311 , n73310 , n72742 );
not ( n73312 , n73311 );
not ( n73313 , n72700 );
nor ( n73314 , n73313 , n73172 );
not ( n73315 , n73314 );
not ( n73316 , n70813 );
or ( n73317 , n73315 , n73316 );
not ( n73318 , n72700 );
not ( n73319 , n73178 );
or ( n73320 , n73318 , n73319 );
nand ( n73321 , n73320 , n72740 );
not ( n73322 , n73321 );
nand ( n73323 , n73317 , n73322 );
not ( n73324 , n73323 );
or ( n73325 , n73312 , n73324 );
or ( n73326 , n73323 , n73311 );
nand ( n73327 , n73325 , n73326 );
and ( n73328 , n72018 , n73327 );
and ( n73329 , n72792 , n69890 );
not ( n73330 , n72792 );
and ( n73331 , n73330 , n69891 );
nor ( n73332 , n73329 , n73331 );
or ( n73333 , n72007 , n73332 );
not ( n73334 , n72479 );
not ( n73335 , n72489 );
nand ( n73336 , n73335 , n72812 );
nor ( n73337 , n70836 , n73336 );
not ( n73338 , n73337 );
or ( n73339 , n73334 , n73338 );
or ( n73340 , n73337 , n72479 );
nand ( n73341 , n73339 , n73340 );
and ( n73342 , n73341 , n72021 );
nor ( n73343 , n69890 , n72075 );
nor ( n73344 , n73342 , n73343 );
nand ( n73345 , n72003 , n72479 );
nand ( n73346 , n73333 , n73344 , n73345 );
nor ( n73347 , n73328 , n73346 );
and ( n73348 , n73309 , n73347 );
nand ( n73349 , n73294 , n73348 );
buf ( n73350 , n73349 );
buf ( n7208 , 1'b0 );
not ( n73352 , n68842 );
buf ( n73353 , n73352 );
buf ( n73354 , n68638 );
and ( n73355 , n71276 , n71062 );
not ( n73356 , n71276 );
not ( n73357 , n71063 );
nand ( n73358 , n73357 , n71041 );
not ( n73359 , n71873 );
and ( n73360 , n73358 , n73359 );
not ( n73361 , n73358 );
and ( n73362 , n73361 , n71873 );
nor ( n73363 , n73360 , n73362 );
and ( n73364 , n73356 , n73363 );
nor ( n73365 , n73355 , n73364 );
or ( n73366 , n73365 , n71990 );
not ( n73367 , n72477 );
not ( n73368 , n70557 );
or ( n73369 , n73367 , n73368 );
not ( n73370 , n72589 );
nand ( n73371 , n73369 , n73370 );
nand ( n73372 , n73299 , n73303 );
xnor ( n73373 , n73371 , n73372 );
nand ( n73374 , n73373 , n72015 );
nand ( n73375 , n72700 , n72740 );
not ( n73376 , n73375 );
not ( n73377 , n72727 );
not ( n73378 , n70813 );
or ( n73379 , n73377 , n73378 );
not ( n73380 , n73178 );
nand ( n73381 , n73379 , n73380 );
not ( n73382 , n73381 );
or ( n73383 , n73376 , n73382 );
or ( n73384 , n73381 , n73375 );
nand ( n73385 , n73383 , n73384 );
and ( n73386 , n73385 , n72018 );
and ( n73387 , n72790 , n69855 );
not ( n73388 , n72790 );
and ( n73389 , n73388 , n72791 );
nor ( n73390 , n73387 , n73389 );
or ( n73391 , n72007 , n73390 );
not ( n73392 , n72489 );
not ( n73393 , n72812 );
nor ( n73394 , n70836 , n73393 );
not ( n73395 , n73394 );
or ( n73396 , n73392 , n73395 );
or ( n73397 , n73394 , n72489 );
nand ( n73398 , n73396 , n73397 );
and ( n73399 , n73398 , n72021 );
nor ( n73400 , n72791 , n72075 );
nor ( n73401 , n73399 , n73400 );
nand ( n73402 , n72003 , n72489 );
nand ( n73403 , n73391 , n73401 , n73402 );
nor ( n73404 , n73386 , n73403 );
and ( n73405 , n73374 , n73404 );
nand ( n73406 , n73366 , n73405 );
buf ( n73407 , n73406 );
buf ( n73408 , 1'b0 );
not ( n73409 , n68842 );
buf ( n73410 , n73409 );
buf ( n73411 , n68638 );
and ( n73412 , n71276 , n69971 );
not ( n73413 , n71276 );
not ( n73414 , n70077 );
not ( n73415 , n72335 );
or ( n73416 , n73414 , n73415 );
or ( n73417 , n72335 , n70077 );
nand ( n73418 , n73416 , n73417 );
and ( n73419 , n73413 , n73418 );
nor ( n73420 , n73412 , n73419 );
or ( n73421 , n73420 , n71990 );
and ( n73422 , n72390 , n70045 );
not ( n73423 , n70528 );
not ( n73424 , n73423 );
not ( n73425 , n70511 );
nand ( n73426 , n73425 , n70522 );
not ( n73427 , n73426 );
or ( n73428 , n73424 , n73427 );
or ( n73429 , n73426 , n73423 );
nand ( n73430 , n73428 , n73429 );
nand ( n73431 , n73430 , n72015 );
xor ( n73432 , n70726 , n70729 );
nand ( n73433 , n72018 , n73432 );
nand ( n73434 , n72003 , n70507 );
not ( n73435 , n70833 );
not ( n73436 , n70526 );
or ( n73437 , n73435 , n73436 );
or ( n73438 , n70526 , n70833 );
nand ( n73439 , n73437 , n73438 );
nand ( n73440 , n72021 , n73439 );
nand ( n73441 , n73431 , n73433 , n73434 , n73440 );
nor ( n73442 , n73422 , n73441 );
nand ( n73443 , n73421 , n73442 );
buf ( n73444 , n73443 );
buf ( n73445 , 1'b0 );
not ( n73446 , n68842 );
buf ( n73447 , n73446 );
buf ( n73448 , n68638 );
not ( n73449 , n71071 );
or ( n73450 , n73449 , n71990 );
nand ( n73451 , n71138 , n72015 );
and ( n73452 , n71192 , n72018 );
not ( n73453 , n69806 );
and ( n73454 , n72789 , n73453 );
not ( n73455 , n72789 );
and ( n73456 , n73455 , n69806 );
nor ( n73457 , n73454 , n73456 );
or ( n73458 , n72007 , n73457 );
and ( n73459 , n71204 , n72021 );
nor ( n73460 , n73453 , n72075 );
nor ( n73461 , n73459 , n73460 );
nand ( n73462 , n72003 , n71126 );
nand ( n73463 , n73458 , n73461 , n73462 );
nor ( n73464 , n73452 , n73463 );
and ( n73465 , n73451 , n73464 );
nand ( n73466 , n73450 , n73465 );
buf ( n7324 , n73466 );
buf ( n73468 , 1'b0 );
not ( n73469 , n68842 );
buf ( n7327 , n73469 );
buf ( n7328 , n68638 );
not ( n73472 , n71229 );
or ( n73473 , n73472 , n71990 );
nand ( n73474 , n71237 , n72015 );
and ( n73475 , n71252 , n72018 );
and ( n73476 , n72787 , n69822 );
not ( n73477 , n72787 );
and ( n73478 , n73477 , n72788 );
nor ( n73479 , n73476 , n73478 );
or ( n73480 , n72007 , n73479 );
and ( n73481 , n71260 , n72021 );
nor ( n73482 , n72788 , n72075 );
nor ( n73483 , n73481 , n73482 );
nand ( n73484 , n72003 , n71096 );
nand ( n73485 , n73480 , n73483 , n73484 );
nor ( n73486 , n73475 , n73485 );
and ( n73487 , n73474 , n73486 );
nand ( n73488 , n73473 , n73487 );
buf ( n7346 , n73488 );
buf ( n73490 , 1'b0 );
not ( n73491 , n68842 );
buf ( n73492 , n73491 );
buf ( n7350 , n68638 );
or ( n73494 , n71285 , n71990 );
nand ( n73495 , n71295 , n72015 );
and ( n73496 , n71308 , n72018 );
not ( n73497 , n3514 );
and ( n73498 , n72786 , n73497 );
not ( n73499 , n72786 );
and ( n73500 , n73499 , n3514 );
nor ( n73501 , n73498 , n73500 );
or ( n73502 , n72007 , n73501 );
and ( n73503 , n71316 , n72021 );
nor ( n73504 , n73497 , n72075 );
nor ( n73505 , n73503 , n73504 );
nand ( n73506 , n72003 , n71078 );
nand ( n73507 , n73502 , n73505 , n73506 );
nor ( n73508 , n73496 , n73507 );
and ( n73509 , n73495 , n73508 );
nand ( n73510 , n73494 , n73509 );
buf ( n73511 , n73510 );
buf ( n73512 , 1'b0 );
not ( n73513 , n68842 );
buf ( n73514 , n73513 );
buf ( n73515 , n68638 );
or ( n73516 , n70113 , n71990 );
not ( n73517 , n70561 );
not ( n73518 , n73517 );
not ( n73519 , n71995 );
and ( n73520 , n73518 , n73519 );
nand ( n73521 , n70816 , n72018 );
nand ( n73522 , n72061 , n70902 );
nand ( n73523 , n70841 , n72021 );
nand ( n73524 , n72003 , n70229 );
nor ( n73525 , n70898 , n72075 );
not ( n73526 , n73525 );
and ( n73527 , n73523 , n73524 , n73526 );
nand ( n73528 , n73521 , n73522 , n73527 );
nor ( n73529 , n73520 , n73528 );
nand ( n73530 , n73516 , n73529 );
buf ( n7388 , n73530 );
buf ( n7389 , 1'b0 );
not ( n73533 , n68842 );
buf ( n73534 , n73533 );
buf ( n7392 , n68638 );
not ( n73536 , n71368 );
or ( n73537 , n73536 , n71990 );
not ( n73538 , n72007 );
not ( n73539 , n69607 );
and ( n73540 , n70896 , n73539 );
not ( n73541 , n70896 );
and ( n73542 , n73541 , n69607 );
nor ( n73543 , n73540 , n73542 );
not ( n73544 , n73543 );
and ( n73545 , n73538 , n73544 );
and ( n73546 , n71394 , n72015 );
nor ( n73547 , n73545 , n73546 );
and ( n73548 , n72018 , n71420 );
nand ( n73549 , n71432 , n72021 );
nand ( n73550 , n72003 , n70242 );
nand ( n73551 , n69607 , n70863 );
nand ( n73552 , n73549 , n73550 , n73551 );
nor ( n73553 , n73548 , n73552 );
and ( n73554 , n73547 , n73553 );
nand ( n73555 , n73537 , n73554 );
buf ( n73556 , n73555 );
buf ( n73557 , 1'b0 );
not ( n73558 , n68842 );
buf ( n73559 , n73558 );
buf ( n73560 , n68638 );
not ( n73561 , n71461 );
or ( n73562 , n73561 , n71990 );
not ( n73563 , n72007 );
and ( n73564 , n70894 , n3454 );
not ( n73565 , n70894 );
and ( n73566 , n73565 , n70895 );
nor ( n73567 , n73564 , n73566 );
not ( n73568 , n73567 );
and ( n73569 , n73563 , n73568 );
and ( n73570 , n71479 , n72015 );
nor ( n73571 , n73569 , n73570 );
and ( n73572 , n72018 , n71495 );
nand ( n73573 , n71505 , n72021 );
nand ( n73574 , n72003 , n70331 );
nand ( n73575 , n3454 , n70863 );
nand ( n73576 , n73573 , n73574 , n73575 );
nor ( n73577 , n73572 , n73576 );
and ( n73578 , n73571 , n73577 );
nand ( n73579 , n73562 , n73578 );
buf ( n73580 , n73579 );
buf ( n73581 , 1'b0 );
not ( n73582 , n68842 );
buf ( n73583 , n73582 );
buf ( n73584 , n68638 );
not ( n73585 , n69362 );
not ( n73586 , n69985 );
not ( n73587 , n71451 );
or ( n73588 , n73586 , n73587 );
or ( n73589 , n71451 , n69985 );
nand ( n73590 , n73588 , n73589 );
not ( n73591 , n73590 );
or ( n73592 , n73585 , n73591 );
nand ( n73593 , n69994 , n69363 );
nand ( n73594 , n73592 , n73593 );
not ( n73595 , n73594 );
or ( n73596 , n73595 , n71990 );
not ( n73597 , n72007 );
not ( n73598 , n69571 );
and ( n73599 , n70893 , n73598 );
not ( n73600 , n70893 );
and ( n73601 , n73600 , n69571 );
nor ( n73602 , n73599 , n73601 );
not ( n73603 , n73602 );
and ( n73604 , n73597 , n73603 );
nand ( n73605 , n70358 , n70361 );
not ( n73606 , n73605 );
nor ( n73607 , n71376 , n70324 );
not ( n73608 , n73607 );
not ( n73609 , n70961 );
or ( n73610 , n73608 , n73609 );
or ( n73611 , n71381 , n70324 );
nand ( n73612 , n73611 , n70355 );
not ( n73613 , n73612 );
nand ( n73614 , n73610 , n73613 );
not ( n73615 , n73614 );
or ( n73616 , n73606 , n73615 );
or ( n73617 , n73614 , n73605 );
nand ( n73618 , n73616 , n73617 );
and ( n73619 , n73618 , n72015 );
nor ( n73620 , n73604 , n73619 );
not ( n73621 , n70674 );
nand ( n73622 , n73621 , n70790 );
not ( n73623 , n73622 );
nor ( n73624 , n71401 , n70683 );
not ( n73625 , n73624 );
not ( n73626 , n70988 );
or ( n73627 , n73625 , n73626 );
not ( n73628 , n71406 );
not ( n73629 , n70683 );
and ( n73630 , n73628 , n73629 );
not ( n73631 , n70788 );
nor ( n73632 , n73630 , n73631 );
nand ( n73633 , n73627 , n73632 );
not ( n73634 , n73633 );
or ( n73635 , n73623 , n73634 );
or ( n73636 , n73633 , n73622 );
nand ( n73637 , n73635 , n73636 );
and ( n73638 , n72018 , n73637 );
not ( n73639 , n70300 );
not ( n73640 , n73639 );
and ( n73641 , n70831 , n71565 );
nand ( n73642 , n71007 , n73641 );
not ( n73643 , n73642 );
or ( n73644 , n73640 , n73643 );
or ( n73645 , n73642 , n73639 );
nand ( n73646 , n73644 , n73645 );
nand ( n73647 , n73646 , n72021 );
nand ( n73648 , n72003 , n70300 );
nand ( n73649 , n69571 , n70863 );
nand ( n73650 , n73647 , n73648 , n73649 );
nor ( n73651 , n73638 , n73650 );
and ( n73652 , n73620 , n73651 );
nand ( n73653 , n73596 , n73652 );
buf ( n73654 , n73653 );
buf ( n73655 , 1'b0 );
not ( n73656 , n68842 );
buf ( n73657 , n73656 );
buf ( n73658 , n68638 );
not ( n73659 , n71536 );
or ( n73660 , n73659 , n71990 );
not ( n73661 , n72007 );
not ( n73662 , n3442 );
and ( n73663 , n70892 , n73662 );
not ( n73664 , n70892 );
and ( n73665 , n73664 , n3442 );
nor ( n73666 , n73663 , n73665 );
not ( n73667 , n73666 );
and ( n73668 , n73661 , n73667 );
and ( n73669 , n71549 , n72015 );
nor ( n73670 , n73668 , n73669 );
and ( n73671 , n71562 , n72018 );
nand ( n73672 , n71571 , n72021 );
nand ( n73673 , n72003 , n70312 );
nand ( n73674 , n3442 , n70863 );
nand ( n73675 , n73672 , n73673 , n73674 );
nor ( n73676 , n73671 , n73675 );
and ( n73677 , n73670 , n73676 );
nand ( n73678 , n73660 , n73677 );
buf ( n7536 , n73678 );
buf ( n7537 , 1'b0 );
not ( n73681 , n68842 );
buf ( n73682 , n73681 );
buf ( n7540 , n68638 );
not ( n73684 , n71602 );
or ( n73685 , n73684 , n71990 );
not ( n73686 , n72007 );
and ( n73687 , n70890 , n69516 );
not ( n73688 , n70890 );
and ( n73689 , n73688 , n70891 );
nor ( n73690 , n73687 , n73689 );
not ( n73691 , n73690 );
and ( n73692 , n73686 , n73691 );
and ( n73693 , n71622 , n72015 );
nor ( n73694 , n73692 , n73693 );
and ( n73695 , n72018 , n71642 );
nand ( n73696 , n71651 , n72021 );
nand ( n73697 , n72003 , n70277 );
nand ( n73698 , n69516 , n70863 );
nand ( n73699 , n73696 , n73697 , n73698 );
nor ( n73700 , n73695 , n73699 );
and ( n73701 , n73694 , n73700 );
nand ( n73702 , n73685 , n73701 );
buf ( n73703 , n73702 );
buf ( n73704 , 1'b0 );
not ( n73705 , n68842 );
buf ( n73706 , n73705 );
buf ( n73707 , n68638 );
not ( n73708 , n71676 );
or ( n73709 , n73708 , n71990 );
not ( n73710 , n72007 );
not ( n73711 , n69524 );
and ( n73712 , n70889 , n73711 );
not ( n73713 , n70889 );
and ( n73714 , n73713 , n69524 );
nor ( n73715 , n73712 , n73714 );
not ( n73716 , n73715 );
and ( n73717 , n73710 , n73716 );
and ( n73718 , n71689 , n72015 );
nor ( n73719 , n73717 , n73718 );
and ( n73720 , n72018 , n71703 );
nand ( n73721 , n71711 , n72021 );
nand ( n73722 , n72003 , n70257 );
nand ( n73723 , n69524 , n70863 );
nand ( n73724 , n73721 , n73722 , n73723 );
nor ( n73725 , n73720 , n73724 );
and ( n73726 , n73719 , n73725 );
nand ( n73727 , n73709 , n73726 );
buf ( n73728 , n73727 );
buf ( n73729 , 1'b0 );
not ( n73730 , n68842 );
buf ( n73731 , n73730 );
buf ( n73732 , n68638 );
not ( n73733 , n70057 );
not ( n73734 , n69974 );
or ( n73735 , n73733 , n73734 );
not ( n73736 , n70057 );
nand ( n73737 , n73736 , n69975 );
nand ( n73738 , n73735 , n73737 );
nand ( n73739 , n73738 , n69362 );
or ( n73740 , n73739 , n71990 );
nand ( n73741 , n72390 , n69954 );
not ( n73742 , n70526 );
nor ( n73743 , n73742 , n72006 );
not ( n73744 , n70527 );
not ( n73745 , n69971 );
or ( n73746 , n73744 , n73745 );
not ( n73747 , n70527 );
nand ( n73748 , n73747 , n70523 );
nand ( n73749 , n73746 , n73748 );
not ( n73750 , n73749 );
not ( n73751 , n72015 );
or ( n73752 , n73750 , n73751 );
not ( n73753 , n70728 );
not ( n73754 , n69971 );
or ( n73755 , n73753 , n73754 );
or ( n73756 , n69971 , n70728 );
nand ( n73757 , n73755 , n73756 );
nand ( n73758 , n72018 , n73757 );
nand ( n73759 , n73752 , n73758 );
nor ( n73760 , n73743 , n73759 );
nand ( n73761 , n73740 , n73741 , n73760 );
buf ( n7619 , n73761 );
buf ( n7620 , 1'b0 );
not ( n73764 , n68842 );
buf ( n73765 , n73764 );
buf ( n7623 , n68638 );
or ( n73767 , n71985 , n70214 );
and ( n73768 , n70577 , n70996 );
not ( n73769 , n70844 );
not ( n73770 , n73769 );
nand ( n73771 , n71012 , n73770 );
not ( n73772 , n70879 );
not ( n73773 , n72012 );
and ( n73774 , n73772 , n73773 );
and ( n73775 , n70853 , n70267 );
nor ( n73776 , n73774 , n73775 );
nand ( n73777 , n70874 , n69537 );
nand ( n73778 , n73771 , n73776 , n73777 );
nor ( n73779 , n73768 , n73778 );
nand ( n73780 , n70969 , n70572 );
and ( n73781 , n73779 , n73780 );
nand ( n73782 , n73767 , n73781 );
buf ( n73783 , n73782 );
buf ( n7641 , 1'b0 );
not ( n73785 , n68842 );
buf ( n73786 , n73785 );
buf ( n73787 , n68638 );
or ( n73788 , n72045 , n70214 );
nand ( n73789 , n72052 , n70577 );
nand ( n73790 , n72059 , n70572 );
not ( n73791 , n72073 );
not ( n73792 , n70844 );
or ( n73793 , n73791 , n73792 );
and ( n73794 , n70874 , n3405 );
and ( n73795 , n70880 , n72066 );
nor ( n73796 , n73794 , n73795 );
nand ( n73797 , n73793 , n73796 );
not ( n73798 , n70382 );
nor ( n73799 , n70852 , n73798 );
nor ( n73800 , n73797 , n73799 );
and ( n73801 , n73789 , n73790 , n73800 );
nand ( n73802 , n73788 , n73801 );
buf ( n73803 , n73802 );
buf ( n73804 , 1'b0 );
not ( n73805 , n68842 );
buf ( n73806 , n73805 );
buf ( n73807 , n68638 );
or ( n73808 , n72098 , n70214 );
nand ( n73809 , n72116 , n70572 );
nand ( n73810 , n72134 , n70577 );
and ( n73811 , n70853 , n70392 );
and ( n73812 , n70880 , n72139 );
nor ( n73813 , n73811 , n73812 );
nand ( n73814 , n70844 , n72154 );
nand ( n73815 , n70874 , n3320 );
and ( n73816 , n73813 , n73814 , n73815 );
and ( n73817 , n73809 , n73810 , n73816 );
nand ( n73818 , n73808 , n73817 );
buf ( n7676 , n73818 );
buf ( n7677 , 1'b0 );
not ( n73821 , n68842 );
buf ( n73822 , n73821 );
buf ( n73823 , n68638 );
or ( n73824 , n72173 , n70214 );
nand ( n73825 , n72182 , n70577 );
nand ( n73826 , n72195 , n70572 );
and ( n73827 , n70853 , n70481 );
and ( n73828 , n70880 , n72201 );
nor ( n73829 , n73827 , n73828 );
nand ( n73830 , n70844 , n72211 );
nand ( n73831 , n70874 , n3276 );
and ( n73832 , n73829 , n73830 , n73831 );
and ( n73833 , n73825 , n73826 , n73832 );
nand ( n73834 , n73824 , n73833 );
buf ( n73835 , n73834 );
buf ( n7693 , 1'b0 );
not ( n73837 , n68842 );
buf ( n73838 , n73837 );
buf ( n73839 , n68638 );
or ( n73840 , n72234 , n70214 );
nand ( n73841 , n72246 , n70572 );
nand ( n73842 , n72258 , n70577 );
and ( n73843 , n70853 , n70436 );
and ( n73844 , n70880 , n72263 );
nor ( n73845 , n73843 , n73844 );
nand ( n73846 , n70844 , n72273 );
not ( n73847 , n70874 );
not ( n73848 , n73847 );
nand ( n73849 , n73848 , n3350 );
and ( n73850 , n73845 , n73846 , n73849 );
and ( n73851 , n73841 , n73842 , n73850 );
nand ( n73852 , n73840 , n73851 );
buf ( n73853 , n73852 );
buf ( n73854 , 1'b0 );
not ( n73855 , n68842 );
buf ( n73856 , n73855 );
buf ( n73857 , n68638 );
or ( n73858 , n72294 , n70214 );
and ( n73859 , n72304 , n70577 );
not ( n73860 , n3346 );
nor ( n73861 , n73847 , n73860 );
nor ( n73862 , n73859 , n73861 );
nand ( n73863 , n72297 , n70572 );
not ( n73864 , n72306 );
not ( n73865 , n70853 );
or ( n73866 , n73864 , n73865 );
not ( n73867 , n70880 );
or ( n73868 , n73867 , n72323 );
nand ( n73869 , n73866 , n73868 );
not ( n73870 , n70844 );
not ( n73871 , n72311 );
nor ( n73872 , n73870 , n73871 );
nor ( n73873 , n73869 , n73872 );
and ( n73874 , n73862 , n73863 , n73873 );
nand ( n73875 , n73858 , n73874 );
buf ( n73876 , n73875 );
buf ( n73877 , 1'b0 );
not ( n73878 , n68842 );
buf ( n73879 , n73878 );
buf ( n73880 , n68638 );
or ( n73881 , n72344 , n70214 );
nand ( n73882 , n72349 , n70572 );
nand ( n73883 , n72360 , n70577 );
nand ( n73884 , n73770 , n72369 );
and ( n73885 , n70853 , n70424 );
and ( n73886 , n70880 , n72321 );
nor ( n73887 , n73885 , n73886 );
nand ( n73888 , n70874 , n69441 );
and ( n73889 , n73884 , n73887 , n73888 );
and ( n73890 , n73882 , n73883 , n73889 );
nand ( n73891 , n73881 , n73890 );
buf ( n73892 , n73891 );
buf ( n7750 , 1'b0 );
not ( n73894 , n68842 );
buf ( n7752 , n73894 );
buf ( n73896 , n68638 );
and ( n73897 , n70874 , n69944 );
not ( n73898 , n70874 );
not ( n73899 , n69951 );
nand ( n73900 , n72458 , n72467 );
not ( n73901 , n73900 );
not ( n73902 , n71754 );
nor ( n73903 , n72453 , n69748 );
nand ( n73904 , n73902 , n72451 , n73903 );
not ( n73905 , n69912 );
xor ( n73906 , n73904 , n73905 );
nand ( n73907 , n73901 , n73906 );
not ( n73908 , n73907 );
or ( n73909 , n73899 , n73908 );
or ( n73910 , n69951 , n73907 );
nand ( n73911 , n73909 , n73910 );
or ( n73912 , n71276 , n4012 );
nand ( n73913 , n73912 , n70226 );
and ( n73914 , n70200 , n73913 );
nand ( n73915 , n73911 , n73914 );
and ( n73916 , n70226 , n68640 );
not ( n73917 , n73916 );
and ( n73918 , n70226 , n2498 );
not ( n73919 , n73918 );
and ( n73920 , n70226 , n2499 );
nor ( n73921 , n72630 , n73920 );
nand ( n73922 , n73919 , n72816 , n73921 , n72821 );
nor ( n73923 , n70836 , n73922 );
not ( n73924 , n73923 );
or ( n73925 , n73917 , n73924 );
or ( n73926 , n73923 , n73916 );
nand ( n73927 , n73925 , n73926 );
and ( n73928 , n73927 , n70999 );
not ( n73929 , n73916 );
nor ( n73930 , n73929 , n70850 );
nor ( n73931 , n73928 , n73930 );
nand ( n73932 , n73915 , n73931 );
and ( n73933 , n73898 , n73932 );
or ( n73934 , n73897 , n73933 );
buf ( n73935 , n73934 );
buf ( n73936 , 1'b0 );
not ( n73937 , n68842 );
buf ( n7795 , n73937 );
buf ( n73939 , n68638 );
and ( n73940 , n70874 , n69906 );
not ( n73941 , n70874 );
and ( n73942 , n70851 , n73918 );
not ( n73943 , n73918 );
nand ( n73944 , n72816 , n72821 , n73921 );
nor ( n73945 , n70836 , n73944 );
not ( n73946 , n73945 );
or ( n73947 , n73943 , n73946 );
or ( n73948 , n73945 , n73918 );
nand ( n73949 , n73947 , n73948 );
and ( n73950 , n73949 , n70999 );
nor ( n73951 , n73942 , n73950 );
nand ( n73952 , n73915 , n73951 );
and ( n73953 , n73941 , n73952 );
or ( n73954 , n73940 , n73953 );
buf ( n73955 , n73954 );
buf ( n73956 , 1'b0 );
not ( n73957 , n68842 );
buf ( n73958 , n73957 );
buf ( n73959 , n68638 );
or ( n73960 , n72388 , n70214 );
nand ( n73961 , n72409 , n70572 );
nand ( n73962 , n70577 , n72422 );
nand ( n73963 , n70880 , n70058 );
nand ( n73964 , n73961 , n73962 , n73963 );
or ( n73965 , n73769 , n72398 );
not ( n73966 , n70062 );
or ( n73967 , n73847 , n73966 );
or ( n73968 , n70852 , n72414 );
nand ( n73969 , n73965 , n73967 , n73968 );
nor ( n73970 , n73964 , n73969 );
nand ( n73971 , n73960 , n73970 );
buf ( n73972 , n73971 );
buf ( n7830 , 1'b0 );
not ( n73974 , n68842 );
buf ( n7832 , n73974 );
buf ( n7833 , n68638 );
not ( n73977 , n73906 );
not ( n73978 , n73977 );
not ( n73979 , n73901 );
or ( n73980 , n73978 , n73979 );
or ( n73981 , n73977 , n73901 );
nand ( n73982 , n73980 , n73981 );
and ( n73983 , n73982 , n73913 );
and ( n73984 , n72456 , n69363 );
nor ( n73985 , n73983 , n73984 );
or ( n73986 , n73985 , n70214 );
nor ( n73987 , n72637 , n72630 );
not ( n73988 , n73987 );
not ( n73989 , n73920 );
not ( n73990 , n69747 );
or ( n73991 , n73989 , n73990 );
or ( n73992 , n69747 , n73920 );
nand ( n73993 , n73991 , n73992 );
not ( n73994 , n73993 );
or ( n73995 , n73988 , n73994 );
or ( n73996 , n73987 , n73993 );
nand ( n73997 , n73995 , n73996 );
not ( n73998 , n73997 );
nor ( n73999 , n72574 , n72642 );
not ( n74000 , n73999 );
nor ( n74001 , n74000 , n72526 );
not ( n74002 , n74001 );
not ( n74003 , n70557 );
or ( n74004 , n74002 , n74003 );
not ( n74005 , n73999 );
not ( n74006 , n72608 );
or ( n74007 , n74005 , n74006 );
not ( n74008 , n72643 );
not ( n74009 , n72624 );
or ( n74010 , n74008 , n74009 );
nand ( n74011 , n74010 , n72644 );
not ( n74012 , n74011 );
nand ( n74013 , n74007 , n74012 );
not ( n74014 , n74013 );
nand ( n74015 , n74004 , n74014 );
not ( n74016 , n74015 );
or ( n74017 , n73998 , n74016 );
or ( n74018 , n74015 , n73997 );
nand ( n74019 , n74017 , n74018 );
nand ( n74020 , n74019 , n70572 );
xor ( n74021 , n73920 , n69747 );
not ( n74022 , n74021 );
and ( n74023 , n72630 , n69733 );
not ( n74024 , n74023 );
or ( n74025 , n74022 , n74024 );
or ( n74026 , n74023 , n74021 );
nand ( n74027 , n74025 , n74026 );
not ( n74028 , n74027 );
nand ( n74029 , n72678 , n72775 );
nor ( n74030 , n74029 , n72728 );
not ( n74031 , n74030 );
not ( n74032 , n70813 );
or ( n74033 , n74031 , n74032 );
not ( n74034 , n72753 );
not ( n74035 , n74029 );
and ( n74036 , n74034 , n74035 );
not ( n74037 , n72775 );
not ( n74038 , n72770 );
or ( n74039 , n74037 , n74038 );
nand ( n74040 , n74039 , n72776 );
nor ( n74041 , n74036 , n74040 );
nand ( n74042 , n74033 , n74041 );
not ( n74043 , n74042 );
or ( n74044 , n74028 , n74043 );
or ( n74045 , n74042 , n74027 );
nand ( n74046 , n74044 , n74045 );
and ( n74047 , n74046 , n70577 );
nand ( n74048 , n72801 , n70880 , n69725 );
not ( n74049 , n73920 );
not ( n74050 , n72630 );
nand ( n74051 , n74050 , n72816 , n72821 );
nor ( n74052 , n70836 , n74051 );
not ( n74053 , n74052 );
or ( n74054 , n74049 , n74053 );
or ( n74055 , n74052 , n73920 );
nand ( n74056 , n74054 , n74055 );
nand ( n74057 , n74056 , n73770 );
nand ( n74058 , n70853 , n73920 );
nand ( n74059 , n70874 , n69745 );
nand ( n74060 , n74048 , n74057 , n74058 , n74059 );
nor ( n74061 , n74047 , n74060 );
nand ( n74062 , n73986 , n74020 , n74061 );
buf ( n7920 , n74062 );
buf ( n7921 , 1'b0 );
not ( n74065 , n68842 );
buf ( n74066 , n74065 );
buf ( n74067 , n68638 );
or ( n74068 , n72474 , n70214 );
nand ( n74069 , n72650 , n70572 );
and ( n74070 , n72782 , n70577 );
nand ( n74071 , n72805 , n70880 );
nand ( n74072 , n72827 , n70844 );
nand ( n74073 , n70853 , n72630 );
nand ( n74074 , n70874 , n69714 );
nand ( n74075 , n74071 , n74072 , n74073 , n74074 );
nor ( n74076 , n74070 , n74075 );
and ( n74077 , n74069 , n74076 );
nand ( n74078 , n74068 , n74077 );
buf ( n74079 , n74078 );
buf ( n7937 , 1'b0 );
not ( n74081 , n68842 );
buf ( n74082 , n74081 );
buf ( n74083 , n68638 );
or ( n74084 , n72849 , n70214 );
nand ( n74085 , n72870 , n70572 );
and ( n74086 , n72893 , n70577 );
not ( n74087 , n72898 );
nand ( n74088 , n74087 , n70880 );
nand ( n74089 , n72910 , n73770 );
nand ( n74090 , n70853 , n72819 );
nand ( n74091 , n70874 , n69692 );
nand ( n74092 , n74088 , n74089 , n74090 , n74091 );
nor ( n74093 , n74086 , n74092 );
and ( n74094 , n74085 , n74093 );
nand ( n74095 , n74084 , n74094 );
buf ( n7953 , n74095 );
buf ( n7954 , 1'b0 );
not ( n74098 , n68842 );
buf ( n74099 , n74098 );
buf ( n74100 , n68638 );
or ( n74101 , n72937 , n70214 );
nand ( n74102 , n72956 , n70572 );
and ( n74103 , n72971 , n70577 );
nor ( n74104 , n72976 , n73867 );
not ( n74105 , n72538 );
nor ( n74106 , n74105 , n70852 );
nor ( n74107 , n74104 , n74106 );
nand ( n74108 , n72986 , n70844 );
nand ( n74109 , n70874 , n69674 );
nand ( n74110 , n74107 , n74108 , n74109 );
nor ( n74111 , n74103 , n74110 );
and ( n74112 , n74102 , n74111 );
nand ( n74113 , n74101 , n74112 );
buf ( n74114 , n74113 );
buf ( n7972 , 1'b0 );
not ( n74116 , n68842 );
buf ( n7974 , n74116 );
buf ( n74118 , n68638 );
or ( n74119 , n73011 , n70214 );
nand ( n74120 , n73026 , n70572 );
and ( n74121 , n73044 , n70577 );
nand ( n74122 , n73060 , n73770 );
and ( n74123 , n70853 , n72548 );
nor ( n74124 , n73049 , n73867 );
nor ( n74125 , n74123 , n74124 );
nand ( n74126 , n70874 , n69835 );
nand ( n74127 , n74122 , n74125 , n74126 );
nor ( n74128 , n74121 , n74127 );
and ( n74129 , n74120 , n74128 );
nand ( n74130 , n74119 , n74129 );
buf ( n74131 , n74130 );
buf ( n7989 , 1'b0 );
not ( n74133 , n68842 );
buf ( n74134 , n74133 );
buf ( n74135 , n68638 );
or ( n74136 , n73083 , n70214 );
nand ( n74137 , n73096 , n70572 );
and ( n74138 , n73108 , n70577 );
nand ( n74139 , n73121 , n73770 );
not ( n74140 , n73113 );
not ( n74141 , n70879 );
and ( n74142 , n74140 , n74141 );
and ( n74143 , n70853 , n72561 );
nor ( n74144 , n74142 , n74143 );
nand ( n74145 , n70874 , n69920 );
nand ( n74146 , n74139 , n74144 , n74145 );
nor ( n74147 , n74138 , n74146 );
and ( n74148 , n74137 , n74147 );
nand ( n74149 , n74136 , n74148 );
buf ( n74150 , n74149 );
buf ( n74151 , 1'b0 );
not ( n74152 , n68842 );
buf ( n74153 , n74152 );
buf ( n8011 , n68638 );
or ( n74155 , n73147 , n70214 );
nand ( n74156 , n73165 , n70572 );
and ( n74157 , n73193 , n70577 );
nand ( n74158 , n73206 , n73770 );
not ( n74159 , n73198 );
not ( n74160 , n70879 );
and ( n74161 , n74159 , n74160 );
and ( n74162 , n70853 , n72514 );
nor ( n74163 , n74161 , n74162 );
nand ( n74164 , n70874 , n69753 );
nand ( n74165 , n74158 , n74163 , n74164 );
nor ( n74166 , n74157 , n74165 );
and ( n74167 , n74156 , n74166 );
nand ( n74168 , n74155 , n74167 );
buf ( n74169 , n74168 );
buf ( n8027 , 1'b0 );
not ( n74171 , n68842 );
buf ( n74172 , n74171 );
buf ( n74173 , n68638 );
or ( n74174 , n73228 , n70214 );
nand ( n74175 , n73243 , n70572 );
and ( n74176 , n73257 , n70577 );
nand ( n74177 , n73270 , n73770 );
not ( n74178 , n73262 );
not ( n74179 , n70879 );
and ( n74180 , n74178 , n74179 );
and ( n74181 , n70853 , n72503 );
nor ( n74182 , n74180 , n74181 );
nand ( n74183 , n70874 , n69787 );
nand ( n74184 , n74177 , n74182 , n74183 );
nor ( n74185 , n74176 , n74184 );
and ( n74186 , n74175 , n74185 );
nand ( n74187 , n74174 , n74186 );
buf ( n74188 , n74187 );
buf ( n8046 , 1'b0 );
not ( n74190 , n68842 );
buf ( n8048 , n74190 );
buf ( n74192 , n68638 );
or ( n74193 , n73293 , n70214 );
nand ( n74194 , n73308 , n70572 );
and ( n74195 , n73327 , n70577 );
nand ( n74196 , n73341 , n73770 );
not ( n74197 , n70879 );
not ( n74198 , n73332 );
and ( n74199 , n74197 , n74198 );
and ( n74200 , n70853 , n72479 );
nor ( n74201 , n74199 , n74200 );
nand ( n74202 , n70874 , n69880 );
nand ( n74203 , n74196 , n74201 , n74202 );
nor ( n74204 , n74195 , n74203 );
and ( n74205 , n74194 , n74204 );
nand ( n74206 , n74193 , n74205 );
buf ( n8064 , n74206 );
buf ( n74208 , 1'b0 );
not ( n74209 , n68842 );
buf ( n8067 , n74209 );
buf ( n8068 , n68638 );
or ( n74212 , n73365 , n70214 );
nand ( n74213 , n73373 , n70572 );
and ( n74214 , n70577 , n73385 );
nand ( n74215 , n73398 , n73770 );
not ( n74216 , n70879 );
not ( n74217 , n73390 );
and ( n74218 , n74216 , n74217 );
and ( n74219 , n70853 , n72489 );
nor ( n74220 , n74218 , n74219 );
nand ( n74221 , n70874 , n69866 );
nand ( n74222 , n74215 , n74220 , n74221 );
nor ( n74223 , n74214 , n74222 );
and ( n74224 , n74213 , n74223 );
nand ( n74225 , n74212 , n74224 );
buf ( n74226 , n74225 );
buf ( n74227 , 1'b0 );
not ( n74228 , n68842 );
buf ( n8086 , n74228 );
buf ( n74230 , n68638 );
or ( n74231 , n73420 , n70214 );
not ( n74232 , n73439 );
or ( n74233 , n73769 , n74232 );
not ( n74234 , n70055 );
or ( n74235 , n73847 , n74234 );
not ( n74236 , n70507 );
or ( n74237 , n70852 , n74236 );
nand ( n74238 , n74233 , n74235 , n74237 );
not ( n74239 , n73430 );
not ( n74240 , n70572 );
or ( n74241 , n74239 , n74240 );
nand ( n74242 , n70577 , n73432 );
nand ( n74243 , n70880 , n70045 );
nand ( n74244 , n74241 , n74242 , n74243 );
nor ( n74245 , n74238 , n74244 );
nand ( n74246 , n74231 , n74245 );
buf ( n74247 , n74246 );
buf ( n74248 , 1'b0 );
not ( n74249 , n68842 );
buf ( n74250 , n74249 );
buf ( n74251 , n68638 );
or ( n74252 , n73449 , n70214 );
nand ( n74253 , n71138 , n70572 );
and ( n74254 , n71192 , n70577 );
nand ( n74255 , n71204 , n73770 );
not ( n74256 , n70879 );
not ( n74257 , n73457 );
and ( n74258 , n74256 , n74257 );
and ( n74259 , n70853 , n71126 );
nor ( n74260 , n74258 , n74259 );
nand ( n74261 , n70874 , n69802 );
nand ( n74262 , n74255 , n74260 , n74261 );
nor ( n74263 , n74254 , n74262 );
and ( n74264 , n74253 , n74263 );
nand ( n74265 , n74252 , n74264 );
buf ( n74266 , n74265 );
buf ( n74267 , 1'b0 );
not ( n74268 , n68842 );
buf ( n8126 , n74268 );
buf ( n8127 , n68638 );
or ( n74271 , n73472 , n70214 );
nand ( n74272 , n71237 , n70572 );
and ( n74273 , n71252 , n70577 );
nand ( n74274 , n71260 , n70844 );
not ( n74275 , n70879 );
not ( n74276 , n73479 );
and ( n74277 , n74275 , n74276 );
and ( n74278 , n70853 , n71096 );
nor ( n74279 , n74277 , n74278 );
nand ( n74280 , n70874 , n69810 );
nand ( n74281 , n74274 , n74279 , n74280 );
nor ( n74282 , n74273 , n74281 );
and ( n74283 , n74272 , n74282 );
nand ( n74284 , n74271 , n74283 );
buf ( n8142 , n74284 );
buf ( n8143 , 1'b0 );
not ( n74287 , n68842 );
buf ( n74288 , n74287 );
buf ( n74289 , n68638 );
or ( n74290 , n71285 , n70214 );
nand ( n74291 , n71295 , n70572 );
and ( n74292 , n71308 , n70577 );
nand ( n74293 , n71316 , n70844 );
not ( n74294 , n70879 );
not ( n74295 , n73501 );
and ( n74296 , n74294 , n74295 );
and ( n74297 , n70853 , n71078 );
nor ( n74298 , n74296 , n74297 );
nand ( n74299 , n73848 , n69655 );
nand ( n74300 , n74293 , n74298 , n74299 );
nor ( n74301 , n74292 , n74300 );
nand ( n74302 , n74290 , n74291 , n74301 );
buf ( n8160 , n74302 );
buf ( n74304 , 1'b0 );
not ( n74305 , n68842 );
buf ( n74306 , n74305 );
buf ( n8164 , n68638 );
or ( n74308 , n73536 , n70214 );
and ( n74309 , n70577 , n71420 );
nand ( n74310 , n71432 , n70844 );
not ( n74311 , n73867 );
not ( n74312 , n73543 );
and ( n74313 , n74311 , n74312 );
and ( n74314 , n70853 , n70242 );
nor ( n74315 , n74313 , n74314 );
nand ( n74316 , n73848 , n3466 );
nand ( n74317 , n74310 , n74315 , n74316 );
nor ( n74318 , n74309 , n74317 );
nand ( n74319 , n71394 , n70572 );
and ( n74320 , n74318 , n74319 );
nand ( n74321 , n74308 , n74320 );
buf ( n74322 , n74321 );
buf ( n74323 , 1'b0 );
not ( n74324 , n68842 );
buf ( n74325 , n74324 );
buf ( n74326 , n68638 );
or ( n74327 , n73561 , n70214 );
and ( n74328 , n70577 , n71495 );
nand ( n74329 , n71505 , n73770 );
not ( n74330 , n70879 );
not ( n74331 , n73567 );
and ( n74332 , n74330 , n74331 );
and ( n74333 , n70853 , n70331 );
nor ( n74334 , n74332 , n74333 );
nand ( n74335 , n73848 , n3450 );
nand ( n74336 , n74329 , n74334 , n74335 );
nor ( n74337 , n74328 , n74336 );
nand ( n74338 , n71479 , n70572 );
and ( n74339 , n74337 , n74338 );
nand ( n74340 , n74327 , n74339 );
buf ( n74341 , n74340 );
buf ( n74342 , 1'b0 );
not ( n74343 , n68842 );
buf ( n8201 , n74343 );
buf ( n8202 , n68638 );
or ( n74346 , n73595 , n70214 );
and ( n74347 , n70577 , n73637 );
nand ( n74348 , n73646 , n70844 );
not ( n74349 , n70879 );
not ( n74350 , n73602 );
and ( n74351 , n74349 , n74350 );
and ( n74352 , n70853 , n70300 );
nor ( n74353 , n74351 , n74352 );
nand ( n74354 , n73848 , n69562 );
nand ( n74355 , n74348 , n74353 , n74354 );
nor ( n74356 , n74347 , n74355 );
nand ( n74357 , n73618 , n70572 );
and ( n74358 , n74356 , n74357 );
nand ( n74359 , n74346 , n74358 );
buf ( n8217 , n74359 );
buf ( n8218 , 1'b0 );
not ( n74362 , n68842 );
buf ( n74363 , n74362 );
buf ( n74364 , n68638 );
or ( n74365 , n73659 , n70214 );
and ( n74366 , n70577 , n71562 );
nand ( n74367 , n71571 , n73770 );
not ( n74368 , n70879 );
not ( n74369 , n73666 );
and ( n74370 , n74368 , n74369 );
and ( n74371 , n70853 , n70312 );
nor ( n74372 , n74370 , n74371 );
nand ( n74373 , n73848 , n69581 );
nand ( n74374 , n74367 , n74372 , n74373 );
nor ( n74375 , n74366 , n74374 );
nand ( n74376 , n71549 , n70572 );
and ( n74377 , n74375 , n74376 );
nand ( n74378 , n74365 , n74377 );
buf ( n74379 , n74378 );
buf ( n74380 , 1'b0 );
not ( n74381 , n68842 );
buf ( n8239 , n74381 );
buf ( n74383 , n68638 );
or ( n74384 , n73684 , n70214 );
and ( n74385 , n70577 , n71642 );
nand ( n74386 , n71651 , n70844 );
not ( n74387 , n70879 );
not ( n74388 , n73690 );
and ( n74389 , n74387 , n74388 );
and ( n74390 , n70853 , n70277 );
nor ( n74391 , n74389 , n74390 );
nand ( n74392 , n73848 , n69511 );
nand ( n74393 , n74386 , n74391 , n74392 );
nor ( n74394 , n74385 , n74393 );
nand ( n74395 , n71622 , n70572 );
and ( n74396 , n74394 , n74395 );
nand ( n74397 , n74384 , n74396 );
buf ( n74398 , n74397 );
buf ( n74399 , 1'b0 );
not ( n74400 , n68842 );
buf ( n74401 , n74400 );
buf ( n74402 , n68638 );
or ( n74403 , n73708 , n70214 );
and ( n74404 , n70577 , n71703 );
nand ( n74405 , n71711 , n70844 );
not ( n74406 , n73867 );
not ( n74407 , n73715 );
and ( n74408 , n74406 , n74407 );
and ( n74409 , n70853 , n70257 );
nor ( n74410 , n74408 , n74409 );
nand ( n74411 , n73848 , n69526 );
nand ( n74412 , n74405 , n74410 , n74411 );
nor ( n74413 , n74404 , n74412 );
nand ( n74414 , n71689 , n70572 );
and ( n74415 , n74413 , n74414 );
nand ( n74416 , n74403 , n74415 );
buf ( n8274 , n74416 );
buf ( n8275 , 1'b0 );
not ( n74419 , n68842 );
buf ( n8277 , n74419 );
buf ( n8278 , n68638 );
or ( n74422 , n73739 , n70214 );
not ( n74423 , n3815 );
not ( n74424 , n70874 );
or ( n74425 , n74423 , n74424 );
or ( n74426 , n70844 , n70853 );
nand ( n74427 , n74426 , n70526 );
nand ( n74428 , n74425 , n74427 );
nand ( n74429 , n70572 , n73749 );
nand ( n74430 , n70577 , n73757 );
nand ( n74431 , n70880 , n69954 );
nand ( n74432 , n74429 , n74430 , n74431 );
nor ( n74433 , n74428 , n74432 );
nand ( n74434 , n74422 , n74433 );
buf ( n8292 , n74434 );
buf ( n74436 , 1'b0 );
not ( n74437 , n68842 );
buf ( n74438 , n74437 );
buf ( n8296 , n68638 );
and ( n74440 , n72044 , n70200 );
nand ( n74441 , n72059 , n70933 );
nand ( n74442 , n72052 , n70575 );
not ( n74443 , n73798 );
not ( n74444 , n70850 );
and ( n74445 , n74443 , n74444 );
and ( n74446 , n72073 , n70999 );
nor ( n74447 , n74445 , n74446 );
nand ( n74448 , n74441 , n74442 , n74447 );
nor ( n74449 , n74440 , n74448 );
or ( n74450 , n74449 , n71020 );
nand ( n74451 , n71020 , n69550 );
nand ( n74452 , n74450 , n74451 );
buf ( n74453 , n74452 );
buf ( n74454 , 1'b0 );
not ( n74455 , n68842 );
buf ( n8313 , n74455 );
buf ( n74457 , n68638 );
not ( n74458 , n72098 );
and ( n74459 , n74458 , n70927 );
not ( n74460 , n70933 );
not ( n74461 , n72116 );
or ( n74462 , n74460 , n74461 );
and ( n74463 , n72134 , n70575 );
not ( n74464 , n70851 );
not ( n74465 , n70392 );
or ( n74466 , n74464 , n74465 );
nand ( n74467 , n72154 , n70999 );
nand ( n74468 , n74466 , n74467 );
nor ( n74469 , n74463 , n74468 );
nand ( n74470 , n74462 , n74469 );
nor ( n74471 , n74459 , n74470 );
or ( n74472 , n74471 , n71020 );
not ( n74473 , n71020 );
not ( n74474 , n74473 );
nand ( n74475 , n74474 , n3316 );
nand ( n74476 , n74472 , n74475 );
buf ( n74477 , n74476 );
buf ( n74478 , 1'b0 );
not ( n74479 , n68842 );
buf ( n74480 , n74479 );
buf ( n74481 , n68638 );
not ( n74482 , n72173 );
and ( n74483 , n74482 , n70927 );
nand ( n74484 , n72195 , n70935 );
nand ( n74485 , n72182 , n70575 );
and ( n74486 , n70481 , n70851 );
and ( n74487 , n72211 , n70999 );
nor ( n74488 , n74486 , n74487 );
nand ( n74489 , n74484 , n74485 , n74488 );
nor ( n74490 , n74483 , n74489 );
or ( n74491 , n74490 , n71020 );
not ( n74492 , n71347 );
nand ( n74493 , n74492 , n3282 );
nand ( n74494 , n74491 , n74493 );
buf ( n8352 , n74494 );
buf ( n74496 , 1'b0 );
not ( n74497 , n68842 );
buf ( n8355 , n74497 );
buf ( n74499 , n68638 );
not ( n74500 , n72234 );
and ( n74501 , n74500 , n70927 );
not ( n74502 , n70933 );
not ( n74503 , n72246 );
or ( n74504 , n74502 , n74503 );
and ( n74505 , n72258 , n70575 );
not ( n74506 , n70851 );
not ( n74507 , n70436 );
or ( n74508 , n74506 , n74507 );
nand ( n74509 , n72273 , n70999 );
nand ( n74510 , n74508 , n74509 );
nor ( n74511 , n74505 , n74510 );
nand ( n74512 , n74504 , n74511 );
nor ( n74513 , n74501 , n74512 );
or ( n74514 , n74513 , n71020 );
nand ( n74515 , n74474 , n69496 );
nand ( n74516 , n74514 , n74515 );
buf ( n74517 , n74516 );
buf ( n74518 , 1'b0 );
not ( n74519 , n68842 );
buf ( n74520 , n74519 );
buf ( n74521 , n68638 );
and ( n74522 , n72293 , n70927 );
not ( n74523 , n70933 );
not ( n74524 , n72297 );
or ( n74525 , n74523 , n74524 );
and ( n74526 , n72304 , n70575 );
not ( n74527 , n72306 );
not ( n74528 , n70851 );
or ( n74529 , n74527 , n74528 );
not ( n74530 , n70999 );
or ( n74531 , n73871 , n74530 );
nand ( n74532 , n74529 , n74531 );
nor ( n74533 , n74526 , n74532 );
nand ( n74534 , n74525 , n74533 );
nor ( n74535 , n74522 , n74534 );
or ( n74536 , n74535 , n71348 );
nand ( n74537 , n74492 , n3342 );
nand ( n74538 , n74536 , n74537 );
buf ( n74539 , n74538 );
buf ( n8397 , 1'b0 );
not ( n74541 , n68842 );
buf ( n74542 , n74541 );
buf ( n74543 , n68638 );
not ( n74544 , n74473 );
or ( n74545 , n72344 , n70199 );
and ( n74546 , n72360 , n70575 );
not ( n74547 , n70424 );
not ( n74548 , n70851 );
or ( n74549 , n74547 , n74548 );
nand ( n74550 , n72369 , n70999 );
nand ( n74551 , n74549 , n74550 );
nor ( n74552 , n74546 , n74551 );
nand ( n74553 , n72349 , n70933 );
and ( n74554 , n74552 , n74553 );
nand ( n74555 , n74545 , n74554 );
not ( n74556 , n74555 );
or ( n74557 , n74544 , n74556 );
nand ( n74558 , n71348 , n3301 );
nand ( n74559 , n74557 , n74558 );
buf ( n8417 , n74559 );
buf ( n8418 , 1'b0 );
not ( n74562 , n68842 );
buf ( n74563 , n74562 );
buf ( n74564 , n68638 );
and ( n74565 , n71020 , n69940 );
not ( n74566 , n71020 );
and ( n74567 , n74566 , n73932 );
or ( n74568 , n74565 , n74567 );
buf ( n8426 , n74568 );
buf ( n74570 , 1'b0 );
not ( n74571 , n68842 );
buf ( n8429 , n74571 );
buf ( n74573 , n68638 );
not ( n74574 , n73952 );
or ( n74575 , n74574 , n74474 );
or ( n74576 , n71347 , n69902 );
nand ( n74577 , n74575 , n74576 );
buf ( n74578 , n74577 );
buf ( n74579 , 1'b0 );
not ( n74580 , n68842 );
buf ( n8438 , n74580 );
buf ( n8439 , n68638 );
not ( n74583 , n72388 );
and ( n74584 , n74583 , n70200 );
not ( n74585 , n70933 );
not ( n74586 , n72409 );
or ( n74587 , n74585 , n74586 );
and ( n74588 , n72422 , n70575 );
or ( n74589 , n72414 , n70850 );
or ( n74590 , n72398 , n74530 );
nand ( n74591 , n74589 , n74590 );
nor ( n74592 , n74588 , n74591 );
nand ( n74593 , n74587 , n74592 );
nor ( n74594 , n74584 , n74593 );
or ( n74595 , n74594 , n71020 );
nand ( n74596 , n71348 , n70073 );
nand ( n74597 , n74595 , n74596 );
buf ( n8455 , n74597 );
buf ( n8456 , 1'b0 );
not ( n74600 , n68842 );
buf ( n74601 , n74600 );
buf ( n74602 , n68638 );
not ( n74603 , n73985 );
and ( n74604 , n74603 , n70200 );
not ( n74605 , n70933 );
not ( n74606 , n74019 );
or ( n74607 , n74605 , n74606 );
and ( n74608 , n74046 , n70575 );
not ( n74609 , n70999 );
not ( n74610 , n74056 );
or ( n74611 , n74609 , n74610 );
nand ( n74612 , n70851 , n73920 );
nand ( n74613 , n74611 , n74612 );
nor ( n74614 , n74608 , n74613 );
nand ( n74615 , n74607 , n74614 );
nor ( n74616 , n74604 , n74615 );
or ( n74617 , n74616 , n74492 );
nand ( n74618 , n71348 , n69741 );
nand ( n74619 , n74617 , n74618 );
buf ( n74620 , n74619 );
buf ( n74621 , 1'b0 );
not ( n74622 , n68842 );
buf ( n74623 , n74622 );
buf ( n74624 , n68638 );
not ( n74625 , n72474 );
not ( n74626 , n70927 );
not ( n74627 , n74626 );
and ( n74628 , n74625 , n74627 );
nand ( n74629 , n72650 , n70933 );
and ( n74630 , n72782 , n70575 );
not ( n74631 , n70999 );
not ( n74632 , n72827 );
or ( n74633 , n74631 , n74632 );
nand ( n74634 , n70851 , n72630 );
nand ( n74635 , n74633 , n74634 );
nor ( n74636 , n74630 , n74635 );
nand ( n74637 , n74629 , n74636 );
nor ( n74638 , n74628 , n74637 );
or ( n74639 , n74638 , n74492 );
nand ( n74640 , n74474 , n69719 );
nand ( n74641 , n74639 , n74640 );
buf ( n8499 , n74641 );
buf ( n8500 , 1'b0 );
not ( n74644 , n68842 );
buf ( n8502 , n74644 );
buf ( n8503 , n68638 );
not ( n74647 , n72849 );
and ( n74648 , n74647 , n74627 );
and ( n74649 , n72893 , n70575 );
not ( n74650 , n70999 );
not ( n74651 , n72910 );
or ( n74652 , n74650 , n74651 );
nand ( n74653 , n70851 , n72819 );
nand ( n74654 , n74652 , n74653 );
nor ( n74655 , n74649 , n74654 );
nand ( n74656 , n72870 , n70933 );
nand ( n74657 , n74655 , n74656 );
nor ( n74658 , n74648 , n74657 );
or ( n74659 , n74658 , n74492 );
nand ( n74660 , n74474 , n69697 );
nand ( n74661 , n74659 , n74660 );
buf ( n8519 , n74661 );
buf ( n8520 , 1'b0 );
not ( n74664 , n68842 );
buf ( n74665 , n74664 );
buf ( n74666 , n68638 );
not ( n74667 , n72937 );
and ( n74668 , n74667 , n70200 );
nand ( n74669 , n72956 , n70933 );
and ( n74670 , n72971 , n70575 );
not ( n74671 , n70999 );
not ( n74672 , n72986 );
or ( n74673 , n74671 , n74672 );
nand ( n74674 , n70851 , n72538 );
nand ( n74675 , n74673 , n74674 );
nor ( n74676 , n74670 , n74675 );
nand ( n74677 , n74669 , n74676 );
nor ( n74678 , n74668 , n74677 );
or ( n74679 , n74678 , n71020 );
nand ( n74680 , n71348 , n69669 );
nand ( n74681 , n74679 , n74680 );
buf ( n74682 , n74681 );
buf ( n8540 , 1'b0 );
not ( n74684 , n68842 );
buf ( n74685 , n74684 );
buf ( n74686 , n68638 );
not ( n74687 , n73011 );
and ( n74688 , n74687 , n74627 );
nand ( n74689 , n73026 , n70933 );
and ( n74690 , n70575 , n73044 );
not ( n74691 , n70999 );
not ( n74692 , n73060 );
or ( n74693 , n74691 , n74692 );
nand ( n74694 , n70851 , n72548 );
nand ( n74695 , n74693 , n74694 );
nor ( n74696 , n74690 , n74695 );
nand ( n74697 , n74689 , n74696 );
nor ( n74698 , n74688 , n74697 );
or ( n74699 , n74698 , n71348 );
nand ( n74700 , n74474 , n69841 );
nand ( n74701 , n74699 , n74700 );
buf ( n74702 , n74701 );
buf ( n74703 , 1'b0 );
not ( n74704 , n68842 );
buf ( n74705 , n74704 );
buf ( n74706 , n68638 );
not ( n74707 , n73083 );
and ( n74708 , n74707 , n70927 );
nand ( n74709 , n73096 , n70933 );
and ( n74710 , n73108 , n70575 );
not ( n74711 , n70999 );
not ( n74712 , n73121 );
or ( n74713 , n74711 , n74712 );
nand ( n74714 , n70851 , n72561 );
nand ( n74715 , n74713 , n74714 );
nor ( n74716 , n74710 , n74715 );
nand ( n74717 , n74709 , n74716 );
nor ( n74718 , n74708 , n74717 );
or ( n74719 , n74718 , n74474 );
nand ( n74720 , n74474 , n69916 );
nand ( n74721 , n74719 , n74720 );
buf ( n74722 , n74721 );
buf ( n74723 , 1'b0 );
not ( n74724 , n68842 );
buf ( n8582 , n74724 );
buf ( n74726 , n68638 );
not ( n74727 , n73147 );
and ( n74728 , n74727 , n70927 );
nand ( n74729 , n73165 , n70933 );
and ( n74730 , n73193 , n70575 );
not ( n74731 , n70999 );
not ( n74732 , n73206 );
or ( n74733 , n74731 , n74732 );
nand ( n74734 , n70851 , n72514 );
nand ( n74735 , n74733 , n74734 );
nor ( n74736 , n74730 , n74735 );
nand ( n74737 , n74729 , n74736 );
nor ( n74738 , n74728 , n74737 );
or ( n74739 , n74738 , n71348 );
nand ( n74740 , n74492 , n69759 );
nand ( n74741 , n74739 , n74740 );
buf ( n74742 , n74741 );
buf ( n74743 , 1'b0 );
not ( n74744 , n68842 );
buf ( n74745 , n74744 );
buf ( n8603 , n68638 );
not ( n74747 , n73228 );
and ( n74748 , n74747 , n70927 );
nand ( n74749 , n73243 , n70933 );
and ( n74750 , n73257 , n70575 );
not ( n74751 , n70999 );
not ( n74752 , n73270 );
or ( n74753 , n74751 , n74752 );
nand ( n74754 , n70851 , n72503 );
nand ( n74755 , n74753 , n74754 );
nor ( n74756 , n74750 , n74755 );
nand ( n74757 , n74749 , n74756 );
nor ( n74758 , n74748 , n74757 );
or ( n74759 , n74758 , n71348 );
nand ( n74760 , n74492 , n69781 );
nand ( n74761 , n74759 , n74760 );
buf ( n8619 , n74761 );
buf ( n8620 , 1'b0 );
not ( n74764 , n68842 );
buf ( n74765 , n74764 );
buf ( n74766 , n68638 );
not ( n74767 , n73293 );
and ( n74768 , n74767 , n70927 );
nand ( n74769 , n73308 , n70933 );
and ( n74770 , n73327 , n70575 );
not ( n74771 , n70999 );
not ( n74772 , n73341 );
or ( n74773 , n74771 , n74772 );
nand ( n74774 , n70851 , n72479 );
nand ( n74775 , n74773 , n74774 );
nor ( n74776 , n74770 , n74775 );
nand ( n74777 , n74769 , n74776 );
nor ( n74778 , n74768 , n74777 );
or ( n74779 , n74778 , n74474 );
nand ( n74780 , n74492 , n69886 );
nand ( n74781 , n74779 , n74780 );
buf ( n8639 , n74781 );
buf ( n8640 , 1'b0 );
not ( n74784 , n68842 );
buf ( n74785 , n74784 );
buf ( n74786 , n68638 );
not ( n74787 , n73365 );
and ( n74788 , n74787 , n74627 );
not ( n74789 , n70933 );
not ( n74790 , n73373 );
or ( n74791 , n74789 , n74790 );
and ( n74792 , n73385 , n70575 );
not ( n74793 , n70999 );
not ( n74794 , n73398 );
or ( n74795 , n74793 , n74794 );
nand ( n74796 , n70851 , n72489 );
nand ( n74797 , n74795 , n74796 );
nor ( n74798 , n74792 , n74797 );
nand ( n74799 , n74791 , n74798 );
nor ( n74800 , n74788 , n74799 );
or ( n74801 , n74800 , n71348 );
nand ( n74802 , n74474 , n69860 );
nand ( n74803 , n74801 , n74802 );
buf ( n8661 , n74803 );
buf ( n8662 , 1'b0 );
not ( n74806 , n68842 );
buf ( n74807 , n74806 );
buf ( n74808 , n68638 );
not ( n74809 , n73420 );
and ( n74810 , n74809 , n70200 );
not ( n74811 , n70933 );
not ( n74812 , n73430 );
or ( n74813 , n74811 , n74812 );
and ( n74814 , n73432 , n70575 );
and ( n74815 , n70851 , n70507 );
and ( n74816 , n73439 , n70999 );
nor ( n74817 , n74814 , n74815 , n74816 );
nand ( n74818 , n74813 , n74817 );
nor ( n74819 , n74810 , n74818 );
or ( n74820 , n74819 , n71020 );
nand ( n74821 , n71348 , n70053 );
nand ( n74822 , n74820 , n74821 );
buf ( n74823 , n74822 );
buf ( n74824 , 1'b0 );
not ( n74825 , n68842 );
buf ( n8683 , n74825 );
buf ( n74827 , n68638 );
and ( n74828 , n73594 , n70927 );
not ( n74829 , n70935 );
not ( n74830 , n73618 );
or ( n74831 , n74829 , n74830 );
and ( n74832 , n73637 , n70575 );
not ( n74833 , n70999 );
not ( n74834 , n73646 );
or ( n74835 , n74833 , n74834 );
nand ( n74836 , n70300 , n70851 );
nand ( n74837 , n74835 , n74836 );
nor ( n74838 , n74832 , n74837 );
nand ( n74839 , n74831 , n74838 );
nor ( n74840 , n74828 , n74839 );
or ( n74841 , n74840 , n71020 );
nand ( n74842 , n71020 , n69566 );
nand ( n74843 , n74841 , n74842 );
buf ( n74844 , n74843 );
buf ( n74845 , 1'b0 );
not ( n74846 , n68842 );
buf ( n74847 , n74846 );
buf ( n74848 , n68638 );
not ( n74849 , n73739 );
not ( n74850 , n70199 );
and ( n74851 , n74849 , n74850 );
not ( n74852 , n70575 );
not ( n74853 , n73757 );
or ( n74854 , n74852 , n74853 );
and ( n74855 , n73749 , n70933 );
nand ( n74856 , n70850 , n74530 );
and ( n74857 , n74856 , n70526 );
nor ( n74858 , n74855 , n74857 );
nand ( n74859 , n74854 , n74858 );
nor ( n74860 , n74851 , n74859 );
or ( n74861 , n74860 , n71020 );
nand ( n74862 , n71020 , n69961 );
nand ( n74863 , n74861 , n74862 );
buf ( n8721 , n74863 );
buf ( n8722 , 1'b0 );
not ( n74866 , n68842 );
buf ( n8724 , n74866 );
buf ( n8725 , n68638 );
not ( n74869 , n70168 );
and ( n74870 , n70152 , n74869 , n70185 , n70858 );
not ( n74871 , n74870 );
or ( n74872 , n71019 , n74871 );
nand ( n74873 , n74871 , n69545 );
nand ( n74874 , n74872 , n74873 );
buf ( n74875 , n74874 );
buf ( n8733 , 1'b0 );
not ( n74877 , n68842 );
buf ( n8735 , n74877 );
buf ( n8736 , n68638 );
or ( n74880 , n74449 , n74871 );
nand ( n74881 , n74871 , n3412 );
nand ( n74882 , n74880 , n74881 );
buf ( n8740 , n74882 );
buf ( n8741 , 1'b0 );
not ( n74885 , n68842 );
buf ( n8743 , n74885 );
buf ( n74887 , n68638 );
or ( n74888 , n74471 , n74871 );
nand ( n74889 , n74871 , n69472 );
nand ( n74890 , n74888 , n74889 );
buf ( n74891 , n74890 );
buf ( n74892 , 1'b0 );
not ( n74893 , n68842 );
buf ( n8751 , n74893 );
buf ( n8752 , n68638 );
or ( n74896 , n74490 , n74871 );
nand ( n74897 , n74871 , n69437 );
nand ( n74898 , n74896 , n74897 );
buf ( n8756 , n74898 );
buf ( n8757 , 1'b0 );
not ( n74901 , n68842 );
buf ( n74902 , n74901 );
buf ( n74903 , n68638 );
or ( n74904 , n74513 , n74871 );
nand ( n74905 , n74871 , n69504 );
nand ( n74906 , n74904 , n74905 );
buf ( n74907 , n74906 );
buf ( n74908 , 1'b0 );
not ( n74909 , n68842 );
buf ( n8767 , n74909 );
buf ( n8768 , n68638 );
or ( n74912 , n74535 , n74871 );
nand ( n74913 , n74871 , n69481 );
nand ( n74914 , n74912 , n74913 );
buf ( n74915 , n74914 );
buf ( n74916 , 1'b0 );
not ( n74917 , n68842 );
buf ( n74918 , n74917 );
buf ( n74919 , n68638 );
not ( n74920 , n74555 );
or ( n74921 , n74920 , n74871 );
or ( n74922 , n74870 , n69452 );
nand ( n74923 , n74921 , n74922 );
buf ( n74924 , n74923 );
buf ( n74925 , 1'b0 );
not ( n74926 , n68842 );
buf ( n74927 , n74926 );
buf ( n74928 , n68638 );
and ( n74929 , n74871 , n3799 );
not ( n74930 , n74871 );
and ( n74931 , n74930 , n73932 );
or ( n74932 , n74929 , n74931 );
buf ( n74933 , n74932 );
buf ( n74934 , 1'b0 );
not ( n74935 , n68842 );
buf ( n8793 , n74935 );
buf ( n8794 , n68638 );
or ( n74938 , n74574 , n74871 );
or ( n74939 , n74870 , n69909 );
nand ( n74940 , n74938 , n74939 );
buf ( n8798 , n74940 );
buf ( n8799 , 1'b0 );
not ( n74943 , n68842 );
buf ( n74944 , n74943 );
buf ( n74945 , n68638 );
or ( n74946 , n74594 , n74871 );
nand ( n74947 , n74871 , n70067 );
nand ( n74948 , n74946 , n74947 );
buf ( n74949 , n74948 );
buf ( n8807 , 1'b0 );
not ( n74951 , n68842 );
buf ( n8809 , n74951 );
buf ( n8810 , n68638 );
or ( n74954 , n74616 , n74871 );
nand ( n74955 , n74871 , n69736 );
nand ( n74956 , n74954 , n74955 );
buf ( n8814 , n74956 );
buf ( n8815 , 1'b0 );
not ( n74959 , n68842 );
buf ( n8817 , n74959 );
buf ( n74961 , n68638 );
or ( n74962 , n74638 , n74871 );
nand ( n74963 , n74871 , n69729 );
nand ( n74964 , n74962 , n74963 );
buf ( n74965 , n74964 );
buf ( n74966 , 1'b0 );
not ( n74967 , n68842 );
buf ( n8825 , n74967 );
buf ( n8826 , n68638 );
not ( n74970 , n69701 );
and ( n74971 , n74871 , n74970 );
not ( n74972 , n74871 );
and ( n74973 , n74972 , n74658 );
nor ( n74974 , n74971 , n74973 );
buf ( n74975 , n74974 );
buf ( n74976 , 1'b0 );
not ( n74977 , n68842 );
buf ( n74978 , n74977 );
buf ( n8836 , n68638 );
or ( n74980 , n74678 , n74871 );
nand ( n74981 , n74871 , n69685 );
nand ( n74982 , n74980 , n74981 );
buf ( n74983 , n74982 );
buf ( n8841 , 1'b0 );
not ( n74985 , n68842 );
buf ( n74986 , n74985 );
buf ( n74987 , n68638 );
or ( n74988 , n74698 , n74871 );
nand ( n74989 , n74871 , n69846 );
nand ( n74990 , n74988 , n74989 );
buf ( n74991 , n74990 );
buf ( n74992 , 1'b0 );
not ( n74993 , n68842 );
buf ( n74994 , n74993 );
buf ( n74995 , n68638 );
or ( n74996 , n74718 , n74871 );
nand ( n74997 , n74871 , n69927 );
nand ( n74998 , n74996 , n74997 );
buf ( n74999 , n74998 );
buf ( n75000 , 1'b0 );
not ( n75001 , n68842 );
buf ( n75002 , n75001 );
buf ( n8860 , n68638 );
or ( n75004 , n74738 , n74871 );
nand ( n75005 , n74871 , n69765 );
nand ( n75006 , n75004 , n75005 );
buf ( n75007 , n75006 );
buf ( n75008 , 1'b0 );
not ( n75009 , n68842 );
buf ( n8867 , n75009 );
buf ( n8868 , n68638 );
or ( n75012 , n74758 , n74871 );
nand ( n75013 , n74871 , n69792 );
nand ( n75014 , n75012 , n75013 );
buf ( n8872 , n75014 );
buf ( n8873 , 1'b0 );
not ( n75017 , n68842 );
buf ( n75018 , n75017 );
buf ( n75019 , n68638 );
or ( n75020 , n74778 , n74871 );
nand ( n75021 , n74871 , n69896 );
nand ( n75022 , n75020 , n75021 );
buf ( n75023 , n75022 );
buf ( n8881 , 1'b0 );
not ( n75025 , n68842 );
buf ( n8883 , n75025 );
buf ( n8884 , n68638 );
or ( n75028 , n74800 , n74871 );
nand ( n75029 , n74871 , n69871 );
nand ( n75030 , n75028 , n75029 );
buf ( n8888 , n75030 );
buf ( n8889 , 1'b0 );
not ( n75033 , n68842 );
buf ( n8891 , n75033 );
buf ( n75035 , n68638 );
or ( n75036 , n74819 , n74871 );
nand ( n75037 , n74871 , n70049 );
nand ( n75038 , n75036 , n75037 );
buf ( n75039 , n75038 );
buf ( n75040 , 1'b0 );
not ( n75041 , n68842 );
buf ( n8899 , n75041 );
buf ( n8900 , n68638 );
or ( n75044 , n71211 , n74871 );
nand ( n75045 , n74871 , n69800 );
nand ( n75046 , n75044 , n75045 );
buf ( n8904 , n75046 );
buf ( n8905 , 1'b0 );
not ( n75049 , n68842 );
buf ( n75050 , n75049 );
buf ( n75051 , n68638 );
or ( n75052 , n71267 , n74871 );
nand ( n75053 , n74871 , n69819 );
nand ( n75054 , n75052 , n75053 );
buf ( n75055 , n75054 );
buf ( n75056 , 1'b0 );
not ( n75057 , n68842 );
buf ( n8915 , n75057 );
buf ( n8916 , n68638 );
or ( n75060 , n71323 , n74871 );
nand ( n75061 , n74871 , n69649 );
nand ( n75062 , n75060 , n75061 );
buf ( n75063 , n75062 );
buf ( n75064 , 1'b0 );
not ( n75065 , n68842 );
buf ( n75066 , n75065 );
buf ( n75067 , n68638 );
or ( n75068 , n71345 , n74871 );
nand ( n75069 , n74871 , n69634 );
nand ( n75070 , n75068 , n75069 );
buf ( n75071 , n75070 );
buf ( n75072 , 1'b0 );
not ( n75073 , n68842 );
buf ( n75074 , n75073 );
buf ( n75075 , n68638 );
or ( n75076 , n71439 , n74871 );
nand ( n75077 , n74871 , n69615 );
nand ( n75078 , n75076 , n75077 );
buf ( n8936 , n75078 );
buf ( n75080 , 1'b0 );
not ( n75081 , n68842 );
buf ( n75082 , n75081 );
buf ( n8940 , n68638 );
or ( n75084 , n71512 , n74871 );
nand ( n75085 , n74871 , n69601 );
nand ( n75086 , n75084 , n75085 );
buf ( n8944 , n75086 );
buf ( n75088 , 1'b0 );
not ( n75089 , n68842 );
buf ( n8947 , n75089 );
buf ( n75091 , n68638 );
or ( n75092 , n74840 , n74871 );
nand ( n75093 , n74871 , n69576 );
nand ( n75094 , n75092 , n75093 );
buf ( n8952 , n75094 );
buf ( n75096 , 1'b0 );
not ( n75097 , n68842 );
buf ( n8955 , n75097 );
buf ( n8956 , n68638 );
or ( n75100 , n71578 , n74871 );
nand ( n75101 , n74871 , n69589 );
nand ( n75102 , n75100 , n75101 );
buf ( n75103 , n75102 );
buf ( n75104 , 1'b0 );
not ( n75105 , n68842 );
buf ( n8963 , n75105 );
buf ( n8964 , n68638 );
or ( n75108 , n71658 , n74871 );
nand ( n75109 , n74871 , n69521 );
nand ( n75110 , n75108 , n75109 );
buf ( n75111 , n75110 );
buf ( n75112 , 1'b0 );
not ( n75113 , n68842 );
buf ( n75114 , n75113 );
buf ( n75115 , n68638 );
or ( n75116 , n71718 , n74871 );
nand ( n75117 , n74871 , n69533 );
nand ( n75118 , n75116 , n75117 );
buf ( n75119 , n75118 );
buf ( n75120 , 1'b0 );
not ( n75121 , n68842 );
buf ( n8979 , n75121 );
buf ( n75123 , n68638 );
or ( n75124 , n74860 , n74871 );
or ( n75125 , n74870 , n69966 );
nand ( n75126 , n75124 , n75125 );
buf ( n8984 , n75126 );
buf ( n8985 , 1'b0 );
not ( n75129 , n68842 );
buf ( n75130 , n75129 );
buf ( n75131 , n68638 );
and ( n75132 , n71847 , n2669 );
not ( n75133 , n71847 );
and ( n75134 , n75133 , n70086 );
or ( n75135 , n75132 , n75134 );
buf ( n75136 , n75135 );
buf ( n75137 , 1'b0 );
not ( n75138 , n68842 );
buf ( n75139 , n75138 );
buf ( n75140 , n68638 );
and ( n75141 , n71847 , n68814 );
not ( n75142 , n71847 );
and ( n75143 , n75142 , n70094 );
or ( n75144 , n75141 , n75143 );
buf ( n75145 , n75144 );
buf ( n75146 , 1'b0 );
not ( n75147 , n68842 );
buf ( n75148 , n75147 );
buf ( n75149 , n68638 );
and ( n75150 , n71847 , n2673 );
not ( n75151 , n71847 );
and ( n75152 , n75151 , n70035 );
or ( n75153 , n75150 , n75152 );
buf ( n75154 , n75153 );
buf ( n75155 , 1'b0 );
not ( n75156 , n68842 );
buf ( n9014 , n75156 );
buf ( n9015 , n68638 );
and ( n75159 , n71847 , n68818 );
not ( n75160 , n71847 );
and ( n75161 , n75160 , n70028 );
or ( n75162 , n75159 , n75161 );
buf ( n9020 , n75162 );
buf ( n9021 , 1'b0 );
not ( n75165 , n68842 );
buf ( n75166 , n75165 );
buf ( n75167 , n68638 );
and ( n75168 , n71729 , n68822 );
not ( n75169 , n71729 );
and ( n75170 , n75169 , n70042 );
or ( n75171 , n75168 , n75170 );
buf ( n9029 , n75171 );
buf ( n9030 , 1'b0 );
not ( n75174 , n68842 );
buf ( n9032 , n75174 );
buf ( n75176 , n68638 );
not ( n75177 , n71729 );
not ( n75178 , n75177 );
not ( n75179 , n70044 );
or ( n75180 , n75178 , n75179 );
nand ( n75181 , n71847 , n68827 );
nand ( n75182 , n75180 , n75181 );
buf ( n75183 , n75182 );
buf ( n75184 , 1'b0 );
not ( n75185 , n68842 );
buf ( n75186 , n75185 );
buf ( n75187 , n68638 );
and ( n75188 , n71729 , n68768 );
not ( n75189 , n71729 );
and ( n75190 , n75189 , n73906 );
or ( n75191 , n75188 , n75190 );
buf ( n75192 , n75191 );
buf ( n75193 , 1'b0 );
not ( n75194 , n68842 );
buf ( n9052 , n75194 );
buf ( n9053 , n68638 );
not ( n75197 , n70077 );
not ( n75198 , n71729 );
not ( n75199 , n75198 );
or ( n75200 , n75197 , n75199 );
not ( n75201 , n68830 );
or ( n75202 , n71846 , n75201 );
nand ( n75203 , n75200 , n75202 );
buf ( n75204 , n75203 );
buf ( n75205 , 1'b0 );
not ( n75206 , n68842 );
buf ( n9064 , n75206 );
buf ( n75208 , n68638 );
and ( n75209 , n71729 , n68770 );
not ( n75210 , n71729 );
and ( n75211 , n75210 , n72467 );
or ( n75212 , n75209 , n75211 );
buf ( n75213 , n75212 );
buf ( n75214 , 1'b0 );
not ( n75215 , n68842 );
buf ( n75216 , n75215 );
buf ( n75217 , n68638 );
and ( n75218 , n71729 , n2629 );
not ( n75219 , n71729 );
and ( n75220 , n75219 , n72456 );
or ( n75221 , n75218 , n75220 );
buf ( n75222 , n75221 );
buf ( n75223 , 1'b0 );
not ( n75224 , n68842 );
buf ( n9082 , n75224 );
buf ( n9083 , n68638 );
not ( n75227 , n70057 );
not ( n75228 , n75198 );
or ( n75229 , n75227 , n75228 );
not ( n75230 , n71729 );
not ( n75231 , n2689 );
or ( n75232 , n75230 , n75231 );
nand ( n75233 , n75229 , n75232 );
buf ( n9091 , n75233 );
buf ( n9092 , 1'b0 );
not ( n75236 , n68842 );
buf ( n75237 , n75236 );
buf ( n75238 , n68638 );
not ( n75239 , n69971 );
not ( n75240 , n71729 );
not ( n75241 , n75240 );
or ( n75242 , n75239 , n75241 );
not ( n75243 , n68834 );
or ( n75244 , n75230 , n75243 );
nand ( n75245 , n75242 , n75244 );
buf ( n75246 , n75245 );
buf ( n75247 , 1'b0 );
not ( n75248 , n68842 );
buf ( n75249 , n75248 );
buf ( n75250 , n68638 );
nor ( n75251 , n70865 , n70151 );
not ( n75252 , n75251 );
or ( n75253 , n75252 , n70185 );
or ( n75254 , n75251 , n70174 );
nand ( n75255 , n75253 , n75254 );
buf ( n75256 , n75255 );
buf ( n75257 , 1'b0 );
not ( n75258 , n68842 );
buf ( n75259 , n75258 );
buf ( n75260 , n68638 );
or ( n75261 , n75252 , n74869 );
not ( n75262 , n4022 );
or ( n75263 , n75251 , n75262 );
nand ( n75264 , n75261 , n75263 );
buf ( n75265 , n75264 );
buf ( n75266 , 1'b0 );
not ( n75267 , n68842 );
buf ( n9125 , n75267 );
buf ( n9126 , n68638 );
not ( n75270 , n70199 );
not ( n75271 , n70144 );
or ( n75272 , n75270 , n75271 );
nand ( n75273 , n70151 , n70143 );
nand ( n75274 , n75272 , n75273 );
not ( n75275 , n70221 );
and ( n75276 , n69362 , n75275 );
and ( n75277 , n75274 , n75276 );
nand ( n75278 , n75277 , n69127 );
and ( n75279 , n69361 , n75275 );
nand ( n75280 , n75274 , n75279 );
not ( n75281 , n75280 );
nor ( n75282 , n69127 , n69537 );
not ( n75283 , n75282 );
nand ( n75284 , n69127 , n69537 );
nand ( n75285 , n75283 , n75284 );
not ( n75286 , n75285 );
or ( n75287 , n3276 , n69063 );
not ( n75288 , n75287 );
not ( n75289 , n69014 );
not ( n75290 , n75289 );
nor ( n75291 , n75290 , n3320 );
nor ( n75292 , n75288 , n75291 );
not ( n75293 , n69029 );
not ( n75294 , n75293 );
nor ( n75295 , n75294 , n3350 );
nand ( n75296 , n69087 , n3346 );
or ( n75297 , n75295 , n75296 );
nand ( n75298 , n75294 , n3350 );
nand ( n75299 , n75297 , n75298 );
and ( n75300 , n75292 , n75299 );
nand ( n75301 , n69063 , n3276 );
or ( n75302 , n75291 , n75301 );
nand ( n75303 , n75290 , n3320 );
nand ( n75304 , n75302 , n75303 );
nor ( n75305 , n75300 , n75304 );
nor ( n75306 , n69087 , n3346 );
nor ( n75307 , n75295 , n75306 );
nor ( n75308 , n69076 , n69441 );
nand ( n75309 , n69099 , n70062 );
or ( n75310 , n75308 , n75309 );
nand ( n75311 , n69076 , n69441 );
nand ( n75312 , n75310 , n75311 );
or ( n75313 , n70062 , n69099 );
and ( n75314 , n3815 , n2728 );
xor ( n75315 , n70055 , n75314 );
and ( n75316 , n75315 , n69110 );
and ( n75317 , n70055 , n75314 );
or ( n75318 , n75316 , n75317 );
nand ( n75319 , n75313 , n75318 );
nor ( n75320 , n75308 , n75319 );
or ( n75321 , n75312 , n75320 );
nand ( n75322 , n75292 , n75307 , n75321 );
nand ( n75323 , n75305 , n75322 );
not ( n75324 , n75323 );
nor ( n75325 , n68992 , n3405 );
or ( n75326 , n75324 , n75325 );
nand ( n75327 , n68992 , n3405 );
nand ( n75328 , n75326 , n75327 );
not ( n75329 , n75328 );
or ( n75330 , n75286 , n75329 );
or ( n75331 , n75328 , n75285 );
nand ( n75332 , n75330 , n75331 );
nand ( n75333 , n75281 , n75332 );
not ( n75334 , n69361 );
nor ( n75335 , n75334 , n75275 );
and ( n75336 , n75274 , n75335 );
nor ( n75337 , n69127 , n69539 );
not ( n75338 , n75337 );
nand ( n75339 , n69127 , n69539 );
nand ( n75340 , n75338 , n75339 );
not ( n75341 , n75340 );
or ( n75342 , n3282 , n69063 );
not ( n75343 , n75342 );
not ( n75344 , n75289 );
nor ( n75345 , n75344 , n3316 );
nor ( n75346 , n75343 , n75345 );
not ( n75347 , n75293 );
nor ( n75348 , n75347 , n69496 );
nand ( n75349 , n69087 , n3342 );
or ( n75350 , n75348 , n75349 );
nand ( n75351 , n75347 , n69496 );
nand ( n75352 , n75350 , n75351 );
and ( n75353 , n75346 , n75352 );
nand ( n75354 , n69063 , n3282 );
or ( n75355 , n75345 , n75354 );
nand ( n75356 , n75344 , n3316 );
nand ( n75357 , n75355 , n75356 );
nor ( n75358 , n75353 , n75357 );
nor ( n75359 , n69087 , n3342 );
nor ( n75360 , n75348 , n75359 );
nor ( n75361 , n69076 , n3301 );
nand ( n75362 , n69099 , n70073 );
or ( n75363 , n75361 , n75362 );
nand ( n75364 , n69076 , n3301 );
nand ( n75365 , n75363 , n75364 );
or ( n75366 , n70073 , n69099 );
and ( n75367 , n69961 , n2728 );
xor ( n75368 , n70053 , n75367 );
and ( n75369 , n75368 , n69110 );
and ( n75370 , n70053 , n75367 );
or ( n75371 , n75369 , n75370 );
nand ( n75372 , n75366 , n75371 );
nor ( n75373 , n75361 , n75372 );
or ( n75374 , n75365 , n75373 );
nand ( n75375 , n75346 , n75360 , n75374 );
nand ( n75376 , n75358 , n75375 );
not ( n75377 , n75376 );
nor ( n75378 , n68992 , n69550 );
or ( n75379 , n75377 , n75378 );
nand ( n75380 , n68992 , n69550 );
nand ( n75381 , n75379 , n75380 );
not ( n75382 , n75381 );
or ( n75383 , n75341 , n75382 );
or ( n75384 , n75381 , n75340 );
nand ( n75385 , n75383 , n75384 );
nand ( n75386 , n75336 , n75385 );
nor ( n75387 , n70140 , n70151 );
not ( n75388 , n70199 );
and ( n75389 , n75388 , n70867 );
nor ( n75390 , n69361 , n75275 );
nor ( n75391 , n75389 , n75390 );
or ( n75392 , n75387 , n75391 , n71996 );
not ( n75393 , n75392 );
and ( n75394 , n75393 , n68724 );
not ( n75395 , n72024 );
nor ( n75396 , n75394 , n75395 );
nand ( n75397 , n75278 , n75333 , n75386 , n75396 );
buf ( n75398 , n75397 );
buf ( n75399 , 1'b0 );
not ( n75400 , n68842 );
buf ( n9258 , n75400 );
buf ( n9259 , n68638 );
nand ( n75403 , n75277 , n68992 );
not ( n75404 , n75325 );
nand ( n75405 , n75404 , n75327 );
not ( n75406 , n75405 );
not ( n75407 , n75323 );
or ( n75408 , n75406 , n75407 );
or ( n75409 , n75323 , n75405 );
nand ( n75410 , n75408 , n75409 );
nand ( n75411 , n75281 , n75410 );
not ( n75412 , n75378 );
nand ( n75413 , n75412 , n75380 );
not ( n75414 , n75413 );
not ( n75415 , n75376 );
or ( n75416 , n75414 , n75415 );
or ( n75417 , n75376 , n75413 );
nand ( n75418 , n75416 , n75417 );
nand ( n75419 , n75336 , n75418 );
and ( n75420 , n75393 , n68729 );
nor ( n75421 , n75420 , n72076 );
nand ( n75422 , n75403 , n75411 , n75419 , n75421 );
buf ( n75423 , n75422 );
buf ( n75424 , 1'b0 );
not ( n75425 , n68842 );
buf ( n75426 , n75425 );
buf ( n9284 , n68638 );
nand ( n75428 , n75277 , n69014 );
not ( n75429 , n75303 );
nor ( n75430 , n75429 , n75291 );
not ( n75431 , n75430 );
and ( n75432 , n75307 , n75321 , n75287 );
not ( n75433 , n75287 );
not ( n75434 , n75299 );
or ( n75435 , n75433 , n75434 );
nand ( n75436 , n75435 , n75301 );
nor ( n75437 , n75432 , n75436 );
not ( n75438 , n75437 );
or ( n75439 , n75431 , n75438 );
or ( n75440 , n75437 , n75430 );
nand ( n75441 , n75439 , n75440 );
nand ( n75442 , n75281 , n75441 );
not ( n75443 , n75356 );
nor ( n75444 , n75443 , n75345 );
not ( n75445 , n75444 );
and ( n75446 , n75360 , n75374 , n75342 );
not ( n75447 , n75342 );
not ( n75448 , n75352 );
or ( n75449 , n75447 , n75448 );
nand ( n75450 , n75449 , n75354 );
nor ( n75451 , n75446 , n75450 );
not ( n75452 , n75451 );
or ( n75453 , n75445 , n75452 );
or ( n75454 , n75451 , n75444 );
nand ( n75455 , n75453 , n75454 );
nand ( n75456 , n75336 , n75455 );
and ( n75457 , n75393 , n68734 );
nor ( n75458 , n75457 , n72142 );
nand ( n75459 , n75428 , n75442 , n75456 , n75458 );
buf ( n9317 , n75459 );
buf ( n9318 , 1'b0 );
not ( n75462 , n68842 );
buf ( n75463 , n75462 );
buf ( n75464 , n68638 );
nand ( n75465 , n75277 , n69063 );
and ( n75466 , n75287 , n75301 );
not ( n75467 , n75466 );
and ( n75468 , n75307 , n75321 );
nor ( n75469 , n75468 , n75299 );
not ( n75470 , n75469 );
or ( n75471 , n75467 , n75470 );
or ( n75472 , n75469 , n75466 );
nand ( n75473 , n75471 , n75472 );
nand ( n75474 , n75281 , n75473 );
and ( n75475 , n75342 , n75354 );
not ( n75476 , n75475 );
and ( n75477 , n75360 , n75374 );
nor ( n75478 , n75477 , n75352 );
not ( n75479 , n75478 );
or ( n75480 , n75476 , n75479 );
or ( n75481 , n75478 , n75475 );
nand ( n75482 , n75480 , n75481 );
nand ( n75483 , n75336 , n75482 );
and ( n75484 , n75393 , n68739 );
nor ( n75485 , n75484 , n72204 );
nand ( n75486 , n75465 , n75474 , n75483 , n75485 );
buf ( n75487 , n75486 );
buf ( n75488 , 1'b0 );
not ( n75489 , n68842 );
buf ( n75490 , n75489 );
buf ( n75491 , n68638 );
nand ( n75492 , n75277 , n69029 );
not ( n75493 , n75295 );
nand ( n75494 , n75493 , n75298 );
not ( n75495 , n75494 );
not ( n75496 , n75321 );
or ( n75497 , n75496 , n75306 );
nand ( n75498 , n75497 , n75296 );
not ( n75499 , n75498 );
or ( n75500 , n75495 , n75499 );
or ( n75501 , n75498 , n75494 );
nand ( n75502 , n75500 , n75501 );
nand ( n75503 , n75281 , n75502 );
not ( n75504 , n75348 );
nand ( n75505 , n75504 , n75351 );
not ( n75506 , n75505 );
not ( n75507 , n75374 );
or ( n75508 , n75507 , n75359 );
nand ( n75509 , n75508 , n75349 );
not ( n75510 , n75509 );
or ( n75511 , n75506 , n75510 );
or ( n75512 , n75509 , n75505 );
nand ( n75513 , n75511 , n75512 );
nand ( n75514 , n75336 , n75513 );
and ( n75515 , n75393 , n68744 );
nor ( n75516 , n75515 , n72266 );
nand ( n75517 , n75492 , n75503 , n75514 , n75516 );
buf ( n75518 , n75517 );
buf ( n75519 , 1'b0 );
not ( n75520 , n68842 );
buf ( n75521 , n75520 );
buf ( n75522 , n68638 );
nand ( n75523 , n75277 , n69087 );
not ( n75524 , n75296 );
nor ( n75525 , n75524 , n75306 );
not ( n75526 , n75525 );
not ( n75527 , n75496 );
or ( n75528 , n75526 , n75527 );
or ( n75529 , n75496 , n75525 );
nand ( n75530 , n75528 , n75529 );
nand ( n75531 , n75281 , n75530 );
not ( n75532 , n75349 );
nor ( n75533 , n75532 , n75359 );
not ( n75534 , n75533 );
not ( n75535 , n75507 );
or ( n75536 , n75534 , n75535 );
or ( n75537 , n75507 , n75533 );
nand ( n75538 , n75536 , n75537 );
nand ( n75539 , n75336 , n75538 );
not ( n75540 , n75392 );
not ( n75541 , n2604 );
not ( n75542 , n75541 );
and ( n75543 , n75540 , n75542 );
not ( n75544 , n3815 );
not ( n75545 , n75279 );
or ( n75546 , n75544 , n75545 );
nand ( n75547 , n75335 , n69961 );
nand ( n75548 , n75546 , n75547 );
xnor ( n75549 , n75548 , n2728 );
or ( n75550 , n71729 , n75549 );
nand ( n75551 , n75550 , n72315 );
nor ( n75552 , n75543 , n75551 );
nand ( n75553 , n75523 , n75531 , n75539 , n75552 );
buf ( n75554 , n75553 );
buf ( n75555 , 1'b0 );
not ( n75556 , n68842 );
buf ( n75557 , n75556 );
buf ( n75558 , n68638 );
nand ( n75559 , n75277 , n69076 );
nand ( n75560 , n75319 , n75309 );
not ( n75561 , n75560 );
not ( n75562 , n75308 );
nand ( n75563 , n75562 , n75311 );
not ( n75564 , n75563 );
or ( n75565 , n75561 , n75564 );
or ( n75566 , n75563 , n75560 );
nand ( n75567 , n75565 , n75566 );
nand ( n75568 , n75281 , n75567 );
nand ( n75569 , n75372 , n75362 );
not ( n75570 , n75569 );
not ( n75571 , n75361 );
nand ( n75572 , n75571 , n75364 );
not ( n75573 , n75572 );
or ( n75574 , n75570 , n75573 );
or ( n75575 , n75572 , n75569 );
nand ( n75576 , n75574 , n75575 );
nand ( n75577 , n75336 , n75576 );
and ( n75578 , n75393 , n68751 );
nor ( n75579 , n75578 , n72372 );
nand ( n75580 , n75559 , n75568 , n75577 , n75579 );
buf ( n75581 , n75580 );
buf ( n75582 , 1'b0 );
not ( n75583 , n68842 );
buf ( n75584 , n75583 );
buf ( n75585 , n68638 );
not ( n75586 , n75318 );
nand ( n75587 , n75309 , n75313 );
not ( n75588 , n75587 );
or ( n75589 , n75586 , n75588 );
or ( n75590 , n75587 , n75318 );
nand ( n75591 , n75589 , n75590 );
nand ( n75592 , n75281 , n75591 );
nand ( n75593 , n75277 , n69099 );
not ( n75594 , n75371 );
nand ( n75595 , n75362 , n75366 );
not ( n75596 , n75595 );
or ( n75597 , n75594 , n75596 );
or ( n75598 , n75595 , n75371 );
nand ( n75599 , n75597 , n75598 );
nand ( n75600 , n75336 , n75599 );
not ( n75601 , n75392 );
not ( n75602 , n68754 );
not ( n75603 , n75602 );
and ( n75604 , n75601 , n75603 );
not ( n75605 , n70863 );
not ( n75606 , n70058 );
or ( n75607 , n75605 , n75606 );
nand ( n75608 , n75607 , n75550 );
nor ( n75609 , n75604 , n75608 );
nand ( n75610 , n75592 , n75593 , n75600 , n75609 );
buf ( n75611 , n75610 );
buf ( n75612 , 1'b0 );
not ( n75613 , n68842 );
buf ( n75614 , n75613 );
buf ( n75615 , n68638 );
nand ( n75616 , n75277 , n69110 );
xor ( n75617 , n70055 , n75314 );
xor ( n75618 , n75617 , n69110 );
nand ( n75619 , n75281 , n75618 );
xor ( n75620 , n70053 , n75367 );
xor ( n75621 , n75620 , n69110 );
nand ( n75622 , n75336 , n75621 );
and ( n75623 , n75393 , n68758 );
and ( n75624 , n70045 , n70863 );
nor ( n75625 , n75623 , n75624 );
nand ( n75626 , n75616 , n75619 , n75622 , n75625 );
buf ( n9484 , n75626 );
buf ( n75628 , 1'b0 );
not ( n75629 , n68842 );
buf ( n75630 , n75629 );
buf ( n9488 , n68638 );
nand ( n75632 , n75277 , n69244 );
not ( n75633 , n69244 );
not ( n75634 , n69802 );
and ( n75635 , n75633 , n75634 );
and ( n75636 , n69244 , n69802 );
nor ( n75637 , n75635 , n75636 );
not ( n75638 , n75637 );
or ( n75639 , n69049 , n69526 );
not ( n75640 , n75639 );
nor ( n75641 , n68981 , n69511 );
nor ( n75642 , n75640 , n75641 );
or ( n75643 , n75282 , n75327 );
nand ( n75644 , n75643 , n75284 );
and ( n75645 , n75642 , n75644 );
nand ( n75646 , n69049 , n69526 );
or ( n75647 , n75641 , n75646 );
nand ( n75648 , n68981 , n69511 );
nand ( n75649 , n75647 , n75648 );
nor ( n75650 , n75645 , n75649 );
nor ( n75651 , n75282 , n75325 );
and ( n75652 , n75642 , n75651 );
nand ( n75653 , n75652 , n75323 );
nand ( n75654 , n75650 , n75653 );
nor ( n75655 , n68938 , n3466 );
nor ( n75656 , n68965 , n3450 );
nor ( n75657 , n75655 , n75656 );
nor ( n75658 , n68951 , n69562 );
nor ( n75659 , n68912 , n69581 );
nor ( n75660 , n75658 , n75659 );
nand ( n75661 , n75657 , n75660 );
not ( n75662 , n75661 );
nor ( n75663 , n69161 , n69810 );
not ( n75664 , n75663 );
nor ( n75665 , n69180 , n69655 );
nor ( n75666 , n69191 , n2697 );
nor ( n75667 , n75665 , n75666 );
nand ( n75668 , n75664 , n75667 );
not ( n75669 , n75668 );
and ( n75670 , n75654 , n75662 , n75669 );
nand ( n75671 , n68912 , n69581 );
or ( n75672 , n75658 , n75671 );
nand ( n75673 , n68951 , n69562 );
nand ( n75674 , n75672 , n75673 );
and ( n75675 , n75657 , n75674 );
nand ( n75676 , n68965 , n3450 );
or ( n75677 , n75655 , n75676 );
nand ( n75678 , n68938 , n3466 );
nand ( n75679 , n75677 , n75678 );
nor ( n75680 , n75675 , n75679 );
or ( n75681 , n75680 , n75668 );
nand ( n75682 , n69191 , n2697 );
or ( n75683 , n75665 , n75682 );
nand ( n75684 , n69180 , n69655 );
nand ( n75685 , n75683 , n75684 );
not ( n75686 , n75685 );
or ( n75687 , n75663 , n75686 );
nand ( n75688 , n69161 , n69810 );
nand ( n75689 , n75681 , n75687 , n75688 );
nor ( n75690 , n75670 , n75689 );
not ( n75691 , n75690 );
or ( n75692 , n75638 , n75691 );
or ( n75693 , n75690 , n75637 );
nand ( n75694 , n75692 , n75693 );
nand ( n75695 , n75281 , n75694 );
not ( n75696 , n69244 );
not ( n75697 , n69804 );
and ( n75698 , n75696 , n75697 );
and ( n75699 , n69244 , n69804 );
nor ( n75700 , n75698 , n75699 );
not ( n75701 , n75700 );
or ( n75702 , n69049 , n69528 );
not ( n75703 , n75702 );
nor ( n75704 , n68981 , n69513 );
nor ( n75705 , n75703 , n75704 );
or ( n75706 , n75337 , n75380 );
nand ( n75707 , n75706 , n75339 );
and ( n75708 , n75705 , n75707 );
nand ( n75709 , n69049 , n69528 );
or ( n75710 , n75704 , n75709 );
nand ( n75711 , n68981 , n69513 );
nand ( n75712 , n75710 , n75711 );
nor ( n75713 , n75708 , n75712 );
nor ( n75714 , n75337 , n75378 );
and ( n75715 , n75705 , n75714 );
nand ( n75716 , n75715 , n75376 );
nand ( n75717 , n75713 , n75716 );
nor ( n75718 , n68938 , n69611 );
nor ( n75719 , n68965 , n69595 );
nor ( n75720 , n75718 , n75719 );
nor ( n75721 , n68951 , n69566 );
nor ( n75722 , n68912 , n69583 );
nor ( n75723 , n75721 , n75722 );
nand ( n75724 , n75720 , n75723 );
not ( n75725 , n75724 );
nor ( n75726 , n69161 , n69814 );
not ( n75727 , n75726 );
nor ( n75728 , n69180 , n3510 );
nor ( n75729 , n69191 , n3498 );
nor ( n75730 , n75728 , n75729 );
nand ( n75731 , n75727 , n75730 );
not ( n75732 , n75731 );
and ( n75733 , n75717 , n75725 , n75732 );
nand ( n75734 , n68912 , n69583 );
or ( n75735 , n75721 , n75734 );
nand ( n75736 , n68951 , n69566 );
nand ( n75737 , n75735 , n75736 );
and ( n75738 , n75720 , n75737 );
nand ( n75739 , n68965 , n69595 );
or ( n75740 , n75718 , n75739 );
nand ( n75741 , n68938 , n69611 );
nand ( n75742 , n75740 , n75741 );
nor ( n75743 , n75738 , n75742 );
or ( n75744 , n75743 , n75731 );
nand ( n75745 , n69191 , n3498 );
or ( n75746 , n75728 , n75745 );
nand ( n75747 , n69180 , n3510 );
nand ( n75748 , n75746 , n75747 );
not ( n75749 , n75748 );
or ( n75750 , n75726 , n75749 );
nand ( n75751 , n69161 , n69814 );
nand ( n75752 , n75744 , n75750 , n75751 );
nor ( n75753 , n75733 , n75752 );
not ( n75754 , n75753 );
or ( n75755 , n75701 , n75754 );
or ( n75756 , n75753 , n75700 );
nand ( n75757 , n75755 , n75756 );
nand ( n75758 , n75336 , n75757 );
and ( n75759 , n75393 , n68674 );
nor ( n75760 , n75759 , n73460 );
nand ( n75761 , n75632 , n75695 , n75758 , n75760 );
buf ( n75762 , n75761 );
buf ( n9620 , 1'b0 );
not ( n75764 , n68842 );
buf ( n9622 , n75764 );
buf ( n9623 , n68638 );
nand ( n75767 , n75277 , n69161 );
not ( n75768 , n75688 );
nor ( n75769 , n75768 , n75663 );
not ( n75770 , n75769 );
and ( n75771 , n75654 , n75662 , n75667 );
not ( n75772 , n75685 );
not ( n75773 , n75680 );
nand ( n75774 , n75773 , n75667 );
nand ( n75775 , n75772 , n75774 );
nor ( n75776 , n75771 , n75775 );
not ( n75777 , n75776 );
or ( n75778 , n75770 , n75777 );
or ( n75779 , n75776 , n75769 );
nand ( n75780 , n75778 , n75779 );
nand ( n75781 , n75281 , n75780 );
not ( n75782 , n75751 );
nor ( n75783 , n75782 , n75726 );
not ( n75784 , n75783 );
and ( n75785 , n75717 , n75725 , n75730 );
not ( n75786 , n75748 );
not ( n75787 , n75743 );
nand ( n75788 , n75787 , n75730 );
nand ( n75789 , n75786 , n75788 );
nor ( n75790 , n75785 , n75789 );
not ( n75791 , n75790 );
or ( n75792 , n75784 , n75791 );
or ( n75793 , n75790 , n75783 );
nand ( n75794 , n75792 , n75793 );
nand ( n75795 , n75336 , n75794 );
and ( n75796 , n75393 , n68679 );
nor ( n75797 , n75796 , n73482 );
nand ( n75798 , n75767 , n75781 , n75795 , n75797 );
buf ( n9656 , n75798 );
buf ( n9657 , 1'b0 );
not ( n75801 , n68842 );
buf ( n75802 , n75801 );
buf ( n75803 , n68638 );
nand ( n75804 , n75277 , n69180 );
not ( n75805 , n75665 );
nand ( n75806 , n75805 , n75684 );
not ( n75807 , n75806 );
or ( n75808 , n75680 , n75666 );
not ( n75809 , n75666 );
nand ( n75810 , n75809 , n75654 , n75662 );
nand ( n75811 , n75808 , n75810 , n75682 );
not ( n75812 , n75811 );
or ( n75813 , n75807 , n75812 );
or ( n75814 , n75811 , n75806 );
nand ( n75815 , n75813 , n75814 );
nand ( n75816 , n75281 , n75815 );
not ( n75817 , n75728 );
nand ( n75818 , n75817 , n75747 );
not ( n75819 , n75818 );
or ( n75820 , n75743 , n75729 );
not ( n75821 , n75729 );
nand ( n75822 , n75821 , n75717 , n75725 );
nand ( n75823 , n75820 , n75822 , n75745 );
not ( n75824 , n75823 );
or ( n75825 , n75819 , n75824 );
or ( n75826 , n75823 , n75818 );
nand ( n75827 , n75825 , n75826 );
nand ( n75828 , n75336 , n75827 );
and ( n75829 , n75393 , n68684 );
nor ( n75830 , n75829 , n73504 );
nand ( n75831 , n75804 , n75816 , n75828 , n75830 );
buf ( n9689 , n75831 );
buf ( n9690 , 1'b0 );
not ( n75834 , n68842 );
buf ( n75835 , n75834 );
buf ( n75836 , n68638 );
nand ( n75837 , n75277 , n69191 );
not ( n75838 , n75666 );
nand ( n75839 , n75838 , n75682 );
not ( n75840 , n75839 );
or ( n75841 , n75653 , n75661 );
or ( n75842 , n75661 , n75650 );
nand ( n75843 , n75841 , n75842 , n75680 );
not ( n75844 , n75843 );
or ( n75845 , n75840 , n75844 );
or ( n75846 , n75843 , n75839 );
nand ( n75847 , n75845 , n75846 );
nand ( n75848 , n75281 , n75847 );
not ( n75849 , n75729 );
nand ( n75850 , n75849 , n75745 );
not ( n75851 , n75850 );
or ( n75852 , n75716 , n75724 );
or ( n75853 , n75724 , n75713 );
nand ( n75854 , n75852 , n75853 , n75743 );
not ( n75855 , n75854 );
or ( n75856 , n75851 , n75855 );
or ( n75857 , n75854 , n75850 );
nand ( n75858 , n75856 , n75857 );
nand ( n75859 , n75336 , n75858 );
and ( n75860 , n75393 , n68689 );
nor ( n75861 , n75860 , n73525 );
nand ( n75862 , n75837 , n75848 , n75859 , n75861 );
buf ( n9720 , n75862 );
buf ( n9721 , 1'b0 );
not ( n75865 , n68842 );
buf ( n9723 , n75865 );
buf ( n75867 , n68638 );
nand ( n75868 , n75277 , n68938 );
not ( n75869 , n75678 );
nor ( n75870 , n75869 , n75655 );
not ( n75871 , n75870 );
not ( n75872 , n75656 );
and ( n75873 , n75660 , n75872 );
and ( n75874 , n75652 , n75873 , n75323 );
not ( n75875 , n75873 );
not ( n75876 , n75650 );
not ( n75877 , n75876 );
or ( n75878 , n75875 , n75877 );
and ( n75879 , n75674 , n75872 );
not ( n75880 , n75676 );
nor ( n75881 , n75879 , n75880 );
nand ( n75882 , n75878 , n75881 );
nor ( n75883 , n75874 , n75882 );
not ( n75884 , n75883 );
or ( n75885 , n75871 , n75884 );
or ( n75886 , n75883 , n75870 );
nand ( n75887 , n75885 , n75886 );
nand ( n75888 , n75281 , n75887 );
not ( n75889 , n75741 );
nor ( n75890 , n75889 , n75718 );
not ( n75891 , n75890 );
not ( n75892 , n75719 );
and ( n75893 , n75723 , n75892 );
and ( n75894 , n75715 , n75893 , n75376 );
not ( n75895 , n75893 );
not ( n75896 , n75713 );
not ( n75897 , n75896 );
or ( n75898 , n75895 , n75897 );
and ( n75899 , n75737 , n75892 );
not ( n75900 , n75739 );
nor ( n75901 , n75899 , n75900 );
nand ( n75902 , n75898 , n75901 );
nor ( n75903 , n75894 , n75902 );
not ( n75904 , n75903 );
or ( n75905 , n75891 , n75904 );
or ( n75906 , n75903 , n75890 );
nand ( n75907 , n75905 , n75906 );
nand ( n75908 , n75336 , n75907 );
and ( n75909 , n75393 , n68694 );
not ( n75910 , n73551 );
nor ( n75911 , n75909 , n75910 );
nand ( n75912 , n75868 , n75888 , n75908 , n75911 );
buf ( n75913 , n75912 );
buf ( n75914 , 1'b0 );
not ( n75915 , n68842 );
buf ( n75916 , n75915 );
buf ( n75917 , n68638 );
nand ( n75918 , n75277 , n68965 );
and ( n75919 , n75872 , n75676 );
not ( n75920 , n75919 );
and ( n75921 , n75876 , n75660 );
and ( n75922 , n75652 , n75323 , n75660 );
nor ( n75923 , n75921 , n75922 , n75674 );
not ( n75924 , n75923 );
or ( n75925 , n75920 , n75924 );
or ( n75926 , n75923 , n75919 );
nand ( n75927 , n75925 , n75926 );
nand ( n75928 , n75281 , n75927 );
and ( n75929 , n75892 , n75739 );
not ( n75930 , n75929 );
and ( n75931 , n75896 , n75723 );
and ( n75932 , n75715 , n75376 , n75723 );
nor ( n75933 , n75931 , n75932 , n75737 );
not ( n75934 , n75933 );
or ( n75935 , n75930 , n75934 );
or ( n75936 , n75933 , n75929 );
nand ( n75937 , n75935 , n75936 );
nand ( n75938 , n75336 , n75937 );
and ( n75939 , n75393 , n68699 );
not ( n75940 , n73575 );
nor ( n75941 , n75939 , n75940 );
nand ( n75942 , n75918 , n75928 , n75938 , n75941 );
buf ( n75943 , n75942 );
buf ( n75944 , 1'b0 );
not ( n75945 , n68842 );
buf ( n75946 , n75945 );
buf ( n75947 , n68638 );
nand ( n75948 , n75277 , n68951 );
not ( n75949 , n75658 );
nand ( n75950 , n75949 , n75673 );
not ( n75951 , n75950 );
or ( n75952 , n75650 , n75659 );
not ( n75953 , n75659 );
nand ( n75954 , n75953 , n75652 , n75323 );
nand ( n75955 , n75952 , n75954 , n75671 );
not ( n75956 , n75955 );
or ( n75957 , n75951 , n75956 );
or ( n75958 , n75955 , n75950 );
nand ( n75959 , n75957 , n75958 );
nand ( n75960 , n75281 , n75959 );
not ( n75961 , n75721 );
nand ( n75962 , n75961 , n75736 );
not ( n75963 , n75962 );
or ( n75964 , n75713 , n75722 );
not ( n75965 , n75722 );
nand ( n75966 , n75965 , n75715 , n75376 );
nand ( n75967 , n75964 , n75966 , n75734 );
not ( n75968 , n75967 );
or ( n75969 , n75963 , n75968 );
or ( n75970 , n75967 , n75962 );
nand ( n75971 , n75969 , n75970 );
nand ( n75972 , n75336 , n75971 );
and ( n75973 , n75393 , n68704 );
not ( n75974 , n73649 );
nor ( n75975 , n75973 , n75974 );
nand ( n75976 , n75948 , n75960 , n75972 , n75975 );
buf ( n75977 , n75976 );
buf ( n75978 , 1'b0 );
not ( n75979 , n68842 );
buf ( n75980 , n75979 );
buf ( n75981 , n68638 );
nand ( n75982 , n75277 , n68912 );
not ( n75983 , n75659 );
nand ( n75984 , n75983 , n75671 );
not ( n75985 , n75984 );
not ( n75986 , n75654 );
or ( n75987 , n75985 , n75986 );
or ( n75988 , n75654 , n75984 );
nand ( n75989 , n75987 , n75988 );
nand ( n75990 , n75281 , n75989 );
not ( n75991 , n75722 );
nand ( n75992 , n75991 , n75734 );
not ( n75993 , n75992 );
not ( n75994 , n75717 );
or ( n75995 , n75993 , n75994 );
or ( n75996 , n75717 , n75992 );
nand ( n75997 , n75995 , n75996 );
nand ( n75998 , n75336 , n75997 );
and ( n75999 , n75393 , n68709 );
not ( n76000 , n73674 );
nor ( n76001 , n75999 , n76000 );
nand ( n76002 , n75982 , n75990 , n75998 , n76001 );
buf ( n76003 , n76002 );
buf ( n76004 , 1'b0 );
not ( n76005 , n68842 );
buf ( n76006 , n76005 );
buf ( n76007 , n68638 );
nand ( n76008 , n75277 , n68981 );
not ( n76009 , n75648 );
nor ( n76010 , n76009 , n75641 );
not ( n76011 , n76010 );
and ( n76012 , n75323 , n75651 , n75639 );
not ( n76013 , n75639 );
not ( n76014 , n75644 );
or ( n76015 , n76013 , n76014 );
nand ( n76016 , n76015 , n75646 );
nor ( n76017 , n76012 , n76016 );
not ( n76018 , n76017 );
or ( n76019 , n76011 , n76018 );
or ( n76020 , n76017 , n76010 );
nand ( n76021 , n76019 , n76020 );
nand ( n76022 , n75281 , n76021 );
not ( n76023 , n75711 );
nor ( n76024 , n76023 , n75704 );
not ( n76025 , n76024 );
and ( n76026 , n75376 , n75714 , n75702 );
not ( n76027 , n75702 );
not ( n76028 , n75707 );
or ( n76029 , n76027 , n76028 );
nand ( n76030 , n76029 , n75709 );
nor ( n76031 , n76026 , n76030 );
not ( n76032 , n76031 );
or ( n76033 , n76025 , n76032 );
or ( n76034 , n76031 , n76024 );
nand ( n76035 , n76033 , n76034 );
nand ( n76036 , n75336 , n76035 );
and ( n76037 , n75393 , n68714 );
not ( n76038 , n73698 );
nor ( n76039 , n76037 , n76038 );
nand ( n76040 , n76008 , n76022 , n76036 , n76039 );
buf ( n76041 , n76040 );
buf ( n76042 , 1'b0 );
not ( n76043 , n68842 );
buf ( n76044 , n76043 );
buf ( n76045 , n68638 );
nand ( n76046 , n75277 , n69049 );
and ( n76047 , n75639 , n75646 );
not ( n76048 , n76047 );
and ( n76049 , n75323 , n75651 );
nor ( n76050 , n76049 , n75644 );
not ( n76051 , n76050 );
or ( n76052 , n76048 , n76051 );
or ( n76053 , n76050 , n76047 );
nand ( n76054 , n76052 , n76053 );
nand ( n76055 , n75281 , n76054 );
and ( n76056 , n75702 , n75709 );
not ( n76057 , n76056 );
and ( n76058 , n75376 , n75714 );
nor ( n76059 , n76058 , n75707 );
not ( n76060 , n76059 );
or ( n76061 , n76057 , n76060 );
or ( n76062 , n76059 , n76056 );
nand ( n76063 , n76061 , n76062 );
nand ( n76064 , n75336 , n76063 );
and ( n76065 , n75393 , n68719 );
not ( n76066 , n73723 );
nor ( n76067 , n76065 , n76066 );
nand ( n76068 , n76046 , n76055 , n76064 , n76067 );
buf ( n76069 , n76068 );
buf ( n76070 , 1'b0 );
not ( n76071 , n68842 );
buf ( n76072 , n76071 );
buf ( n76073 , n68638 );
nand ( n76074 , n75277 , n2728 );
xor ( n76075 , n3815 , n2728 );
nand ( n76076 , n75281 , n76075 );
xor ( n76077 , n69961 , n2728 );
nand ( n76078 , n75336 , n76077 );
and ( n76079 , n75393 , n68763 );
and ( n76080 , n69954 , n70863 );
nor ( n76081 , n76079 , n76080 );
nand ( n76082 , n76074 , n76076 , n76078 , n76081 );
buf ( n76083 , n76082 );
buf ( n76084 , 1'b0 );
not ( n76085 , n68842 );
buf ( n76086 , n76085 );
buf ( n9944 , n68638 );
not ( n76088 , n69127 );
or ( n76089 , n71996 , n76088 );
nand ( n76090 , n70863 , n2519 );
nand ( n76091 , n76089 , n76090 );
buf ( n76092 , n76091 );
buf ( n9950 , 1'b0 );
not ( n76094 , n68842 );
buf ( n9952 , n76094 );
buf ( n9953 , n68638 );
not ( n76097 , n68992 );
or ( n76098 , n71996 , n76097 );
not ( n76099 , n68663 );
or ( n76100 , n72075 , n76099 );
nand ( n76101 , n76098 , n76100 );
buf ( n76102 , n76101 );
buf ( n76103 , 1'b0 );
not ( n76104 , n68842 );
buf ( n76105 , n76104 );
buf ( n76106 , n68638 );
not ( n76107 , n69014 );
not ( n76108 , n70143 );
or ( n76109 , n76107 , n76108 );
nand ( n76110 , n70863 , n68664 );
nand ( n76111 , n76109 , n76110 );
buf ( n76112 , n76111 );
buf ( n76113 , 1'b0 );
not ( n76114 , n68842 );
buf ( n76115 , n76114 );
buf ( n76116 , n68638 );
not ( n76117 , n69063 );
not ( n76118 , n70143 );
or ( n76119 , n76117 , n76118 );
nand ( n76120 , n70863 , n68665 );
nand ( n76121 , n76119 , n76120 );
buf ( n9979 , n76121 );
buf ( n76123 , 1'b0 );
not ( n76124 , n68842 );
buf ( n76125 , n76124 );
buf ( n9983 , n68638 );
not ( n76127 , n69029 );
not ( n76128 , n70143 );
or ( n76129 , n76127 , n76128 );
nand ( n76130 , n70863 , n2523 );
nand ( n76131 , n76129 , n76130 );
buf ( n76132 , n76131 );
buf ( n76133 , 1'b0 );
not ( n76134 , n68842 );
buf ( n76135 , n76134 );
buf ( n76136 , n68638 );
not ( n76137 , n69087 );
not ( n76138 , n70143 );
or ( n76139 , n76137 , n76138 );
nand ( n76140 , n70863 , n2524 );
nand ( n76141 , n76139 , n76140 );
buf ( n76142 , n76141 );
buf ( n76143 , 1'b0 );
not ( n76144 , n68842 );
buf ( n76145 , n76144 );
buf ( n76146 , n68638 );
not ( n76147 , n69076 );
not ( n76148 , n70143 );
or ( n76149 , n76147 , n76148 );
nand ( n76150 , n70863 , n68668 );
nand ( n76151 , n76149 , n76150 );
buf ( n76152 , n76151 );
buf ( n10010 , 1'b0 );
not ( n76154 , n68842 );
buf ( n10012 , n76154 );
buf ( n76156 , n68638 );
not ( n76157 , n69234 );
or ( n76158 , n71996 , n76157 );
nand ( n76159 , n70863 , n68640 );
nand ( n76160 , n76158 , n76159 );
buf ( n10018 , n76160 );
buf ( n10019 , 1'b0 );
not ( n76163 , n68842 );
buf ( n76164 , n76163 );
buf ( n76165 , n68638 );
not ( n76166 , n69404 );
or ( n76167 , n76166 , n71996 );
nand ( n76168 , n70863 , n2498 );
nand ( n76169 , n76167 , n76168 );
buf ( n76170 , n76169 );
buf ( n76171 , 1'b0 );
not ( n76172 , n68842 );
buf ( n76173 , n76172 );
buf ( n76174 , n68638 );
not ( n76175 , n69099 );
not ( n76176 , n70143 );
or ( n76177 , n76175 , n76176 );
nand ( n76178 , n70863 , n68669 );
nand ( n76179 , n76177 , n76178 );
buf ( n76180 , n76179 );
buf ( n76181 , 1'b0 );
not ( n76182 , n68842 );
buf ( n76183 , n76182 );
buf ( n76184 , n68638 );
not ( n76185 , n69413 );
or ( n76186 , n71996 , n76185 );
nand ( n76187 , n70863 , n2499 );
nand ( n76188 , n76186 , n76187 );
buf ( n76189 , n76188 );
buf ( n76190 , 1'b0 );
not ( n76191 , n68842 );
buf ( n10049 , n76191 );
buf ( n10050 , n68638 );
not ( n76194 , n69356 );
or ( n76195 , n71996 , n76194 );
not ( n76196 , n2500 );
or ( n76197 , n72075 , n76196 );
nand ( n76198 , n76195 , n76197 );
buf ( n76199 , n76198 );
buf ( n76200 , 1'b0 );
not ( n76201 , n68842 );
buf ( n10059 , n76201 );
buf ( n10060 , n68638 );
not ( n76204 , n69342 );
or ( n76205 , n71996 , n76204 );
not ( n76206 , n2501 );
or ( n76207 , n72075 , n76206 );
nand ( n76208 , n76205 , n76207 );
buf ( n76209 , n76208 );
buf ( n10067 , 1'b0 );
not ( n76211 , n68842 );
buf ( n10069 , n76211 );
buf ( n10070 , n68638 );
not ( n76214 , n69328 );
or ( n76215 , n71996 , n76214 );
not ( n76216 , n2502 );
or ( n76217 , n72075 , n76216 );
nand ( n76218 , n76215 , n76217 );
buf ( n10076 , n76218 );
buf ( n76220 , 1'b0 );
not ( n76221 , n68842 );
buf ( n76222 , n76221 );
buf ( n76223 , n68638 );
not ( n76224 , n69302 );
not ( n76225 , n70143 );
or ( n76226 , n76224 , n76225 );
nand ( n76227 , n70863 , n2503 );
nand ( n76228 , n76226 , n76227 );
buf ( n76229 , n76228 );
buf ( n76230 , 1'b0 );
not ( n76231 , n68842 );
buf ( n10089 , n76231 );
buf ( n10090 , n68638 );
not ( n76234 , n69315 );
or ( n76235 , n71996 , n76234 );
not ( n76236 , n2504 );
or ( n76237 , n72075 , n76236 );
nand ( n76238 , n76235 , n76237 );
buf ( n10096 , n76238 );
buf ( n76240 , 1'b0 );
not ( n76241 , n68842 );
buf ( n76242 , n76241 );
buf ( n10100 , n68638 );
not ( n76244 , n69293 );
not ( n76245 , n70143 );
or ( n76246 , n76244 , n76245 );
nand ( n76247 , n70863 , n68648 );
nand ( n76248 , n76246 , n76247 );
buf ( n76249 , n76248 );
buf ( n76250 , 1'b0 );
not ( n76251 , n68842 );
buf ( n76252 , n76251 );
buf ( n76253 , n68638 );
not ( n76254 , n69281 );
or ( n76255 , n71996 , n76254 );
not ( n76256 , n68649 );
or ( n76257 , n72075 , n76256 );
nand ( n76258 , n76255 , n76257 );
buf ( n76259 , n76258 );
buf ( n76260 , 1'b0 );
not ( n76261 , n68842 );
buf ( n10119 , n76261 );
buf ( n10120 , n68638 );
not ( n76264 , n69269 );
or ( n76265 , n71996 , n76264 );
not ( n76266 , n68650 );
or ( n76267 , n72075 , n76266 );
nand ( n76268 , n76265 , n76267 );
buf ( n10126 , n76268 );
buf ( n10127 , 1'b0 );
not ( n76271 , n68842 );
buf ( n10129 , n76271 );
buf ( n10130 , n68638 );
not ( n76274 , n69260 );
or ( n76275 , n71996 , n76274 );
not ( n76276 , n2508 );
or ( n76277 , n72075 , n76276 );
nand ( n76278 , n76275 , n76277 );
buf ( n76279 , n76278 );
buf ( n10137 , 1'b0 );
not ( n76281 , n68842 );
buf ( n10139 , n76281 );
buf ( n76283 , n68638 );
not ( n76284 , n69110 );
not ( n76285 , n70143 );
or ( n76286 , n76284 , n76285 );
nand ( n76287 , n70863 , n68670 );
nand ( n76288 , n76286 , n76287 );
buf ( n76289 , n76288 );
buf ( n76290 , 1'b0 );
not ( n76291 , n68842 );
buf ( n76292 , n76291 );
buf ( n76293 , n68638 );
not ( n76294 , n69244 );
or ( n76295 , n71996 , n76294 );
not ( n76296 , n2509 );
or ( n76297 , n72075 , n76296 );
nand ( n76298 , n76295 , n76297 );
buf ( n10156 , n76298 );
buf ( n10157 , 1'b0 );
not ( n76301 , n68842 );
buf ( n76302 , n76301 );
buf ( n76303 , n68638 );
not ( n76304 , n68653 );
not ( n76305 , n70863 );
or ( n76306 , n76304 , n76305 );
not ( n76307 , n69161 );
or ( n76308 , n71996 , n76307 );
nand ( n76309 , n76306 , n76308 );
buf ( n76310 , n76309 );
buf ( n76311 , 1'b0 );
not ( n76312 , n68842 );
buf ( n76313 , n76312 );
buf ( n76314 , n68638 );
not ( n76315 , n69180 );
or ( n76316 , n71996 , n76315 );
not ( n76317 , n68654 );
or ( n76318 , n72075 , n76317 );
nand ( n76319 , n76316 , n76318 );
buf ( n76320 , n76319 );
buf ( n76321 , 1'b0 );
not ( n76322 , n68842 );
buf ( n76323 , n76322 );
buf ( n76324 , n68638 );
not ( n76325 , n69191 );
not ( n76326 , n70143 );
or ( n76327 , n76325 , n76326 );
nand ( n76328 , n70863 , n68655 );
nand ( n76329 , n76327 , n76328 );
buf ( n76330 , n76329 );
buf ( n76331 , 1'b0 );
not ( n76332 , n68842 );
buf ( n10190 , n76332 );
buf ( n10191 , n68638 );
not ( n76335 , n68938 );
or ( n76336 , n76335 , n71996 );
nand ( n76337 , n70863 , n2513 );
nand ( n76338 , n76336 , n76337 );
buf ( n10196 , n76338 );
buf ( n10197 , 1'b0 );
not ( n76341 , n68842 );
buf ( n10199 , n76341 );
buf ( n76343 , n68638 );
not ( n76344 , n68965 );
or ( n76345 , n71996 , n76344 );
nand ( n76346 , n70863 , n2514 );
nand ( n76347 , n76345 , n76346 );
buf ( n76348 , n76347 );
buf ( n76349 , 1'b0 );
not ( n76350 , n68842 );
buf ( n76351 , n76350 );
buf ( n76352 , n68638 );
not ( n76353 , n68951 );
or ( n76354 , n71996 , n76353 );
nand ( n76355 , n70863 , n2515 );
nand ( n76356 , n76354 , n76355 );
buf ( n76357 , n76356 );
buf ( n76358 , 1'b0 );
not ( n76359 , n68842 );
buf ( n76360 , n76359 );
buf ( n76361 , n68638 );
not ( n76362 , n68912 );
or ( n76363 , n71996 , n76362 );
nand ( n76364 , n70863 , n2516 );
nand ( n76365 , n76363 , n76364 );
buf ( n76366 , n76365 );
buf ( n10224 , 1'b0 );
not ( n76368 , n68842 );
buf ( n10226 , n76368 );
buf ( n76370 , n68638 );
not ( n76371 , n68981 );
or ( n76372 , n71996 , n76371 );
nand ( n76373 , n70863 , n2517 );
nand ( n76374 , n76372 , n76373 );
buf ( n10232 , n76374 );
buf ( n10233 , 1'b0 );
not ( n76377 , n68842 );
buf ( n76378 , n76377 );
buf ( n76379 , n68638 );
not ( n76380 , n69049 );
or ( n76381 , n71996 , n76380 );
nand ( n76382 , n70863 , n2518 );
nand ( n76383 , n76381 , n76382 );
buf ( n76384 , n76383 );
buf ( n76385 , 1'b0 );
not ( n76386 , n68842 );
buf ( n76387 , n76386 );
buf ( n76388 , n68638 );
not ( n76389 , n2728 );
not ( n76390 , n70143 );
or ( n76391 , n76389 , n76390 );
nand ( n76392 , n70863 , n2528 );
nand ( n76393 , n76391 , n76392 );
buf ( n76394 , n76393 );
buf ( n76395 , 1'b0 );
not ( n76396 , n68842 );
buf ( n76397 , n76396 );
buf ( n76398 , n68638 );
not ( n76399 , n69623 );
not ( n76400 , n76399 );
not ( n76401 , n69951 );
nand ( n76402 , n76401 , n73906 );
not ( n76403 , n76402 );
or ( n76404 , n76400 , n76403 );
not ( n76405 , n76402 );
not ( n76406 , n76405 );
and ( n76407 , n69557 , n69547 );
and ( n76408 , n76407 , n69535 , n69523 );
nand ( n76409 , n69474 , n69455 , n69439 , n69475 );
nand ( n76410 , n69491 , n69506 );
nor ( n76411 , n76409 , n76410 );
nand ( n76412 , n76408 , n76411 );
not ( n76413 , n76412 );
and ( n76414 , n69591 , n69580 );
and ( n76415 , n76414 , n69603 );
nand ( n76416 , n76413 , n76415 );
not ( n76417 , n69617 );
xor ( n76418 , n76416 , n76417 );
not ( n76419 , n76418 );
or ( n76420 , n76406 , n76419 );
nand ( n76421 , n76404 , n76420 );
not ( n76422 , n70242 );
nor ( n76423 , n76421 , n76422 );
not ( n76424 , n69603 );
nand ( n76425 , n76408 , n76411 , n76414 );
not ( n76426 , n76425 );
or ( n76427 , n76424 , n76426 );
or ( n76428 , n76425 , n69603 );
nand ( n76429 , n76427 , n76428 );
not ( n76430 , n76429 );
or ( n76431 , n76402 , n76430 );
nand ( n76432 , n76402 , n69985 );
nand ( n76433 , n76431 , n76432 );
not ( n76434 , n70331 );
nor ( n76435 , n76433 , n76434 );
nor ( n76436 , n76423 , n76435 );
not ( n76437 , n70300 );
and ( n76438 , n76407 , n69535 , n69523 );
nand ( n76439 , n76438 , n76411 , n69591 );
xnor ( n76440 , n76439 , n69580 );
not ( n76441 , n76440 );
or ( n76442 , n76402 , n76441 );
nand ( n76443 , n76402 , n70102 );
nand ( n76444 , n76442 , n76443 );
nor ( n76445 , n76437 , n76444 );
not ( n76446 , n70312 );
not ( n76447 , n69994 );
not ( n76448 , n76402 );
not ( n76449 , n76448 );
not ( n76450 , n76449 );
or ( n76451 , n76447 , n76450 );
not ( n76452 , n69591 );
not ( n76453 , n76412 );
or ( n76454 , n76452 , n76453 );
or ( n76455 , n76412 , n69591 );
nand ( n76456 , n76454 , n76455 );
not ( n76457 , n76456 );
or ( n76458 , n76402 , n76457 );
nand ( n76459 , n76451 , n76458 );
nor ( n76460 , n76446 , n76459 );
nor ( n76461 , n76445 , n76460 );
and ( n76462 , n76436 , n76461 );
not ( n76463 , n70382 );
not ( n76464 , n76463 );
not ( n76465 , n70086 );
not ( n76466 , n76402 );
or ( n76467 , n76465 , n76466 );
not ( n76468 , n76405 );
xor ( n76469 , n69557 , n76411 );
not ( n76470 , n76469 );
or ( n76471 , n76468 , n76470 );
nand ( n76472 , n76467 , n76471 );
not ( n76473 , n76472 );
or ( n76474 , n76464 , n76473 );
not ( n76475 , n70267 );
not ( n76476 , n69547 );
nand ( n76477 , n76411 , n69557 );
not ( n76478 , n76477 );
or ( n76479 , n76476 , n76478 );
or ( n76480 , n76477 , n69547 );
nand ( n76481 , n76479 , n76480 );
not ( n76482 , n76481 );
or ( n76483 , n76402 , n76482 );
nand ( n76484 , n76402 , n70011 );
nand ( n76485 , n76483 , n76484 );
nand ( n76486 , n76475 , n76485 );
nand ( n76487 , n76474 , n76486 );
not ( n76488 , n76485 );
nand ( n76489 , n76488 , n70267 );
nand ( n76490 , n76487 , n76489 );
not ( n76491 , n70257 );
not ( n76492 , n70017 );
not ( n76493 , n76402 );
or ( n76494 , n76492 , n76493 );
not ( n76495 , n69535 );
nand ( n76496 , n76411 , n76407 );
not ( n76497 , n76496 );
or ( n76498 , n76495 , n76497 );
or ( n76499 , n76496 , n69535 );
nand ( n76500 , n76498 , n76499 );
not ( n76501 , n76500 );
or ( n76502 , n76406 , n76501 );
nand ( n76503 , n76494 , n76502 );
not ( n76504 , n76503 );
not ( n76505 , n76504 );
or ( n76506 , n76491 , n76505 );
not ( n76507 , n69523 );
nand ( n76508 , n76411 , n76407 , n69535 );
not ( n76509 , n76508 );
or ( n76510 , n76507 , n76509 );
or ( n76511 , n76508 , n69523 );
nand ( n76512 , n76510 , n76511 );
not ( n76513 , n76512 );
or ( n76514 , n76402 , n76513 );
not ( n76515 , n76402 );
not ( n76516 , n76515 );
not ( n76517 , n71533 );
nand ( n76518 , n76516 , n76517 );
nand ( n76519 , n76514 , n76518 );
not ( n76520 , n70277 );
nor ( n76521 , n76519 , n76520 );
not ( n76522 , n76521 );
nand ( n76523 , n76506 , n76522 );
or ( n76524 , n76490 , n76523 );
not ( n76525 , n70257 );
nand ( n76526 , n76525 , n76503 );
or ( n76527 , n76521 , n76526 );
not ( n76528 , n76519 );
or ( n76529 , n76528 , n70277 );
nand ( n76530 , n76527 , n76529 );
not ( n76531 , n76530 );
nand ( n76532 , n76524 , n76531 );
and ( n76533 , n76462 , n76532 );
not ( n76534 , n76436 );
not ( n76535 , n70312 );
nand ( n76536 , n76535 , n76459 );
or ( n76537 , n76445 , n76536 );
not ( n76538 , n76444 );
or ( n76539 , n76538 , n70300 );
nand ( n76540 , n76537 , n76539 );
not ( n76541 , n76540 );
or ( n76542 , n76534 , n76541 );
not ( n76543 , n76423 );
nand ( n76544 , n76433 , n76434 );
not ( n76545 , n76544 );
and ( n76546 , n76543 , n76545 );
and ( n76547 , n76421 , n76422 );
nor ( n76548 , n76546 , n76547 );
nand ( n76549 , n76542 , n76548 );
nor ( n76550 , n76533 , n76549 );
not ( n76551 , n70382 );
not ( n76552 , n76472 );
not ( n76553 , n76552 );
or ( n76554 , n76551 , n76553 );
nand ( n76555 , n76554 , n76489 );
nor ( n76556 , n76555 , n76523 );
not ( n76557 , n70028 );
not ( n76558 , n76402 );
or ( n76559 , n76557 , n76558 );
not ( n76560 , n76402 );
not ( n76561 , n69506 );
nand ( n76562 , n69455 , n69475 );
not ( n76563 , n76562 );
nand ( n76564 , n76563 , n69491 );
not ( n76565 , n76564 );
or ( n76566 , n76561 , n76565 );
or ( n76567 , n76564 , n69506 );
nand ( n76568 , n76566 , n76567 );
nand ( n76569 , n76560 , n76568 );
nand ( n76570 , n76559 , n76569 );
not ( n76571 , n70436 );
nor ( n76572 , n76570 , n76571 );
not ( n76573 , n72306 );
not ( n76574 , n69491 );
not ( n76575 , n76562 );
or ( n76576 , n76574 , n76575 );
or ( n76577 , n76562 , n69491 );
nand ( n76578 , n76576 , n76577 );
not ( n76579 , n76578 );
or ( n76580 , n76402 , n76579 );
nand ( n76581 , n76516 , n70042 );
nand ( n76582 , n76580 , n76581 );
nor ( n76583 , n76573 , n76582 );
nor ( n76584 , n76572 , n76583 );
not ( n76585 , n69474 );
not ( n76586 , n76410 );
nand ( n76587 , n76586 , n76563 , n69439 );
not ( n76588 , n76587 );
or ( n76589 , n76585 , n76588 );
or ( n76590 , n76587 , n69474 );
nand ( n76591 , n76589 , n76590 );
not ( n76592 , n76591 );
or ( n76593 , n76402 , n76592 );
nand ( n76594 , n76516 , n70094 );
nand ( n76595 , n76593 , n76594 );
not ( n76596 , n70392 );
nor ( n76597 , n76595 , n76596 );
not ( n76598 , n70035 );
not ( n76599 , n76402 );
or ( n76600 , n76598 , n76599 );
not ( n76601 , n76448 );
not ( n76602 , n69439 );
or ( n76603 , n76562 , n76410 );
not ( n76604 , n76603 );
or ( n76605 , n76602 , n76604 );
or ( n76606 , n76603 , n69439 );
nand ( n76607 , n76605 , n76606 );
not ( n76608 , n76607 );
or ( n76609 , n76601 , n76608 );
nand ( n76610 , n76600 , n76609 );
not ( n76611 , n70481 );
nor ( n76612 , n76610 , n76611 );
nor ( n76613 , n76597 , n76612 );
not ( n76614 , n70424 );
not ( n76615 , n76614 );
not ( n76616 , n69455 );
not ( n76617 , n69475 );
and ( n76618 , n76616 , n76617 );
nor ( n76619 , n76618 , n76563 );
not ( n76620 , n76619 );
or ( n76621 , n76402 , n76620 );
nand ( n76622 , n76516 , n70044 );
nand ( n76623 , n76621 , n76622 );
not ( n76624 , n76623 );
or ( n76625 , n76615 , n76624 );
or ( n76626 , n76623 , n76614 );
not ( n76627 , n70057 );
nand ( n76628 , n76627 , n70507 );
not ( n76629 , n69971 );
nand ( n76630 , n76629 , n70526 );
and ( n76631 , n76628 , n76630 );
not ( n76632 , n70507 );
and ( n76633 , n70057 , n76632 );
nor ( n76634 , n76631 , n76633 );
not ( n76635 , n70077 );
and ( n76636 , n76635 , n70463 );
or ( n76637 , n76634 , n76636 );
or ( n76638 , n76635 , n70463 );
nand ( n76639 , n76637 , n76638 );
nand ( n76640 , n76626 , n76639 );
nand ( n76641 , n76625 , n76640 );
nand ( n76642 , n76584 , n76613 , n76641 );
not ( n76643 , n72306 );
nand ( n76644 , n76643 , n76582 );
not ( n76645 , n70436 );
nand ( n76646 , n76645 , n76570 );
and ( n76647 , n76644 , n76646 );
nor ( n76648 , n76647 , n76572 );
nand ( n76649 , n76648 , n76613 );
nand ( n76650 , n76610 , n76611 );
nor ( n76651 , n76597 , n76650 );
and ( n76652 , n76595 , n76596 );
nor ( n76653 , n76651 , n76652 );
nand ( n76654 , n76642 , n76649 , n76653 );
nand ( n76655 , n76556 , n76462 , n76654 );
nand ( n76656 , n76550 , n76655 );
and ( n76657 , n69603 , n69617 );
nand ( n76658 , n76414 , n76657 );
nor ( n76659 , n76412 , n76658 );
nand ( n76660 , n69659 , n69645 );
nand ( n76661 , n69900 , n69773 );
nor ( n76662 , n76660 , n76661 );
and ( n76663 , n69826 , n69875 , n69808 , n69796 );
nand ( n76664 , n76662 , n76663 );
nand ( n76665 , n69936 , n69854 );
nand ( n76666 , n69689 , n69710 );
nor ( n76667 , n76665 , n76666 );
not ( n76668 , n72632 );
nand ( n76669 , n76667 , n76668 );
nor ( n76670 , n76664 , n76669 );
nand ( n76671 , n76659 , n76670 );
not ( n76672 , n69747 );
and ( n76673 , n76671 , n76672 );
not ( n76674 , n76671 );
and ( n76675 , n76674 , n69747 );
nor ( n76676 , n76673 , n76675 );
not ( n76677 , n76676 );
or ( n76678 , n76449 , n76677 );
nand ( n76679 , n76402 , n72467 );
nand ( n76680 , n76678 , n76679 );
not ( n76681 , n76680 );
nand ( n76682 , n76681 , n73920 );
not ( n76683 , n76667 );
nand ( n76684 , n76662 , n76663 );
nor ( n76685 , n76683 , n76684 );
nand ( n76686 , n76659 , n76685 );
not ( n76687 , n76668 );
and ( n76688 , n76686 , n76687 );
not ( n76689 , n76686 );
and ( n76690 , n76689 , n76668 );
nor ( n76691 , n76688 , n76690 );
not ( n76692 , n76691 );
or ( n76693 , n76402 , n76692 );
nand ( n76694 , n76516 , n72456 );
nand ( n76695 , n76693 , n76694 );
not ( n76696 , n76695 );
nand ( n76697 , n76696 , n72630 );
nand ( n76698 , n76682 , n76697 );
not ( n76699 , n73918 );
nand ( n76700 , n76668 , n69747 );
not ( n76701 , n76700 );
nand ( n76702 , n76701 , n76667 );
nor ( n76703 , n76684 , n76702 );
nand ( n76704 , n76659 , n76703 );
and ( n76705 , n76704 , n69912 );
not ( n76706 , n76704 );
not ( n76707 , n69912 );
and ( n76708 , n76706 , n76707 );
nor ( n76709 , n76705 , n76708 );
not ( n76710 , n76709 );
or ( n76711 , n76402 , n76710 );
nand ( n76712 , n76402 , n73906 );
nand ( n76713 , n76711 , n76712 );
not ( n76714 , n76713 );
not ( n76715 , n76714 );
or ( n76716 , n76699 , n76715 );
nor ( n76717 , n76700 , n69912 );
nand ( n76718 , n76667 , n76717 );
nor ( n76719 , n76684 , n76718 );
nand ( n76720 , n76659 , n76719 );
not ( n76721 , n69946 );
and ( n76722 , n76721 , n76707 );
not ( n76723 , n76721 );
and ( n76724 , n76723 , n69912 );
nor ( n76725 , n76722 , n76724 );
xor ( n76726 , n76720 , n76725 );
not ( n76727 , n76726 );
not ( n76728 , n76402 );
not ( n76729 , n76728 );
or ( n76730 , n76727 , n76729 );
not ( n76731 , n69951 );
nand ( n76732 , n76730 , n76731 );
not ( n76733 , n73916 );
nand ( n76734 , n76732 , n76733 );
nand ( n76735 , n76716 , n76734 );
nor ( n76736 , n76698 , n76735 );
not ( n76737 , n76665 );
nand ( n76738 , n76737 , n69689 );
nor ( n76739 , n76664 , n76738 );
nand ( n76740 , n76659 , n76739 );
not ( n76741 , n69710 );
and ( n76742 , n76740 , n76741 );
not ( n76743 , n76740 );
and ( n76744 , n76743 , n69710 );
nor ( n76745 , n76742 , n76744 );
not ( n76746 , n76745 );
or ( n76747 , n76601 , n76746 );
nand ( n76748 , n76402 , n71767 );
nand ( n76749 , n76747 , n76748 );
not ( n76750 , n72819 );
nor ( n76751 , n76749 , n76750 );
not ( n76752 , n71783 );
not ( n76753 , n76752 );
not ( n76754 , n76516 );
or ( n76755 , n76753 , n76754 );
nor ( n76756 , n76664 , n76665 );
nand ( n76757 , n76659 , n76756 );
not ( n76758 , n69689 );
and ( n76759 , n76757 , n76758 );
not ( n76760 , n76757 );
and ( n76761 , n76760 , n69689 );
nor ( n76762 , n76759 , n76761 );
not ( n76763 , n76762 );
or ( n76764 , n76601 , n76763 );
nand ( n76765 , n76755 , n76764 );
not ( n76766 , n72538 );
nor ( n76767 , n76765 , n76766 );
nor ( n76768 , n76751 , n76767 );
not ( n76769 , n76768 );
not ( n76770 , n72561 );
not ( n76771 , n76684 );
nand ( n76772 , n76771 , n76659 );
not ( n76773 , n69936 );
and ( n76774 , n76772 , n76773 );
not ( n76775 , n76772 );
and ( n76776 , n76775 , n69936 );
nor ( n76777 , n76774 , n76776 );
not ( n76778 , n76777 );
or ( n76779 , n76402 , n76778 );
nand ( n76780 , n76402 , n71818 );
nand ( n76781 , n76779 , n76780 );
not ( n76782 , n76781 );
not ( n76783 , n76782 );
or ( n76784 , n76770 , n76783 );
not ( n76785 , n71802 );
not ( n76786 , n76785 );
not ( n76787 , n76402 );
or ( n76788 , n76786 , n76787 );
nor ( n76789 , n76664 , n76773 );
nand ( n76790 , n76659 , n76789 );
not ( n76791 , n69854 );
and ( n76792 , n76790 , n76791 );
not ( n76793 , n76790 );
and ( n76794 , n76793 , n69854 );
nor ( n76795 , n76792 , n76794 );
not ( n76796 , n76795 );
or ( n76797 , n76402 , n76796 );
nand ( n76798 , n76788 , n76797 );
not ( n76799 , n72548 );
nor ( n76800 , n76798 , n76799 );
not ( n76801 , n76800 );
nand ( n76802 , n76784 , n76801 );
nor ( n76803 , n76769 , n76802 );
nand ( n76804 , n76736 , n76803 );
nand ( n76805 , n69808 , n69826 );
nor ( n76806 , n76660 , n76805 );
nand ( n76807 , n69900 , n69875 );
not ( n76808 , n69796 );
nor ( n76809 , n76807 , n76808 );
and ( n76810 , n76806 , n76809 );
nand ( n76811 , n76659 , n76810 );
not ( n76812 , n69773 );
and ( n76813 , n76811 , n76812 );
not ( n76814 , n76811 );
and ( n76815 , n76814 , n69773 );
nor ( n76816 , n76813 , n76815 );
not ( n76817 , n76816 );
or ( n76818 , n76601 , n76817 );
not ( n76819 , n71837 );
nand ( n76820 , n76402 , n76819 );
nand ( n76821 , n76818 , n76820 );
not ( n76822 , n72514 );
nor ( n76823 , n76821 , n76822 );
not ( n76824 , n72503 );
not ( n76825 , n71856 );
not ( n76826 , n76449 );
or ( n76827 , n76825 , n76826 );
not ( n76828 , n76807 );
and ( n76829 , n76806 , n76828 );
nand ( n76830 , n76659 , n76829 );
and ( n76831 , n76830 , n76808 );
not ( n76832 , n76830 );
and ( n76833 , n76832 , n69796 );
nor ( n76834 , n76831 , n76833 );
not ( n76835 , n76834 );
or ( n76836 , n76402 , n76835 );
nand ( n76837 , n76827 , n76836 );
nor ( n76838 , n76824 , n76837 );
nor ( n76839 , n76823 , n76838 );
not ( n76840 , n71873 );
not ( n76841 , n76402 );
or ( n76842 , n76840 , n76841 );
and ( n76843 , n76806 , n69875 );
nand ( n76844 , n76659 , n76843 );
not ( n76845 , n69900 );
and ( n76846 , n76844 , n76845 );
not ( n76847 , n76844 );
and ( n76848 , n76847 , n69900 );
nor ( n76849 , n76846 , n76848 );
not ( n76850 , n76849 );
or ( n76851 , n76468 , n76850 );
nand ( n76852 , n76842 , n76851 );
not ( n76853 , n72479 );
nor ( n76854 , n76852 , n76853 );
not ( n76855 , n71041 );
not ( n76856 , n76402 );
or ( n76857 , n76855 , n76856 );
nand ( n76858 , n76659 , n76806 );
not ( n76859 , n69875 );
and ( n76860 , n76858 , n76859 );
not ( n76861 , n76858 );
and ( n76862 , n76861 , n69875 );
nor ( n76863 , n76860 , n76862 );
not ( n76864 , n76863 );
or ( n76865 , n76406 , n76864 );
nand ( n76866 , n76857 , n76865 );
not ( n76867 , n72489 );
nor ( n76868 , n76866 , n76867 );
nor ( n76869 , n76854 , n76868 );
and ( n76870 , n76839 , n76869 );
not ( n76871 , n70229 );
not ( n76872 , n69981 );
not ( n76873 , n76402 );
or ( n76874 , n76872 , n76873 );
xor ( n76875 , n69645 , n76659 );
not ( n76876 , n76875 );
or ( n76877 , n76402 , n76876 );
nand ( n76878 , n76874 , n76877 );
not ( n76879 , n76878 );
not ( n76880 , n76879 );
or ( n76881 , n76871 , n76880 );
nand ( n76882 , n76659 , n69645 );
not ( n76883 , n69659 );
and ( n76884 , n76882 , n76883 );
not ( n76885 , n76882 );
and ( n76886 , n76885 , n69659 );
nor ( n76887 , n76884 , n76886 );
not ( n76888 , n76887 );
or ( n76889 , n76402 , n76888 );
nand ( n76890 , n76449 , n69664 );
nand ( n76891 , n76889 , n76890 );
not ( n76892 , n76891 );
nand ( n76893 , n76892 , n71078 );
nand ( n76894 , n76881 , n76893 );
not ( n76895 , n71096 );
not ( n76896 , n71051 );
not ( n76897 , n76402 );
or ( n76898 , n76896 , n76897 );
not ( n76899 , n76660 );
nand ( n76900 , n76899 , n76659 );
not ( n76901 , n69826 );
and ( n76902 , n76900 , n76901 );
not ( n76903 , n76900 );
and ( n76904 , n76903 , n69826 );
nor ( n76905 , n76902 , n76904 );
not ( n76906 , n76905 );
or ( n76907 , n76406 , n76906 );
nand ( n76908 , n76898 , n76907 );
not ( n76909 , n76908 );
not ( n76910 , n76909 );
or ( n76911 , n76895 , n76910 );
nor ( n76912 , n76660 , n76901 );
nand ( n76913 , n76659 , n76912 );
xnor ( n76914 , n76913 , n69808 );
not ( n76915 , n76914 );
not ( n76916 , n76405 );
or ( n76917 , n76915 , n76916 );
not ( n76918 , n76402 );
not ( n76919 , n71062 );
or ( n76920 , n76918 , n76919 );
nand ( n76921 , n76917 , n76920 );
not ( n76922 , n71126 );
nor ( n76923 , n76921 , n76922 );
not ( n76924 , n76923 );
nand ( n76925 , n76911 , n76924 );
nor ( n76926 , n76894 , n76925 );
nand ( n76927 , n76870 , n76926 );
nor ( n76928 , n76804 , n76927 );
and ( n76929 , n76656 , n76928 );
not ( n76930 , n71078 );
nand ( n76931 , n76930 , n76891 );
not ( n76932 , n76931 );
not ( n76933 , n70229 );
nand ( n76934 , n76933 , n76878 );
not ( n76935 , n76934 );
or ( n76936 , n76932 , n76935 );
nand ( n76937 , n76936 , n76893 );
or ( n76938 , n76925 , n76937 );
not ( n76939 , n71096 );
nand ( n76940 , n76939 , n76908 );
or ( n76941 , n76923 , n76940 );
nand ( n76942 , n76921 , n76922 );
nand ( n76943 , n76941 , n76942 );
not ( n76944 , n76943 );
nand ( n76945 , n76938 , n76944 );
and ( n76946 , n76870 , n76945 );
not ( n76947 , n76839 );
nand ( n76948 , n76866 , n76867 );
or ( n76949 , n76854 , n76948 );
nand ( n76950 , n76852 , n76853 );
nand ( n76951 , n76949 , n76950 );
not ( n76952 , n76951 );
or ( n76953 , n76947 , n76952 );
not ( n76954 , n76823 );
not ( n76955 , n72503 );
nand ( n76956 , n76955 , n76837 );
not ( n76957 , n76956 );
and ( n76958 , n76954 , n76957 );
and ( n76959 , n76821 , n76822 );
nor ( n76960 , n76958 , n76959 );
nand ( n76961 , n76953 , n76960 );
nor ( n76962 , n76946 , n76961 );
or ( n76963 , n76962 , n76804 );
not ( n76964 , n76768 );
not ( n76965 , n72561 );
nand ( n76966 , n76965 , n76781 );
or ( n76967 , n76800 , n76966 );
nand ( n76968 , n76798 , n76799 );
nand ( n76969 , n76967 , n76968 );
not ( n76970 , n76969 );
or ( n76971 , n76964 , n76970 );
not ( n76972 , n76751 );
nand ( n76973 , n76765 , n76766 );
not ( n76974 , n76973 );
and ( n76975 , n76972 , n76974 );
and ( n76976 , n76749 , n76750 );
nor ( n76977 , n76975 , n76976 );
nand ( n76978 , n76971 , n76977 );
and ( n76979 , n76978 , n76736 );
not ( n76980 , n76695 );
nor ( n76981 , n76980 , n72630 );
and ( n76982 , n76682 , n76981 );
not ( n76983 , n76680 );
nor ( n76984 , n76983 , n73920 );
nor ( n76985 , n76982 , n76984 );
or ( n76986 , n76985 , n76735 );
nor ( n76987 , n76714 , n73918 );
and ( n76988 , n76987 , n76734 );
nor ( n76989 , n76732 , n76733 );
nor ( n76990 , n76988 , n76989 );
nand ( n76991 , n76986 , n76990 );
nor ( n76992 , n76979 , n76991 );
nand ( n76993 , n76963 , n76992 );
nor ( n76994 , n76929 , n76993 );
not ( n76995 , n76994 );
not ( n76996 , n72503 );
not ( n76997 , n76996 );
not ( n76998 , n71856 );
or ( n76999 , n76997 , n76998 );
not ( n77000 , n72514 );
nand ( n77001 , n76819 , n77000 );
nand ( n77002 , n76999 , n77001 );
not ( n77003 , n72489 );
not ( n77004 , n77003 );
not ( n77005 , n71041 );
or ( n77006 , n77004 , n77005 );
not ( n77007 , n72479 );
nand ( n77008 , n71873 , n77007 );
nand ( n77009 , n77006 , n77008 );
nor ( n77010 , n77002 , n77009 );
not ( n77011 , n71096 );
not ( n77012 , n77011 );
not ( n77013 , n71051 );
or ( n77014 , n77012 , n77013 );
not ( n77015 , n71126 );
nand ( n77016 , n71062 , n77015 );
nand ( n77017 , n77014 , n77016 );
not ( n77018 , n71078 );
not ( n77019 , n69664 );
not ( n77020 , n77019 );
or ( n77021 , n77018 , n77020 );
not ( n77022 , n69981 );
nand ( n77023 , n77022 , n70229 );
nand ( n77024 , n77021 , n77023 );
not ( n77025 , n71078 );
nand ( n77026 , n77025 , n69664 );
nand ( n77027 , n77024 , n77026 );
or ( n77028 , n77017 , n77027 );
nor ( n77029 , n71051 , n77011 );
and ( n77030 , n77016 , n77029 );
nor ( n77031 , n71062 , n77015 );
nor ( n77032 , n77030 , n77031 );
nand ( n77033 , n77028 , n77032 );
and ( n77034 , n77010 , n77033 );
nor ( n77035 , n71041 , n77003 );
and ( n77036 , n77008 , n77035 );
nor ( n77037 , n71873 , n77007 );
nor ( n77038 , n77036 , n77037 );
or ( n77039 , n77038 , n77002 );
nor ( n77040 , n71856 , n76996 );
and ( n77041 , n77001 , n77040 );
nor ( n77042 , n76819 , n77000 );
nor ( n77043 , n77041 , n77042 );
nand ( n77044 , n77039 , n77043 );
nor ( n77045 , n77034 , n77044 );
not ( n77046 , n72630 );
not ( n77047 , n77046 );
not ( n77048 , n72456 );
or ( n77049 , n77047 , n77048 );
not ( n77050 , n73920 );
nand ( n77051 , n77050 , n72467 );
nand ( n77052 , n77049 , n77051 );
not ( n77053 , n73918 );
not ( n77054 , n77053 );
not ( n77055 , n73906 );
or ( n77056 , n77054 , n77055 );
not ( n77057 , n69951 );
nand ( n77058 , n77057 , n73916 );
nand ( n77059 , n77056 , n77058 );
nor ( n77060 , n77052 , n77059 );
not ( n77061 , n72538 );
not ( n77062 , n77061 );
not ( n77063 , n76752 );
or ( n77064 , n77062 , n77063 );
not ( n77065 , n72819 );
nand ( n77066 , n71767 , n77065 );
nand ( n77067 , n77064 , n77066 );
not ( n77068 , n72561 );
not ( n77069 , n77068 );
not ( n77070 , n71818 );
or ( n77071 , n77069 , n77070 );
not ( n77072 , n72548 );
nand ( n77073 , n76785 , n77072 );
nand ( n77074 , n77071 , n77073 );
nor ( n77075 , n77067 , n77074 );
nand ( n77076 , n77060 , n77075 );
or ( n77077 , n77045 , n77076 );
nor ( n77078 , n76785 , n77072 );
nor ( n77079 , n71818 , n77068 );
or ( n77080 , n77078 , n77079 );
nand ( n77081 , n77080 , n77073 );
or ( n77082 , n77067 , n77081 );
nor ( n77083 , n76752 , n77061 );
and ( n77084 , n77066 , n77083 );
nor ( n77085 , n71767 , n77065 );
nor ( n77086 , n77084 , n77085 );
nand ( n77087 , n77082 , n77086 );
and ( n77088 , n77060 , n77087 );
not ( n77089 , n72467 );
not ( n77090 , n73920 );
not ( n77091 , n77090 );
and ( n77092 , n77089 , n77091 );
nor ( n77093 , n72456 , n77046 );
and ( n77094 , n77051 , n77093 );
nor ( n77095 , n77092 , n77094 );
or ( n77096 , n77095 , n77059 );
nor ( n77097 , n73906 , n77053 );
and ( n77098 , n77058 , n77097 );
not ( n77099 , n69951 );
nor ( n77100 , n77099 , n73916 );
nor ( n77101 , n77098 , n77100 );
nand ( n77102 , n77096 , n77101 );
nor ( n77103 , n77088 , n77102 );
nand ( n77104 , n77077 , n77103 );
not ( n77105 , n70229 );
not ( n77106 , n77105 );
not ( n77107 , n69981 );
or ( n77108 , n77106 , n77107 );
nand ( n77109 , n77108 , n77026 );
nor ( n77110 , n77017 , n77109 );
nand ( n77111 , n77010 , n77110 );
not ( n77112 , n70331 );
not ( n77113 , n77112 );
not ( n77114 , n69985 );
or ( n77115 , n77113 , n77114 );
not ( n77116 , n70242 );
nand ( n77117 , n77116 , n76399 );
nand ( n77118 , n77115 , n77117 );
not ( n77119 , n70312 );
not ( n77120 , n77119 );
not ( n77121 , n69994 );
or ( n77122 , n77120 , n77121 );
not ( n77123 , n70300 );
nand ( n77124 , n77123 , n70102 );
nand ( n77125 , n77122 , n77124 );
nor ( n77126 , n77118 , n77125 );
not ( n77127 , n70257 );
not ( n77128 , n77127 );
not ( n77129 , n70017 );
or ( n77130 , n77128 , n77129 );
not ( n77131 , n71533 );
not ( n77132 , n70277 );
nand ( n77133 , n77131 , n77132 );
nand ( n77134 , n77130 , n77133 );
not ( n77135 , n70382 );
not ( n77136 , n77135 );
not ( n77137 , n70086 );
or ( n77138 , n77136 , n77137 );
not ( n77139 , n70267 );
nand ( n77140 , n77139 , n70011 );
nand ( n77141 , n77138 , n77140 );
nor ( n77142 , n77134 , n77141 );
not ( n77143 , n70392 );
nand ( n77144 , n70094 , n77143 );
not ( n77145 , n70481 );
nand ( n77146 , n77145 , n70035 );
and ( n77147 , n77144 , n77146 );
not ( n77148 , n70436 );
nand ( n77149 , n77148 , n70028 );
not ( n77150 , n70821 );
not ( n77151 , n77150 );
nand ( n77152 , n77151 , n70042 );
and ( n77153 , n77149 , n77152 );
not ( n77154 , n70424 );
nand ( n77155 , n77154 , n70044 );
not ( n77156 , n69971 );
nor ( n77157 , n77156 , n70526 );
not ( n77158 , n70057 );
nor ( n77159 , n77158 , n70507 );
or ( n77160 , n77157 , n77159 );
not ( n77161 , n70507 );
or ( n77162 , n70057 , n77161 );
nand ( n77163 , n77160 , n77162 );
not ( n77164 , n70463 );
nand ( n77165 , n77164 , n70077 );
nand ( n77166 , n77155 , n77163 , n77165 );
not ( n77167 , n70463 );
nor ( n77168 , n77167 , n70077 );
nand ( n77169 , n77155 , n77168 );
not ( n77170 , n70044 );
nand ( n77171 , n77170 , n70424 );
nand ( n77172 , n77166 , n77169 , n77171 );
nand ( n77173 , n77147 , n77153 , n77172 );
not ( n77174 , n77150 );
nor ( n77175 , n77174 , n70042 );
not ( n77176 , n77175 );
not ( n77177 , n77149 );
or ( n77178 , n77176 , n77177 );
not ( n77179 , n70028 );
nand ( n77180 , n77179 , n70436 );
nand ( n77181 , n77178 , n77180 );
nand ( n77182 , n77147 , n77181 );
not ( n77183 , n70481 );
nor ( n77184 , n77183 , n70035 );
and ( n77185 , n77144 , n77184 );
nor ( n77186 , n70094 , n77143 );
nor ( n77187 , n77185 , n77186 );
nand ( n77188 , n77173 , n77182 , n77187 );
and ( n77189 , n77126 , n77142 , n77188 );
not ( n77190 , n77126 );
nor ( n77191 , n70086 , n77135 );
and ( n77192 , n77140 , n77191 );
not ( n77193 , n70011 );
and ( n77194 , n77193 , n70267 );
nor ( n77195 , n77192 , n77194 );
or ( n77196 , n77195 , n77134 );
nor ( n77197 , n70017 , n77127 );
and ( n77198 , n77133 , n77197 );
nor ( n77199 , n77131 , n77132 );
nor ( n77200 , n77198 , n77199 );
nand ( n77201 , n77196 , n77200 );
not ( n77202 , n77201 );
or ( n77203 , n77190 , n77202 );
not ( n77204 , n77118 );
nor ( n77205 , n69994 , n77119 );
not ( n77206 , n77205 );
not ( n77207 , n77124 );
or ( n77208 , n77206 , n77207 );
not ( n77209 , n70102 );
nand ( n77210 , n77209 , n70300 );
nand ( n77211 , n77208 , n77210 );
and ( n77212 , n77204 , n77211 );
nor ( n77213 , n69985 , n77112 );
not ( n77214 , n77213 );
not ( n77215 , n77117 );
or ( n77216 , n77214 , n77215 );
not ( n77217 , n76399 );
nand ( n77218 , n77217 , n70242 );
nand ( n77219 , n77216 , n77218 );
nor ( n77220 , n77212 , n77219 );
nand ( n77221 , n77203 , n77220 );
nor ( n77222 , n77189 , n77221 );
nor ( n77223 , n77111 , n77222 , n77076 );
nor ( n77224 , n77104 , n77223 );
nand ( n77225 , n70200 , n70151 );
or ( n77226 , n77224 , n77225 );
or ( n77227 , n77225 , n70156 );
nand ( n77228 , n77226 , n77227 );
nand ( n77229 , n77228 , n71987 );
not ( n77230 , n70198 );
nor ( n77231 , n77230 , n70192 );
nand ( n77232 , n77231 , n70151 );
nand ( n77233 , n77225 , n77232 );
not ( n77234 , n77233 );
not ( n77235 , n77224 );
or ( n77236 , n77234 , n77235 );
nand ( n77237 , n77236 , n77227 );
nand ( n77238 , n77237 , n70878 );
not ( n77239 , n77224 );
not ( n77240 , n77232 );
nand ( n77241 , n77240 , n71987 );
not ( n77242 , n77241 );
and ( n77243 , n77239 , n77242 );
and ( n77244 , n70206 , n70210 , n70143 );
not ( n77245 , n77244 );
not ( n77246 , n70229 );
nand ( n77247 , n77246 , n69645 );
not ( n77248 , n69645 );
nand ( n77249 , n77248 , n70229 );
nand ( n77250 , n77247 , n77249 );
not ( n77251 , n70242 );
nand ( n77252 , n77251 , n69617 );
and ( n77253 , n77250 , n77252 );
not ( n77254 , n77250 );
not ( n77255 , n77252 );
and ( n77256 , n77254 , n77255 );
nor ( n77257 , n77253 , n77256 );
not ( n77258 , n72561 );
nand ( n77259 , n77258 , n69936 );
not ( n77260 , n69936 );
nand ( n77261 , n77260 , n72561 );
nand ( n77262 , n77259 , n77261 );
not ( n77263 , n72514 );
nand ( n77264 , n77263 , n69773 );
xor ( n77265 , n77262 , n77264 );
nand ( n77266 , n77257 , n77265 );
not ( n77267 , n72630 );
nand ( n77268 , n77267 , n69733 );
not ( n77269 , n69733 );
nand ( n77270 , n77269 , n72630 );
nand ( n77271 , n77268 , n77270 );
not ( n77272 , n72818 );
not ( n77273 , n77272 );
nand ( n77274 , n77273 , n69710 );
xor ( n77275 , n77271 , n77274 );
not ( n77276 , n73920 );
nand ( n77277 , n77276 , n69747 );
not ( n77278 , n77277 );
not ( n77279 , n77278 );
not ( n77280 , n73918 );
nand ( n77281 , n77280 , n69912 );
not ( n77282 , n69912 );
nand ( n77283 , n77282 , n73918 );
nand ( n77284 , n77281 , n77283 );
not ( n77285 , n77284 );
or ( n77286 , n77279 , n77285 );
or ( n77287 , n77284 , n77278 );
nand ( n77288 , n77286 , n77287 );
not ( n77289 , n77281 );
not ( n77290 , n77289 );
xor ( n77291 , n69946 , n73916 );
not ( n77292 , n77291 );
or ( n77293 , n77290 , n77292 );
or ( n77294 , n77291 , n77289 );
nand ( n77295 , n77293 , n77294 );
nand ( n77296 , n77275 , n77288 , n77295 );
nor ( n77297 , n77266 , n77296 );
not ( n77298 , n71126 );
not ( n77299 , n69808 );
not ( n77300 , n77299 );
or ( n77301 , n77298 , n77300 );
not ( n77302 , n71126 );
nand ( n77303 , n77302 , n69808 );
nand ( n77304 , n77301 , n77303 );
not ( n77305 , n77304 );
not ( n77306 , n71096 );
nand ( n77307 , n77306 , n69826 );
not ( n77308 , n77307 );
and ( n77309 , n77305 , n77308 );
and ( n77310 , n77304 , n77307 );
nor ( n77311 , n77309 , n77310 );
not ( n77312 , n71096 );
not ( n77313 , n69826 );
not ( n77314 , n77313 );
or ( n77315 , n77312 , n77314 );
nand ( n77316 , n77315 , n77307 );
not ( n77317 , n71078 );
nand ( n77318 , n77317 , n69659 );
and ( n77319 , n77316 , n77318 );
not ( n77320 , n77316 );
not ( n77321 , n77318 );
and ( n77322 , n77320 , n77321 );
nor ( n77323 , n77319 , n77322 );
not ( n77324 , n69580 );
not ( n77325 , n77324 );
not ( n77326 , n70300 );
or ( n77327 , n77325 , n77326 );
not ( n77328 , n70300 );
nand ( n77329 , n77328 , n69580 );
nand ( n77330 , n77327 , n77329 );
not ( n77331 , n70312 );
nand ( n77332 , n77331 , n69591 );
xor ( n77333 , n77330 , n77332 );
not ( n77334 , n72503 );
nand ( n77335 , n77334 , n69796 );
not ( n77336 , n69796 );
nand ( n77337 , n77336 , n72503 );
nand ( n77338 , n77335 , n77337 );
not ( n77339 , n72479 );
nand ( n77340 , n77339 , n69900 );
xor ( n77341 , n77338 , n77340 );
nand ( n77342 , n77311 , n77323 , n77333 , n77341 );
not ( n77343 , n72548 );
nand ( n77344 , n77343 , n69854 );
not ( n77345 , n69854 );
nand ( n77346 , n77345 , n72548 );
nand ( n77347 , n77344 , n77346 );
xor ( n77348 , n77347 , n77259 );
not ( n77349 , n69591 );
not ( n77350 , n77349 );
not ( n77351 , n70312 );
or ( n77352 , n77350 , n77351 );
nand ( n77353 , n77352 , n77332 );
not ( n77354 , n70277 );
nand ( n77355 , n77354 , n69523 );
xor ( n77356 , n77353 , n77355 );
not ( n77357 , n69710 );
nand ( n77358 , n77357 , n77272 );
nand ( n77359 , n77274 , n77358 );
not ( n77360 , n72538 );
nand ( n77361 , n77360 , n69689 );
xor ( n77362 , n77359 , n77361 );
not ( n77363 , n69689 );
nand ( n77364 , n77363 , n72538 );
nand ( n77365 , n77361 , n77364 );
xor ( n77366 , n77365 , n77344 );
nand ( n77367 , n77348 , n77356 , n77362 , n77366 );
nor ( n77368 , n77342 , n77367 );
not ( n77369 , n69659 );
nand ( n77370 , n77369 , n71078 );
nand ( n77371 , n77318 , n77370 );
and ( n77372 , n77371 , n77247 );
not ( n77373 , n77371 );
not ( n77374 , n77247 );
and ( n77375 , n77373 , n77374 );
nor ( n77376 , n77372 , n77375 );
not ( n77377 , n69900 );
nand ( n77378 , n77377 , n72479 );
nand ( n77379 , n77340 , n77378 );
not ( n77380 , n72489 );
nand ( n77381 , n77380 , n69875 );
xor ( n77382 , n77379 , n77381 );
not ( n77383 , n70277 );
not ( n77384 , n69523 );
not ( n77385 , n77384 );
or ( n77386 , n77383 , n77385 );
nand ( n77387 , n77386 , n77355 );
not ( n77388 , n70257 );
nand ( n77389 , n77388 , n69535 );
xor ( n77390 , n77387 , n77389 );
not ( n77391 , n69439 );
not ( n77392 , n77391 );
not ( n77393 , n70481 );
or ( n77394 , n77392 , n77393 );
not ( n77395 , n70481 );
nand ( n77396 , n77395 , n69439 );
nand ( n77397 , n77394 , n77396 );
not ( n77398 , n70436 );
nand ( n77399 , n77398 , n69506 );
xor ( n77400 , n77397 , n77399 );
nand ( n77401 , n77376 , n77382 , n77390 , n77400 );
not ( n77402 , n70331 );
not ( n77403 , n69603 );
not ( n77404 , n77403 );
or ( n77405 , n77402 , n77404 );
not ( n77406 , n70331 );
nand ( n77407 , n77406 , n69603 );
nand ( n77408 , n77405 , n77407 );
xor ( n77409 , n77408 , n77329 );
not ( n77410 , n70242 );
not ( n77411 , n69617 );
not ( n77412 , n77411 );
or ( n77413 , n77410 , n77412 );
nand ( n77414 , n77413 , n77252 );
xor ( n77415 , n77414 , n77407 );
not ( n77416 , n69875 );
nand ( n77417 , n77416 , n72489 );
nand ( n77418 , n77381 , n77417 );
xor ( n77419 , n77418 , n77303 );
not ( n77420 , n69773 );
nand ( n77421 , n77420 , n72514 );
nand ( n77422 , n77264 , n77421 );
xor ( n77423 , n77422 , n77335 );
nand ( n77424 , n77409 , n77415 , n77419 , n77423 );
nor ( n77425 , n77401 , n77424 );
not ( n77426 , n69747 );
nand ( n77427 , n77426 , n73920 );
nand ( n77428 , n77277 , n77427 );
xor ( n77429 , n77428 , n77268 );
not ( n77430 , n69491 );
not ( n77431 , n77430 );
not ( n77432 , n70821 );
not ( n77433 , n77432 );
or ( n77434 , n77431 , n77433 );
not ( n77435 , n77432 );
nand ( n77436 , n77435 , n69491 );
nand ( n77437 , n77434 , n77436 );
not ( n77438 , n70424 );
nand ( n77439 , n77438 , n69475 );
xor ( n77440 , n77437 , n77439 );
not ( n77441 , n69474 );
not ( n77442 , n77441 );
not ( n77443 , n70392 );
or ( n77444 , n77442 , n77443 );
not ( n77445 , n70392 );
nand ( n77446 , n77445 , n69474 );
nand ( n77447 , n77444 , n77446 );
xor ( n77448 , n77447 , n77396 );
not ( n77449 , n69547 );
not ( n77450 , n77449 );
not ( n77451 , n70267 );
or ( n77452 , n77450 , n77451 );
not ( n77453 , n70267 );
nand ( n77454 , n77453 , n69547 );
nand ( n77455 , n77452 , n77454 );
not ( n77456 , n70382 );
nand ( n77457 , n77456 , n69557 );
xor ( n77458 , n77455 , n77457 );
nand ( n77459 , n77429 , n77440 , n77448 , n77458 );
not ( n77460 , n70257 );
not ( n77461 , n69535 );
not ( n77462 , n77461 );
or ( n77463 , n77460 , n77462 );
nand ( n77464 , n77463 , n77389 );
xor ( n77465 , n77464 , n77454 );
not ( n77466 , n69506 );
not ( n77467 , n77466 );
not ( n77468 , n70436 );
or ( n77469 , n77467 , n77468 );
nand ( n77470 , n77469 , n77399 );
and ( n77471 , n77470 , n77436 );
not ( n77472 , n77470 );
not ( n77473 , n77436 );
and ( n77474 , n77472 , n77473 );
nor ( n77475 , n77471 , n77474 );
not ( n77476 , n69557 );
not ( n77477 , n77476 );
not ( n77478 , n70382 );
or ( n77479 , n77477 , n77478 );
nand ( n77480 , n77479 , n77457 );
xor ( n77481 , n77480 , n77446 );
xnor ( n77482 , n70077 , n70463 );
not ( n77483 , n69971 );
and ( n77484 , n70526 , n77483 );
not ( n77485 , n70526 );
and ( n77486 , n77485 , n69971 );
nor ( n77487 , n77484 , n77486 );
xnor ( n77488 , n70507 , n70057 );
nand ( n77489 , n77482 , n77487 , n77488 );
xor ( n77490 , n69475 , n69455 );
xor ( n77491 , n77490 , n70424 );
nor ( n77492 , n77489 , n77491 );
nand ( n77493 , n77465 , n77475 , n77481 , n77492 );
nor ( n77494 , n77459 , n77493 );
and ( n77495 , n77297 , n77368 , n77425 , n77494 );
not ( n77496 , n70192 );
nor ( n77497 , n77496 , n70867 , n70198 );
not ( n77498 , n77497 );
or ( n77499 , n77495 , n77498 );
nand ( n77500 , n77497 , n4012 );
nand ( n77501 , n77499 , n77500 );
not ( n77502 , n77501 );
or ( n77503 , n77245 , n77502 );
nor ( n77504 , n70564 , n70867 );
nand ( n77505 , n77504 , n77244 );
nor ( n77506 , n77495 , n77505 );
not ( n77507 , n71987 );
nand ( n77508 , n70206 , n70869 , n70143 );
and ( n77509 , n70877 , n77507 , n77508 );
nor ( n77510 , n77509 , n77500 );
nor ( n77511 , n77506 , n77510 );
nand ( n77512 , n77503 , n77511 );
nor ( n77513 , n77243 , n77512 );
and ( n77514 , n77229 , n77238 , n77513 );
not ( n77515 , n71126 );
nor ( n77516 , n71062 , n77515 );
not ( n77517 , n71096 );
nor ( n77518 , n71051 , n77517 );
nor ( n77519 , n77516 , n77518 );
not ( n77520 , n71078 );
nand ( n77521 , n77520 , n69664 );
not ( n77522 , n70229 );
nand ( n77523 , n77522 , n69981 );
and ( n77524 , n77521 , n77523 );
not ( n77525 , n71078 );
nor ( n77526 , n77525 , n69664 );
nor ( n77527 , n77524 , n77526 );
and ( n77528 , n77519 , n77527 );
not ( n77529 , n71096 );
nand ( n77530 , n77529 , n71051 );
or ( n77531 , n77516 , n77530 );
nand ( n77532 , n71062 , n77515 );
nand ( n77533 , n77531 , n77532 );
nor ( n77534 , n77528 , n77533 );
not ( n77535 , n71837 );
not ( n77536 , n72514 );
nor ( n77537 , n77535 , n77536 );
not ( n77538 , n72503 );
nor ( n77539 , n71856 , n77538 );
nor ( n77540 , n77537 , n77539 );
not ( n77541 , n72479 );
nor ( n77542 , n71873 , n77541 );
not ( n77543 , n72489 );
nor ( n77544 , n77543 , n71041 );
nor ( n77545 , n77542 , n77544 );
nand ( n77546 , n77540 , n77545 );
or ( n77547 , n77534 , n77546 );
not ( n77548 , n71873 );
not ( n77549 , n77541 );
or ( n77550 , n77548 , n77549 );
not ( n77551 , n72489 );
nand ( n77552 , n77551 , n71041 );
or ( n77553 , n77542 , n77552 );
nand ( n77554 , n77550 , n77553 );
and ( n77555 , n77554 , n77540 );
nand ( n77556 , n71856 , n77538 );
or ( n77557 , n77537 , n77556 );
nand ( n77558 , n77535 , n77536 );
nand ( n77559 , n77557 , n77558 );
nor ( n77560 , n77555 , n77559 );
nand ( n77561 , n77547 , n77560 );
not ( n77562 , n77561 );
not ( n77563 , n73918 );
not ( n77564 , n73906 );
not ( n77565 , n77564 );
or ( n77566 , n77563 , n77565 );
not ( n77567 , n73916 );
nand ( n77568 , n69951 , n77567 );
nand ( n77569 , n77566 , n77568 );
not ( n77570 , n77569 );
not ( n77571 , n73920 );
nor ( n77572 , n72467 , n77571 );
not ( n77573 , n72630 );
nor ( n77574 , n77573 , n72456 );
nor ( n77575 , n77572 , n77574 );
nand ( n77576 , n77570 , n77575 );
not ( n77577 , n72819 );
nor ( n77578 , n77577 , n71767 );
not ( n77579 , n72538 );
nor ( n77580 , n77579 , n76752 );
nor ( n77581 , n77578 , n77580 );
not ( n77582 , n72548 );
nor ( n77583 , n76785 , n77582 );
not ( n77584 , n72561 );
nor ( n77585 , n71818 , n77584 );
nor ( n77586 , n77583 , n77585 );
nand ( n77587 , n77581 , n77586 );
nor ( n77588 , n77576 , n77587 );
not ( n77589 , n77588 );
or ( n77590 , n77562 , n77589 );
not ( n77591 , n77576 );
nand ( n77592 , n76785 , n77582 );
nand ( n77593 , n71818 , n77584 );
and ( n77594 , n77592 , n77593 );
nor ( n77595 , n77594 , n77583 );
not ( n77596 , n77595 );
not ( n77597 , n77581 );
or ( n77598 , n77596 , n77597 );
not ( n77599 , n77578 );
not ( n77600 , n76752 );
nor ( n77601 , n77600 , n72538 );
and ( n77602 , n77599 , n77601 );
not ( n77603 , n71767 );
nor ( n77604 , n77603 , n72819 );
nor ( n77605 , n77602 , n77604 );
nand ( n77606 , n77598 , n77605 );
and ( n77607 , n77591 , n77606 );
not ( n77608 , n72467 );
not ( n77609 , n77608 );
not ( n77610 , n73920 );
and ( n77611 , n77609 , n77610 );
not ( n77612 , n77572 );
not ( n77613 , n72456 );
nor ( n77614 , n77613 , n72630 );
and ( n77615 , n77612 , n77614 );
nor ( n77616 , n77611 , n77615 );
or ( n77617 , n77616 , n77569 );
not ( n77618 , n73906 );
nor ( n77619 , n77618 , n73918 );
and ( n77620 , n77568 , n77619 );
nor ( n77621 , n69951 , n77567 );
nor ( n77622 , n77620 , n77621 );
nand ( n77623 , n77617 , n77622 );
nor ( n77624 , n77607 , n77623 );
nand ( n77625 , n77590 , n77624 );
not ( n77626 , n76399 );
nand ( n77627 , n77626 , n70242 );
not ( n77628 , n69985 );
nand ( n77629 , n77628 , n70331 );
nand ( n77630 , n77627 , n77629 );
not ( n77631 , n70102 );
nand ( n77632 , n77631 , n70300 );
not ( n77633 , n69994 );
nand ( n77634 , n77633 , n70312 );
nand ( n77635 , n77632 , n77634 );
nor ( n77636 , n77630 , n77635 );
not ( n77637 , n70277 );
nor ( n77638 , n77637 , n76517 );
not ( n77639 , n70257 );
nor ( n77640 , n77639 , n70017 );
nor ( n77641 , n77638 , n77640 );
not ( n77642 , n77641 );
not ( n77643 , n70382 );
not ( n77644 , n70086 );
not ( n77645 , n77644 );
or ( n77646 , n77643 , n77645 );
not ( n77647 , n70267 );
nor ( n77648 , n77647 , n70011 );
not ( n77649 , n77648 );
nand ( n77650 , n77646 , n77649 );
nor ( n77651 , n77642 , n77650 );
not ( n77652 , n70392 );
nor ( n77653 , n77652 , n70094 );
not ( n77654 , n70481 );
nor ( n77655 , n77654 , n70035 );
nor ( n77656 , n77653 , n77655 );
not ( n77657 , n70436 );
nor ( n77658 , n70028 , n77657 );
not ( n77659 , n72306 );
nor ( n77660 , n77659 , n70042 );
nor ( n77661 , n77658 , n77660 );
not ( n77662 , n70044 );
nand ( n77663 , n77662 , n70424 );
not ( n77664 , n70526 );
nor ( n77665 , n77664 , n69971 );
not ( n77666 , n70057 );
and ( n77667 , n77666 , n70507 );
or ( n77668 , n77665 , n77667 );
or ( n77669 , n77666 , n70507 );
nand ( n77670 , n77668 , n77669 );
not ( n77671 , n70077 );
nand ( n77672 , n77671 , n70463 );
nand ( n77673 , n77663 , n77670 , n77672 );
not ( n77674 , n70077 );
nor ( n77675 , n77674 , n70463 );
nand ( n77676 , n77663 , n77675 );
not ( n77677 , n70424 );
nand ( n77678 , n77677 , n70044 );
nand ( n77679 , n77673 , n77676 , n77678 );
nand ( n77680 , n77656 , n77661 , n77679 );
not ( n77681 , n72306 );
nand ( n77682 , n77681 , n70042 );
or ( n77683 , n77658 , n77682 );
nand ( n77684 , n70028 , n77657 );
nand ( n77685 , n77683 , n77684 );
nand ( n77686 , n77656 , n77685 );
not ( n77687 , n77653 );
not ( n77688 , n70035 );
nor ( n77689 , n77688 , n70481 );
and ( n77690 , n77687 , n77689 );
not ( n77691 , n70094 );
nor ( n77692 , n77691 , n70392 );
nor ( n77693 , n77690 , n77692 );
nand ( n77694 , n77680 , n77686 , n77693 );
nand ( n77695 , n77636 , n77651 , n77694 );
not ( n77696 , n77641 );
not ( n77697 , n70382 );
nand ( n77698 , n77697 , n70086 );
or ( n77699 , n77648 , n77698 );
not ( n77700 , n70011 );
or ( n77701 , n77700 , n70267 );
nand ( n77702 , n77699 , n77701 );
not ( n77703 , n77702 );
or ( n77704 , n77696 , n77703 );
not ( n77705 , n77638 );
not ( n77706 , n70017 );
nor ( n77707 , n77706 , n70257 );
and ( n77708 , n77705 , n77707 );
not ( n77709 , n76517 );
nor ( n77710 , n77709 , n70277 );
nor ( n77711 , n77708 , n77710 );
nand ( n77712 , n77704 , n77711 );
nand ( n77713 , n77712 , n77636 );
not ( n77714 , n77632 );
not ( n77715 , n70312 );
nand ( n77716 , n77715 , n69994 );
or ( n77717 , n77714 , n77716 );
not ( n77718 , n70300 );
nand ( n77719 , n77718 , n70102 );
nand ( n77720 , n77717 , n77719 );
not ( n77721 , n77630 );
and ( n77722 , n77720 , n77721 );
not ( n77723 , n77627 );
not ( n77724 , n70331 );
nand ( n77725 , n77724 , n69985 );
or ( n77726 , n77723 , n77725 );
not ( n77727 , n70242 );
nand ( n77728 , n77727 , n76399 );
nand ( n77729 , n77726 , n77728 );
nor ( n77730 , n77722 , n77729 );
nand ( n77731 , n77695 , n77713 , n77730 );
not ( n77732 , n70229 );
nor ( n77733 , n77732 , n69981 );
nor ( n77734 , n77526 , n77733 );
nand ( n77735 , n77519 , n77734 );
nor ( n77736 , n77546 , n77735 );
not ( n77737 , n77587 );
and ( n77738 , n77591 , n77731 , n77736 , n77737 );
nor ( n77739 , n77625 , n77738 );
or ( n77740 , n77739 , n70877 );
not ( n77741 , n77508 );
nand ( n77742 , n77495 , n77741 );
nand ( n77743 , n77740 , n77742 );
not ( n77744 , n77743 );
nand ( n77745 , n77739 , n71987 );
nand ( n77746 , n77744 , n77745 );
nand ( n77747 , n77746 , n77497 );
nand ( n77748 , n77746 , n77504 );
and ( n77749 , n77233 , n77741 );
not ( n77750 , n77227 );
and ( n77751 , n77750 , n77244 );
nor ( n77752 , n77749 , n77751 );
and ( n77753 , n77514 , n77747 , n77748 , n77752 );
or ( n77754 , n76995 , n77753 );
nand ( n77755 , n77514 , n77747 , n77748 );
not ( n77756 , n77244 );
not ( n77757 , n77233 );
or ( n77758 , n77756 , n77757 );
or ( n77759 , n77227 , n77508 );
nand ( n77760 , n77758 , n77759 );
nor ( n77761 , n77755 , n77760 );
or ( n77762 , n77761 , n76994 );
not ( n77763 , n75279 );
nor ( n77764 , n70145 , n70212 , n77763 );
not ( n77765 , n77764 );
nand ( n77766 , n70151 , n70864 );
nand ( n77767 , n77765 , n77766 , n4012 );
nand ( n77768 , n77754 , n77762 , n77767 );
buf ( n77769 , n77768 );
buf ( n77770 , 1'b0 );
not ( n77771 , n68639 );
not ( n77772 , n77771 );
buf ( n77773 , n77772 );
buf ( n77774 , n68638 );
buf ( n77775 , n71728 );
buf ( n77776 , 1'b0 );
not ( n77777 , n77771 );
buf ( n77778 , n77777 );
buf ( n77779 , n68638 );
nand ( n77780 , n70192 , n70198 );
and ( n77781 , n70140 , n77780 );
nor ( n77782 , n77781 , n70151 );
not ( n77783 , n70226 );
or ( n77784 , n77782 , n77783 );
nand ( n77785 , n77784 , n70864 );
buf ( n77786 , n77785 );
endmodule

