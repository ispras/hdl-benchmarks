module GTECH_NOT(Z, A);

output Z;
input A;

not U(Z,A);

endmodule
