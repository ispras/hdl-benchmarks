// IWLS benchmark module "t481" printed on Wed May 29 17:29:17 2002
module t481(v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14, v15, \v16.0 );
input
  v10,
  v11,
  v12,
  v13,
  v14,
  v15,
  v0,
  v1,
  v2,
  v3,
  v4,
  v5,
  v6,
  v7,
  v8,
  v9;
output
  \v16.0 ;
wire
  \[60] ,
  \[338] ,
  \[145] ,
  \[13028] ,
  \[61] ,
  \[146] ,
  \[62] ,
  \[13963] ,
  \[147] ,
  \[63] ,
  \[148] ,
  \[64] ,
  \[13412] ,
  \[149] ,
  \[436] ,
  \[65] ,
  \[12664] ,
  \[8397] ,
  \[66] ,
  \[1182] ,
  \[8415] ,
  \[438] ,
  \[67] ,
  \[439] ,
  \[68] ,
  \[69] ,
  \[13129] ,
  \[343] ,
  \[0] ,
  \[344] ,
  \[1] ,
  \[345] ,
  \[2] ,
  \[13592] ,
  \[153] ,
  \[3] ,
  \[440] ,
  \[5649] ,
  \[12961] ,
  \[1478] ,
  \[154] ,
  \[4] ,
  \[441] ,
  \[70] ,
  \[155] ,
  \[5] ,
  \[442] ,
  \[71] ,
  \[156] ,
  \[6] ,
  \[443] ,
  \[72] ,
  \[7] ,
  \[73] ,
  \[11753] ,
  \[8] ,
  \[74] ,
  \[2687] ,
  \[159] ,
  \[9] ,
  \[75] ,
  \[11472] ,
  \[2705] ,
  \[76] ,
  \[448] ,
  \[77] ,
  \[449] ,
  \[78] ,
  \[256] ,
  \[79] ,
  \[6571] ,
  \[259] ,
  \[10079] ,
  \[13694] ,
  \[163] ,
  \[1581] ,
  \[164] ,
  \[80] ,
  \[11190] ,
  \[165] ,
  \[81] ,
  \[453] ,
  \[82] ,
  \[260] ,
  \[454] ,
  \[83] ,
  \[261] ,
  \[455] ,
  \[84] ,
  \[262] ,
  \[8433] ,
  \[169] ,
  \[456] ,
  \[85] ,
  \[263] ,
  \[86] ,
  \[458] ,
  \[87] ,
  \[11576] ,
  \[13525] ,
  \[88] ,
  \[13627] ,
  \[12494] ,
  \[89] ,
  \[361] ,
  \[268] ,
  \[362] ,
  \[1030] ,
  \[269] ,
  \[12784] ,
  \[363] ,
  \[364] ,
  \[171] ,
  \[14256] ,
  \[10] ,
  \[5667] ,
  \[365] ,
  \[172] ,
  \[11] ,
  \[1033] ,
  \[173] ,
  \[12] ,
  \[1514] ,
  \[367] ,
  \[174] ,
  \[13] ,
  \[368] ,
  \[14] ,
  \[91] ,
  \[13244] ,
  \[15] ,
  \[463] ,
  \[92] ,
  \[270] ,
  \[464] ,
  \[93] ,
  \[10110] ,
  \[2723] ,
  \[17] ,
  \[465] ,
  \[13348] ,
  \[94] ,
  \[18] ,
  \[95] ,
  \[96] ,
  \[97] ,
  \[98] ,
  \[100] ,
  \[99] ,
  \[101] ,
  \[102] ,
  \[373] ,
  \[103] ,
  \[374] ,
  \[104] ,
  \[181] ,
  \[375] ,
  \[105] ,
  \[106] ,
  \[183] ,
  \[10095] ,
  \[107] ,
  \[184] ,
  \[23] ,
  \[108] ,
  \[185] ,
  \[24] ,
  \[109] ,
  \[187] ,
  \[26] ,
  \[474] ,
  \[27] ,
  \[475] ,
  \[12822] ,
  \[28] ,
  \[476] ,
  \[300] ,
  \[29] ,
  \[13063] ,
  \[477] ,
  \[301] ,
  \[302] ,
  \[303] ,
  \[110] ,
  \[1241] ,
  \[287] ,
  \[304] ,
  \[111] ,
  \[288] ,
  \[305] ,
  \[112] ,
  \[289] ,
  \[10319] ,
  \[113] ,
  \[307] ,
  \[114] ,
  \[308] ,
  \[115] ,
  \[672] ,
  \[403] ,
  \[193] ,
  \[32] ,
  \[5689] ,
  \[117] ,
  \[404] ,
  \[194] ,
  \[33] ,
  \[118] ,
  \[10123] ,
  \[405] ,
  \[195] ,
  \[34] ,
  \[119] ,
  \[35] ,
  \[1537] ,
  \[213] ,
  \[36] ,
  \[214] ,
  \[215] ,
  \[216] ,
  \[293] ,
  \[39] ,
  \[218] ,
  \[313] ,
  \[120] ,
  \[314] ,
  \[121] ,
  \[298] ,
  \[5711] ,
  \[315] ,
  \[299] ,
  \[10516] ,
  \[393] ,
  \[123] ,
  \[394] ,
  \[124] ,
  \[40] ,
  \[395] ,
  \[125] ,
  \[12359] ,
  \[41] ,
  \[1063] ,
  \[396] ,
  \[127] ,
  \[971] ,
  \[43] ,
  \[11539] ,
  \[129] ,
  \[45] ,
  \[223] ,
  \[46] ,
  \[224] ,
  \[10693] ,
  \[47] ,
  \[48] ,
  \[49] ,
  \[130] ,
  \[14213] ,
  \[13103] ,
  \[131] ,
  \[132] ,
  \[12848] ,
  \[12745] ,
  \[133] ,
  \[10795] ,
  \[134] ,
  \[50] ,
  \[135] ,
  \[51] ,
  \[136] ,
  \[52] ,
  \[11641] ,
  \[53] ,
  \[54] ,
  \[10626] ,
  \[55] ,
  \[10728] ,
  \[56] ,
  \[2669] ,
  \[57] ,
  \[1559] ,
  \[58] ,
  \[59] ,
  \[794] ,
  \[14132] ,
  \[333] ,
  \[1464] ,
  \[334] ,
  \[13386] ,
  \[335] ,
  \[1273] ,
  \[336] ,
  \[143] ,
  \[13311] ;
assign
  \[60]  = \[12]  | \[10] ,
  \[338]  = 0,
  \[145]  = \[53]  | (\[52]  | \[8433] ),
  \[13028]  = \[109]  & \[53] ,
  \[61]  = \[33]  & \[11] ,
  \[146]  = \[129]  & ~\[6] ,
  \[62]  = \[45]  & ~\[15] ,
  \[13963]  = \[85]  & \[61] ,
  \[147]  = \[45]  & ~v6,
  \[63]  = v2 | ~v0,
  \[148]  = ~\[1581]  & \[5649] ,
  \[64]  = \[62]  & \[47] ,
  \[13412]  = \[118]  & \[65] ,
  \[149]  = v7 & ~v5,
  \[436]  = \[84]  & ~\[58] ,
  \[65]  = \[11]  & ~\[10] ,
  \[12664]  = \[77]  & \[67] ,
  \[8397]  = \[169]  & \[159] ,
  \[66]  = \[5711]  & ~v7,
  \[1182]  = (~\[132]  & (~\[55]  & (~\[53]  & ~\[50] ))) | \[71] ,
  \[8415]  = \[174]  & \[159] ,
  \[438]  = 0,
  \[67]  = \[33]  & ~\[12] ,
  \[439]  = \[120]  & ~\[58] ,
  \[68]  = \[5]  | v9,
  \[69]  = (~\[7]  & \[5] ) | (\[7]  & ~\[5] ),
  \[13129]  = (\[101]  & \[56] ) | (\[89]  & \[11] ),
  \[343]  = \[109]  & \[64] ,
  \[0]  = ~\[794]  | (~\[1033]  | (~\[1273]  | ~\[1514] )),
  \[344]  = \[109]  & ~\[13] ,
  \[1]  = ~v13 | v12,
  \[345]  = \[109]  & \[2723] ,
  \[2]  = v15 | ~v14,
  \[13592]  = \[82]  & \[53] ,
  \[153]  = \[75]  & ~\[54] ,
  \[3]  = \[1]  | v14,
  \[440]  = \[100]  & ~\[58] ,
  \[5649]  = \[169]  & \[149] ,
  \[12961]  = \[59]  & \[11] ,
  \[1478]  = (~\[114]  & \[48] ) | \[63] ,
  \[154]  = \[73]  & ~\[54] ,
  \[4]  = v3 | ~v2,
  \[441]  = \[101]  & \[61] ,
  \[70]  = \[7]  | v10,
  \[155]  = \[66]  & ~\[54] ,
  \[5]  = v11 | ~v10,
  \[442]  = \[102]  & \[61] ,
  \[71]  = \[9]  | \[3] ,
  \[156]  = \[84]  & ~\[54] ,
  \[6]  = ~v1 | v0,
  \[443]  = \[64]  & \[61] ,
  \[72]  = \[23]  & \[11] ,
  \[7]  = ~v9 | v8,
  \[73]  = \[36]  & v0,
  \[11753]  = \[59]  & ~\[12] ,
  \[8]  = \[2]  | ~v12,
  \[74]  = ~\[6]  & v3,
  \[2687]  = \[47]  & (~v6 & v4),
  \[159]  = ~v6 & ~v5,
  \[9]  = v10 | v9,
  \[75]  = \[36]  & ~v1,
  \[11472]  = \[77]  & \[57] ,
  \[2705]  = \[159]  & \[74] ,
  \[76]  = \[17]  | \[12] ,
  \[448]  = \[61]  & \[2669] ,
  \[77]  = \[41]  | \[6571] ,
  \[449]  = \[61]  & \[6571] ,
  \[78]  = (v15 & v12) | \[49] ,
  \[256]  = \[84]  & ~\[60] ,
  \[79]  = \[23]  & ~\[8] ,
  \[6571]  = \[149]  & \[47] ,
  \[259]  = \[101]  & ~\[18] ,
  \[10079]  = \[108]  & (~v2 & ~v1),
  \[13694]  = (\[101]  & ~\[58] ) | ((\[88]  & \[82] ) | (\[82]  & \[55] )),
  \[163]  = ~\[71]  & \[64] ,
  \[1581]  = \[5649]  & ~v8,
  \v16.0  = \[0] ,
  \[164]  = ~\[71]  & ~\[13] ,
  \[80]  = \[23]  & ~\[12] ,
  \[11190]  = (\[146]  & ~\[71] ) | (\[110]  & ~\[54] ),
  \[165]  = ~\[71]  & \[2723] ,
  \[81]  = \[33]  & ~\[8] ,
  \[453]  = \[75]  & \[61] ,
  \[82]  = \[23]  & ~\[3] ,
  \[260]  = \[120]  & ~\[60] ,
  \[454]  = \[73]  & \[61] ,
  \[83]  = ~\[14]  & ~\[7] ,
  \[261]  = \[100]  & ~\[60] ,
  \[455]  = \[66]  & \[61] ,
  \[84]  = \[5689]  & ~v7,
  \[262]  = \[102]  & ~\[18] ,
  \[8433]  = \[149]  & \[74] ,
  \[169]  = ~\[4]  & v0,
  \[456]  = \[84]  & \[61] ,
  \[85]  = \[52]  | \[40] ,
  \[263]  = \[64]  & ~\[18] ,
  \[86]  = ~\[5]  & v9,
  \[458]  = 0,
  \[87]  = ~\[70]  | ~\[68] ,
  \[11576]  = (\[115]  & \[80] ) | (\[100]  & \[57] ),
  \[13525]  = (\[146]  & \[82] ) | (\[110]  & \[65] ),
  \[88]  = \[120]  | \[5649] ,
  \[13627]  = \[82]  & \[50] ,
  \[12494]  = \[81]  & \[55] ,
  \[89]  = \[88]  & ~\[17] ,
  \[361]  = \[109]  & \[100] ,
  \[268]  = ~\[18]  & \[2669] ,
  \[362]  = \[102]  & \[56] ,
  \[1030]  = (~\[117]  & (~\[115]  & (~\[77]  & (~\[52]  & (~\[40]  & ~\[2669] ))))) | \[60] ,
  \[269]  = ~\[18]  & \[6571] ,
  \[12784]  = (\[86]  & (~\[12]  & \[1537] )) | (\[115]  & \[72] ),
  \[363]  = \[64]  & \[56] ,
  \[364]  = \[56]  & ~\[13] ,
  \[171]  = \[45]  & v6,
  \[14256]  = \[83]  & \[50] ,
  \[10]  = ~v11 | v9,
  \[5667]  = \[174]  & \[149] ,
  \[365]  = \[56]  & \[2723] ,
  \[172]  = \[148]  & v11,
  \[11]  = ~\[1]  & v15,
  \[1033]  = (\[28]  & (~\[2705]  & (~\[336]  & (~\[335]  & (~\[334]  & (~\[333]  & (~\[344]  & (~\[343]  & (~\[345]  & (~\[12961]  & (~\[13129]  & (~\[13103]  & (~\[13063]  & (~\[13028]  & (~\[308]  & (~\[307]  & (~\[305]  & (~\[304]  & (~\[303]  & (~\[302]  & (~\[301]  & (~\[314]  & (~\[313]  & (~\[315]  & (~\[12664]  & (~\[12848]  & (~\[12822]  & (~\[12784]  & (~\[12745]  & (~\[293]  & (~\[289]  & (~\[288]  & (~\[287]  & (~\[299]  & (~\[300]  & (~\[12494]  & (\[971]  & (~\[5649]  & (~\[5667]  & (~\[263]  & (~\[262]  & (~\[261]  & (~\[260]  & (~\[259]  & (~\[256]  & (~\[269]  & (~\[268]  & (\[1030]  & (~\[8397]  & (~\[8415]  & ~\[8433] )))))))))))))))))))))))))))))))))))))))))))))))))) | (~\[81]  & (~\[72]  & (~\[67]  & (\[60]  & (\[28]  & (~\[344]  & (~\[343]  & (~\[345]  & (~\[12961]  & (~\[13129]  & (~\[13103]  & (~\[13063]  & (~\[13028]  & (\[971]  & (~\[263]  & (~\[262]  & (~\[259]  & (~\[269]  & (~\[268]  & ~\[270] ))))))))))))))))))),
  \[173]  = \[86]  & ~\[8] ,
  \[12]  = \[2]  | v13,
  \[1514]  = (\[32]  & (~\[98]  & (~\[97]  & (~\[96]  & (~\[95]  & (~\[94]  & (~\[93]  & (~\[92]  & (~\[91]  & (~\[104]  & (~\[103]  & (~\[105]  & (~\[10626]  & (~\[10728]  & (~\[10693]  & (~\[10795]  & (~\[10516]  & (~\[10319]  & (\[1478]  & (\[1464]  & (~\[10123]  & (~\[10110]  & (~\[10095]  & ~\[10079] ))))))))))))))))))))))) | ((\[99]  & (\[34]  & (~\[32]  & (\[5]  & (\[1464]  & ~v15))))) | ((\[99]  & (~\[34]  & (~\[5]  & (\[1464]  & ~v15)))) | ((\[34]  & (~\[32]  & (\[5]  & (\[1464]  & v13)))) | (~\[34]  & (~\[5]  & (\[1464]  & v13)))))),
  \[367]  = \[56]  & \[2687] ,
  \[174]  = ~\[4]  & ~v1,
  \[13]  = ~\[171]  | (~\[74]  | v7),
  \[368]  = \[56]  & \[2669] ,
  \[14]  = \[5]  | \[3] ,
  \[91]  = \[79]  & \[8415] ,
  \[13244]  = \[77]  & \[56] ,
  \[15]  = v7 | ~v6,
  \[463]  = \[83]  & \[64] ,
  \[92]  = \[79]  & \[8397] ,
  \[270]  = ~\[18]  & \[8433] ,
  \[464]  = \[83]  & ~\[13] ,
  \[93]  = \[79]  & \[75] ,
  \[10110]  = (~\[119]  & ~v2) | ((~\[99]  & ~\[63] ) | (\[87]  & ~\[63] )),
  \[2723]  = \[159]  & \[47] ,
  \[17]  = v10 | ~v8,
  \[465]  = \[83]  & \[2723] ,
  \[13348]  = (\[115]  & \[65] ) | (\[100]  & \[56] ),
  \[94]  = \[79]  & \[73] ,
  \[18]  = \[10]  | \[3] ,
  \[95]  = \[79]  & \[66] ,
  \[96]  = \[84]  & \[79] ,
  \[97]  = \[79]  & \[5667] ,
  \[98]  = \[172]  & ~\[8] ,
  \[100]  = \[46]  & v0,
  \[99]  = v14 | v13,
  \[101]  = \[51]  & \[47] ,
  \[102]  = \[74]  & \[51] ,
  \[373]  = \[75]  & \[56] ,
  \[103]  = \[111]  & \[64] ,
  \[374]  = \[73]  & \[56] ,
  \[104]  = \[111]  & ~\[13] ,
  \[181]  = \[101]  & \[57] ,
  \[375]  = \[66]  & \[56] ,
  \[105]  = \[111]  & \[2723] ,
  \[106]  = (\[2]  & \[1] ) | \[69] ,
  \[183]  = \[64]  & \[57] ,
  \[10095]  = \[107]  & (~v2 & ~v1),
  \[107]  = \[114]  | \[78] ,
  \[184]  = \[57]  & ~\[13] ,
  \[23]  = v11 & v8,
  \[108]  = (\[2]  & ~v13) | \[87] ,
  \[185]  = 0,
  \[24]  = \[9]  | \[8] ,
  \[109]  = ~\[17]  & \[11] ,
  \[187]  = \[57]  & \[2687] ,
  \[26]  = (~\[131]  & ~\[1537] ) | (\[14]  | ~v9),
  \[474]  = \[83]  & \[73] ,
  \[27]  = ~\[4]  & v4,
  \[475]  = \[83]  & \[66] ,
  \[12822]  = \[85]  & \[72] ,
  \[28]  = ~\[85]  | \[18] ,
  \[476]  = \[84]  & \[83] ,
  \[300]  = \[173]  & \[1559] ,
  \[29]  = ~\[77]  | \[24] ,
  \[13063]  = \[109]  & \[50] ,
  \[477]  = \[83]  & \[5667] ,
  \[301]  = \[173]  & \[1537] ,
  \[302]  = \[102]  & \[67] ,
  \[303]  = \[67]  & \[64] ,
  \[110]  = \[46]  & \[6] ,
  \[1241]  = (~\[136]  & (~\[118]  & (~\[101]  & (~\[85]  & ~\[54] )))) | ((~\[132]  & (\[54]  & ~\[35] )) | (\[54]  & \[24] )),
  \[287]  = \[81]  & \[2687] ,
  \[304]  = \[67]  & ~\[13] ,
  \[111]  = ~\[17]  & ~\[8] ,
  \[288]  = \[81]  & \[2669] ,
  \[305]  = \[67]  & \[2723] ,
  \[112]  = ~v3 | v1,
  \[289]  = \[81]  & \[6571] ,
  \[10319]  = (\[114]  & (~\[15]  & ~v5)) | ((\[106]  & (~\[15]  & ~v5)) | ((\[147]  & \[113] ) | ((\[147]  & ~\[99] ) | ((\[147]  & \[69] ) | ((~\[130]  & \[114] ) | (~\[130]  & \[106] )))))),
  \[113]  = (\[1]  & v15) | \[49] ,
  \[307]  = \[67]  & \[2687] ,
  \[114]  = ~\[2]  & ~\[1] ,
  \[308]  = \[67]  & \[2669] ,
  \[115]  = (\[62]  & \[47] ) | \[146] ,
  \[672]  = (~\[136]  & (~\[117]  & (~\[100]  & (~\[77]  & (~\[52]  & (~\[40]  & ~\[2669] )))))) | ((~\[100]  & \[58] ) | (~\[82]  & \[58] )),
  \[403]  = \[82]  & \[64] ,
  \[193]  = \[75]  & \[57] ,
  \[32]  = \[15]  | ~v4,
  \[5689]  = \[171]  & \[169] ,
  \[117]  = (\[36]  & \[6] ) | \[66] ,
  \[404]  = \[82]  & ~\[13] ,
  \[194]  = \[73]  & \[57] ,
  \[33]  = ~\[7]  & ~\[5] ,
  \[118]  = \[43]  | \[8433] ,
  \[10123]  = \[113]  & ~\[63] ,
  \[405]  = \[82]  & \[2723] ,
  \[195]  = \[66]  & \[57] ,
  \[34]  = \[32]  | \[7] ,
  \[119]  = \[48]  | v1,
  \[35]  = \[84]  | \[5667] ,
  \[1537]  = \[100]  & ~v8,
  \[213]  = \[80]  & \[75] ,
  \[36]  = \[27]  & ~v6,
  \[214]  = \[80]  & \[73] ,
  \[215]  = \[80]  & \[66] ,
  \[216]  = \[84]  & \[80] ,
  \[293]  = \[81]  & \[75] ,
  \[39]  = \[8397]  | \[8415] ,
  \[218]  = 0,
  \[313]  = \[75]  & \[67] ,
  \[120]  = \[46]  & ~v1,
  \[314]  = \[73]  & \[67] ,
  \[121]  = \[111]  & \[100] ,
  \[298]  = 0,
  \[5711]  = \[174]  & \[171] ,
  \[315]  = \[67]  & \[66] ,
  \[299]  = \[101]  & \[67] ,
  \[10516]  = (\[114]  & (~\[62]  & \[45] )) | ((\[107]  & (~\[6]  & ~\[4] )) | ((\[106]  & (~\[62]  & \[45] )) | ((\[106]  & (~\[6]  & ~\[4] )) | ((\[145]  & \[79] ) | (\[115]  & \[79] ))))),
  \[393]  = \[75]  & \[65] ,
  \[123]  = \[64]  & ~\[24] ,
  \[394]  = \[73]  & \[65] ,
  \[124]  = ~\[24]  & ~\[13] ,
  \[40]  = \[2687]  | \[2705] ,
  \[395]  = \[66]  & \[65] ,
  \[125]  = 0,
  \[12359]  = (\[115]  & \[81] ) | ((\[110]  & ~\[18] ) | (\[81]  & \[52] )),
  \[41]  = \[39]  | \[8433] ,
  \[1063]  = (~\[132]  & (~\[55]  & (~\[53]  & ~\[50] ))) | \[76] ,
  \[396]  = \[84]  & \[65] ,
  \[127]  = ~\[24]  & \[2687] ,
  \[971]  = (~\[39]  & (~\[36]  & (~\[5649]  & (~\[5667]  & (~\[5689]  & (~\[5711]  & ~\[12359] )))))) | ((~\[39]  & (~\[6]  & (~\[5649]  & (~\[5667]  & (~\[5689]  & (~\[5711]  & ~\[12359] )))))) | ((~\[39]  & (~\[36]  & (~\[5649]  & (~\[5667]  & (~\[12359]  & v7))))) | ((~\[39]  & (~\[6]  & (~\[5649]  & (~\[5667]  & (~\[12359]  & v7))))) | (\[18]  & ~\[12359] )))),
  \[43]  = \[2669]  | \[6571] ,
  \[11539]  = \[143]  & \[57] ,
  \[129]  = \[51]  & \[4] ,
  \[45]  = v5 & ~v4,
  \[223]  = ~\[76]  & \[64] ,
  \[46]  = \[27]  & v7,
  \[224]  = ~\[76]  & ~\[13] ,
  \[10693]  = \[111]  & \[53] ,
  \[47]  = ~\[6]  & ~v2,
  \[48]  = v14 | ~v12,
  \[49]  = (~\[7]  & v11) | (~\[5]  & v8),
  \[130]  = ~\[6]  | ~v3,
  \[14213]  = \[83]  & \[53] ,
  \[13103]  = \[109]  & \[55] ,
  \[131]  = \[1559]  | \[1581] ,
  \[132]  = \[110]  | \[5649] ,
  \[12848]  = \[118]  & \[72] ,
  \[12745]  = (\[131]  & \[67] ) | (\[67]  & \[35] ),
  \[133]  = \[75]  & ~\[24] ,
  \[10795]  = (\[111]  & \[55] ) | ((\[101]  & ~\[24] ) | (\[89]  & ~\[8] )),
  \[134]  = \[73]  & ~\[24] ,
  \[50]  = \[75]  | \[41] ,
  \[135]  = \[66]  & ~\[24] ,
  \[51]  = v7 & v4,
  \[136]  = \[102]  | \[64] ,
  \[52]  = ~\[13]  | \[2723] ,
  \[11641]  = \[145]  & \[80] ,
  \[53]  = \[43]  | \[40] ,
  \[54]  = \[12]  | \[9] ,
  \[10626]  = \[59]  & ~\[8] ,
  \[55]  = \[73]  | (\[66]  | \[35] ),
  \[10728]  = \[111]  & \[50] ,
  \[56]  = \[11]  & ~\[9] ,
  \[2669]  = \[74]  & (~v6 & v4),
  \[57]  = ~\[10]  & ~\[8] ,
  \[1559]  = \[120]  & ~v8,
  \[58]  = \[17]  | \[3] ,
  \[59]  = (\[146]  & ~\[17] ) | (\[110]  & \[23] ),
  \[794]  = (\[26]  & (~\[456]  & (~\[455]  & (~\[454]  & (~\[453]  & (~\[464]  & (~\[463]  & (~\[465]  & (~\[14132]  & (~\[14256]  & (~\[14213]  & (~\[476]  & (~\[475]  & (~\[474]  & (~\[443]  & (~\[442]  & (~\[441]  & (~\[440]  & (~\[439]  & (~\[436]  & (~\[449]  & (~\[448]  & (~\[13963]  & (\[672]  & (~\[2705]  & (~\[396]  & (~\[395]  & (~\[394]  & (~\[393]  & (~\[404]  & (~\[403]  & (~\[405]  & (~\[13525]  & (~\[13627]  & (~\[13592]  & (~\[13694]  & (~\[368]  & (~\[367]  & (~\[365]  & (~\[364]  & (~\[363]  & (~\[362]  & (~\[361]  & (~\[374]  & (~\[373]  & (~\[375]  & (~\[13244]  & (~\[13412]  & (~\[13386]  & (~\[13348]  & (~\[13311]  & (~\[5649]  & (~\[5667]  & (~\[8397]  & (~\[8415]  & ~\[8433] ))))))))))))))))))))))))))))))))))))))))))))))))))))))) | (~\[65]  & (~\[61]  & (\[58]  & (~\[56]  & (\[26]  & (~\[464]  & (~\[463]  & (~\[465]  & (~\[14132]  & (~\[14256]  & (~\[14213]  & (~\[477]  & (~\[476]  & (~\[475]  & (~\[474]  & (\[672]  & (~\[404]  & (~\[403]  & (~\[405]  & (~\[13525]  & (~\[13627]  & (~\[13592]  & (~\[13694]  & ~\[361] ))))))))))))))))))))))),
  \[14132]  = (\[86]  & (\[11]  & \[1559] )) | ((\[86]  & (\[11]  & \[1537] )) | (\[146]  & \[83] )),
  \[333]  = \[75]  & \[72] ,
  \[1464]  = (~\[114]  & (~\[87]  & ~\[2] )) | ((~\[87]  & (\[32]  & v13)) | ((~\[32]  & (\[2]  & ~\[1] )) | (\[112]  & \[32] ))),
  \[334]  = \[73]  & \[72] ,
  \[13386]  = \[85]  & \[65] ,
  \[335]  = \[72]  & \[66] ,
  \[1273]  = (~\[102]  & (\[29]  & (~\[2669]  & (~\[2705]  & (~\[2723]  & (~\[5649]  & (~\[5667]  & (~\[216]  & (~\[215]  & (~\[214]  & (~\[213]  & (~\[224]  & (~\[223]  & (~\[11753]  & (\[1063]  & (~\[187]  & (~\[184]  & (~\[183]  & (~\[181]  & (~\[194]  & (~\[193]  & (~\[195]  & (~\[11472]  & (~\[11576]  & (~\[11539]  & (~\[11641]  & (~\[156]  & (~\[155]  & (~\[154]  & (~\[153]  & (~\[164]  & (~\[163]  & (~\[11190]  & (\[1182]  & (~\[127]  & (~\[124]  & (~\[123]  & (~\[121]  & (~\[134]  & (~\[133]  & (~\[135]  & (~\[8397]  & (~\[8415]  & \[1241] ))))))))))))))))))))))))))))))))))))))))))) | (~\[80]  & (\[76]  & (~\[57]  & (\[54]  & (\[24]  & (~\[164]  & (~\[163]  & (~\[165]  & (~\[11190]  & (\[1182]  & ~\[121] )))))))))),
  \[336]  = \[84]  & \[72] ,
  \[143]  = \[88]  | \[35] ,
  \[13311]  = \[143]  & \[56] ;
endmodule

