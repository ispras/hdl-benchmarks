// IWLS benchmark module "cht" printed on Wed May 29 16:31:27 2002
module cht(a, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, \x , y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, r0, s0, t0, u0, v0, w0, x0, y0, z0, a1, b1, c1, d1, e1, f1, g1, h1, i1, j1, k1, l1, m1, n1, o1, p1, q1, r1, s1, t1, u1, v1, w1, x1, y1, z1, a2, b2, c2, d2, e2, f2);
input
  a,
  c,
  d,
  e,
  f,
  g,
  h,
  i,
  j,
  k,
  l,
  m,
  n,
  o,
  p,
  q,
  r,
  s,
  t,
  u,
  v,
  w,
  \x ,
  y,
  z,
  a0,
  b0,
  c0,
  d0,
  e0,
  f0,
  g0,
  h0,
  i0,
  j0,
  k0,
  l0,
  m0,
  n0,
  o0,
  p0,
  q0,
  r0,
  s0,
  t0,
  u0,
  v0;
output
  a1,
  a2,
  b1,
  b2,
  c1,
  c2,
  d1,
  d2,
  e1,
  e2,
  f1,
  f2,
  g1,
  h1,
  i1,
  j1,
  k1,
  l1,
  m1,
  n1,
  o1,
  p1,
  q1,
  r1,
  s1,
  t1,
  u1,
  v1,
  w0,
  w1,
  x0,
  x1,
  y0,
  y1,
  z0,
  z1;
wire
  \[5] ,
  \[6] ,
  \[7] ,
  \[8] ,
  \[9] ,
  \[20] ,
  \[21] ,
  \[22] ,
  \[23] ,
  \[24] ,
  \[25] ,
  \[26] ,
  \[27] ,
  \[28] ,
  \[29] ,
  \[30] ,
  \[31] ,
  \[32] ,
  \[33] ,
  \[34] ,
  \[35] ,
  \[10] ,
  \[11] ,
  \[12] ,
  \[13] ,
  \[14] ,
  \[15] ,
  \[0] ,
  \[16] ,
  \[1] ,
  \[17] ,
  \[2] ,
  \[18] ,
  \[3] ,
  \[19] ,
  \[4] ;
assign
  \[5]  = (e & (r & ~l)) | ((e & (~l & i)) | (r & (~l & ~i))),
  \[6]  = (s & (t & ~l)) | ((s & (~l & ~j)) | (t & (~l & j))),
  \[7]  = (t & (u & ~l)) | ((t & (~l & ~j)) | (u & (~l & j))),
  \[8]  = (u & (v & ~l)) | ((u & (~l & ~j)) | (v & (~l & j))),
  \[9]  = (v & (w & ~l)) | ((v & (~l & ~j)) | (w & (~l & j))),
  \[20]  = (g0 & (h0 & ~l)) | ((g0 & (~l & ~k)) | (h0 & (~l & k))),
  \[21]  = (h0 & (i0 & ~l)) | ((h0 & (~l & ~k)) | (i0 & (~l & k))),
  \[22]  = (i0 & (j0 & ~l)) | ((i0 & (~l & ~k)) | (j0 & (~l & k))),
  \[23]  = (j0 & (k0 & ~l)) | ((j0 & (~l & ~k)) | (k0 & (~l & k))),
  \[24]  = (k0 & (l0 & ~l)) | ((k0 & (~l & ~k)) | (l0 & (~l & k))),
  \[25]  = (l0 & (m0 & ~l)) | ((l0 & (~l & ~k)) | (m0 & (~l & k))),
  \[26]  = (m0 & (n0 & ~l)) | ((m0 & (~l & ~k)) | (n0 & (~l & k))),
  \[27]  = (o0 & (n0 & (~p & ~l))) | ((o0 & (n0 & (~l & a))) | ((o0 & (~p & (~l & k))) | ((o0 & (~l & (k & a))) | ((n0 & (p & (~l & a))) | ((p & (~l & (k & a))) | (n0 & (~l & ~k))))))),
  \[28]  = (p0 & (~p & (~l & k))) | ((p0 & (o0 & ~l)) | ((o0 & (p & ~l)) | (o0 & (~l & ~k)))),
  \[29]  = (q0 & (~p & (~l & k))) | ((q0 & (p0 & ~l)) | ((p0 & (p & ~l)) | (p0 & (~l & ~k)))),
  a1 = \[4] ,
  a2 = \[30] ,
  b1 = \[5] ,
  b2 = \[31] ,
  c1 = \[6] ,
  c2 = \[32] ,
  d1 = \[7] ,
  d2 = \[33] ,
  e1 = \[8] ,
  e2 = \[34] ,
  f1 = \[9] ,
  f2 = \[35] ,
  g1 = \[10] ,
  \[30]  = (r0 & (~p & (~l & k))) | ((r0 & (q0 & ~l)) | ((q0 & (p & ~l)) | (q0 & (~l & ~k)))),
  h1 = \[11] ,
  \[31]  = (s0 & (~p & (~l & k))) | ((s0 & (r0 & ~l)) | ((r0 & (p & ~l)) | (r0 & (~l & ~k)))),
  i1 = \[12] ,
  \[32]  = (t0 & (~p & (~l & k))) | ((t0 & (s0 & ~l)) | ((s0 & (p & ~l)) | (s0 & (~l & ~k)))),
  j1 = \[13] ,
  \[33]  = (u0 & (~p & (~l & k))) | ((u0 & (t0 & ~l)) | ((t0 & (p & ~l)) | (t0 & (~l & ~k)))),
  k1 = \[14] ,
  \[34]  = (v0 & (~p & (~l & k))) | ((v0 & (u0 & ~l)) | ((u0 & (p & ~l)) | (u0 & (~l & ~k)))),
  l1 = \[15] ,
  \[35]  = (~p & (~l & (k & a))) | ((v0 & (p & ~l)) | ((v0 & (~l & ~k)) | (v0 & (~l & a)))),
  m1 = \[16] ,
  n1 = \[17] ,
  o1 = \[18] ,
  p1 = \[19] ,
  q1 = \[20] ,
  \[10]  = (w & (\x  & ~l)) | ((w & (~l & ~j)) | (\x  & (~l & j))),
  r1 = \[21] ,
  \[11]  = (\x  & (y & ~l)) | ((\x  & (~l & ~j)) | (y & (~l & j))),
  s1 = \[22] ,
  \[12]  = (y & (z & ~l)) | ((y & (~l & ~j)) | (z & (~l & j))),
  t1 = \[23] ,
  \[13]  = (z & (a0 & ~l)) | ((z & (~l & ~j)) | (a0 & (~l & j))),
  u1 = \[24] ,
  \[14]  = (a0 & (b0 & ~l)) | ((a0 & (~l & ~j)) | (b0 & (~l & j))),
  v1 = \[25] ,
  \[15]  = (b0 & (c0 & ~l)) | ((b0 & (~l & ~j)) | (c0 & (~l & j))),
  \[0]  = (f & (m & ~l)) | ((f & (~l & i)) | (m & (~l & ~i))),
  w0 = \[0] ,
  w1 = \[26] ,
  \[16]  = (c0 & (d0 & ~l)) | ((c0 & (~l & ~j)) | (d0 & (~l & j))),
  \[1]  = (g & (n & ~l)) | ((g & (~l & i)) | (n & (~l & ~i))),
  x0 = \[1] ,
  x1 = \[27] ,
  \[17]  = (d0 & (e0 & ~l)) | ((d0 & (~l & ~j)) | (e0 & (~l & j))),
  \[2]  = (h & (o & ~l)) | ((h & (~l & i)) | (o & (~l & ~i))),
  y0 = \[2] ,
  y1 = \[28] ,
  \[18]  = (e0 & (f0 & ~l)) | ((e0 & (~l & ~j)) | (f0 & (~l & j))),
  \[3]  = (c & (p & ~l)) | ((c & (~l & i)) | (p & (~l & ~i))),
  z0 = \[3] ,
  z1 = \[29] ,
  \[19]  = (a & (f0 & ~l)) | ((a & (~l & j)) | (f0 & (~l & ~j))),
  \[4]  = (d & (q & ~l)) | ((d & (~l & i)) | (q & (~l & ~i)));
endmodule

