//NOTE: no-implementation module stub

module GTECH_AND3 (
    output Z,
    input A,
    input B,
    input C
);

endmodule
