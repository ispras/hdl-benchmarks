// IWLS benchmark module "dalu" printed on Wed May 29 16:31:30 2002
module dalu(inA15, inA14, inA13, inA12, inA11, inA10, inA9, inA8, inA7, inA6, inA5, inA4, inA3, inA2, inA1, inA0, inB15, inB14, inB13, inB12, inB11, inB10, inB9, inB8, inB7, inB6, inB5, inB4, inB3, inB2, inB1, inB0, inC15, inC14, inC13, inC12, inC11, inC10, inC9, inC8, inC7, inC6, inC5, inC4, inC3, inC2, inC1, inC0, inD15, inD14, inD13, inD12, inD11, inD10, inD9, inD8, inD7, inD6, inD5, inD4, inD3, inD2, inD1, inD0, opsel3, opsel2, opsel1, opsel0, musel4, musel3, musel2, musel1, sh2, sh1, sh0, O15, O14, O13, O12, O11, O10, O9, O8, O7, O6, O5, O4, O3, O2, O1, O0);
input
  inA10,
  inA11,
  inA12,
  inA13,
  inA14,
  inA15,
  inB10,
  inB11,
  inB12,
  inB13,
  inB14,
  inB15,
  inC10,
  inC11,
  inC12,
  inC13,
  inC14,
  inC15,
  inD10,
  inD11,
  inD12,
  inD13,
  inD14,
  inD15,
  inA0,
  inA1,
  inA2,
  inA3,
  inA4,
  inA5,
  inA6,
  inA7,
  inA8,
  inA9,
  inB0,
  inB1,
  inB2,
  inB3,
  inB4,
  inB5,
  inB6,
  inB7,
  inB8,
  inB9,
  inC0,
  inC1,
  inC2,
  inC3,
  inC4,
  inC5,
  inC6,
  inC7,
  inC8,
  inC9,
  inD0,
  inD1,
  inD2,
  inD3,
  inD4,
  inD5,
  inD6,
  inD7,
  inD8,
  inD9,
  sh0,
  sh1,
  sh2,
  musel1,
  musel2,
  musel3,
  musel4,
  opsel0,
  opsel1,
  opsel2,
  opsel3;
output
  O0,
  O1,
  O2,
  O3,
  O4,
  O5,
  O6,
  O7,
  O8,
  O9,
  O10,
  O11,
  O12,
  O13,
  O14,
  O15;
wire
  \[5893] ,
  \[378] ,
  \[189] ,
  \[5894] ,
  \[569] ,
  \[8520] ,
  \[8521] ,
  \[6055] ,
  \[9880] ,
  \[6056] ,
  \[4349] ,
  \[5897] ,
  \[5898] ,
  \[10744] ,
  \[8714] ,
  \[8335] ,
  \[9883] ,
  \[8905] ,
  \[10556] ,
  \[190] ,
  \[8337] ,
  \[570] ,
  \[950] ,
  \[381] ,
  \[9886] ,
  \[8908] ,
  \[382] ,
  \[11100] ,
  \[2642] ,
  \[10372] ,
  \[193] ,
  \[383] ,
  \[4540] ,
  \[194] ,
  \[384] ,
  \[4352] ,
  \[2645] ,
  \[575] ,
  \[576] ,
  \[6061] ,
  \[197] ,
  \[6062] ,
  \[198] ,
  \[6063] ,
  \[199] ,
  \[8530] ,
  \[8911] ,
  \[6065] ,
  \[6066] ,
  \[10944] ,
  \[8914] ,
  \[0] ,
  \[10946] ,
  \[1] ,
  \[8726] ,
  \[2] ,
  \[8917] ,
  \[10570] ,
  \[391] ,
  \[581] ,
  \[3] ,
  \[8349] ,
  \[582] ,
  \[4] ,
  \[1105] ,
  \[5] ,
  \[11302] ,
  \[6] ,
  \[1107] ,
  \[7] ,
  \[8] ,
  \[6071] ,
  \[587] ,
  \[9] ,
  \[6072] ,
  \[588] ,
  \[6073] ,
  \[399] ,
  \[8540] ,
  \[969] ,
  \[8920] ,
  \[6074] ,
  \[11308] ,
  \[8541] ,
  \[6075] ,
  \[8923] ,
  \[10764] ,
  \[8926] ,
  \[10960] ,
  \[11310] ,
  \[8549] ,
  \[782] ,
  \[8929] ,
  \[1115] ,
  \[593] ,
  \[594] ,
  \[6080] ,
  \[6081] ,
  \[6082] ,
  \[10588] ,
  \[8360] ,
  \[599] ,
  \[8361] ,
  \[11318] ,
  \[8741] ,
  \[8932] ,
  \[6086] ,
  \[6087] ,
  \[8935] ,
  \[10396] ,
  \[1501] ,
  \[1312] ,
  \[11316] ,
  \[1502] ,
  \[11506] ,
  \[8938] ,
  \[3404] ,
  \[4954] ,
  \[6092] ,
  \[5304] ,
  \[6093] ,
  \[10978] ,
  \[799] ,
  \[6094] ,
  \[8181] ,
  \[8941] ,
  \[8372] ,
  \[8562] ,
  \[9101] ,
  \[8563] ,
  \[6097] ,
  \[8754] ,
  \[8944] ,
  \[6098] ,
  \[8185] ,
  \[1130] ,
  \[11324] ,
  \[10786] ,
  \[1511] ,
  \[2490] ,
  \[11326] ,
  \[1512] ,
  \[8947] ,
  \[3600] ,
  G3,
  \[2493] ,
  \[1136] ,
  \[11332] ,
  \[4392] ,
  \[1517] ,
  \[1329] ,
  \[1519] ,
  \[4965] ,
  \[3228] ,
  \[8570] ,
  \[8950] ,
  \[11908] ,
  \[4968] ,
  \[9301] ,
  \[8952] ,
  \[8953] ,
  \[8195] ,
  \[11334] ,
  \[1520] ,
  \[8955] ,
  \[1331] ,
  \[8956] ,
  \[11146] ,
  \[1332] ,
  \[8767] ,
  \[8388] ,
  \[9117] ,
  \[8389] ,
  \[3231] ,
  \[11340] ,
  \[8959] ,
  \[11910] ,
  \[4780] ,
  \[1525] ,
  \[9119] ,
  \[11342] ,
  \[1526] ,
  \[1337] ,
  \[5701] ,
  \[1338] ,
  \[5514] ,
  \[5704] ,
  \[10998] ,
  \[5705] ,
  \[11348] ,
  \[11728] ,
  \[8961] ,
  \[5517] ,
  \[8962] ,
  \[9312] ,
  \[5708] ,
  b0,
  b1,
  b2,
  b3,
  b4,
  b5,
  b6,
  b7,
  b8,
  b9,
  \[8964] ,
  \[9314] ,
  \[8965] ,
  \[1910] ,
  \[8586] ,
  e0,
  e1,
  e2,
  e3,
  e5,
  \[8587] ,
  e6,
  e7,
  \[8777] ,
  e9,
  \[11726] ,
  \[8967] ,
  \[8968] ,
  \[1913] ,
  \[9507] ,
  \[11350] ,
  \[11920] ,
  \[1535] ,
  \[11922] ,
  \[5900] ,
  \[1347] ,
  \[1537] ,
  \[1538] ,
  \[5712] ,
  \[1349] ,
  \[3626] ,
  \[5523] ,
  \[5713] ,
  \[5903] ,
  \[5524] ,
  \[5904] ,
  \[5525] ,
  \[5905] ,
  \[11358] ,
  \[9130] ,
  \[8781] ,
  \[3629] ,
  \[8971] ,
  \[9511] ,
  \[8593] ,
  \[9132] ,
  \[5528] ,
  \[8973] ,
  \[5908] ,
  \[5529] ,
  \[8974] ,
  \[5719] ,
  \[9513] ,
  \[5909] ,
  \[1350] ,
  \[11544] ,
  \[8976] ,
  \[11166] ,
  \[11356] ,
  \[11546] ,
  \[8977] ,
  \[1353] ,
  \[1543] ,
  \[202] ,
  \[9707] ,
  \[1354] ,
  \[1544] ,
  \[8979] ,
  \[203] ,
  \[204] ,
  \[1356] ,
  \[1167] ,
  \[5911] ,
  \[5722] ,
  \[207] ,
  \[5533] ,
  \[5723] ,
  \[208] ,
  \[5913] ,
  \[5534] ,
  \[209] ,
  \[8790] ,
  \[5535] ,
  \[8980] ,
  \[5156] ,
  \[5536] ,
  \[5726] ,
  \[5916] ,
  \[5537] ,
  \[9331] ,
  \[5917] ,
  \[9711] ,
  \[9901] ,
  b10,
  b11,
  b12,
  \[8983] ,
  b13,
  b14,
  b15,
  \[5918] ,
  \[9143] ,
  \[9523] ,
  \[9713] ,
  \[11364] ,
  \[8985] ,
  \[1361] ,
  \[9145] ,
  \[9335] ,
  \[8986] ,
  \[210] ,
  \[9905] ,
  \[11366] ,
  \[1363] ,
  \[1553] ,
  \[9337] ,
  \[8988] ,
  \[9527] ,
  \[11180] ,
  \[1364] ,
  \[8989] ,
  \[213] ,
  \[1555] ,
  \[9529] ,
  \[214] ,
  \[9719] ,
  \[11372] ,
  \[1556] ,
  \[5730] ,
  \[5731] ,
  \[5921] ,
  \[5542] ,
  \[217] ,
  \[5922] ,
  \[3076] ,
  \[1369] ,
  \[5543] ,
  \[218] ,
  \[219] ,
  \[5924] ,
  \[3079] ,
  \[8991] ,
  \[8992] ,
  \[5737] ,
  \[5927] ,
  \[9721] ,
  \[9911] ,
  \[10204] ,
  \[5928] ,
  \[10013] ,
  \[5549] ,
  \[8994] ,
  \[5929] ,
  \[9913] ,
  \[1370] ,
  \[11374] ,
  \[10015] ,
  \[1561] ,
  \[600] ,
  \[1562] ,
  \[9156] ,
  \[10400] ,
  \[411] ,
  \[3270] ,
  \[9347] ,
  \[222] ,
  \[11380] ,
  \[11760] ,
  \[223] ,
  \[9728] ,
  \[9539] ,
  \[224] ,
  \[11382] ,
  \[5550] ,
  \[11762] ,
  \[5740] ,
  \[605] ,
  \[1567] ,
  \[5551] ,
  \[5741] ,
  \[606] ,
  \[1568] ,
  \[227] ,
  \[5932] ,
  \[1379] ,
  \[228] ,
  \[5933] ,
  \[5554] ,
  \[5744] ,
  \[229] ,
  \[5555] ,
  \[5935] ,
  \[11388] ,
  \[11578] ,
  \[5556] ,
  \[9920] ,
  \[10029] ,
  \[9161] ,
  \[9351] ,
  \[5937] ,
  \[9731] ,
  \[5748] ,
  \[5559] ,
  \[9353] ,
  \[5749] ,
  \[9543] ,
  \[5939] ,
  \[1190] ,
  \[9923] ,
  \[1381] ,
  \[10025] ,
  \[9165] ,
  \[9545] ,
  \[230] ,
  \[11196] ,
  \[1382] ,
  \[611] ,
  \[612] ,
  \[11390] ,
  \[11580] ,
  \[233] ,
  \[423] ,
  \[10031] ,
  \[9169] ,
  \[234] ,
  \[424] ,
  \[11772] ,
  \[425] ,
  \[1387] ,
  \[1577] ,
  \[426] ,
  \[1388] ,
  \[237] ,
  \[617] ,
  \[1579] ,
  \[5563] ,
  \[238] ,
  \[618] ,
  \[5564] ,
  \[6103] ,
  \[239] ,
  \[10608] ,
  \[6104] ,
  \[5755] ,
  \[5945] ,
  \[11398] ,
  \[6105] ,
  \[5946] ,
  \[9740] ,
  \[9171] ,
  \[5947] ,
  \[9741] ,
  \[5378] ,
  e10,
  \[10224] ,
  e11,
  e13,
  \[6107] ,
  \[10414] ,
  e14,
  \[5758] ,
  e15,
  \[5948] ,
  \[9932] ,
  \[9363] ,
  \[6108] ,
  \[9743] ,
  \[9933] ,
  \[1580] ,
  \[11774] ,
  \[9555] ,
  \[9935] ,
  \[11396] ,
  \[1772] ,
  \[9367] ,
  \[242] ,
  \[432] ,
  \[243] ,
  \[623] ,
  \[1775] ,
  \[9369] ,
  \[9559] ,
  \[244] ,
  \[9749] ,
  \[624] ,
  \[5570] ,
  \[5760] ,
  \[5950] ,
  \[1397] ,
  \[5951] ,
  \[247] ,
  \[5952] ,
  \[1399] ,
  \[1589] ,
  \[5573] ,
  \[5763] ,
  \[248] ,
  \[438] ,
  \[10048] ,
  \[5574] ,
  \[6113] ,
  \[5764] ,
  \[249] ,
  \[6114] ,
  \[5955] ,
  \[6115] ,
  \[11978] ,
  \[5956] ,
  \[5577] ,
  \[5767] ,
  \[9561] ,
  \[5957] ,
  \[9941] ,
  \[10044] ,
  \[9182] ,
  \[6117] ,
  \[9753] ,
  \[10046] ,
  \[9184] ,
  pgx3,
  \[1591] ,
  \[9755] ,
  \[9945] ,
  \[10050] ,
  \[1592] ,
  \[11976] ,
  \[441] ,
  \[631] ,
  \[252] ,
  \[9757] ,
  \[9947] ,
  \[10432] ,
  \[9379] ,
  \[9759] ,
  \[9949] ,
  \[4222] ,
  \[255] ,
  \[1597] ,
  \[5581] ,
  \[5771] ,
  \[256] ,
  \[1598] ,
  \[5582] ,
  \[5772] ,
  \[5962] ,
  \[258] ,
  \[5963] ,
  \[10058] ,
  \[11988] ,
  \[5966] ,
  \[9760] ,
  \[9571] ,
  \[5967] ,
  \[9951] ,
  \[10244] ,
  \[5588] ,
  \[5778] ,
  \[9952] ,
  \[9383] ,
  \[5969] ,
  \[9763] ,
  \[8405] ,
  \[10056] ,
  \[9195] ,
  \[9385] ,
  \[9575] ,
  \[9955] ,
  \[10060] ,
  \[10630] ,
  \[9766] ,
  \[9197] ,
  \[9577] ,
  \[10062] ,
  \[11990] ,
  \[263] ,
  \[10632] ,
  \[9958] ,
  \[264] ,
  \[5970] ,
  \[835] ,
  \[5591] ,
  \[5781] ,
  \[266] ,
  \[5592] ,
  \[5782] ,
  \[10068] ,
  \[10258] ,
  \[5595] ,
  \[5785] ,
  \[5975] ,
  \[5976] ,
  \[5977] ,
  \[5978] ,
  \[9772] ,
  \[5599] ,
  \[5789] ,
  \[5979] ,
  \[9964] ,
  \[9395] ,
  \[10070] ,
  \[271] ,
  \[9776] ,
  \[8418] ,
  \[10830] ,
  \[272] ,
  \[8419] ,
  \[10072] ,
  \[10452] ,
  \[9778] ,
  \[9968] ,
  \[9399] ,
  \[274] ,
  \[9779] ,
  \[464] ,
  \[5790] ,
  \[5980] ,
  \[465] ,
  \[5981] ,
  \[466] ,
  \[5982] ,
  \[467] ,
  \[468] ,
  \[279] ,
  \[8611] ,
  \[5796] ,
  \[9970] ,
  \[8612] ,
  \[8802] ,
  \[5987] ,
  \[9971] ,
  \[10074] ,
  \[5988] ,
  \[9782] ,
  \[5799] ,
  \[10646] ,
  \[9974] ,
  \[280] ,
  \[10080] ,
  \[661] ,
  \[2352] ,
  \[282] ,
  \[8619] ,
  \[10082] ,
  \[2355] ,
  \[5990] ,
  \[287] ,
  \[5992] ,
  \[667] ,
  \[288] ,
  \[5993] ,
  \[10468] ,
  \[5994] ,
  \[8430] ,
  \[10084] ,
  \[5998] ,
  \[10086] ,
  \[10276] ,
  \[290] ,
  \[480] ,
  \[8817] ,
  \[10850] ,
  \[8628] ,
  \[10092] ,
  \[1005] ,
  \[483] ,
  \[4640] ,
  \[484] ,
  \[295] ,
  \[865] ,
  \[296] ,
  \[298] ,
  \[2938] ,
  \[10098] ,
  \[489] ,
  \[8440] ,
  \[11018] ,
  \[8441] ,
  \[10094] ,
  \[10474] ,
  \[8254] ,
  \[10664] ,
  \[11014] ,
  \[1200] ,
  \[11204] ,
  \[10096] ,
  \[10476] ,
  \[2941] ,
  \[11022] ,
  \[875] ,
  \[496] ,
  \[4466] ,
  \[10868] ,
  \[8640] ,
  \[8830] ,
  \[8451] ,
  \[8263] ,
  \[5008] ,
  \[11024] ,
  \[1400] ,
  \[11404] ,
  \[10296] ,
  \[11026] ,
  \[11406] ,
  \[10870] ,
  \[1405] ,
  \[1406] ,
  \[11412] ,
  \[4663] ,
  \[697] ,
  \[4854] ,
  \[8270] ,
  \[4666] ,
  \[8271] ,
  \[11228] ,
  \[8274] ,
  \[10684] ,
  \[8464] ,
  \[8465] ,
  \[8655] ,
  \[1221] ,
  \[1411] ,
  \[11226] ,
  \[1412] ,
  \[1603] ,
  \[11040] ,
  \[11420] ,
  \[1604] ,
  \[8849] ,
  \[1035] ,
  \[11612] ,
  \[9012] ,
  \[10884] ,
  \[8475] ,
  \[11424] ,
  \[11614] ,
  \[8855] ,
  \[8286] ,
  \[1421] ,
  \[8287] ,
  \[11806] ,
  \[1423] ,
  \[1613] ,
  \[1424] ,
  \[9208] ,
  \[1045] ,
  \[1235] ,
  \[1615] ,
  \[3512] ,
  \[11242] ,
  \[12790] ,
  \[1616] ,
  \[5600] ,
  \[3515] ,
  \[10] ,
  \[11] ,
  \[12] ,
  \[13] ,
  \[8861] ,
  \[5606] ,
  \[14] ,
  \[9401] ,
  \[15] ,
  \[8673] ,
  \[9213] ,
  \[5609] ,
  \[11434] ,
  \[11624] ,
  \[12799] ,
  \[1431] ,
  \[1432] ,
  \[11626] ,
  \[8298] ,
  \[12793] ,
  \[9217] ,
  \[12796] ,
  \[1434] ,
  \[5610] ,
  \[5800] ,
  \[1627] ,
  \[1439] ,
  \[1629] ,
  \[5613] ,
  \[5803] ,
  \[8870] ,
  \[11068] ,
  \[8491] ,
  \[8492] ,
  \[9221] ,
  \[5617] ,
  \[9411] ,
  \[5807] ,
  \[5618] ,
  \[5808] ,
  \[9223] ,
  \[11254] ,
  \[1630] ,
  \[1441] ,
  \[9415] ,
  \[9605] ,
  \[1442] ,
  \[9417] ,
  \[1635] ,
  \[9609] ,
  \[11262] ,
  \[1636] ,
  \[1447] ,
  \[1448] ,
  \[5624] ,
  \[5814] ,
  \[3348] ,
  \[9040] ,
  \[5627] ,
  \[5817] ,
  \[9611] ,
  \[8693] ,
  \[5628] ,
  \[5818] ,
  \[8884] ,
  \[9234] ,
  \[9615] ,
  \[11456] ,
  \[9236] ,
  \[9427] ,
  \[9617] ,
  \[9807] ,
  \[11840] ,
  \[303] ,
  \[1075] ,
  \[304] ,
  \[11842] ,
  \[1457] ,
  \[5631] ,
  \[5821] ,
  \[306] ,
  \[1459] ,
  \[3736] ,
  \[10108] ,
  \[5635] ,
  \[5825] ,
  \[5256] ,
  \[5636] ,
  \[5826] ,
  \[9431] ,
  \[9621] ,
  \[10104] ,
  \[9433] ,
  \[9623] ,
  \[1460] ,
  \[10106] ,
  \[11654] ,
  \[9815] ,
  \[10110] ,
  \[311] ,
  \[9247] ,
  \[312] ,
  \[11090] ,
  \[9817] ,
  \[8899] ,
  \[503] ,
  \[1465] ,
  \[9249] ,
  \[9629] ,
  \[314] ,
  \[11282] ,
  \[1466] ,
  \[506] ,
  \[5642] ,
  \[5832] ,
  \[1089] ,
  \[507] ,
  \[508] ,
  \[10118] ,
  \[319] ,
  \[509] ,
  \[5645] ,
  \[5835] ,
  \[11288] ,
  \[5456] ,
  \[5646] ,
  \[9630] ,
  \[5837] ,
  \[5649] ,
  \[9443] ,
  \[9823] ,
  \[10116] ,
  \[9635] ,
  \[320] ,
  \[9825] ,
  \[11286] ,
  \[10120] ,
  \[511] ,
  \[9447] ,
  \[322] ,
  \[11290] ,
  \[10122] ,
  \[9638] ,
  \[1475] ,
  \[12020] ,
  \[9449] ,
  \[514] ,
  \[5840] ,
  \[1477] ,
  \[6000] ,
  \[5082] ,
  \[1478] ,
  \[6001] ,
  \[327] ,
  \[517] ,
  \[707] ,
  \[5653] ,
  \[5843] ,
  \[328] ,
  \[10128] ,
  \[10318] ,
  \[5654] ,
  \[5844] ,
  \[11298] ,
  \[11488] ,
  \[9260] ,
  \[5846] ,
  \[6006] ,
  \[9641] ,
  \[6007] ,
  \[9832] ,
  \[9073] ,
  \[6008] ,
  \[5849] ,
  \[10316] ,
  \[9265] ,
  \[330] ,
  \[9835] ,
  \[10130] ,
  \[10320] ,
  \[1483] ,
  \[9647] ,
  \[1484] ,
  \[11490] ,
  \[10132] ,
  \[9079] ,
  \[9269] ,
  \[3762] ,
  \[9459] ,
  \[5660] ,
  \[5850] ,
  \[335] ,
  \[905] ,
  \[336] ,
  \[6011] ,
  \[3765] ,
  \[1489] ,
  \[6012] ,
  \[5663] ,
  \[5853] ,
  \[338] ,
  \[5664] ,
  \[5854] ,
  \[10708] ,
  \[3388] ,
  \[5855] ,
  \[4308] ,
  \[5667] ,
  \[10134] ,
  \[6017] ,
  \[5858] ,
  \[10704] ,
  \[9273] ,
  \[6018] ,
  \[9463] ,
  \[5859] ,
  \[9653] ,
  \[1490] ,
  \[6019] ,
  \[11874] ,
  \[10516] ,
  \[9844] ,
  \[9275] ,
  \[9465] ,
  \[9655] ,
  \[11496] ,
  \[10140] ,
  \[11876] ,
  \[10710] ,
  \[9847] ,
  \[3391] ,
  \[10142] ,
  \[343] ,
  \[10712] ,
  \[10902] ,
  \[344] ,
  \[11692] ,
  \[5671] ,
  \[5861] ,
  \[346] ,
  \[12802] ,
  \[6021] ,
  \[5672] ,
  \[1499] ,
  \[2228] ,
  \[6022] ,
  \[5864] ,
  \[919] ,
  \[5865] ,
  \[5866] ,
  \[12048] ,
  \[9661] ,
  \[12808] ,
  \[10144] ,
  \[6027] ,
  \[10334] ,
  \[5678] ,
  \[6028] ,
  \[5869] ,
  \[9663] ,
  \[9853] ,
  \[10146] ,
  \[11694] ,
  \[6029] ,
  \[9664] ,
  \[9475] ,
  \[9286] ,
  \[2231] ,
  \[351] ,
  \[352] ,
  \[9857] ,
  \[10152] ,
  \[9288] ,
  \[12805] ,
  \[12050] ,
  \[3592] ,
  \[9479] ,
  \[354] ,
  \[9859] ,
  \[5870] ,
  \[6030] ,
  \[5681] ,
  \[5871] ,
  \[6031] ,
  \[5682] ,
  \[12811] ,
  \[737] ,
  \[10158] ,
  \[5874] ,
  \[359] ,
  \[4706] ,
  \[5875] ,
  \[9670] ,
  \[8502] ,
  \[6036] ,
  \[5687] ,
  \[9481] ,
  \[5877] ,
  \[8313] ,
  \[9861] ,
  \[10154] ,
  \[6037] ,
  \[8314] ,
  \[6038] ,
  \[10156] ,
  \[6039] ,
  \[10536] ,
  \[9674] ,
  \[10726] ,
  \[9864] ,
  \[360] ,
  \[9677] ,
  \[362] ,
  \[9867] ,
  \[10352] ,
  \[173] ,
  \[10922] ,
  \[9299] ,
  \[2814] ,
  \[5690] ,
  \[5880] ,
  \[555] ,
  \[5881] ,
  \[556] ,
  \[177] ,
  \[5882] ,
  \[367] ,
  \[2817] ,
  \[6042] ,
  \[178] ,
  \[368] ,
  \[10168] ,
  \[5694] ,
  \[179] ,
  \[6044] ,
  \[5695] ,
  \[5885] ,
  \[6045] ,
  \[4338] ,
  \[5886] ,
  \[9870] ,
  \[9491] ,
  \[10164] ,
  \[5888] ,
  \[5889] ,
  \[8705] ,
  \[10166] ,
  \[9495] ,
  \[370] ,
  \[10170] ,
  \[8328] ,
  \[9876] ,
  \[561] ,
  \[751] ,
  \[2062] ,
  \[9497] ,
  \[182] ,
  \[562] ,
  \[10172] ,
  \[183] ,
  \[563] ,
  \[184] ,
  \[564] ,
  \[2065] ,
  \[375] ,
  \[6050] ,
  \[376] ,
  \[6051] ,
  \[187] ,
  \[5892] ,
  \[6052] ,
  \[188] ;
assign
  \[5893]  = (~\[5892]  & ~\[8195] ) | ~\[11358] ,
  \[378]  = (~inB0 & ~\[1772] ) | ((~inB0 & ~musel1) | ((~\[9575]  & ~\[1772] ) | (~\[9575]  & ~musel1))),
  \[189]  = (~\[8911]  & ~opsel2) | ((~\[8911]  & ~\[8956] ) | ((~\[5550]  & ~opsel2) | (~\[5550]  & ~\[8956] ))),
  \[5894]  = ~inC10 | ~musel2,
  \[569]  = (~\[10060]  & ~sh1) | ((~\[10060]  & ~\[10056] ) | ((~\[5947]  & ~sh1) | (~\[5947]  & ~\[10056] ))),
  \[8520]  = (~\[6071]  & ~\[346] ) | ~\[10536] ,
  \[8521]  = ~\[8520] ,
  \[6055]  = ~\[5886]  | (~\[5881]  | ~\[12790] ),
  \[9880]  = \[5671]  | \[8817] ,
  \[6056]  = ~opsel2 | ~\[8929] ,
  \[4349]  = (~\[8655]  & ~\[8640] ) | ((~\[8655]  & ~\[5807] ) | ((~\[5825]  & ~\[8640] ) | (~\[5825]  & ~\[5807] ))),
  \[5897]  = ~musel4 | (~\[5523]  | ~\[9417] ),
  \[5898]  = (~\[5897]  & ~\[8195] ) | ~\[11350] ,
  \[10744]  = ~sh2 | ~\[8440] ,
  \[8714]  = ~\[5722] ,
  \[8335]  = (~\[5987]  & ~\[290] ) | ~\[11068] ,
  \[9883]  = ~\[8817]  | ~\[5671] ,
  \[8905]  = (~\[5955]  & ~\[5854] ) | ~\[11242] ,
  \[10556]  = ~opsel3 | (~\[5550]  | ~\[9249] ),
  \[190]  = (~\[9165]  & ~\[9161] ) | ((~\[9165]  & ~\[8956] ) | ((~\[8899]  & ~\[9161] ) | (~\[8899]  & ~\[8956] ))),
  \[8337]  = ~\[8335] ,
  \[570]  = (~\[10062]  & ~sh1) | ((~\[10062]  & ~\[10058] ) | ((~\[5947]  & ~sh1) | (~\[5947]  & ~\[10058] ))),
  \[950]  = (~\[6038]  & ~\[10786] ) | (~\[6038]  & ~\[9740] ),
  \[381]  = ~\[1421]  & (~opsel0 & ~\[5778] ),
  \[9886]  = ~\[6029] ,
  \[8908]  = (~\[5969]  & ~\[5859] ) | ~\[11180] ,
  \[382]  = ~\[1397]  & (~opsel0 & ~\[5796] ),
  \[11100]  = ~\[8781]  | ~\[8328] ,
  \[2642]  = ~\[5708]  & ~\[5528] ,
  \[10372]  = ~inD2 | (~musel4 | (~\[5523]  | ~\[2065] )),
  \[193]  = (~\[1089]  & ~\[9169] ) | (~\[1089]  & ~\[5992] ),
  \[383]  = ~\[1379]  & (~opsel0 & ~\[5814] ),
  \[4540]  = ~\[5782]  & ~\[5528] ,
  \[194]  = (~\[8914]  & ~opsel2) | ((~\[8914]  & ~\[8959] ) | ((~\[5550]  & ~opsel2) | (~\[5550]  & ~\[8959] ))),
  \[384]  = ~\[1361]  & (~opsel0 & ~\[5832] ),
  \[4352]  = (~\[8628]  & ~\[8619] ) | ((~\[8628]  & ~\[5771] ) | ((~\[5789]  & ~\[8619] ) | (~\[5789]  & ~\[5771] ))),
  \[2645]  = ~musel1 & ~musel2,
  \[575]  = (~\[10072]  & ~sh1) | ((~\[10072]  & ~\[10068] ) | ((~\[5947]  & ~sh1) | (~\[5947]  & ~\[10068] ))),
  \[576]  = (~\[10074]  & ~sh1) | ((~\[10074]  & ~\[10070] ) | ((~\[5947]  & ~sh1) | (~\[5947]  & ~\[10070] ))),
  \[6061]  = ~musel3 | ~\[5525] ,
  \[197]  = (~opsel0 & ~opsel1) | ((~opsel0 & ~\[5535] ) | ((~\[5534]  & ~opsel1) | (~\[5534]  & ~\[5535] ))),
  \[6062]  = ~\[5535]  | ~\[5534] ,
  \[198]  = (~\[1045]  & ~\[9182] ) | (~\[1045]  & ~\[6007] ),
  \[6063]  = (~\[8726]  & ~\[8475] ) | (~\[5740]  & ~\[5730] ),
  \[199]  = (~\[8917]  & ~opsel2) | ((~\[8917]  & ~\[8962] ) | ((~\[5550]  & ~opsel2) | (~\[5550]  & ~\[8962] ))),
  \[8530]  = ~\[5771] ,
  \[8911]  = (~\[5937]  & ~\[5865] ) | (~pgx3 & ~\[9101] ),
  \[6065]  = ~\[12790]  | ~\[5886] ,
  \[6066]  = ~opsel2 | ~\[8932] ,
  \[10944]  = ~\[9883]  | ~\[5994] ,
  \[8914]  = (~\[6000]  & ~\[5893] ) | ~\[11040] ,
  \[0]  = (~\[173]  & ~opsel3) | ~\[11290] ,
  \[10946]  = ~opsel3 | (~\[5550]  | ~\[9184] ),
  \[1]  = (~\[178]  & ~opsel3) | ~\[11228] ,
  \[8726]  = ~\[5740] ,
  \[2]  = (~\[183]  & ~opsel3) | ~\[11166] ,
  \[8917]  = (~\[6011]  & ~\[5898] ) | ~\[10960] ,
  \[10570]  = ~\[6065]  | ~\[5881] ,
  \[391]  = (~\[1356]  & ~\[4338] ) | (~\[1356]  & ~\[9605] ),
  \[581]  = (~\[10084]  & ~sh1) | ((~\[10084]  & ~\[10080] ) | ((~\[5947]  & ~sh1) | (~\[5947]  & ~\[10080] ))),
  \[3]  = (~\[188]  & ~opsel3) | (~\[5981]  & ~\[190] ),
  \[8349]  = ~\[5635] ,
  \[582]  = (~\[10086]  & ~sh1) | ((~\[10086]  & ~\[10082] ) | ((~\[5947]  & ~sh1) | (~\[5947]  & ~\[10082] ))),
  \[4]  = (~\[193]  & ~opsel3) | ~\[11026] ,
  \[1105]  = ~\[5947]  & ~\[8287] ,
  \[5]  = (~\[198]  & ~opsel3) | ~\[10946] ,
  \[11302]  = ~\[8195]  | ~\[5932] ,
  \[6]  = (~\[203]  & ~opsel3) | ~\[10870] ,
  \[1107]  = ~\[8270]  & ~sh2,
  \[7]  = (~\[208]  & ~opsel3) | (~\[6030]  & ~\[210] ),
  \[8]  = (~\[213]  & ~opsel3) | ~\[10712] ,
  \[6071]  = ~musel3 | ~\[5525] ,
  \[587]  = (~\[10096]  & ~sh1) | ((~\[10096]  & ~\[10092] ) | ((~\[5947]  & ~sh1) | (~\[5947]  & ~\[10092] ))),
  \[9]  = (~\[218]  & ~opsel3) | ~\[10632] ,
  \[6072]  = ~\[5535]  | ~\[5534] ,
  \[588]  = (~\[10098]  & ~sh1) | ((~\[10098]  & ~\[10094] ) | ((~\[5947]  & ~sh1) | (~\[5947]  & ~\[10094] ))),
  \[6073]  = (~\[5758]  & ~\[5748] ) | (~\[8741]  & ~\[8502] ),
  \[399]  = (~\[12799]  & ~\[9623] ) | (~\[12799]  & ~\[5840] ),
  \[8540]  = (~\[6080]  & ~\[354] ) | ~\[10452] ,
  \[969]  = ~\[6031]  & ~\[6028] ,
  \[8920]  = (~\[6021]  & ~\[5904] ) | ~\[10884] ,
  \[6074]  = ~opsel3 | ~\[5550] ,
  \[11308]  = ~inA0 | (~\[5528]  | ~musel1),
  \[8541]  = ~\[8540] ,
  \[6075]  = ~opsel2 | ~\[8935] ,
  \[8923]  = (~\[5998]  & ~\[5909] ) | (~\[9079]  & ~\[9073] ),
  \[10764]  = ~inD7 | (~musel4 | (~\[5523]  | ~\[2817] )),
  \[8926]  = (~\[6044]  & ~\[5870] ) | ~\[10726] ,
  \[10960]  = ~\[6011]  | ~\[5898] ,
  \[11310]  = ~\[8195]  | ~\[5927] ,
  \[8549]  = ~\[5789] ,
  \[782]  = (~\[6082]  & ~\[10474] ) | (~\[6082]  & ~\[9638] ),
  \[8929]  = (~\[6055]  & ~\[5875] ) | ~\[10646] ,
  \[1115]  = (~\[5993]  & ~\[11090] ) | (~\[5993]  & ~\[9844] ),
  \[593]  = (~\[10108]  & ~sh1) | ((~\[10108]  & ~\[10104] ) | ((~\[5947]  & ~sh1) | (~\[5947]  & ~\[10104] ))),
  \[594]  = (~\[10110]  & ~sh1) | ((~\[10110]  & ~\[10106] ) | ((~\[5947]  & ~sh1) | (~\[5947]  & ~\[10106] ))),
  \[6080]  = ~musel3 | ~\[5525] ,
  \[6081]  = ~\[5535]  | ~\[5534] ,
  \[6082]  = (~\[8619]  & ~\[8530] ) | (~\[5781]  & ~\[5771] ),
  \[10588]  = ~sh2 | ~\[8491] ,
  \[8360]  = (~\[6006]  & ~\[298] ) | ~\[10998] ,
  \[599]  = (~\[10120]  & ~sh1) | ((~\[10120]  & ~\[10116] ) | ((~\[5947]  & ~sh1) | (~\[5947]  & ~\[10116] ))),
  \[8361]  = ~\[8360] ,
  \[11318]  = ~\[8195]  | ~\[5921] ,
  \[8741]  = ~\[5758] ,
  \[8932]  = (~\[6065]  & ~\[5881] ) | ~\[10570] ,
  \[6086]  = ~\[8195]  | (~\[5933]  | (~\[5928]  | ~\[5922] )),
  \[6087]  = ~opsel2 | ~\[8938] ,
  \[8935]  = (~\[6042]  & ~\[5886] ) | (~\[12790]  & ~\[9040] ),
  \[10396]  = ~\[9653]  | ~\[9664] ,
  \[1501]  = ~musel1 & (~musel2 & (~\[5695]  & ~musel3)),
  \[1312]  = (~\[5555]  & ~\[11456] ) | (~\[5555]  & ~\[9932] ),
  \[11316]  = ~inA1 | (~\[5528]  | ~musel1),
  \[1502]  = ~\[5523]  & (~musel4 & ~\[320] ),
  \[11506]  = (~\[1354]  & ~\[1353] ) | ~\[9609] ,
  \[8938]  = (~\[6086]  & ~\[5917] ) | ~\[10414] ,
  \[3404]  = ~\[5946]  & ~\[8185] ,
  \[4954]  = ~\[5687]  & ~\[5528] ,
  \[6092]  = ~musel3 | ~\[5525] ,
  \[5304]  = ~\[5574]  & ~\[5528] ,
  \[6093]  = ~\[5535]  | ~\[5534] ,
  \[10978]  = ~sh2 | ~\[8360] ,
  \[799]  = ~\[6075]  & ~\[6072] ,
  \[6094]  = (~\[8628]  & ~\[8549] ) | (~\[5799]  & ~\[5789] ),
  \[8181]  = (~\[5533]  & ~\[258] ) | ~\[11434] ,
  \[8941]  = (~\[6097]  & ~\[5922] ) | ~\[10334] ,
  \[8372]  = ~\[5653] ,
  \[8562]  = (~\[6092]  & ~\[362] ) | ~\[10372] ,
  \[9101]  = ~\[5865] ,
  \[8563]  = ~\[8562] ,
  \[6097]  = ~\[5933]  | (~\[5928]  | ~\[8195] ),
  \[8754]  = ~\[6039] ,
  \[8944]  = (~\[6107]  & ~\[5928] ) | ~\[10258] ,
  \[6098]  = ~opsel2 | ~\[8941] ,
  \[8185]  = ~\[8181] ,
  \[1130]  = ~\[5843]  & ~\[5840] ,
  \[11324]  = ~inA2 | (~\[5528]  | ~musel1),
  \[10786]  = ~\[9719]  | ~\[9743] ,
  \[1511]  = (~\[5682]  & ~\[8802] ) | (~\[5682]  & ~\[5653] ),
  \[2490]  = ~\[5726]  & ~\[5528] ,
  \[11326]  = ~\[8195]  | ~\[5916] ,
  \[1512]  = ~\[5653]  & ~\[8802] ,
  \[8947]  = (~\[5933]  & ~\[5849] ) | (~\[9012]  & ~\[8195] ),
  \[3600]  = ~sh1 & ~sh2,
  G3 = (~\[8328]  & ~\[9807] ) | ((~\[8328]  & ~\[9815] ) | ((~\[5627]  & ~\[9807] ) | (~\[5627]  & ~\[9815] ))),
  \[2493]  = ~musel1 & ~musel2,
  \[1136]  = ~\[5982]  & ~\[5979] ,
  \[11332]  = ~inA3 | (~\[5528]  | ~musel1),
  \[4392]  = ~\[5818]  & ~\[5528] ,
  \[1517]  = ~\[5550]  & ~\[5549] ,
  \[1329]  = ~\[5550]  & ~\[5549] ,
  \[1519]  = ~musel1 & (~musel2 & (~\[5672]  & ~musel3)),
  \[4965]  = (~\[8817]  & ~\[8802] ) | ((~\[8817]  & ~\[5653] ) | ((~\[5671]  & ~\[8802] ) | (~\[5671]  & ~\[5653] ))),
  \[3228]  = ~\[5631]  & ~\[5528] ,
  \[8570]  = ~\[5807] ,
  \[8950]  = (~\[5950]  & ~\[8270] ) | ~\[11254] ,
  O0 = \[15] ,
  O1 = \[14] ,
  O2 = \[13] ,
  O3 = \[12] ,
  O4 = \[11] ,
  O5 = \[10] ,
  O6 = \[9] ,
  O7 = \[8] ,
  O8 = \[7] ,
  O9 = \[6] ,
  \[11908]  = ~inD10 | (~musel3 | ~\[5528] ),
  \[4968]  = (~\[8790]  & ~\[8781] ) | ((~\[8790]  & ~\[5617] ) | ((~\[5635]  & ~\[8781] ) | (~\[5635]  & ~\[5617] ))),
  \[9301]  = (~\[247]  & ~e1) | (~\[6104]  & ~\[8991] ),
  \[8952]  = ~\[8950] ,
  \[8953]  = (~\[5963]  & ~\[5957] ) | ~\[3592] ,
  \[8195]  = ~\[5849] ,
  \[11334]  = ~\[8195]  | ~\[5908] ,
  \[1520]  = ~\[5523]  & (~musel4 & ~\[312] ),
  \[8955]  = ~\[8953] ,
  \[1331]  = ~musel1 & (~musel2 & (~\[5600]  & ~musel3)),
  \[8956]  = (~\[556]  & ~sh2) | (~\[5946]  & ~\[555] ),
  \[11146]  = ~inD12 | (~musel4 | (~\[5523]  | ~\[3515] )),
  \[1332]  = ~\[5523]  & (~musel4 & ~\[280] ),
  \[8767]  = ~\[5760] ,
  \[8388]  = (~\[6017]  & ~\[306] ) | ~\[10922] ,
  \[9117]  = (~\[5939]  & ~opsel2) | ~\[11298] ,
  \[8389]  = ~\[8388] ,
  \[3231]  = ~musel1 & ~musel2,
  \[11340]  = ~inA8 | (~\[5528]  | ~musel1),
  \[8959]  = (~\[5988]  & ~\[561] ) | ~\[3348] ,
  \[11910]  = ~inB10 | (~\[5523]  | ~musel2),
  \[4780]  = ~\[5723]  & ~\[5528] ,
  \[1525]  = ~\[5529]  & (~musel3 & ~\[311] ),
  \[9119]  = (~\[177]  & ~e15) | (~\[5536]  & ~\[8185] ),
  \[11342]  = ~\[8195]  | ~\[5903] ,
  \[1526]  = (~musel1 & ~\[11842] ) | (~musel1 & ~\[11840] ),
  \[1337]  = ~\[5529]  & (~musel3 & ~\[279] ),
  \[5701]  = (~\[5534]  & ~opsel2) | (~opsel1 & ~opsel3),
  \[1338]  = (~musel1 & ~\[11490] ) | (~musel1 & ~\[11488] ),
  \[5514]  = ~\[5528]  & ~\[5524] ,
  \[5704]  = (~\[423]  & ~b7) | (\[423]  & b7),
  \[10998]  = ~inD10 | (~musel4 | (~\[5523]  | ~\[3231] )),
  \[5705]  = ~inC6,
  \[11348]  = ~inA9 | (~\[5528]  | ~musel1),
  \[11728]  = ~inB5 | (~\[5523]  | ~musel2),
  \[8961]  = ~\[8959] ,
  \[5517]  = ~musel1 & ~musel2,
  \[8962]  = (~\[564]  & ~sh0) | (~\[5948]  & ~\[563] ),
  \[9312]  = ~\[249] ,
  \[5708]  = ~inD6,
  b0 = ~\[1364]  & ~\[1363] ,
  b1 = ~\[1382]  & ~\[1381] ,
  b2 = ~\[1400]  & ~\[1399] ,
  b3 = ~\[1424]  & ~\[1423] ,
  b4 = ~\[1442]  & ~\[1441] ,
  b5 = ~\[1460]  & ~\[1459] ,
  b6 = ~\[1478]  & ~\[1477] ,
  b7 = ~\[1502]  & ~\[1501] ,
  b8 = ~\[1520]  & ~\[1519] ,
  b9 = ~\[1538]  & ~\[1537] ,
  \[8964]  = ~\[8962] ,
  \[9314]  = (~\[252]  & ~e0) | (~\[6114]  & ~\[8994] ),
  \[8965]  = (~\[570]  & ~sh0) | (~\[5948]  & ~\[569] ),
  \[1910]  = ~\[5803]  & ~\[5528] ,
  \[8586]  = (~\[6103]  & ~\[370] ) | ~\[10296] ,
  e0 = (~\[661]  & ~\[6115] ) | (~\[661]  & ~\[5840] ),
  e1 = (~\[697]  & ~\[6105] ) | (~\[697]  & ~\[9670] ),
  e2 = (~\[737]  & ~\[6094] ) | (~\[737]  & ~\[9647] ),
  e3 = (~\[782]  & ~\[9611] ) | (~\[782]  & ~\[6082] ),
  e5 = (~\[865]  & ~\[6063] ) | (~\[865]  & ~\[9772] ),
  \[8587]  = ~\[8586] ,
  e6 = (~\[905]  & ~\[6052] ) | (~\[905]  & ~\[9749] ),
  e7 = (~\[950]  & ~\[9713] ) | (~\[950]  & ~\[6038] ),
  \[8777]  = (~\[6039]  & ~\[9782] ) | (~\[6073]  & ~\[8754] ),
  e9 = (~\[1035]  & ~\[6019] ) | (~\[1035]  & ~\[9876] ),
  \[11726]  = ~inD5 | (~musel3 | ~\[5528] ),
  \[8967]  = ~\[8965] ,
  \[8968]  = (~\[576]  & ~sh0) | (~\[5948]  & ~\[575] ),
  \[1913]  = ~musel1 & ~musel2,
  \[9507]  = (~\[5529]  & ~musel2) | (~\[5528]  & ~musel1),
  \[11350]  = ~\[8195]  | ~\[5897] ,
  \[11920]  = ~inD11 | (~musel3 | ~\[5528] ),
  \[1535]  = ~\[5550]  & ~\[5549] ,
  \[11922]  = ~inB11 | (~\[5523]  | ~musel2),
  \[5900]  = ~inC9 | ~musel2,
  \[1347]  = ~\[5843]  & ~\[5840] ,
  \[1537]  = ~musel1 & (~musel2 & (~\[5654]  & ~musel3)),
  \[1538]  = ~\[5523]  & (~musel4 & ~\[304] ),
  \[5712]  = (~\[1484]  & ~\[1483] ) | ~\[5525] ,
  \[1349]  = ~\[5549]  & (~opsel2 & ~opsel1),
  \[3626]  = ~\[5577]  & ~\[5528] ,
  \[5523]  = ~musel3,
  \[5713]  = ~inC6 | ~musel4,
  \[5903]  = ~musel4 | (~\[5523]  | ~\[9433] ),
  \[5524]  = ~inD15,
  \[5904]  = (~\[5903]  & ~\[8195] ) | ~\[11342] ,
  \[5525]  = ~musel4,
  \[5905]  = ~inC8 | ~musel2,
  \[11358]  = ~\[8195]  | ~\[5892] ,
  \[9130]  = ~\[179] ,
  \[8781]  = ~\[5627] ,
  \[3629]  = ~musel1 & ~musel2,
  \[8971]  = (~\[582]  & ~sh0) | (~\[5948]  & ~\[581] ),
  \[9511]  = (~\[5529]  & ~musel2) | (~\[5528]  & ~musel1),
  \[8593]  = ~\[5825] ,
  \[9132]  = (~\[182]  & ~e14) | (~\[5951]  & ~\[8952] ),
  \[5528]  = ~musel2,
  \[8973]  = ~\[8971] ,
  \[5908]  = ~musel4 | (~\[5523]  | ~\[9449] ),
  \[5529]  = ~musel1,
  \[8974]  = (~\[588]  & ~sh0) | (~\[5948]  & ~\[587] ),
  \[5719]  = (~\[5534]  & ~opsel2) | (~opsel1 & ~opsel3),
  \[9513]  = (~\[5882]  & ~musel1) | ~\[11372] ,
  \[5909]  = (~\[5908]  & ~\[8195] ) | ~\[11334] ,
  \[1350]  = ~\[5550]  & (~opsel3 & ~\[5534] ),
  \[11544]  = ~inD0 | (~musel3 | ~\[5528] ),
  \[8976]  = ~\[8974] ,
  \[11166]  = ~opsel3 | (~\[5550]  | ~\[9145] ),
  \[11356]  = ~inA10 | (~\[5528]  | ~musel1),
  \[11546]  = ~inB0 | (~\[5523]  | ~musel2),
  \[8977]  = (~\[594]  & ~sh0) | (~\[5948]  & ~\[593] ),
  \[1353]  = (~\[391]  & ~\[8628] ) | (~\[391]  & ~\[5789] ),
  \[1543]  = ~\[5529]  & (~musel3 & ~\[303] ),
  \[202]  = (~opsel0 & ~opsel1) | ((~opsel0 & ~\[5535] ) | ((~\[5534]  & ~opsel1) | (~\[5534]  & ~\[5535] ))),
  \[9707]  = ~\[8726]  | ~\[5730] ,
  \[1354]  = ~\[5789]  & ~\[8628] ,
  \[1544]  = (~musel1 & ~\[11876] ) | (~musel1 & ~\[11874] ),
  \[8979]  = ~\[8977] ,
  \[203]  = (~\[1005]  & ~\[9195] ) | (~\[1005]  & ~\[6018] ),
  \[204]  = (~\[8920]  & ~opsel2) | ((~\[8920]  & ~\[8965] ) | ((~\[5550]  & ~opsel2) | (~\[5550]  & ~\[8965] ))),
  \[1356]  = ~\[5807]  & ~\[8640] ,
  \[1167]  = ~\[5970]  & ~\[5966] ,
  \[5911]  = ~\[5909]  | (~\[5904]  | (~\[5898]  | ~\[5893] )),
  \[5722]  = (~\[424]  & ~b6) | (\[424]  & b6),
  \[207]  = (~opsel0 & ~opsel1) | ((~opsel0 & ~\[5535] ) | ((~\[5534]  & ~opsel1) | (~\[5534]  & ~\[5535] ))),
  \[5533]  = ~musel3 | ~\[5525] ,
  \[5723]  = ~inC5,
  \[208]  = (~\[969]  & ~\[9208] ) | (~\[969]  & ~\[6028] ),
  \[5913]  = ~inC3 | ~musel2,
  \[5534]  = ~opsel1,
  \[209]  = (~\[8923]  & ~opsel2) | ((~\[8923]  & ~\[8968] ) | ((~\[5550]  & ~opsel2) | (~\[5550]  & ~\[8968] ))),
  \[8790]  = ~\[5645] ,
  \[5535]  = ~opsel0,
  \[8980]  = (~\[600]  & ~sh0) | (~\[5948]  & ~\[599] ),
  \[5156]  = ~\[5628]  & ~\[5528] ,
  \[5536]  = ~\[5535]  | ~\[5534] ,
  \[5726]  = ~inD5,
  \[5916]  = ~musel4 | (~\[5523]  | ~\[9529] ),
  \[5537]  = ~inC15,
  \[9331]  = (~\[5529]  & ~musel2) | (~\[5528]  & ~musel1),
  \[5917]  = (~\[5916]  & ~\[8195] ) | ~\[11326] ,
  \[9711]  = ~\[8705]  | ~\[5694] ,
  \[9901]  = (~\[5763]  & ~\[511] ) | ~\[8767] ,
  b10 = ~\[1556]  & ~\[1555] ,
  b11 = ~\[1580]  & ~\[1579] ,
  b12 = ~\[1332]  & ~\[1331] ,
  \[8983]  = (~\[606]  & ~sh0) | (~\[5948]  & ~\[605] ),
  b13 = ~\[1592]  & ~\[1591] ,
  b14 = ~\[1616]  & ~\[1615] ,
  b15 = ~\[1630]  & ~\[1629] ,
  \[5918]  = ~inC2 | ~musel2,
  \[9143]  = ~\[184] ,
  \[9523]  = (~\[5529]  & ~musel2) | (~\[5528]  & ~musel1),
  \[9713]  = (~\[438]  & ~\[9741] ) | ~\[9743] ,
  \[11364]  = ~inA11 | (~\[5528]  | ~musel1),
  \[8985]  = ~\[8983] ,
  \[1361]  = ~\[5550]  & ~\[5549] ,
  \[9145]  = (~\[187]  & ~e13) | (~\[5966]  & ~\[8955] ),
  \[9335]  = (~\[5529]  & ~musel2) | (~\[5528]  & ~musel1),
  \[8986]  = (~\[612]  & ~sh0) | (~\[5948]  & ~\[611] ),
  \[210]  = (~\[9217]  & ~\[9213] ) | ((~\[9217]  & ~\[8968] ) | ((~\[8849]  & ~\[9213] ) | (~\[8849]  & ~\[8968] ))),
  \[9905]  = (~\[514]  & ~\[9933] ) | ~\[9935] ,
  \[11366]  = ~\[8195]  | ~\[5885] ,
  \[1363]  = ~musel1 & (~musel2 & (~\[5826]  & ~musel3)),
  \[1553]  = ~\[5550]  & ~\[5549] ,
  \[9337]  = (~\[5846]  & ~musel1) | ~\[11424] ,
  \[8988]  = ~\[8986] ,
  \[9527]  = (~\[5529]  & ~musel2) | (~\[5528]  & ~musel1),
  \[11180]  = ~\[5969]  | ~\[5859] ,
  \[1364]  = ~\[5523]  & (~musel4 & ~\[376] ),
  \[8989]  = (~\[618]  & ~sh0) | (~\[5948]  & ~\[617] ),
  \[213]  = (~\[919]  & ~\[9221] ) | (~\[919]  & ~\[6037] ),
  \[1555]  = ~musel1 & (~musel2 & (~\[5636]  & ~musel3)),
  \[9529]  = (~\[5913]  & ~musel1) | ~\[11332] ,
  \[214]  = (~\[8926]  & ~opsel2) | ((~\[8926]  & ~\[8971] ) | ((~\[5550]  & ~opsel2) | (~\[5550]  & ~\[8971] ))),
  \[9719]  = (~\[441]  & ~\[12805] ) | ~\[9731] ,
  \[11372]  = ~inA4 | (~\[5528]  | ~musel1),
  \[1556]  = ~\[5523]  & (~musel4 & ~\[296] ),
  \[5730]  = (~\[1466]  & ~\[1465] ) | ~\[5525] ,
  \[5731]  = ~inC5 | ~musel4,
  \[5921]  = ~musel4 | (~\[5523]  | ~\[9545] ),
  \[5542]  = (~\[1636]  & ~\[1635] ) | ~\[5525] ,
  \[217]  = (~opsel0 & ~opsel1) | ((~opsel0 & ~\[5535] ) | ((~\[5534]  & ~opsel1) | (~\[5534]  & ~\[5535] ))),
  \[5922]  = (~\[5921]  & ~\[8195] ) | ~\[11318] ,
  \[3076]  = ~\[5649]  & ~\[5528] ,
  \[1369]  = ~\[5529]  & (~musel3 & ~\[375] ),
  \[5543]  = ~inC15 | ~musel4,
  \[218]  = (~\[875]  & ~\[9234] ) | (~\[875]  & ~\[6051] ),
  \[219]  = (~\[8929]  & ~opsel2) | ((~\[8929]  & ~\[8974] ) | ((~\[5550]  & ~opsel2) | (~\[5550]  & ~\[8974] ))),
  \[5924]  = ~inC1 | ~musel2,
  \[3079]  = ~musel1 & ~musel2,
  \[8991]  = ~\[8989] ,
  \[8992]  = (~\[624]  & ~sh0) | (~\[5948]  & ~\[623] ),
  \[5737]  = (~\[5534]  & ~opsel2) | (~opsel1 & ~opsel3),
  \[5927]  = ~musel4 | (~\[5523]  | ~\[9561] ),
  \[9721]  = (~\[6039]  & ~\[12808] ) | ~\[9728] ,
  \[9911]  = (~\[517]  & ~\[12793] ) | ~\[9923] ,
  \[10204]  = ~sh2 | ~\[8611] ,
  \[5928]  = (~\[5927]  & ~\[8195] ) | ~\[11310] ,
  \[10013]  = (~\[5946]  & ~sh1) | ~\[11196] ,
  \[5549]  = ~opsel3,
  \[8994]  = ~\[8992] ,
  \[5929]  = ~inC0 | ~musel2,
  \[9913]  = (~\[5844]  & ~\[12796] ) | ~\[9920] ,
  \[1370]  = (~musel1 & ~\[11546] ) | (~musel1 & ~\[11544] ),
  \[11374]  = ~\[8195]  | ~\[5880] ,
  \[10015]  = (~\[5948]  & ~\[8270] ) | (~\[8287]  & ~sh0),
  \[1561]  = ~\[5529]  & (~musel3 & ~\[295] ),
  \[600]  = (~\[10122]  & ~sh1) | ((~\[10122]  & ~\[10118] ) | ((~\[5947]  & ~sh1) | (~\[5947]  & ~\[10118] ))),
  \[1562]  = (~musel1 & ~\[11910] ) | (~musel1 & ~\[11908] ),
  \[9156]  = ~\[189] ,
  \[10400]  = ~opsel3 | (~\[5550]  | ~\[9275] ),
  \[411]  = (~\[12802]  & ~\[9655] ) | (~\[12802]  & ~\[5840] ),
  \[3270]  = ~\[5935]  & ~\[5911] ,
  \[9347]  = (~\[5529]  & ~musel2) | (~\[5528]  & ~musel1),
  \[222]  = (~opsel0 & ~opsel1) | ((~opsel0 & ~\[5535] ) | ((~\[5534]  & ~opsel1) | (~\[5534]  & ~\[5535] ))),
  \[11380]  = ~inA5 | (~\[5528]  | ~musel1),
  \[11760]  = ~inD6 | (~musel3 | ~\[5528] ),
  \[223]  = (~\[835]  & ~\[9247] ) | (~\[835]  & ~\[6062] ),
  \[9728]  = ~\[8741]  | ~\[5748] ,
  \[9539]  = (~\[5529]  & ~musel2) | (~\[5528]  & ~musel1),
  \[224]  = (~\[8932]  & ~opsel2) | ((~\[8932]  & ~\[8977] ) | ((~\[5550]  & ~opsel2) | (~\[5550]  & ~\[8977] ))),
  \[11382]  = ~\[8195]  | ~\[5874] ,
  \[5550]  = ~opsel2,
  \[11762]  = ~inB6 | (~\[5523]  | ~musel2),
  \[5740]  = (~\[425]  & ~b5) | (\[425]  & b5),
  \[605]  = (~\[10132]  & ~sh1) | ((~\[10132]  & ~\[10128] ) | ((~\[5947]  & ~sh1) | (~\[5947]  & ~\[10128] ))),
  \[1567]  = ~\[5529]  & (~musel3 & ~\[287] ),
  \[5551]  = (~\[5534]  & ~opsel2) | (~opsel1 & ~opsel3),
  \[5741]  = ~inC4,
  \[606]  = (~\[10134]  & ~sh1) | ((~\[10134]  & ~\[10130] ) | ((~\[5947]  & ~sh1) | (~\[5947]  & ~\[10130] ))),
  \[1568]  = (~musel1 & ~\[11922] ) | (~musel1 & ~\[11920] ),
  \[227]  = (~opsel0 & ~opsel1) | ((~opsel0 & ~\[5535] ) | ((~\[5534]  & ~opsel1) | (~\[5534]  & ~\[5535] ))),
  \[5932]  = ~musel4 | (~\[5523]  | ~\[9577] ),
  \[1379]  = ~\[5550]  & ~\[5549] ,
  \[228]  = (~\[799]  & ~\[9260] ) | (~\[799]  & ~\[6072] ),
  \[5933]  = (~\[5932]  & ~\[8195] ) | ~\[11302] ,
  \[5554]  = (~\[506]  & ~b15) | (\[506]  & b15),
  \[5744]  = ~inD4,
  \[229]  = (~\[8935]  & ~opsel2) | ((~\[8935]  & ~\[8980] ) | ((~\[5550]  & ~opsel2) | (~\[5550]  & ~\[8980] ))),
  \[5555]  = (~\[5554]  & ~\[5542] ) | ~\[12020] ,
  \[5935]  = ~\[5933]  | (~\[5928]  | (~\[5922]  | ~\[5917] )),
  \[11388]  = ~inA6 | (~\[5528]  | ~musel1),
  \[11578]  = ~inD1 | (~musel3 | ~\[5528] ),
  \[5556]  = ~inC14,
  \[9920]  = ~\[8870]  | ~\[5599] ,
  \[10029]  = (~\[5947]  & ~\[8270] ) | (~\[8314]  & ~sh1),
  \[9161]  = ~\[5979] ,
  \[9351]  = (~\[5529]  & ~musel2) | (~\[5528]  & ~musel1),
  \[5937]  = ~pgx3,
  \[9731]  = \[5730]  | \[8726] ,
  \[5748]  = (~\[1448]  & ~\[1447] ) | ~\[5525] ,
  \[5559]  = ~inD14,
  \[9353]  = (~\[5850]  & ~musel1) | ~\[11420] ,
  \[5749]  = ~inC4 | ~musel4,
  \[9543]  = (~\[5529]  & ~musel2) | (~\[5528]  & ~musel1),
  \[5939]  = ~pgx3 | (~\[5865]  | (~\[5859]  | ~\[5854] )),
  \[1190]  = (~\[5967]  & ~\[11226] ) | (~\[5967]  & ~\[9968] ),
  \[9923]  = \[5581]  | \[8861] ,
  \[1381]  = ~musel1 & (~musel2 & (~\[5808]  & ~musel3)),
  \[10025]  = ~\[5976] ,
  \[9165]  = (~\[5535]  & ~opsel1) | (~\[5534]  & ~opsel0),
  \[9545]  = (~\[5918]  & ~musel1) | ~\[11324] ,
  \[230]  = (~\[9269]  & ~\[9265] ) | ((~\[9269]  & ~\[8980] ) | ((~\[8777]  & ~\[9265] ) | (~\[8777]  & ~\[8980] ))),
  \[11196]  = ~sh1 | ~\[5957] ,
  \[1382]  = ~\[5523]  & (~musel4 & ~\[368] ),
  \[611]  = (~\[10144]  & ~sh1) | ((~\[10144]  & ~\[10140] ) | ((~\[5947]  & ~sh1) | (~\[5947]  & ~\[10140] ))),
  \[612]  = (~\[10146]  & ~sh1) | ((~\[10146]  & ~\[10142] ) | ((~\[5947]  & ~sh1) | (~\[5947]  & ~\[10142] ))),
  \[11390]  = ~\[8195]  | ~\[5869] ,
  \[11580]  = ~inB1 | (~\[5523]  | ~musel2),
  \[233]  = (~\[751]  & ~\[9273] ) | (~\[751]  & ~\[6081] ),
  \[423]  = ~\[1499]  & (~opsel0 & ~\[5701] ),
  \[10031]  = (~\[562]  & ~sh0) | (~\[5990]  & ~\[8314] ),
  \[9169]  = ~\[194] ,
  \[234]  = (~\[8938]  & ~opsel2) | ((~\[8938]  & ~\[8983] ) | ((~\[5550]  & ~opsel2) | (~\[5550]  & ~\[8983] ))),
  \[424]  = ~\[1475]  & (~opsel0 & ~\[5719] ),
  \[11772]  = ~inD7 | (~musel3 | ~\[5528] ),
  \[425]  = ~\[1457]  & (~opsel0 & ~\[5737] ),
  \[1387]  = ~\[5529]  & (~musel3 & ~\[367] ),
  \[1577]  = ~\[5550]  & ~\[5549] ,
  \[426]  = ~\[1439]  & (~opsel0 & ~\[5755] ),
  \[1388]  = (~musel1 & ~\[11580] ) | (~musel1 & ~\[11578] ),
  \[237]  = (~opsel0 & ~opsel1) | ((~opsel0 & ~\[5535] ) | ((~\[5534]  & ~opsel1) | (~\[5534]  & ~\[5535] ))),
  \[617]  = (~\[10156]  & ~sh1) | ((~\[10156]  & ~\[10152] ) | ((~\[5947]  & ~sh1) | (~\[5947]  & ~\[10152] ))),
  \[1579]  = ~musel1 & (~musel2 & (~\[5618]  & ~musel3)),
  \[5563]  = (~\[1604]  & ~\[1603] ) | ~\[5525] ,
  \[238]  = (~\[707]  & ~\[9286] ) | (~\[707]  & ~\[6093] ),
  \[618]  = (~\[10158]  & ~sh1) | ((~\[10158]  & ~\[10154] ) | ((~\[5947]  & ~sh1) | (~\[5947]  & ~\[10154] ))),
  \[5564]  = ~inC14 | ~musel4,
  \[6103]  = ~musel3 | ~\[5525] ,
  \[239]  = (~\[8941]  & ~opsel2) | ((~\[8941]  & ~\[8986] ) | ((~\[5550]  & ~opsel2) | (~\[5550]  & ~\[8986] ))),
  \[10608]  = ~inD5 | (~musel4 | (~\[5523]  | ~\[2493] )),
  \[6104]  = ~\[5535]  | ~\[5534] ,
  \[5755]  = (~\[5534]  & ~opsel2) | (~opsel1 & ~opsel3),
  \[5945]  = ~musel3 | ~\[5525] ,
  \[11398]  = ~\[8195]  | ~\[5864] ,
  \[6105]  = (~\[8640]  & ~\[8570] ) | (~\[5817]  & ~\[5807] ),
  \[5946]  = ~sh2,
  \[9740]  = \[5712]  | \[8714] ,
  \[9171]  = (~\[197]  & ~e11) | (~\[5992]  & ~\[8961] ),
  \[5947]  = ~sh1,
  \[9741]  = ~\[9740] ,
  \[5378]  = ~\[5556]  & ~\[5528] ,
  e10 = (~\[1075]  & ~\[6008] ) | (~\[1075]  & ~\[9853] ),
  \[10224]  = ~inD0 | (~musel4 | (~\[5523]  | ~\[1775] )),
  e11 = (~\[1115]  & ~\[9817] ) | (~\[1115]  & ~\[5993] ),
  e13 = (~\[1190]  & ~\[5967] ) | (~\[1190]  & ~\[9964] ),
  \[6107]  = ~\[8195]  | ~\[5933] ,
  \[10414]  = ~\[6086]  | ~\[5917] ,
  e14 = (~\[1221]  & ~\[5952] ) | (~\[1221]  & ~\[9941] ),
  \[5758]  = (~\[426]  & ~b4) | (\[426]  & b4),
  e15 = (~\[1312]  & ~\[9905] ) | (~\[1312]  & ~\[5555] ),
  \[5948]  = ~sh0,
  \[9932]  = \[5563]  | \[8855] ,
  \[9363]  = (~\[5529]  & ~musel2) | (~\[5528]  & ~musel1),
  \[6108]  = ~opsel2 | ~\[8944] ,
  \[9743]  = ~\[8714]  | ~\[5712] ,
  \[9933]  = ~\[9932] ,
  \[1580]  = ~\[5523]  & (~musel4 & ~\[288] ),
  \[11774]  = ~inB7 | (~\[5523]  | ~musel2),
  \[9555]  = (~\[5529]  & ~musel2) | (~\[5528]  & ~musel1),
  \[9935]  = ~\[8855]  | ~\[5563] ,
  \[11396]  = ~inA7 | (~\[5528]  | ~musel1),
  \[1772]  = ~\[5821]  & ~\[5528] ,
  \[9367]  = (~\[5529]  & ~musel2) | (~\[5528]  & ~musel1),
  \[242]  = (~opsel0 & ~opsel1) | ((~opsel0 & ~\[5535] ) | ((~\[5534]  & ~opsel1) | (~\[5534]  & ~\[5535] ))),
  \[432]  = (~\[1434]  & ~\[4308] ) | (~\[1434]  & ~\[9707] ),
  \[243]  = (~\[667]  & ~\[9299] ) | (~\[667]  & ~\[6104] ),
  \[623]  = (~\[10168]  & ~sh1) | ((~\[10168]  & ~\[10164] ) | ((~\[5947]  & ~sh1) | (~\[5947]  & ~\[10164] ))),
  \[1775]  = ~musel1 & ~musel2,
  \[9369]  = (~\[5855]  & ~musel1) | ~\[11412] ,
  \[9559]  = (~\[5529]  & ~musel2) | (~\[5528]  & ~musel1),
  \[244]  = (~\[8944]  & ~opsel2) | ((~\[8944]  & ~\[8989] ) | ((~\[5550]  & ~opsel2) | (~\[5550]  & ~\[8989] ))),
  \[9749]  = ~\[10704]  | ~\[9766] ,
  \[624]  = (~\[10170]  & ~sh1) | ((~\[10170]  & ~\[10166] ) | ((~\[5947]  & ~sh1) | (~\[5947]  & ~\[10166] ))),
  \[5570]  = (~\[5534]  & ~opsel2) | (~opsel1 & ~opsel3),
  \[5760]  = (~\[5694]  & ~\[8705] ) | ~\[11654] ,
  \[5950]  = (~\[5947]  & ~sh2) | ~\[3736] ,
  \[1397]  = ~\[5550]  & ~\[5549] ,
  \[5951]  = ~\[5535]  | ~\[5534] ,
  \[247]  = (~opsel0 & ~opsel1) | ((~opsel0 & ~\[5535] ) | ((~\[5534]  & ~opsel1) | (~\[5534]  & ~\[5535] ))),
  \[5952]  = (~\[8855]  & ~\[8254] ) | (~\[5573]  & ~\[5563] ),
  \[1399]  = ~musel1 & (~musel2 & (~\[5790]  & ~musel3)),
  \[1589]  = ~\[5550]  & ~\[5549] ,
  \[5573]  = (~\[507]  & ~b14) | (\[507]  & b14),
  \[5763]  = ~\[4663]  | ~\[4666] ,
  \[248]  = (~\[631]  & ~\[9312] ) | (~\[631]  & ~\[6114] ),
  \[438]  = (~\[12805]  & ~\[9721] ) | (~\[12805]  & ~\[9731] ),
  \[10048]  = (~\[5946]  & ~\[8185] ) | (~\[8337]  & ~sh2),
  \[5574]  = ~inC13,
  \[6113]  = ~musel3 | ~\[5525] ,
  \[5764]  = ~inC3,
  \[249]  = (~\[8947]  & ~opsel2) | ((~\[8947]  & ~\[8992] ) | ((~\[5550]  & ~opsel2) | (~\[5550]  & ~\[8992] ))),
  \[6114]  = ~\[5535]  | ~\[5534] ,
  \[5955]  = ~\[5865]  | (~\[5859]  | ~pgx3),
  \[6115]  = (~\[5835]  & ~\[5825] ) | (~\[8655]  & ~\[8593] ),
  \[11978]  = ~inB13 | (~\[5523]  | ~musel2),
  \[5956]  = ~opsel2 | ~\[8905] ,
  \[5577]  = ~inD13,
  \[5767]  = ~inD3,
  \[9561]  = (~\[5924]  & ~musel1) | ~\[11316] ,
  \[5957]  = ~sh0 | ~sh2,
  \[9941]  = ~\[11282]  | ~\[9958] ,
  \[10044]  = (~\[8287]  & ~sh2) | ~\[10978] ,
  \[9182]  = ~\[199] ,
  \[6117]  = ~opsel2 | ~\[8947] ,
  \[9753]  = (~\[6039]  & ~\[9759] ) | ~\[9760] ,
  \[10046]  = (~\[5946]  & ~\[8185] ) | (~\[8314]  & ~sh2),
  \[9184]  = (~\[202]  & ~e10) | (~\[6007]  & ~\[8964] ),
  pgx3 = ~\[5935]  & (~\[5849]  & (~\[5911]  & ~\[5888] )),
  \[1591]  = ~musel1 & (~musel2 & (~\[5582]  & ~musel3)),
  \[9755]  = ~\[10710]  | ~\[9757] ,
  \[9945]  = (~\[5844]  & ~\[9951] ) | ~\[9952] ,
  \[10050]  = (~\[5946]  & ~\[8270] ) | (~\[8361]  & ~sh2),
  \[1592]  = ~\[5523]  & (~musel4 & ~\[272] ),
  \[11976]  = ~inD13 | (~musel3 | ~\[5528] ),
  \[441]  = (~\[12808]  & ~\[9728] ) | (~\[12808]  & ~\[6039] ),
  \[631]  = ~\[6117]  & ~\[6114] ,
  \[252]  = (~opsel0 & ~opsel1) | ((~opsel0 & ~\[5535] ) | ((~\[5534]  & ~opsel1) | (~\[5534]  & ~\[5535] ))),
  \[9757]  = \[5748]  | \[8741] ,
  \[9947]  = ~\[11288]  | ~\[9949] ,
  \[10432]  = ~sh2 | ~\[8540] ,
  \[9379]  = (~\[5529]  & ~musel2) | (~\[5528]  & ~musel1),
  \[9759]  = ~\[9757] ,
  \[9949]  = \[5599]  | \[8870] ,
  \[4222]  = ~\[5592]  & ~\[5528] ,
  \[255]  = (~inA15 & ~inC15) | ((~inA15 & ~musel2) | ((~\[5528]  & ~inC15) | (~\[5528]  & ~musel2))),
  \[1597]  = ~\[5529]  & (~musel3 & ~\[271] ),
  \[5581]  = (~\[1598]  & ~\[1597] ) | ~\[5525] ,
  \[5771]  = (~\[1412]  & ~\[1411] ) | ~\[5525] ,
  \[256]  = (~inA15 & ~\[5456] ) | ((~inA15 & ~musel1) | ((~\[9331]  & ~\[5456] ) | (~\[9331]  & ~musel1))),
  \[1598]  = (~musel1 & ~\[11978] ) | (~musel1 & ~\[11976] ),
  \[5582]  = ~inC13 | ~musel4,
  \[5772]  = ~inC3 | ~musel4,
  \[5962]  = ~musel3 | ~\[5525] ,
  \[258]  = (~inB15 & ~\[5514] ) | ((~inB15 & ~musel1) | ((~\[9335]  & ~\[5514] ) | (~\[9335]  & ~musel1))),
  \[5963]  = ~sh1 | ~\[8286] ,
  \[10058]  = (~\[5946]  & ~\[8185] ) | (~\[8337]  & ~sh2),
  \[11988]  = ~inD14 | (~musel3 | ~\[5528] ),
  \[5966]  = ~\[5535]  | ~\[5534] ,
  \[9760]  = ~\[8741]  | ~\[5748] ,
  \[9571]  = (~\[5529]  & ~musel2) | (~\[5528]  & ~musel1),
  \[5967]  = (~\[8861]  & ~\[8274] ) | (~\[5591]  & ~\[5581] ),
  \[9951]  = ~\[9949] ,
  \[10244]  = ~opsel3 | (~\[5550]  | ~\[9301] ),
  \[5588]  = (~\[5534]  & ~opsel2) | (~opsel1 & ~opsel3),
  \[5778]  = (~\[5534]  & ~opsel2) | (~opsel1 & ~opsel3),
  \[9952]  = ~\[8870]  | ~\[5599] ,
  \[9383]  = (~\[5529]  & ~musel2) | (~\[5528]  & ~musel1),
  \[5969]  = ~pgx3 | ~\[5865] ,
  \[9763]  = \[5730]  | \[8726] ,
  \[8405]  = ~\[5671] ,
  \[10056]  = (~\[8314]  & ~sh2) | ~\[10902] ,
  \[9195]  = ~\[204] ,
  \[9385]  = (~\[5861]  & ~musel1) | ~\[11404] ,
  \[9575]  = (~\[5529]  & ~musel2) | (~\[5528]  & ~musel1),
  \[9955]  = \[5581]  | \[8861] ,
  \[10060]  = (~\[5946]  & ~\[8270] ) | (~\[8361]  & ~sh2),
  \[10630]  = ~\[9779]  | ~\[6039] ,
  \[9766]  = ~\[8726]  | ~\[5730] ,
  \[9197]  = (~\[207]  & ~e9) | (~\[6018]  & ~\[8967] ),
  \[9577]  = (~\[5929]  & ~musel1) | ~\[11308] ,
  \[10062]  = (~\[5946]  & ~\[8287] ) | (~\[8389]  & ~sh2),
  \[11990]  = ~inB14 | (~\[5523]  | ~musel2),
  \[263]  = (~inA14 & ~inC14) | ((~inA14 & ~musel2) | ((~\[5528]  & ~inC14) | (~\[5528]  & ~musel2))),
  \[10632]  = ~opsel3 | (~\[5550]  | ~\[9236] ),
  \[9958]  = ~\[8861]  | ~\[5581] ,
  \[264]  = (~inA14 & ~\[5378] ) | ((~inA14 & ~musel1) | ((~\[9347]  & ~\[5378] ) | (~\[9347]  & ~musel1))),
  \[5970]  = ~opsel2 | ~\[8908] ,
  \[835]  = ~\[6066]  & ~\[6062] ,
  \[5591]  = (~\[508]  & ~b13) | (\[508]  & b13),
  \[5781]  = (~\[381]  & ~b3) | (\[381]  & b3),
  \[266]  = (~inB14 & ~\[3762] ) | ((~inB14 & ~musel1) | ((~\[9351]  & ~\[3762] ) | (~\[9351]  & ~musel1))),
  \[5592]  = ~inC12,
  \[5782]  = ~inC2,
  \[10068]  = (~\[8337]  & ~sh2) | ~\[10830] ,
  \[10258]  = ~\[6107]  | ~\[5928] ,
  \[5595]  = ~inD12,
  \[5785]  = ~inD2,
  \[5975]  = ~musel3 | ~\[5525] ,
  \[5976]  = ~sh0 | ~sh1,
  \[5977]  = ~sh0 | ~\[5947] ,
  \[5978]  = (~\[5976]  & ~\[8185] ) | (~\[5977]  & ~\[8287] ),
  \[9772]  = (~\[6039]  & ~\[9778] ) | ~\[9779] ,
  \[5599]  = (~\[1338]  & ~\[1337] ) | ~\[5525] ,
  \[5789]  = (~\[1406]  & ~\[1405] ) | ~\[5525] ,
  \[5979]  = ~\[5535]  | ~\[5534] ,
  \[9964]  = (~\[5844]  & ~\[9970] ) | ~\[9971] ,
  \[9395]  = (~\[5529]  & ~musel2) | (~\[5528]  & ~musel1),
  \[10070]  = (~\[5946]  & ~\[8185] ) | (~\[8361]  & ~sh2),
  \[271]  = (~inA13 & ~inC13) | ((~inA13 & ~musel2) | ((~\[5528]  & ~inC13) | (~\[5528]  & ~musel2))),
  \[9776]  = \[5748]  | \[8741] ,
  \[8418]  = (~\[6027]  & ~\[314] ) | ~\[10850] ,
  \[10830]  = ~sh2 | ~\[8418] ,
  \[272]  = (~inA13 & ~\[5304] ) | ((~inA13 & ~musel1) | ((~\[9363]  & ~\[5304] ) | (~\[9363]  & ~musel1))),
  \[8419]  = ~\[8418] ,
  \[10072]  = (~\[5946]  & ~\[8287] ) | (~\[8389]  & ~sh2),
  \[10452]  = ~inD3 | (~musel4 | (~\[5523]  | ~\[2231] )),
  \[9778]  = ~\[9776] ,
  \[9968]  = \[5599]  | \[8870] ,
  \[9399]  = (~\[5529]  & ~musel2) | (~\[5528]  & ~musel1),
  \[274]  = (~inB13 & ~\[3626] ) | ((~inB13 & ~musel1) | ((~\[9367]  & ~\[3626] ) | (~\[9367]  & ~musel1))),
  \[9779]  = ~\[8741]  | ~\[5748] ,
  \[464]  = ~\[1577]  & (~opsel0 & ~\[5624] ),
  \[5790]  = ~inC2 | ~musel4,
  \[5980]  = (~\[5609]  & ~\[5599] ) | (~\[8870]  & ~\[8298] ),
  \[465]  = ~\[1553]  & (~opsel0 & ~\[5642] ),
  \[5981]  = ~opsel3 | ~\[5550] ,
  \[466]  = ~\[1535]  & (~opsel0 & ~\[5660] ),
  \[5982]  = ~opsel2 | ~\[8911] ,
  \[467]  = ~\[1517]  & (~opsel0 & ~\[5678] ),
  \[468]  = ~\[5837]  & ~\[1130] ,
  \[279]  = (~inA12 & ~inC12) | ((~inA12 & ~musel2) | ((~\[5528]  & ~inC12) | (~\[5528]  & ~musel2))),
  \[8611]  = (~\[6113]  & ~\[378] ) | ~\[10224] ,
  \[5796]  = (~\[5534]  & ~opsel2) | (~opsel1 & ~opsel3),
  \[9970]  = ~\[9968] ,
  \[8612]  = ~\[8611] ,
  \[8802]  = ~\[5663] ,
  \[5987]  = ~musel3 | ~\[5525] ,
  \[9971]  = ~\[8870]  | ~\[5599] ,
  \[10074]  = (~\[5946]  & ~\[8314] ) | (~\[8419]  & ~sh2),
  \[5988]  = ~sh0 | ~sh1,
  \[9782]  = ~\[6073] ,
  \[5799]  = (~\[382]  & ~b2) | (\[382]  & b2),
  \[10646]  = ~\[6055]  | ~\[5875] ,
  \[9974]  = ~\[5980] ,
  \[280]  = (~inA12 & ~\[4222] ) | ((~inA12 & ~musel1) | ((~\[9379]  & ~\[4222] ) | (~\[9379]  & ~musel1))),
  \[10080]  = (~\[8361]  & ~sh2) | ~\[10744] ,
  \[661]  = ~\[6115]  & ~\[5840] ,
  \[2352]  = ~\[5744]  & ~\[5528] ,
  \[282]  = (~inB12 & ~\[3512] ) | ((~inB12 & ~musel1) | ((~\[9383]  & ~\[3512] ) | (~\[9383]  & ~musel1))),
  \[8619]  = ~\[5781] ,
  \[10082]  = (~\[5946]  & ~\[8185] ) | (~\[8389]  & ~sh2),
  \[2355]  = ~musel1 & ~musel2,
  \[5990]  = ~sh0 | ~\[5947] ,
  \[287]  = (~inA11 & ~inC11) | ((~inA11 & ~musel2) | ((~\[5528]  & ~inC11) | (~\[5528]  & ~musel2))),
  \[5992]  = ~\[5535]  | ~\[5534] ,
  \[667]  = ~\[6108]  & ~\[6104] ,
  \[288]  = (~inA11 & ~\[5256] ) | ((~inA11 & ~musel1) | ((~\[9395]  & ~\[5256] ) | (~\[9395]  & ~musel1))),
  \[5993]  = (~\[8781]  & ~\[8328] ) | ~\[11100] ,
  \[10468]  = ~\[9615]  | ~\[9638] ,
  \[5994]  = (~\[5763]  & ~\[468] ) | ~\[8767] ,
  \[8430]  = ~\[5694] ,
  \[10084]  = (~\[5946]  & ~\[8314] ) | (~\[8419]  & ~sh2),
  \[5998]  = ~\[3270]  | ~\[8195] ,
  \[10086]  = (~\[5946]  & ~\[8337] ) | (~\[8441]  & ~sh2),
  \[10276]  = ~sh2 | ~\[8586] ,
  \[290]  = (~inB11 & ~\[3388] ) | ((~inB11 & ~musel1) | ((~\[9399]  & ~\[3388] ) | (~\[9399]  & ~musel1))),
  \[480]  = (~\[12811]  & ~\[9825] ) | (~\[12811]  & ~\[9835] ),
  \[8817]  = ~\[5681] ,
  \[10850]  = ~inD8 | (~musel4 | (~\[5523]  | ~\[2941] )),
  \[8628]  = ~\[5799] ,
  \[10092]  = (~\[8389]  & ~sh2) | ~\[10664] ,
  \[1005]  = ~\[6022]  & ~\[6018] ,
  \[483]  = (~\[484]  & ~\[9832] ) | (~\[484]  & ~\[5994] ),
  \[4640]  = ~\[5764]  & ~\[5528] ,
  \[484]  = ~\[5671]  & ~\[8817] ,
  \[295]  = (~inA10 & ~inC10) | ((~inA10 & ~musel2) | ((~\[5528]  & ~inC10) | (~\[5528]  & ~musel2))),
  \[865]  = (~\[6063]  & ~\[10630] ) | (~\[6063]  & ~\[9776] ),
  \[296]  = (~inA10 & ~\[5156] ) | ((~inA10 & ~musel1) | ((~\[9411]  & ~\[5156] ) | (~\[9411]  & ~musel1))),
  \[298]  = (~inB10 & ~\[3228] ) | ((~inB10 & ~musel1) | ((~\[9415]  & ~\[3228] ) | (~\[9415]  & ~musel1))),
  \[2938]  = ~\[5667]  & ~\[5528] ,
  \[10098]  = (~\[5946]  & ~\[8361] ) | (~\[8465]  & ~sh2),
  \[489]  = ~\[5635]  & ~\[8790] ,
  \[8440]  = (~\[6036]  & ~\[322] ) | ~\[10764] ,
  \[11018]  = ~\[9857]  | ~\[9867] ,
  \[8441]  = ~\[8440] ,
  \[10094]  = (~\[5946]  & ~\[8270] ) | (~\[8419]  & ~sh2),
  \[10474]  = ~\[9617]  | ~\[9641] ,
  \[8254]  = ~\[5563] ,
  \[10664]  = ~sh2 | ~\[8464] ,
  \[11014]  = ~\[8790]  | ~\[8349] ,
  \[1200]  = ~\[5956]  & ~\[5951] ,
  \[11204]  = ~inD13 | (~musel4 | (~\[5523]  | ~\[3629] )),
  \[10096]  = (~\[5946]  & ~\[8337] ) | (~\[8441]  & ~sh2),
  \[10476]  = ~\[9621]  | ~\[9635] ,
  \[2941]  = ~musel1 & ~musel2,
  \[11022]  = ~\[9859]  | ~\[9870] ,
  \[875]  = ~\[6056]  & ~\[6051] ,
  \[496]  = ~\[5671]  & ~\[8817] ,
  \[4466]  = ~\[5800]  & ~\[5528] ,
  \[10868]  = ~\[8817]  | ~\[8405] ,
  \[8640]  = ~\[5817] ,
  \[8830]  = ~\[5994] ,
  \[8451]  = ~\[5712] ,
  \[8263]  = (~\[5945]  & ~\[266] ) | ~\[11262] ,
  \[5008]  = ~\[5664]  & ~\[5528] ,
  \[11024]  = ~\[9864]  | ~\[5994] ,
  \[1400]  = ~\[5523]  & (~musel4 & ~\[360] ),
  \[11404]  = ~inA12 | (~\[5528]  | ~musel1),
  \[10296]  = ~inD1 | (~musel4 | (~\[5523]  | ~\[1913] )),
  \[11026]  = ~opsel3 | (~\[5550]  | ~\[9171] ),
  \[11406]  = ~\[8195]  | ~\[5858] ,
  \[10870]  = ~opsel3 | (~\[5550]  | ~\[9197] ),
  \[1405]  = ~\[5529]  & (~musel3 & ~\[359] ),
  \[1406]  = (~musel1 & ~\[11614] ) | (~musel1 & ~\[11612] ),
  \[11412]  = ~inA13 | (~\[5528]  | ~musel1),
  \[4663]  = (~\[8741]  & ~\[8726] ) | ((~\[8741]  & ~\[5730] ) | ((~\[5748]  & ~\[8726] ) | (~\[5748]  & ~\[5730] ))),
  \[697]  = (~\[6105]  & ~\[10318] ) | (~\[6105]  & ~\[9674] ),
  \[4854]  = ~\[5705]  & ~\[5528] ,
  \[8270]  = ~\[8263] ,
  \[4666]  = (~\[8714]  & ~\[8705] ) | ((~\[8714]  & ~\[5694] ) | ((~\[5712]  & ~\[8705] ) | (~\[5712]  & ~\[5694] ))),
  \[8271]  = ~\[5853] ,
  \[11228]  = ~opsel3 | (~\[5550]  | ~\[9132] ),
  \[8274]  = ~\[5581] ,
  \[10684]  = ~inD6 | (~musel4 | (~\[5523]  | ~\[2645] )),
  \[8464]  = (~\[6050]  & ~\[330] ) | ~\[10684] ,
  \[8465]  = ~\[8464] ,
  \[8655]  = ~\[5835] ,
  \[1221]  = (~\[5952]  & ~\[11286] ) | (~\[5952]  & ~\[9955] ),
  \[1411]  = ~\[5529]  & (~musel3 & ~\[351] ),
  \[11226]  = ~\[9971]  | ~\[5844] ,
  \[1412]  = (~musel1 & ~\[11626] ) | (~musel1 & ~\[11624] ),
  \[1603]  = ~\[5529]  & (~musel3 & ~\[263] ),
  \[11040]  = ~\[6000]  | ~\[5893] ,
  \[11420]  = ~inA14 | (~\[5528]  | ~musel1),
  \[1604]  = (~musel1 & ~\[11990] ) | (~musel1 & ~\[11988] ),
  \[8849]  = (~\[5994]  & ~\[9886] ) | (~\[6029]  & ~\[8830] ),
  \[1035]  = (~\[6019]  & ~\[10944] ) | (~\[6019]  & ~\[9880] ),
  \[11612]  = ~inD2 | (~musel3 | ~\[5528] ),
  \[9012]  = ~\[5933] ,
  O10 = \[5] ,
  O11 = \[4] ,
  O12 = \[3] ,
  O13 = \[2] ,
  O14 = \[1] ,
  O15 = \[0] ,
  \[10884]  = ~\[6021]  | ~\[5904] ,
  \[8475]  = ~\[5730] ,
  \[11424]  = ~inA15 | (~\[5528]  | ~musel1),
  \[11614]  = ~inB2 | (~\[5523]  | ~musel2),
  \[8855]  = ~\[5573] ,
  \[8286]  = (~\[5962]  & ~\[274] ) | ~\[11204] ,
  \[1421]  = ~\[5550]  & ~\[5549] ,
  \[8287]  = ~\[8286] ,
  \[11806]  = (~\[1512]  & ~\[1511] ) | (~\[5645]  & ~\[8349] ),
  \[1423]  = ~musel1 & (~musel2 & (~\[5772]  & ~musel3)),
  \[1613]  = ~\[5550]  & ~\[5549] ,
  \[1424]  = ~\[5523]  & (~musel4 & ~\[352] ),
  \[9208]  = ~\[209] ,
  \[1045]  = ~\[6012]  & ~\[6007] ,
  \[1235]  = ~\[5939]  & (~\[5550]  & ~\[5536] ),
  \[1615]  = ~musel1 & (~musel2 & (~\[5564]  & ~musel3)),
  \[3512]  = ~\[5595]  & ~\[5528] ,
  \[11242]  = ~\[5955]  | ~\[5854] ,
  \[12790]  = ~\[5935]  & ~\[5849] ,
  \[1616]  = ~\[5523]  & (~musel4 & ~\[264] ),
  \[5600]  = ~inC12 | ~musel4,
  \[3515]  = ~musel1 & ~musel2,
  \[10]  = (~\[223]  & ~opsel3) | ~\[10556] ,
  \[11]  = (~\[228]  & ~opsel3) | (~\[6074]  & ~\[230] ),
  \[12]  = (~\[233]  & ~opsel3) | ~\[10400] ,
  \[13]  = (~\[238]  & ~opsel3) | ~\[10320] ,
  \[8861]  = ~\[5591] ,
  \[5606]  = (~\[5534]  & ~opsel2) | (~opsel1 & ~opsel3),
  \[14]  = (~\[243]  & ~opsel3) | ~\[10244] ,
  \[9401]  = (~\[5889]  & ~musel1) | ~\[11364] ,
  \[15]  = (~\[248]  & ~opsel3) | ~\[10172] ,
  \[8673]  = ~\[5840] ,
  \[9213]  = ~\[6028] ,
  \[5609]  = (~\[509]  & ~b12) | (\[509]  & b12),
  \[11434]  = ~musel4 | (~inD15 | (~\[5523]  | ~\[5517] )),
  \[11624]  = ~inD3 | (~musel3 | ~\[5528] ),
  \[12799]  = ~\[5835]  & ~\[8593] ,
  \[1431]  = (~\[432]  & ~\[8714] ) | (~\[432]  & ~\[5712] ),
  \[1432]  = ~\[5712]  & ~\[8714] ,
  \[11626]  = ~inB3 | (~\[5523]  | ~musel2),
  \[8298]  = ~\[5599] ,
  \[12793]  = ~\[5591]  & ~\[8274] ,
  \[9217]  = (~\[5535]  & ~opsel1) | (~\[5534]  & ~opsel0),
  \[12796]  = \[8298]  & \[5609] ,
  \[1434]  = ~\[5730]  & ~\[8726] ,
  \[5610]  = ~inC11,
  \[5800]  = ~inC1,
  \[1627]  = ~\[5550]  & ~\[5549] ,
  \[1439]  = ~\[5550]  & ~\[5549] ,
  \[1629]  = ~musel1 & (~musel2 & (~\[5543]  & ~musel3)),
  \[5613]  = ~inD11,
  \[5803]  = ~inD1,
  \[8870]  = ~\[5609] ,
  \[11068]  = ~inD11 | (~musel4 | (~\[5523]  | ~\[3391] )),
  \[8491]  = (~\[6061]  & ~\[338] ) | ~\[10608] ,
  \[8492]  = ~\[8491] ,
  \[9221]  = ~\[214] ,
  \[5617]  = (~\[1568]  & ~\[1567] ) | ~\[5525] ,
  \[9411]  = (~\[5529]  & ~musel2) | (~\[5528]  & ~musel1),
  \[5807]  = (~\[1388]  & ~\[1387] ) | ~\[5525] ,
  \[5618]  = ~inC11 | ~musel4,
  \[5808]  = ~inC1 | ~musel4,
  \[9223]  = (~\[217]  & ~e7) | (~\[6037]  & ~\[8973] ),
  \[11254]  = ~\[5950]  | ~\[8181] ,
  \[1630]  = ~\[5523]  & (~musel4 & ~\[256] ),
  \[1441]  = ~musel1 & (~musel2 & (~\[5749]  & ~musel3)),
  \[9415]  = (~\[5529]  & ~musel2) | (~\[5528]  & ~musel1),
  \[9605]  = ~\[8640]  | ~\[5807] ,
  \[1442]  = ~\[5523]  & (~musel4 & ~\[344] ),
  \[9417]  = (~\[5894]  & ~musel1) | ~\[11356] ,
  \[1635]  = ~\[5529]  & (~musel3 & ~\[255] ),
  \[9609]  = ~\[8619]  | ~\[5771] ,
  \[11262]  = ~inD14 | (~musel4 | (~\[5523]  | ~\[3765] )),
  \[1636]  = (~musel1 & ~\[12050] ) | (~musel1 & ~\[12048] ),
  \[1447]  = ~\[5529]  & (~musel3 & ~\[343] ),
  \[1448]  = (~musel1 & ~\[11694] ) | (~musel1 & ~\[11692] ),
  \[5624]  = (~\[5534]  & ~opsel2) | (~opsel1 & ~opsel3),
  \[5814]  = (~\[5534]  & ~opsel2) | (~opsel1 & ~opsel3),
  \[3348]  = (~\[10031]  & ~\[3404] ) | ((~\[10031]  & ~\[5988] ) | ((~\[5946]  & ~\[3404] ) | (~\[5946]  & ~\[5988] ))),
  \[9040]  = ~\[5886] ,
  \[5627]  = (~\[464]  & ~b11) | (\[464]  & b11),
  \[5817]  = (~\[383]  & ~b1) | (\[383]  & b1),
  \[9611]  = ~\[10468]  | ~\[9641] ,
  \[8693]  = ~\[5837] ,
  \[5628]  = ~inC10,
  \[5818]  = ~inC0,
  \[8884]  = ~\[5844] ,
  \[9234]  = ~\[219] ,
  \[9615]  = (~\[399]  & ~\[9630] ) | ~\[9635] ,
  \[11456]  = ~\[9911]  | ~\[9935] ,
  \[9236]  = (~\[222]  & ~e6) | (~\[6051]  & ~\[8976] ),
  \[9427]  = (~\[5529]  & ~musel2) | (~\[5528]  & ~musel1),
  \[9617]  = ~\[10476]  | ~\[9629] ,
  \[9807]  = (~\[5635]  & ~\[8790] ) | ~\[11806] ,
  \[11840]  = ~inD8 | (~musel3 | ~\[5528] ),
  \[303]  = (~inA9 & ~inC9) | ((~inA9 & ~musel2) | ((~\[5528]  & ~inC9) | (~\[5528]  & ~musel2))),
  \[1075]  = (~\[6008]  & ~\[11022] ) | (~\[6008]  & ~\[9867] ),
  \[304]  = (~inA9 & ~\[5082] ) | ((~inA9 & ~musel1) | ((~\[9427]  & ~\[5082] ) | (~\[9427]  & ~musel1))),
  \[11842]  = ~inB8 | (~\[5523]  | ~musel2),
  \[1457]  = ~\[5550]  & ~\[5549] ,
  \[5631]  = ~inD10,
  \[5821]  = ~inD0,
  \[306]  = (~inB9 & ~\[3076] ) | ((~inB9 & ~musel1) | ((~\[9431]  & ~\[3076] ) | (~\[9431]  & ~musel1))),
  \[1459]  = ~musel1 & (~musel2 & (~\[5731]  & ~musel3)),
  \[3736]  = (~sh0 & ~sh2) | ((~sh0 & ~\[5948] ) | ((~\[5947]  & ~sh2) | (~\[5947]  & ~\[5948] ))),
  \[10108]  = (~\[5946]  & ~\[8361] ) | (~\[8465]  & ~sh2),
  \[5635]  = (~\[1562]  & ~\[1561] ) | ~\[5525] ,
  \[5825]  = (~\[1370]  & ~\[1369] ) | ~\[5525] ,
  \[5256]  = ~\[5610]  & ~\[5528] ,
  \[5636]  = ~inC10 | ~musel4,
  \[5826]  = ~inC0 | ~musel4,
  \[9431]  = (~\[5529]  & ~musel2) | (~\[5528]  & ~musel1),
  \[9621]  = (~\[5840]  & ~\[12799] ) | ~\[9623] ,
  \[10104]  = (~\[8419]  & ~sh2) | ~\[10588] ,
  \[9433]  = (~\[5900]  & ~musel1) | ~\[11348] ,
  \[9623]  = \[5825]  | \[8655] ,
  \[1460]  = ~\[5523]  & (~musel4 & ~\[336] ),
  \[10106]  = (~\[5946]  & ~\[8287] ) | (~\[8441]  & ~sh2),
  \[11654]  = (~\[1432]  & ~\[1431] ) | ~\[9711] ,
  \[9815]  = ~\[8781]  | ~\[5617] ,
  \[10110]  = (~\[5946]  & ~\[8389] ) | (~\[8492]  & ~sh2),
  \[311]  = (~inA8 & ~inC8) | ((~inA8 & ~musel2) | ((~\[5528]  & ~inC8) | (~\[5528]  & ~musel2))),
  \[9247]  = ~\[224] ,
  \[312]  = (~inA8 & ~\[5008] ) | ((~inA8 & ~musel1) | ((~\[9443]  & ~\[5008] ) | (~\[9443]  & ~musel1))),
  \[11090]  = ~\[9823]  | ~\[9847] ,
  \[9817]  = (~\[480]  & ~\[489] ) | ~\[9847] ,
  \[8899]  = (~\[5844]  & ~\[9974] ) | (~\[5980]  & ~\[8884] ),
  \[503]  = ~\[5671]  & ~\[8817] ,
  \[1465]  = ~\[5529]  & (~musel3 & ~\[335] ),
  \[9249]  = (~\[227]  & ~e5) | (~\[6062]  & ~\[8979] ),
  \[9629]  = \[5807]  | \[8640] ,
  \[314]  = (~inB8 & ~\[2938] ) | ((~inB8 & ~musel1) | ((~\[9447]  & ~\[2938] ) | (~\[9447]  & ~musel1))),
  \[11282]  = ~\[9945]  | ~\[9955] ,
  \[1466]  = (~musel1 & ~\[11728] ) | (~musel1 & ~\[11726] ),
  \[506]  = ~\[1627]  & (~opsel0 & ~\[5551] ),
  \[5642]  = (~\[5534]  & ~opsel2) | (~opsel1 & ~opsel3),
  \[5832]  = (~\[5534]  & ~opsel2) | (~opsel1 & ~opsel3),
  \[1089]  = ~\[6001]  & ~\[5992] ,
  \[507]  = ~\[1613]  & (~opsel0 & ~\[5570] ),
  \[508]  = ~\[1589]  & (~opsel0 & ~\[5588] ),
  \[10118]  = (~\[5946]  & ~\[8314] ) | (~\[8465]  & ~sh2),
  \[319]  = (~inA7 & ~inC7) | ((~inA7 & ~musel2) | ((~\[5528]  & ~inC7) | (~\[5528]  & ~musel2))),
  \[509]  = ~\[1329]  & (~opsel0 & ~\[5606] ),
  \[5645]  = (~\[465]  & ~b10) | (\[465]  & b10),
  \[5835]  = (~\[384]  & ~b0) | (\[384]  & b0),
  \[11288]  = ~\[9952]  | ~\[5844] ,
  \[5456]  = ~\[5537]  & ~\[5528] ,
  \[5646]  = ~inC9,
  \[9630]  = ~\[9629] ,
  \[5837]  = (~\[5771]  & ~\[8619] ) | ~\[11506] ,
  \[5649]  = ~inD9,
  \[9443]  = (~\[5529]  & ~musel2) | (~\[5528]  & ~musel1),
  \[9823]  = (~\[483]  & ~\[12811] ) | ~\[9835] ,
  \[10116]  = (~\[8441]  & ~sh2) | ~\[10516] ,
  \[9635]  = ~\[8640]  | ~\[5807] ,
  \[320]  = (~inA7 & ~\[4954] ) | ((~inA7 & ~musel1) | ((~\[9459]  & ~\[4954] ) | (~\[9459]  & ~musel1))),
  \[9825]  = (~\[5994]  & ~\[484] ) | ~\[9832] ,
  \[11286]  = ~\[9947]  | ~\[9958] ,
  \[10120]  = (~\[5946]  & ~\[8389] ) | (~\[8492]  & ~sh2),
  \[511]  = ~\[5837]  & ~\[1347] ,
  \[9447]  = (~\[5529]  & ~musel2) | (~\[5528]  & ~musel1),
  \[322]  = (~inB7 & ~\[2814] ) | ((~inB7 & ~musel1) | ((~\[9463]  & ~\[2814] ) | (~\[9463]  & ~musel1))),
  \[11290]  = ~opsel3 | (~\[5550]  | ~\[9119] ),
  \[10122]  = (~\[5946]  & ~\[8419] ) | (~\[8521]  & ~sh2),
  \[9638]  = \[5789]  | \[8628] ,
  \[1475]  = ~\[5550]  & ~\[5549] ,
  \[12020]  = ~\[5554]  | ~\[5542] ,
  \[9449]  = (~\[5905]  & ~musel1) | ~\[11340] ,
  \[514]  = (~\[12793]  & ~\[9913] ) | (~\[12793]  & ~\[9923] ),
  \[5840]  = (~\[1350]  & ~\[1349] ) | ~\[5535] ,
  \[1477]  = ~musel1 & (~musel2 & (~\[5713]  & ~musel3)),
  \[6000]  = ~\[9079]  | (~\[5909]  | (~\[5904]  | ~\[5898] )),
  \[5082]  = ~\[5646]  & ~\[5528] ,
  \[1478]  = ~\[5523]  & (~musel4 & ~\[328] ),
  \[6001]  = ~opsel2 | ~\[8914] ,
  \[327]  = (~inA6 & ~inC6) | ((~inA6 & ~musel2) | ((~\[5528]  & ~inC6) | (~\[5528]  & ~musel2))),
  \[517]  = (~\[12796]  & ~\[9920] ) | (~\[12796]  & ~\[5844] ),
  \[707]  = ~\[6098]  & ~\[6093] ,
  \[5653]  = (~\[1544]  & ~\[1543] ) | ~\[5525] ,
  \[5843]  = ~\[4349]  | ~\[4352] ,
  \[328]  = (~inA6 & ~\[4854] ) | ((~inA6 & ~musel1) | ((~\[9475]  & ~\[4854] ) | (~\[9475]  & ~musel1))),
  \[10128]  = (~\[8465]  & ~sh2) | ~\[10432] ,
  \[10318]  = ~\[8673]  | ~\[9677] ,
  \[5654]  = ~inC9 | ~musel4,
  \[5844]  = ~G3 | ~\[11496] ,
  \[11298]  = ~opsel2 | ~\[8181] ,
  \[11488]  = ~inD12 | (~musel3 | ~\[5528] ),
  \[9260]  = ~\[229] ,
  \[5846]  = ~inC15 | ~musel2,
  \[6006]  = ~musel3 | ~\[5525] ,
  \[9641]  = ~\[8628]  | ~\[5789] ,
  \[6007]  = ~\[5535]  | ~\[5534] ,
  \[9832]  = ~\[8817]  | ~\[5671] ,
  \[9073]  = ~\[5909] ,
  \[6008]  = (~\[8790]  & ~\[8349] ) | ~\[11014] ,
  \[5849]  = ~musel4 | (~\[5523]  | ~\[9337] ),
  \[10316]  = ~\[9674]  | ~\[5840] ,
  \[9265]  = ~\[6072] ,
  \[330]  = (~inB6 & ~\[2642] ) | ((~inB6 & ~musel1) | ((~\[9479]  & ~\[2642] ) | (~\[9479]  & ~musel1))),
  \[9835]  = \[5653]  | \[8802] ,
  \[10130]  = (~\[5946]  & ~\[8337] ) | (~\[8492]  & ~sh2),
  \[10320]  = ~opsel3 | (~\[5550]  | ~\[9288] ),
  \[1483]  = ~\[5529]  & (~musel3 & ~\[327] ),
  \[9647]  = (~\[411]  & ~\[9663] ) | ~\[9664] ,
  \[1484]  = (~musel1 & ~\[11762] ) | (~musel1 & ~\[11760] ),
  \[11490]  = ~inB12 | (~\[5523]  | ~musel2),
  \[10132]  = (~\[5946]  & ~\[8419] ) | (~\[8521]  & ~sh2),
  \[9079]  = ~\[5998] ,
  \[9269]  = (~\[5535]  & ~opsel1) | (~\[5534]  & ~opsel0),
  \[3762]  = ~\[5559]  & ~\[5528] ,
  \[9459]  = (~\[5529]  & ~musel2) | (~\[5528]  & ~musel1),
  \[5660]  = (~\[5534]  & ~opsel2) | (~opsel1 & ~opsel3),
  \[5850]  = ~inC14 | ~musel2,
  \[335]  = (~inA5 & ~inC5) | ((~inA5 & ~musel2) | ((~\[5528]  & ~inC5) | (~\[5528]  & ~musel2))),
  \[905]  = (~\[6052]  & ~\[10708] ) | (~\[6052]  & ~\[9763] ),
  \[336]  = (~inA5 & ~\[4780] ) | ((~inA5 & ~musel1) | ((~\[9491]  & ~\[4780] ) | (~\[9491]  & ~musel1))),
  \[6011]  = ~\[5909]  | (~\[5904]  | ~\[9079] ),
  \[3765]  = ~musel1 & ~musel2,
  \[1489]  = ~\[5529]  & (~musel3 & ~\[319] ),
  \[6012]  = ~opsel2 | ~\[8917] ,
  \[5663]  = (~\[466]  & ~b9) | (\[466]  & b9),
  \[5853]  = ~musel4 | (~\[5523]  | ~\[9353] ),
  \[338]  = (~inB5 & ~\[2490] ) | ((~inB5 & ~musel1) | ((~\[9495]  & ~\[2490] ) | (~\[9495]  & ~musel1))),
  \[5664]  = ~inC8,
  \[5854]  = (~\[5853]  & ~\[8195] ) | (~\[5849]  & ~\[8271] ),
  \[10708]  = ~\[9755]  | ~\[9766] ,
  \[3388]  = ~\[5613]  & ~\[5528] ,
  \[5855]  = ~inC13 | ~musel2,
  \[4308]  = ~\[5748]  & ~\[8741] ,
  \[5667]  = ~inD8,
  \[10134]  = (~\[5946]  & ~\[8441] ) | (~\[8541]  & ~sh2),
  \[6017]  = ~musel3 | ~\[5525] ,
  \[5858]  = ~musel4 | (~\[5523]  | ~\[9369] ),
  \[10704]  = ~\[9753]  | ~\[9763] ,
  \[9273]  = ~\[234] ,
  \[6018]  = ~\[5535]  | ~\[5534] ,
  \[9463]  = (~\[5529]  & ~musel2) | (~\[5528]  & ~musel1),
  \[5859]  = (~\[5858]  & ~\[8195] ) | ~\[11406] ,
  \[9653]  = (~\[5840]  & ~\[12802] ) | ~\[9655] ,
  \[1490]  = (~musel1 & ~\[11774] ) | (~musel1 & ~\[11772] ),
  \[6019]  = (~\[8802]  & ~\[8372] ) | (~\[5663]  & ~\[5653] ),
  \[11874]  = ~inD9 | (~musel3 | ~\[5528] ),
  \[10516]  = ~sh2 | ~\[8520] ,
  \[9844]  = \[5635]  | \[8790] ,
  \[9275]  = (~\[237]  & ~e3) | (~\[6081]  & ~\[8985] ),
  \[9465]  = (~\[5866]  & ~musel1) | ~\[11396] ,
  \[9655]  = \[5825]  | \[8655] ,
  \[11496]  = ~\[4965]  | (~\[4968]  | ~\[9901] ),
  \[10140]  = (~\[8492]  & ~sh2) | ~\[10352] ,
  \[11876]  = ~inB9 | (~\[5523]  | ~musel2),
  \[10710]  = ~\[9760]  | ~\[6039] ,
  \[9847]  = \[5645]  | \[8349] ,
  \[3391]  = ~musel1 & ~musel2,
  \[10142]  = (~\[5946]  & ~\[8361] ) | (~\[8521]  & ~sh2),
  \[343]  = (~inA4 & ~inC4) | ((~inA4 & ~musel2) | ((~\[5528]  & ~inC4) | (~\[5528]  & ~musel2))),
  \[10712]  = ~opsel3 | (~\[5550]  | ~\[9223] ),
  \[10902]  = ~sh2 | ~\[8388] ,
  \[344]  = (~inA4 & ~\[4706] ) | ((~inA4 & ~musel1) | ((~\[9507]  & ~\[4706] ) | (~\[9507]  & ~musel1))),
  \[11692]  = ~inD4 | (~musel3 | ~\[5528] ),
  \[5671]  = (~\[1526]  & ~\[1525] ) | ~\[5525] ,
  \[5861]  = ~inC12 | ~musel2,
  \[346]  = (~inB4 & ~\[2352] ) | ((~inB4 & ~musel1) | ((~\[9511]  & ~\[2352] ) | (~\[9511]  & ~musel1))),
  \[12802]  = ~\[5835]  & ~\[8593] ,
  \[6021]  = ~\[9079]  | ~\[5909] ,
  \[5672]  = ~inC8 | ~musel4,
  \[1499]  = ~\[5550]  & ~\[5549] ,
  \[2228]  = ~\[5767]  & ~\[5528] ,
  \[6022]  = ~opsel2 | ~\[8920] ,
  \[5864]  = ~musel4 | (~\[5523]  | ~\[9385] ),
  \[919]  = ~\[6045]  & ~\[6037] ,
  \[5865]  = (~\[5864]  & ~\[8195] ) | ~\[11398] ,
  \[5866]  = ~inC7 | ~musel2,
  \[12048]  = ~inD15 | (~musel3 | ~\[5528] ),
  \[9661]  = \[5807]  | \[8640] ,
  \[12808]  = \[8502]  & \[5758] ,
  \[10144]  = (~\[5946]  & ~\[8441] ) | (~\[8541]  & ~sh2),
  \[6027]  = ~musel3 | ~\[5525] ,
  \[10334]  = ~\[6097]  | ~\[5922] ,
  \[5678]  = (~\[5534]  & ~opsel2) | (~opsel1 & ~opsel3),
  \[6028]  = ~\[5535]  | ~\[5534] ,
  \[5869]  = ~musel4 | (~\[5523]  | ~\[9465] ),
  \[9663]  = ~\[9661] ,
  \[9853]  = ~\[11018]  | ~\[9870] ,
  \[10146]  = (~\[5946]  & ~\[8465] ) | (~\[8563]  & ~sh2),
  \[11694]  = ~inB4 | (~\[5523]  | ~musel2),
  \[6029]  = (~\[8817]  & ~\[8405] ) | ~\[10868] ,
  \[9664]  = ~\[8640]  | ~\[5807] ,
  \[9475]  = (~\[5529]  & ~musel2) | (~\[5528]  & ~musel1),
  \[9286]  = ~\[239] ,
  \[2231]  = ~musel1 & ~musel2,
  \[351]  = (~inA3 & ~inC3) | ((~inA3 & ~musel2) | ((~\[5528]  & ~inC3) | (~\[5528]  & ~musel2))),
  \[352]  = (~inA3 & ~\[4640] ) | ((~inA3 & ~musel1) | ((~\[9523]  & ~\[4640] ) | (~\[9523]  & ~musel1))),
  \[9857]  = (~\[5994]  & ~\[496] ) | ~\[9864] ,
  \[10152]  = (~\[8521]  & ~sh2) | ~\[10276] ,
  \[9288]  = (~\[242]  & ~e2) | (~\[6093]  & ~\[8988] ),
  \[12805]  = ~\[5740]  & ~\[8475] ,
  \[12050]  = ~inB15 | (~\[5523]  | ~musel2),
  \[3592]  = (~\[3600]  & ~\[10013] ) | ((~\[3600]  & ~\[8181] ) | ((~\[10015]  & ~\[10013] ) | (~\[10015]  & ~\[8181] ))),
  \[9479]  = (~\[5529]  & ~musel2) | (~\[5528]  & ~musel1),
  \[354]  = (~inB3 & ~\[2228] ) | ((~inB3 & ~musel1) | ((~\[9527]  & ~\[2228] ) | (~\[9527]  & ~musel1))),
  \[9859]  = ~\[11024]  | ~\[9861] ,
  \[5870]  = (~\[5869]  & ~\[8195] ) | ~\[11390] ,
  \[6030]  = ~opsel3 | ~\[5550] ,
  \[5681]  = (~\[467]  & ~b8) | (\[467]  & b8),
  \[5871]  = ~inC6 | ~musel2,
  \[6031]  = ~opsel2 | ~\[8923] ,
  \[5682]  = ~\[8405]  | ~\[5681] ,
  \[12811]  = ~\[5663]  & ~\[8372] ,
  \[737]  = (~\[6094]  & ~\[10396] ) | (~\[6094]  & ~\[9661] ),
  \[10158]  = (~\[5946]  & ~\[8492] ) | (~\[8587]  & ~sh2),
  \[5874]  = ~musel4 | (~\[5523]  | ~\[9481] ),
  \[359]  = (~inA2 & ~inC2) | ((~inA2 & ~musel2) | ((~\[5528]  & ~inC2) | (~\[5528]  & ~musel2))),
  \[4706]  = ~\[5741]  & ~\[5528] ,
  \[5875]  = (~\[5874]  & ~\[8195] ) | ~\[11382] ,
  \[9670]  = ~\[10316]  | ~\[9677] ,
  \[8502]  = ~\[5748] ,
  \[6036]  = ~musel3 | ~\[5525] ,
  \[5687]  = ~inC7,
  \[9481]  = (~\[5871]  & ~musel1) | ~\[11388] ,
  \[5877]  = ~inC5 | ~musel2,
  \[8313]  = (~\[5975]  & ~\[282] ) | ~\[11146] ,
  \[9861]  = \[5671]  | \[8817] ,
  \[10154]  = (~\[5946]  & ~\[8389] ) | (~\[8541]  & ~sh2),
  \[6037]  = ~\[5535]  | ~\[5534] ,
  \[8314]  = ~\[8313] ,
  \[6038]  = (~\[8705]  & ~\[8430] ) | (~\[5704]  & ~\[5694] ),
  \[10156]  = (~\[5946]  & ~\[8465] ) | (~\[8563]  & ~sh2),
  \[6039]  = (~\[5843]  & ~\[5840] ) | ~\[8693] ,
  \[10536]  = ~inD4 | (~musel4 | (~\[5523]  | ~\[2355] )),
  \[9674]  = \[5825]  | \[8655] ,
  \[10726]  = ~\[6044]  | ~\[5870] ,
  \[9864]  = ~\[8817]  | ~\[5671] ,
  \[360]  = (~inA2 & ~\[4540] ) | ((~inA2 & ~musel1) | ((~\[9539]  & ~\[4540] ) | (~\[9539]  & ~musel1))),
  \[9677]  = ~\[8655]  | ~\[5825] ,
  \[362]  = (~inB2 & ~\[2062] ) | ((~inB2 & ~musel1) | ((~\[9543]  & ~\[2062] ) | (~\[9543]  & ~musel1))),
  \[9867]  = \[5653]  | \[8802] ,
  \[10352]  = ~sh2 | ~\[8562] ,
  \[173]  = (~\[1235]  & ~\[9117] ) | (~\[1235]  & ~\[5536] ),
  \[10922]  = ~inD9 | (~musel4 | (~\[5523]  | ~\[3079] )),
  \[9299]  = ~\[244] ,
  \[2814]  = ~\[5690]  & ~\[5528] ,
  \[5690]  = ~inD7,
  \[5880]  = ~musel4 | (~\[5523]  | ~\[9497] ),
  \[555]  = (~\[5976]  & ~\[10025] ) | ((~\[5976]  & ~\[8313] ) | ((~\[8181]  & ~\[10025] ) | (~\[8181]  & ~\[8313] ))),
  \[5881]  = (~\[5880]  & ~\[8195] ) | ~\[11374] ,
  \[556]  = (~\[5978]  & ~\[10029] ) | (~\[5978]  & ~\[5948] ),
  \[177]  = (~opsel0 & ~opsel1) | ((~opsel0 & ~\[5535] ) | ((~\[5534]  & ~opsel1) | (~\[5534]  & ~\[5535] ))),
  \[5882]  = ~inC4 | ~musel2,
  \[367]  = (~inA1 & ~inC1) | ((~inA1 & ~musel2) | ((~\[5528]  & ~inC1) | (~\[5528]  & ~musel2))),
  \[2817]  = ~musel1 & ~musel2,
  \[6042]  = ~\[12790] ,
  \[178]  = (~\[1200]  & ~\[9130] ) | (~\[1200]  & ~\[5951] ),
  \[368]  = (~inA1 & ~\[4466] ) | ((~inA1 & ~musel1) | ((~\[9555]  & ~\[4466] ) | (~\[9555]  & ~musel1))),
  \[10168]  = (~\[5946]  & ~\[8492] ) | (~\[8587]  & ~sh2),
  \[5694]  = (~\[1490]  & ~\[1489] ) | ~\[5525] ,
  \[179]  = (~\[8905]  & ~opsel2) | ((~\[8905]  & ~\[8950] ) | ((~\[5550]  & ~opsel2) | (~\[5550]  & ~\[8950] ))),
  \[6044]  = ~\[12790]  | (~\[5886]  | (~\[5881]  | ~\[5875] )),
  \[5695]  = ~inC7 | ~musel4,
  \[5885]  = ~musel4 | (~\[5523]  | ~\[9513] ),
  \[6045]  = ~opsel2 | ~\[8926] ,
  \[4338]  = ~\[5825]  & ~\[8655] ,
  \[5886]  = (~\[5885]  & ~\[8195] ) | ~\[11366] ,
  \[9870]  = ~\[8802]  | ~\[5653] ,
  \[9491]  = (~\[5529]  & ~musel2) | (~\[5528]  & ~musel1),
  \[10164]  = (~\[8541]  & ~sh2) | ~\[10204] ,
  \[5888]  = ~\[5886]  | (~\[5881]  | (~\[5875]  | ~\[5870] )),
  \[5889]  = ~inC11 | ~musel2,
  \[8705]  = ~\[5704] ,
  \[10166]  = (~\[5946]  & ~\[8419] ) | (~\[8563]  & ~sh2),
  \[9495]  = (~\[5529]  & ~musel2) | (~\[5528]  & ~musel1),
  \[370]  = (~inB1 & ~\[1910] ) | ((~inB1 & ~musel1) | ((~\[9559]  & ~\[1910] ) | (~\[9559]  & ~musel1))),
  \[10170]  = (~\[5946]  & ~\[8521] ) | (~\[8612]  & ~sh2),
  \[8328]  = ~\[5617] ,
  \[9876]  = (~\[5994]  & ~\[503] ) | ~\[9883] ,
  \[561]  = (~\[1107]  & ~sh2) | (~\[1107]  & ~\[8335] ),
  \[751]  = ~\[6087]  & ~\[6081] ,
  \[2062]  = ~\[5785]  & ~\[5528] ,
  \[9497]  = (~\[5877]  & ~musel1) | ~\[11380] ,
  \[182]  = (~opsel0 & ~opsel1) | ((~opsel0 & ~\[5535] ) | ((~\[5534]  & ~opsel1) | (~\[5534]  & ~\[5535] ))),
  \[562]  = (~\[1105]  & ~\[8335] ) | (~\[1105]  & ~\[5947] ),
  \[10172]  = ~opsel3 | (~\[5550]  | ~\[9314] ),
  \[183]  = (~\[1167]  & ~\[9143] ) | (~\[1167]  & ~\[5966] ),
  \[563]  = (~\[10048]  & ~sh1) | ((~\[10048]  & ~\[10044] ) | ((~\[5947]  & ~sh1) | (~\[5947]  & ~\[10044] ))),
  \[184]  = (~\[8908]  & ~opsel2) | ((~\[8908]  & ~\[8953] ) | ((~\[5550]  & ~opsel2) | (~\[5550]  & ~\[8953] ))),
  \[564]  = (~\[10050]  & ~sh1) | ((~\[10050]  & ~\[10046] ) | ((~\[5947]  & ~sh1) | (~\[5947]  & ~\[10046] ))),
  \[2065]  = ~musel1 & ~musel2,
  \[375]  = (~inA0 & ~inC0) | ((~inA0 & ~musel2) | ((~\[5528]  & ~inC0) | (~\[5528]  & ~musel2))),
  \[6050]  = ~musel3 | ~\[5525] ,
  \[376]  = (~inA0 & ~\[4392] ) | ((~inA0 & ~musel1) | ((~\[9571]  & ~\[4392] ) | (~\[9571]  & ~musel1))),
  \[6051]  = ~\[5535]  | ~\[5534] ,
  \[187]  = (~opsel0 & ~opsel1) | ((~opsel0 & ~\[5535] ) | ((~\[5534]  & ~opsel1) | (~\[5534]  & ~\[5535] ))),
  \[5892]  = ~musel4 | (~\[5523]  | ~\[9401] ),
  \[6052]  = (~\[8714]  & ~\[8451] ) | (~\[5722]  & ~\[5712] ),
  \[188]  = (~\[1136]  & ~\[9156] ) | (~\[1136]  & ~\[5979] );
endmodule

