//
// Conformal-LEC Version 14.20-d237 ( 26-Mar-2015) ( 64 bit executable)
//
module top ( PI_clock , PI_reset , n0 , n1 , n2 , n3 , n4 , n5 , n6 , 
  n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , 
  n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , 
  n27 , n28 , n29 , n30 , n31 , DFF_state_reg_Q , n32 , n33 , n34 , n35 , 
  n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , 
  n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , 
  n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , 
  n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , 
  n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , 
  n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , 
  n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , 
  n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , 
  n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , 
  n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , 
  n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , 
  n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , 
  n156 , n157 , n158 , DFF_B_reg_Q , n159 , n160 , n161 , n162 , n163 , n164 , 
  n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , 
  n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , 
  n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , 
  n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , 
  n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , 
  n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , 
  n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , 
  n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , DFF_rd_reg_Q , DFF_wr_reg_Q , 
  n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , 
  n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , 
  n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , 
  n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , 
  n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , 
  n293 , n294 , PO_rd , PO_wr , DFF_state_reg_S , DFF_state_reg_R , DFF_state_reg_CK , DFF_state_reg_D , n295 , n296 , 
  n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , 
  n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , 
  n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , 
  n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , 
  n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , 
  n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , 
  n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , 
  n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , 
  n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , 
  n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , 
  n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , 
  n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , 
  n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , 
  n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , 
  n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , 
  n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , 
  n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , 
  n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , 
  n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , 
  n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , 
  n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , 
  n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , 
  n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , 
  n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , 
  n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , 
  n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , 
  n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , 
  n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , 
  n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , 
  n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , 
  n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , 
  n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , 
  n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , 
  n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , 
  n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , 
  n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , 
  n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , 
  n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , 
  n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , 
  n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , 
  n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , 
  n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , 
  n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , 
  n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , 
  n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , 
  n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , 
  n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , 
  n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , 
  n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , 
  n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , 
  n797 , n798 , n799 , n800 , n801 , n802 , DFF_B_reg_S , DFF_B_reg_R , DFF_B_reg_CK , DFF_B_reg_D , 
  n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , 
  n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , 
  n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , 
  n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , 
  n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , 
  n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , 
  n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , 
  n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , 
  n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , 
  n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , 
  n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , 
  n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , 
  n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , 
  n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , 
  n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , 
  n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , 
  n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , 
  n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , 
  n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , 
  n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , 
  n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , 
  n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , 
  n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , 
  n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , 
  n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , 
  n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , 
  n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , 
  n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , 
  n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , 
  n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , 
  n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , 
  n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , 
  n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , 
  n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , DFF_rd_reg_S , DFF_rd_reg_R , DFF_rd_reg_CK , DFF_rd_reg_D , 
  DFF_wr_reg_S , DFF_wr_reg_R , DFF_wr_reg_CK , DFF_wr_reg_D);
input PI_clock , PI_reset , n0 , n1 , n2 , n3 , n4 , n5 , n6 , 
  n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , 
  n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , 
  n27 , n28 , n29 , n30 , n31 , DFF_state_reg_Q , n32 , n33 , n34 , n35 , 
  n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , 
  n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , 
  n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , 
  n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , 
  n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , 
  n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , 
  n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , 
  n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , 
  n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , 
  n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , 
  n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , 
  n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , 
  n156 , n157 , n158 , DFF_B_reg_Q , n159 , n160 , n161 , n162 , n163 , n164 , 
  n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , 
  n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , 
  n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , 
  n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , 
  n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , 
  n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , 
  n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , 
  n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , DFF_rd_reg_Q , DFF_wr_reg_Q;
output n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , 
  n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , 
  n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , 
  n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , 
  n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , 
  n292 , n293 , n294 , PO_rd , PO_wr , DFF_state_reg_S , DFF_state_reg_R , DFF_state_reg_CK , DFF_state_reg_D , n295 , 
  n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , 
  n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , 
  n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , 
  n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , 
  n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , 
  n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , 
  n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , 
  n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , 
  n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , 
  n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , 
  n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , 
  n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , 
  n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , 
  n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , 
  n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , 
  n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , 
  n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , 
  n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , 
  n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , 
  n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , 
  n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , 
  n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , 
  n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , 
  n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , 
  n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , 
  n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , 
  n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , 
  n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , 
  n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , 
  n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , 
  n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , 
  n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , 
  n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , 
  n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , 
  n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , 
  n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , 
  n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , 
  n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , 
  n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , 
  n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , 
  n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , 
  n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , 
  n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , 
  n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , 
  n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , 
  n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , 
  n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , 
  n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , 
  n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , 
  n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , 
  n796 , n797 , n798 , n799 , n800 , n801 , n802 , DFF_B_reg_S , DFF_B_reg_R , DFF_B_reg_CK , 
  DFF_B_reg_D , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , 
  n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , 
  n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , 
  n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , 
  n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , 
  n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , 
  n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , 
  n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , 
  n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , 
  n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , 
  n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , 
  n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , 
  n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , 
  n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , 
  n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , 
  n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , 
  n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , 
  n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , 
  n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , 
  n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , 
  n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , 
  n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , 
  n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , 
  n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , 
  n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , 
  n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , 
  n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , 
  n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , 
  n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , 
  n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , 
  n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , 
  n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , 
  n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , 
  n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , DFF_rd_reg_S , DFF_rd_reg_R , DFF_rd_reg_CK , 
  DFF_rd_reg_D , DFF_wr_reg_S , DFF_wr_reg_R , DFF_wr_reg_CK , DFF_wr_reg_D;

wire n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , 
   n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , 
   n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , 
   n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , 
   n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , 
   n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , 
   n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , 
   n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , 
   n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , 
   n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , 
   n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , 
   n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , 
   n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , 
   n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , 
   n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , 
   n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , 
   n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , 
   n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , 
   n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , 
   n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , 
   n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , 
   n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , 
   n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , 
   n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , 
   n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , 
   n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , 
   n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , 
   n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , 
   n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , 
   n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , 
   n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , 
   n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , 
   n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , 
   n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , 
   n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , 
   n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , 
   n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , 
   n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , 
   n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , 
   n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , 
   n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , 
   n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , 
   n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , 
   n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , 
   n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , 
   n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , 
   n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , 
   n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , 
   n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , 
   n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , 
   n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , 
   n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , 
   n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , 
   n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , 
   n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , 
   n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , 
   n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , 
   n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , 
   n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , 
   n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , 
   n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , 
   n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , 
   n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , 
   n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , 
   n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , 
   n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , 
   n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , 
   n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , 
   n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , 
   n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , 
   n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , 
   n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , 
   n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , 
   n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , 
   n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , 
   n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , 
   n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , 
   n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , 
   n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , 
   n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , 
   n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , 
   n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , 
   n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , 
   n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , 
   n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , 
   n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , 
   n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , 
   n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , 
   n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , 
   n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , 
   n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , 
   n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , 
   n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , 
   n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , 
   n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , 
   n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , 
   n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , 
   n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , 
   n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , 
   n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , 
   n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , 
   n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , 
   n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , 
   n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , 
   n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , 
   n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , 
   n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , 
   n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , 
   n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , 
   n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , 
   n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , 
   n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , 
   n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , 
   n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , 
   n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , 
   n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , 
   n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , 
   n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , 
   n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , 
   n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , 
   n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , 
   n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , 
   n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , 
   n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , 
   n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , 
   n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , 
   n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , 
   n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , 
   n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , 
   n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , 
   n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , 
   n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , 
   n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , 
   n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , 
   n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , 
   n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , 
   n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , 
   n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , 
   n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , 
   n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , 
   n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , 
   n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , 
   n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , 
   n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , 
   n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , 
   n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , 
   n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , 
   n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , 
   n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , 
   n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , 
   n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , 
   n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , 
   n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , 
   n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , 
   n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , 
   n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , 
   n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , 
   n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , 
   n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , 
   n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , 
   n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , 
   n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , 
   n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , 
   n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , 
   n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , 
   n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , 
   n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , 
   n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , 
   n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , 
   n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , 
   n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , 
   n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , 
   n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , 
   n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , 
   n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , 
   n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , 
   n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , 
   n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , 
   n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , 
   n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , 
   n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , 
   n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , 
   n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , 
   n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , 
   n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , 
   n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , 
   n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , 
   n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , 
   n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , 
   n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , 
   n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , 
   n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , 
   n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , 
   n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , 
   n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , 
   n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , 
   n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , 
   n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , 
   n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , 
   n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , 
   n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , 
   n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , 
   n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , 
   n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , 
   n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , 
   n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , 
   n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , 
   n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , 
   n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , 
   n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , 
   n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , 
   n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , 
   n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , 
   n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , 
   n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , 
   n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , 
   n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , 
   n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , 
   n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , 
   n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , 
   n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , 
   n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , 
   n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , 
   n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , 
   n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , 
   n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , 
   n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , 
   n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , 
   n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , 
   n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , 
   n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , 
   n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , 
   n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , 
   n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , 
   n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , 
   n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , 
   n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , 
   n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , 
   n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , 
   n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , 
   n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , 
   n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , 
   n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , 
   n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , 
   n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , 
   n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , 
   n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , 
   n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , 
   n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , 
   n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , 
   n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , 
   n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , 
   n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , 
   n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , 
   n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , 
   n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , 
   n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , 
   n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , 
   n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , 
   n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , 
   n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , 
   n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , 
   n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , 
   n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , 
   n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , 
   n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , 
   n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , 
   n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , 
   n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , 
   n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , 
   n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , 
   n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , 
   n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , 
   n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , 
   n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , 
   n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , 
   n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , 
   n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , 
   n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , 
   n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , 
   n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , 
   n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , 
   n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , 
   n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , 
   n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , 
   n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , 
   n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , 
   n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , 
   n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , 
   n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , 
   n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , 
   n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , 
   n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , 
   n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , 
   n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , 
   n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , 
   n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , 
   n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , 
   n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , 
   n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , 
   n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , 
   n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , 
   n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , 
   n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , 
   n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , 
   n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , 
   n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , 
   n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , 
   n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , 
   n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , 
   n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , 
   n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , 
   n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , 
   n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , 
   n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , 
   n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , 
   n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , 
   n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , 
   n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , 
   n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , 
   n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , 
   n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , 
   n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , 
   n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , 
   n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , 
   n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , 
   n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , 
   n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , 
   n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , 
   n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , 
   n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , 
   n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , 
   n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , 
   n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , 
   n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , 
   n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , 
   n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , 
   n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , 
   n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , 
   n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , 
   n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , 
   n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , 
   n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , 
   n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , 
   n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , 
   n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , 
   n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , 
   n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , 
   n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , 
   n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , 
   n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , 
   n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , 
   n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , 
   n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , 
   n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , 
   n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , 
   n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , 
   n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , 
   n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , 
   n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , 
   n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , 
   n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , 
   n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , 
   n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , 
   n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , 
   n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , 
   n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , 
   n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , 
   n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , 
   n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , 
   n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , 
   n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , 
   n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , 
   n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , 
   n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , 
   n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , 
   n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , 
   n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , 
   n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , 
   n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , 
   n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , 
   n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , 
   n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , 
   n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , 
   n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , 
   n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , 
   n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , 
   n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , 
   n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , 
   n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , 
   n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , 
   n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , 
   n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , 
   n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , 
   n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , 
   n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , 
   n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , 
   n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , 
   n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , 
   n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , 
   n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , 
   n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , 
   n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , 
   n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , 
   n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , 
   n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , 
   n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , 
   n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , 
   n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , 
   n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , 
   n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , 
   n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , 
   n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , 
   n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , 
   n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , 
   n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , 
   n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , 
   n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , 
   n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , 
   n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , 
   n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , 
   n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , 
   n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , 
   n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , 
   n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , 
   n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , 
   n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , 
   n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , 
   n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , 
   n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , 
   n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , 
   n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , 
   n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , 
   n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , 
   n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , 
   n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , 
   n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , 
   n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , 
   n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , 
   n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , 
   n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , 
   n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , 
   n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , 
   n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , 
   n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , 
   n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , 
   n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , 
   n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , 
   n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , 
   n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , 
   n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , 
   n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , 
   n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , 
   n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , 
   n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , 
   n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , 
   n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , 
   n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , 
   n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , 
   n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , 
   n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , 
   n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , 
   n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , 
   n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , 
   n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , 
   n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , 
   n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , 
   n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , 
   n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , 
   n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , 
   n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , 
   n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , 
   n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , 
   n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , 
   n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , 
   n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , 
   n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , 
   n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , 
   n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , 
   n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , 
   n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , 
   n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , 
   n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , 
   n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , 
   n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , 
   n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , 
   n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , 
   n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , 
   n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , 
   n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , 
   n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , 
   n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , 
   n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , 
   n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , 
   n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , 
   n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , 
   n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , 
   n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , 
   n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , 
   n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , 
   n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , 
   n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , 
   n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , 
   n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , 
   n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , 
   n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , 
   n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , 
   n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , 
   n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , 
   n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , 
   n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , 
   n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , 
   n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , 
   n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , 
   n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , 
   n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , 
   n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , 
   n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , 
   n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , 
   n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , 
   n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , 
   n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , 
   n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , 
   n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , 
   n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , 
   n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , 
   n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , 
   n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , 
   n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , 
   n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , 
   n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , 
   n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , 
   n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , 
   n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , 
   n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , 
   n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , 
   n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , 
   n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , 
   n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , 
   n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , 
   n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , 
   n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , 
   n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , 
   n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , 
   n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , 
   n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , 
   n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , 
   n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , 
   n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , 
   n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , 
   n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , 
   n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , 
   n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , 
   n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , 
   n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , 
   n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , 
   n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , 
   n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , 
   n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , 
   n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , 
   n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , 
   n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , 
   n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , 
   n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , 
   n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , 
   n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , 
   n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , 
   n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , 
   n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , 
   n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , 
   n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , 
   n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , 
   n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , 
   n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , 
   n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , 
   n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , 
   n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , 
   n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , 
   n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , 
   n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , 
   n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , 
   n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , 
   n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , 
   n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , 
   n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , 
   n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , 
   n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , 
   n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , 
   n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , 
   n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , 
   n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , 
   n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , 
   n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , 
   n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , 
   n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , 
   n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , 
   n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , 
   n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , 
   n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , 
   n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , 
   n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , 
   n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , 
   n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , 
   n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , 
   n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , 
   n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , 
   n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , 
   n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , 
   n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , 
   n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , 
   n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , 
   n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , 
   n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , 
   n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , 
   n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , 
   n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , 
   n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , 
   n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , 
   n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , 
   n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , 
   n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , 
   n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , 
   n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , 
   n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , 
   n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , 
   n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , 
   n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , 
   n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , 
   n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , 
   n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , 
   n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , 
   n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , 
   n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , 
   n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , 
   n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , 
   n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , 
   n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , 
   n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , 
   n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , 
   n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , 
   n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , 
   n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , 
   n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , 
   n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , 
   n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , 
   n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , 
   n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , 
   n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , 
   n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , 
   n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , 
   n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , 
   n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , 
   n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , 
   n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , 
   n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , 
   n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , 
   n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , 
   n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , 
   n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , 
   n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , 
   n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , 
   n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , 
   n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , 
   n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , 
   n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , 
   n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , 
   n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , 
   n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , 
   n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , 
   n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , 
   n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , 
   n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , 
   n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , 
   n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , 
   n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , 
   n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , 
   n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , 
   n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , 
   n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , 
   n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , 
   n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , 
   n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , 
   n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , 
   n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , 
   n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , 
   n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , 
   n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , 
   n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , 
   n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , 
   n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , 
   n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , 
   n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , 
   n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , 
   n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , 
   n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , 
   n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , 
   n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , 
   n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , 
   n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , 
   n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , 
   n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , 
   n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , 
   n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , 
   n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , 
   n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , 
   n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , 
   n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , 
   n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , 
   n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , 
   n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , 
   n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , 
   n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , 
   n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , 
   n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , 
   n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , 
   n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , 
   n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , 
   n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , 
   n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , 
   n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , 
   n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , 
   n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , 
   n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , 
   n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , 
   n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , 
   n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , 
   n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , 
   n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , 
   n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , 
   n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , 
   n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , 
   n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , 
   n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , 
   n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , 
   n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , 
   n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , 
   n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , 
   n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , 
   n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , 
   n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , 
   n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , 
   n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , 
   n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , 
   n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , 
   n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , 
   n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , 
   n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , 
   n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , 
   n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , 
   n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , 
   n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , 
   n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , 
   n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , 
   n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , 
   n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , 
   n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , 
   n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , 
   n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , 
   n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , 
   n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , 
   n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , 
   n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , 
   n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , 
   n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , 
   n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , 
   n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , 
   n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , 
   n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , 
   n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , 
   n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , 
   n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , 
   n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , 
   n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , 
   n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , 
   n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , 
   n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , 
   n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , 
   n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , 
   n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , 
   n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , 
   n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , 
   n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , 
   n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , 
   n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , 
   n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , 
   n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , 
   n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , 
   n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , 
   n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , 
   n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , 
   n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , 
   n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , 
   n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , 
   n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , 
   n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , 
   n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , 
   n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , 
   n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , 
   n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , 
   n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , 
   n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , 
   n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , 
   n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , 
   n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , 
   n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , 
   n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , 
   n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , 
   n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , 
   n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , 
   n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , 
   n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , 
   n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , 
   n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , 
   n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , 
   n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , 
   n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , 
   n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , 
   n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , 
   n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , 
   n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , 
   n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , 
   n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , 
   n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , 
   n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , 
   n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , 
   n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , 
   n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , 
   n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , 
   n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , 
   n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , 
   n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , 
   n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , 
   n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , 
   n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , 
   n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , 
   n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , 
   n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , 
   n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , 
   n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , 
   n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , 
   n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , 
   n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , 
   n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , 
   n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , 
   n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , 
   n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , 
   n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , 
   n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , 
   n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , 
   n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , 
   n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , 
   n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , 
   n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , 
   n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , 
   n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , 
   n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , 
   n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , 
   n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , 
   n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , 
   n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , 
   n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , 
   n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , 
   n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , 
   n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , 
   n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , 
   n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , 
   n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , 
   n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , 
   n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , 
   n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , 
   n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , 
   n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , 
   n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , 
   n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , 
   n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , 
   n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , 
   n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , 
   n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , 
   n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , 
   n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , 
   n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , 
   n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , 
   n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , 
   n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , 
   n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , 
   n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , 
   n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , 
   n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , 
   n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , 
   n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , 
   n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , 
   n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , 
   n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , 
   n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , 
   n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , 
   n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , 
   n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , 
   n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , 
   n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , 
   n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , 
   n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , 
   n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , 
   n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , 
   n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , 
   n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , 
   n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , 
   n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , 
   n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , 
   n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , 
   n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , 
   n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , 
   n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , 
   n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , 
   n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , 
   n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , 
   n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , 
   n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , 
   n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , 
   n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , 
   n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , 
   n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , 
   n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , 
   n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , 
   n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , 
   n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , 
   n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , 
   n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , 
   n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , 
   n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , 
   n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , 
   n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , 
   n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , 
   n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , 
   n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , 
   n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , 
   n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , 
   n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , 
   n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , 
   n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , 
   n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , 
   n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , 
   n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , 
   n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , 
   n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , 
   n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , 
   n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , 
   n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , 
   n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , 
   n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , 
   n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , 
   n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , 
   n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , 
   n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , 
   n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , 
   n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , 
   n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , 
   n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , 
   n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , 
   n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , 
   n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , 
   n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , 
   n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , 
   n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , 
   n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , 
   n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , 
   n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , 
   n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , 
   n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , 
   n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , 
   n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , 
   n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , 
   n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , 
   n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , 
   n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , 
   n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , 
   n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , 
   n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , 
   n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , 
   n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , 
   n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , 
   n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , 
   n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , 
   n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , 
   n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , 
   n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , 
   n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , 
   n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , 
   n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , 
   n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , 
   n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , 
   n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , 
   n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , 
   n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , 
   n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , 
   n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , 
   n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , 
   n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , 
   n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , 
   n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , 
   n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , 
   n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , 
   n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , 
   n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , 
   n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , 
   n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , 
   n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , 
   n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , 
   n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , 
   n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , 
   n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , 
   n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , 
   n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , 
   n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , 
   n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , 
   n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , 
   n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , 
   n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , 
   n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , 
   n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , 
   n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , 
   n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , 
   n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , 
   n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , 
   n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , 
   n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , 
   n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , 
   n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , 
   n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , 
   n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , 
   n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , 
   n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , 
   n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , 
   n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , 
   n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , 
   n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , 
   n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , 
   n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , 
   n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , 
   n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , 
   n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , 
   n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , 
   n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , 
   n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , 
   n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , 
   n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , 
   n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , 
   n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , 
   n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , 
   n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , 
   n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , 
   n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , 
   n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , 
   n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , 
   n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , 
   n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , 
   n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , 
   n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , 
   n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , 
   n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , 
   n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , 
   n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , 
   n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , 
   n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , 
   n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , 
   n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , 
   n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , 
   n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , 
   n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , 
   n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , 
   n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , 
   n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , 
   n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , 
   n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , 
   n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , 
   n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , 
   n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , 
   n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , 
   n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , 
   n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , 
   n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , 
   n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , 
   n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , 
   n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , 
   n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , 
   n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , 
   n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , 
   n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , 
   n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , 
   n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , 
   n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , 
   n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , 
   n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , 
   n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , 
   n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , 
   n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , 
   n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , 
   n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , 
   n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , 
   n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , 
   n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , 
   n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , 
   n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , 
   n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , 
   n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , 
   n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , 
   n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , 
   n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , 
   n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , 
   n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , 
   n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , 
   n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , 
   n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , 
   n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , 
   n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , 
   n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , 
   n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , 
   n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , 
   n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , 
   n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , 
   n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , 
   n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , 
   n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , 
   n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , 
   n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , 
   n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , 
   n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , 
   n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , 
   n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , 
   n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , 
   n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , 
   n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , 
   n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , 
   n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , 
   n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , 
   n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , 
   n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , 
   n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , 
   n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , 
   n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , 
   n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , 
   n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , 
   n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , 
   n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , 
   n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , 
   n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , 
   n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , 
   n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , 
   n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , 
   n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , 
   n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , 
   n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , 
   n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , 
   n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , 
   n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , 
   n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , 
   n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , 
   n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , 
   n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , 
   n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , 
   n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , 
   n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , 
   n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , 
   n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , 
   n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , 
   n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , 
   n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , 
   n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , 
   n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , 
   n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , 
   n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , 
   n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , 
   n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , 
   n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , 
   n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , 
   n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , 
   n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , 
   n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , 
   n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , 
   n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , 
   n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , 
   n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , 
   n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , 
   n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , 
   n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , 
   n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , 
   n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , 
   n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , 
   n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , 
   n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , 
   n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , 
   n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , 
   n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , 
   n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , 
   n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , 
   n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , 
   n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , 
   n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , 
   n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , 
   n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , 
   n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , 
   n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , 
   n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , 
   n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , 
   n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , 
   n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , 
   n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , 
   n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , 
   n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , 
   n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , 
   n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , 
   n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , 
   n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , 
   n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , 
   n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , 
   n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , 
   n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , 
   n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , 
   n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , 
   n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , 
   n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , 
   n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , 
   n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , 
   n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , 
   n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , 
   n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , 
   n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , 
   n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , 
   n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , 
   n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , 
   n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , 
   n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , 
   n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , 
   n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , 
   n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , 
   n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , 
   n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , 
   n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , 
   n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , 
   n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , 
   n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , 
   n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , 
   n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , 
   n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , 
   n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , 
   n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , 
   n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , 
   n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , 
   n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , 
   n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , 
   n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , 
   n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , 
   n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , 
   n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , 
   n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , 
   n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , 
   n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , 
   n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , 
   n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , 
   n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , 
   n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , 
   n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , 
   n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , 
   n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , 
   n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , 
   n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , 
   n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , 
   n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , 
   n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , 
   n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , 
   n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , 
   n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , 
   n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , 
   n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , 
   n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , 
   n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , 
   n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , 
   n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , 
   n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , 
   n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , 
   n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , 
   n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , 
   n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , 
   n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , 
   n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , 
   n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , 
   n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , 
   n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , 
   n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , 
   n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , 
   n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , 
   n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , 
   n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , 
   n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , 
   n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , 
   n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , 
   n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , 
   n15237 , n15238 , n15239 , n15240 , n15241 , n15242 ;
buf ( n243 , n2315 );
buf ( n244 , n2317 );
buf ( n245 , n2319 );
buf ( n246 , n2321 );
buf ( n247 , n2323 );
buf ( n248 , n2325 );
buf ( n249 , n2327 );
buf ( n250 , n2329 );
buf ( n251 , n2331 );
buf ( n252 , n2333 );
buf ( n253 , n2335 );
buf ( n254 , n2337 );
buf ( n255 , n2339 );
buf ( n256 , n2341 );
buf ( n257 , n2343 );
buf ( n258 , n2345 );
buf ( n259 , n2347 );
buf ( n260 , n2349 );
buf ( n261 , n2351 );
buf ( n262 , n2353 );
buf ( n263 , n2355 );
buf ( n264 , n2357 );
buf ( n265 , n2359 );
buf ( n266 , n2361 );
buf ( n267 , n2363 );
buf ( n268 , n2365 );
buf ( n269 , n2367 );
buf ( n270 , n2369 );
buf ( n271 , n2371 );
buf ( n272 , n2373 );
buf ( n273 , n2375 );
buf ( n274 , n2377 );
buf ( n275 , n2379 );
buf ( n276 , n2381 );
buf ( n277 , n2383 );
buf ( n278 , n2385 );
buf ( n279 , n2387 );
buf ( n280 , n2389 );
buf ( n281 , n2391 );
buf ( n282 , n2393 );
buf ( n283 , n2395 );
buf ( n284 , n2397 );
buf ( n285 , n2399 );
buf ( n286 , n2401 );
buf ( n287 , n2403 );
buf ( n288 , n2405 );
buf ( n289 , n2407 );
buf ( n290 , n2409 );
buf ( n291 , n2411 );
buf ( n292 , n2413 );
buf ( n293 , n2415 );
buf ( n294 , n2417 );
buf ( PO_rd , n2419 );
buf ( PO_wr , n2421 );
buf ( DFF_state_reg_S , n2425 );
buf ( DFF_state_reg_R , n2426 );
buf ( DFF_state_reg_CK , n2427 );
buf ( DFF_state_reg_D , n2429 );
buf ( n295 , n2431 );
buf ( n296 , n2432 );
buf ( n297 , n2433 );
buf ( n298 , n2437 );
buf ( n299 , n2439 );
buf ( n300 , n2440 );
buf ( n301 , n2441 );
buf ( n302 , n2453 );
buf ( n303 , n2455 );
buf ( n304 , n2456 );
buf ( n305 , n2457 );
buf ( n306 , n2468 );
buf ( n307 , n2470 );
buf ( n308 , n2471 );
buf ( n309 , n2472 );
buf ( n310 , n2483 );
buf ( n311 , n2485 );
buf ( n312 , n2486 );
buf ( n313 , n2487 );
buf ( n314 , n2498 );
buf ( n315 , n2500 );
buf ( n316 , n2501 );
buf ( n317 , n2502 );
buf ( n318 , n2513 );
buf ( n319 , n2515 );
buf ( n320 , n2516 );
buf ( n321 , n2517 );
buf ( n322 , n2528 );
buf ( n323 , n2530 );
buf ( n324 , n2531 );
buf ( n325 , n2532 );
buf ( n326 , n2543 );
buf ( n327 , n2545 );
buf ( n328 , n2546 );
buf ( n329 , n2547 );
buf ( n330 , n2558 );
buf ( n331 , n2560 );
buf ( n332 , n2561 );
buf ( n333 , n2562 );
buf ( n334 , n2573 );
buf ( n335 , n2575 );
buf ( n336 , n2576 );
buf ( n337 , n2577 );
buf ( n338 , n2588 );
buf ( n339 , n2590 );
buf ( n340 , n2591 );
buf ( n341 , n2592 );
buf ( n342 , n2603 );
buf ( n343 , n2605 );
buf ( n344 , n2606 );
buf ( n345 , n2607 );
buf ( n346 , n2618 );
buf ( n347 , n2620 );
buf ( n348 , n2621 );
buf ( n349 , n2622 );
buf ( n350 , n2633 );
buf ( n351 , n2635 );
buf ( n352 , n2636 );
buf ( n353 , n2637 );
buf ( n354 , n2648 );
buf ( n355 , n2650 );
buf ( n356 , n2651 );
buf ( n357 , n2652 );
buf ( n358 , n2663 );
buf ( n359 , n2665 );
buf ( n360 , n2666 );
buf ( n361 , n2667 );
buf ( n362 , n2678 );
buf ( n363 , n2680 );
buf ( n364 , n2681 );
buf ( n365 , n2682 );
buf ( n366 , n2693 );
buf ( n367 , n2695 );
buf ( n368 , n2696 );
buf ( n369 , n2697 );
buf ( n370 , n2708 );
buf ( n371 , n2710 );
buf ( n372 , n2711 );
buf ( n373 , n2712 );
buf ( n374 , n2723 );
buf ( n375 , n2725 );
buf ( n376 , n2726 );
buf ( n377 , n2727 );
buf ( n378 , n2738 );
buf ( n379 , n2740 );
buf ( n380 , n2741 );
buf ( n381 , n2742 );
buf ( n382 , n2753 );
buf ( n383 , n2755 );
buf ( n384 , n2756 );
buf ( n385 , n2757 );
buf ( n386 , n2768 );
buf ( n387 , n2770 );
buf ( n388 , n2771 );
buf ( n389 , n2772 );
buf ( n390 , n2783 );
buf ( n391 , n2785 );
buf ( n392 , n2786 );
buf ( n393 , n2787 );
buf ( n394 , n2798 );
buf ( n395 , n2800 );
buf ( n396 , n2801 );
buf ( n397 , n2802 );
buf ( n398 , n2813 );
buf ( n399 , n2815 );
buf ( n400 , n2816 );
buf ( n401 , n2817 );
buf ( n402 , n2828 );
buf ( n403 , n2830 );
buf ( n404 , n2831 );
buf ( n405 , n2832 );
buf ( n406 , n2843 );
buf ( n407 , n2845 );
buf ( n408 , n2846 );
buf ( n409 , n2847 );
buf ( n410 , n2858 );
buf ( n411 , n2860 );
buf ( n412 , n2861 );
buf ( n413 , n2862 );
buf ( n414 , n2873 );
buf ( n415 , n2875 );
buf ( n416 , n2876 );
buf ( n417 , n2877 );
buf ( n418 , n2888 );
buf ( n419 , n2889 );
buf ( n420 , n2890 );
buf ( n421 , n2891 );
buf ( n422 , n2903 );
buf ( n423 , n2905 );
buf ( n424 , n2906 );
buf ( n425 , n2907 );
buf ( n426 , n3311 );
buf ( n427 , n3313 );
buf ( n428 , n3314 );
buf ( n429 , n3315 );
buf ( n430 , n3355 );
buf ( n431 , n3357 );
buf ( n432 , n3358 );
buf ( n433 , n3359 );
buf ( n434 , n6734 );
buf ( n435 , n6735 );
buf ( n436 , n6736 );
buf ( n437 , n6737 );
buf ( n438 , n7090 );
buf ( n439 , n7091 );
buf ( n440 , n7092 );
buf ( n441 , n7093 );
buf ( n442 , n7164 );
buf ( n443 , n7165 );
buf ( n444 , n7166 );
buf ( n445 , n7167 );
buf ( n446 , n7238 );
buf ( n447 , n7239 );
buf ( n448 , n7240 );
buf ( n449 , n7241 );
buf ( n450 , n7312 );
buf ( n451 , n7313 );
buf ( n452 , n7314 );
buf ( n453 , n7315 );
buf ( n454 , n7386 );
buf ( n455 , n7387 );
buf ( n456 , n7388 );
buf ( n457 , n7389 );
buf ( n458 , n7460 );
buf ( n459 , n7461 );
buf ( n460 , n7462 );
buf ( n461 , n7463 );
buf ( n462 , n7534 );
buf ( n463 , n7535 );
buf ( n464 , n7536 );
buf ( n465 , n7537 );
buf ( n466 , n7608 );
buf ( n467 , n7609 );
buf ( n468 , n7610 );
buf ( n469 , n7611 );
buf ( n470 , n7682 );
buf ( n471 , n7683 );
buf ( n472 , n7684 );
buf ( n473 , n7685 );
buf ( n474 , n7756 );
buf ( n475 , n7757 );
buf ( n476 , n7758 );
buf ( n477 , n7759 );
buf ( n478 , n7830 );
buf ( n479 , n7831 );
buf ( n480 , n7832 );
buf ( n481 , n7833 );
buf ( n482 , n7904 );
buf ( n483 , n7905 );
buf ( n484 , n7906 );
buf ( n485 , n7907 );
buf ( n486 , n7978 );
buf ( n487 , n7979 );
buf ( n488 , n7980 );
buf ( n489 , n7981 );
buf ( n490 , n8052 );
buf ( n491 , n8053 );
buf ( n492 , n8054 );
buf ( n493 , n8055 );
buf ( n494 , n8126 );
buf ( n495 , n8127 );
buf ( n496 , n8128 );
buf ( n497 , n8129 );
buf ( n498 , n8200 );
buf ( n499 , n8201 );
buf ( n500 , n8202 );
buf ( n501 , n8203 );
buf ( n502 , n8274 );
buf ( n503 , n8275 );
buf ( n504 , n8276 );
buf ( n505 , n8277 );
buf ( n506 , n8348 );
buf ( n507 , n8349 );
buf ( n508 , n8350 );
buf ( n509 , n8351 );
buf ( n510 , n8422 );
buf ( n511 , n8423 );
buf ( n512 , n8424 );
buf ( n513 , n8425 );
buf ( n514 , n8496 );
buf ( n515 , n8497 );
buf ( n516 , n8498 );
buf ( n517 , n8499 );
buf ( n518 , n8570 );
buf ( n519 , n8571 );
buf ( n520 , n8572 );
buf ( n521 , n8573 );
buf ( n522 , n8644 );
buf ( n523 , n8645 );
buf ( n524 , n8646 );
buf ( n525 , n8647 );
buf ( n526 , n8718 );
buf ( n527 , n8719 );
buf ( n528 , n8720 );
buf ( n529 , n8721 );
buf ( n530 , n8792 );
buf ( n531 , n8793 );
buf ( n532 , n8794 );
buf ( n533 , n8795 );
buf ( n534 , n8866 );
buf ( n535 , n8867 );
buf ( n536 , n8868 );
buf ( n537 , n8869 );
buf ( n538 , n8940 );
buf ( n539 , n8941 );
buf ( n540 , n8942 );
buf ( n541 , n8943 );
buf ( n542 , n9014 );
buf ( n543 , n9015 );
buf ( n544 , n9016 );
buf ( n545 , n9017 );
buf ( n546 , n9088 );
buf ( n547 , n9089 );
buf ( n548 , n9090 );
buf ( n549 , n9091 );
buf ( n550 , n9125 );
buf ( n551 , n9126 );
buf ( n552 , n9127 );
buf ( n553 , n9128 );
buf ( n554 , n9158 );
buf ( n555 , n9159 );
buf ( n556 , n9160 );
buf ( n557 , n9161 );
buf ( n558 , n9191 );
buf ( n559 , n9192 );
buf ( n560 , n9193 );
buf ( n561 , n9194 );
buf ( n562 , n9224 );
buf ( n563 , n9225 );
buf ( n564 , n9226 );
buf ( n565 , n9227 );
buf ( n566 , n9257 );
buf ( n567 , n9258 );
buf ( n568 , n9259 );
buf ( n569 , n9260 );
buf ( n570 , n9290 );
buf ( n571 , n9291 );
buf ( n572 , n9292 );
buf ( n573 , n9293 );
buf ( n574 , n9323 );
buf ( n575 , n9324 );
buf ( n576 , n9325 );
buf ( n577 , n9326 );
buf ( n578 , n9356 );
buf ( n579 , n9357 );
buf ( n580 , n9358 );
buf ( n581 , n9359 );
buf ( n582 , n9389 );
buf ( n583 , n9390 );
buf ( n584 , n9391 );
buf ( n585 , n9392 );
buf ( n586 , n9422 );
buf ( n587 , n9423 );
buf ( n588 , n9424 );
buf ( n589 , n9425 );
buf ( n590 , n9455 );
buf ( n591 , n9456 );
buf ( n592 , n9457 );
buf ( n593 , n9458 );
buf ( n594 , n9488 );
buf ( n595 , n9489 );
buf ( n596 , n9490 );
buf ( n597 , n9491 );
buf ( n598 , n9521 );
buf ( n599 , n9522 );
buf ( n600 , n9523 );
buf ( n601 , n9524 );
buf ( n602 , n9554 );
buf ( n603 , n9555 );
buf ( n604 , n9556 );
buf ( n605 , n9557 );
buf ( n606 , n9587 );
buf ( n607 , n9588 );
buf ( n608 , n9589 );
buf ( n609 , n9590 );
buf ( n610 , n9620 );
buf ( n611 , n9621 );
buf ( n612 , n9622 );
buf ( n613 , n9623 );
buf ( n614 , n9653 );
buf ( n615 , n9654 );
buf ( n616 , n9655 );
buf ( n617 , n9656 );
buf ( n618 , n9686 );
buf ( n619 , n9687 );
buf ( n620 , n9688 );
buf ( n621 , n9689 );
buf ( n622 , n9719 );
buf ( n623 , n9720 );
buf ( n624 , n9721 );
buf ( n625 , n9722 );
buf ( n626 , n9752 );
buf ( n627 , n9753 );
buf ( n628 , n9754 );
buf ( n629 , n9755 );
buf ( n630 , n9785 );
buf ( n631 , n9786 );
buf ( n632 , n9787 );
buf ( n633 , n9788 );
buf ( n634 , n9818 );
buf ( n635 , n9819 );
buf ( n636 , n9820 );
buf ( n637 , n9821 );
buf ( n638 , n9851 );
buf ( n639 , n9852 );
buf ( n640 , n9853 );
buf ( n641 , n9854 );
buf ( n642 , n9884 );
buf ( n643 , n9885 );
buf ( n644 , n9886 );
buf ( n645 , n9887 );
buf ( n646 , n9917 );
buf ( n647 , n9918 );
buf ( n648 , n9919 );
buf ( n649 , n9920 );
buf ( n650 , n9950 );
buf ( n651 , n9951 );
buf ( n652 , n9952 );
buf ( n653 , n9953 );
buf ( n654 , n9983 );
buf ( n655 , n9984 );
buf ( n656 , n9985 );
buf ( n657 , n9986 );
buf ( n658 , n10016 );
buf ( n659 , n10017 );
buf ( n660 , n10018 );
buf ( n661 , n10019 );
buf ( n662 , n10049 );
buf ( n663 , n10050 );
buf ( n664 , n10051 );
buf ( n665 , n10052 );
buf ( n666 , n10125 );
buf ( n667 , n10126 );
buf ( n668 , n10127 );
buf ( n669 , n10128 );
buf ( n670 , n10190 );
buf ( n671 , n10191 );
buf ( n672 , n10192 );
buf ( n673 , n10193 );
buf ( n674 , n10230 );
buf ( n675 , n10231 );
buf ( n676 , n10232 );
buf ( n677 , n10233 );
buf ( n678 , n10266 );
buf ( n679 , n10267 );
buf ( n680 , n10268 );
buf ( n681 , n10269 );
buf ( n682 , n10299 );
buf ( n683 , n10300 );
buf ( n684 , n10301 );
buf ( n685 , n10302 );
buf ( n686 , n10332 );
buf ( n687 , n10333 );
buf ( n688 , n10334 );
buf ( n689 , n10335 );
buf ( n690 , n10365 );
buf ( n691 , n10366 );
buf ( n692 , n10367 );
buf ( n693 , n10368 );
buf ( n694 , n10398 );
buf ( n695 , n10399 );
buf ( n696 , n10400 );
buf ( n697 , n10401 );
buf ( n698 , n10431 );
buf ( n699 , n10432 );
buf ( n700 , n10433 );
buf ( n701 , n10434 );
buf ( n702 , n10464 );
buf ( n703 , n10465 );
buf ( n704 , n10466 );
buf ( n705 , n10467 );
buf ( n706 , n10497 );
buf ( n707 , n10498 );
buf ( n708 , n10499 );
buf ( n709 , n10500 );
buf ( n710 , n10530 );
buf ( n711 , n10531 );
buf ( n712 , n10532 );
buf ( n713 , n10533 );
buf ( n714 , n10563 );
buf ( n715 , n10564 );
buf ( n716 , n10565 );
buf ( n717 , n10566 );
buf ( n718 , n10596 );
buf ( n719 , n10597 );
buf ( n720 , n10598 );
buf ( n721 , n10599 );
buf ( n722 , n10629 );
buf ( n723 , n10630 );
buf ( n724 , n10631 );
buf ( n725 , n10632 );
buf ( n726 , n10662 );
buf ( n727 , n10663 );
buf ( n728 , n10664 );
buf ( n729 , n10665 );
buf ( n730 , n10695 );
buf ( n731 , n10696 );
buf ( n732 , n10697 );
buf ( n733 , n10698 );
buf ( n734 , n10728 );
buf ( n735 , n10729 );
buf ( n736 , n10730 );
buf ( n737 , n10731 );
buf ( n738 , n10761 );
buf ( n739 , n10762 );
buf ( n740 , n10763 );
buf ( n741 , n10764 );
buf ( n742 , n10794 );
buf ( n743 , n10795 );
buf ( n744 , n10796 );
buf ( n745 , n10797 );
buf ( n746 , n10827 );
buf ( n747 , n10828 );
buf ( n748 , n10829 );
buf ( n749 , n10830 );
buf ( n750 , n10860 );
buf ( n751 , n10861 );
buf ( n752 , n10862 );
buf ( n753 , n10863 );
buf ( n754 , n10893 );
buf ( n755 , n10894 );
buf ( n756 , n10895 );
buf ( n757 , n10896 );
buf ( n758 , n10926 );
buf ( n759 , n10927 );
buf ( n760 , n10928 );
buf ( n761 , n10929 );
buf ( n762 , n10959 );
buf ( n763 , n10960 );
buf ( n764 , n10961 );
buf ( n765 , n10962 );
buf ( n766 , n10992 );
buf ( n767 , n10993 );
buf ( n768 , n10994 );
buf ( n769 , n10995 );
buf ( n770 , n11025 );
buf ( n771 , n11026 );
buf ( n772 , n11027 );
buf ( n773 , n11028 );
buf ( n774 , n11058 );
buf ( n775 , n11059 );
buf ( n776 , n11060 );
buf ( n777 , n11061 );
buf ( n778 , n11091 );
buf ( n779 , n11092 );
buf ( n780 , n11093 );
buf ( n781 , n11094 );
buf ( n782 , n11124 );
buf ( n783 , n11125 );
buf ( n784 , n11126 );
buf ( n785 , n11127 );
buf ( n786 , n11157 );
buf ( n787 , n11158 );
buf ( n788 , n11159 );
buf ( n789 , n11160 );
buf ( n790 , n11190 );
buf ( n791 , n11191 );
buf ( n792 , n11192 );
buf ( n793 , n11193 );
buf ( n794 , n11223 );
buf ( n795 , n11224 );
buf ( n796 , n11225 );
buf ( n797 , n11226 );
buf ( n798 , n11256 );
buf ( n799 , n11257 );
buf ( n800 , n11258 );
buf ( n801 , n11259 );
buf ( n802 , n11285 );
buf ( DFF_B_reg_S , n11286 );
buf ( DFF_B_reg_R , n11287 );
buf ( DFF_B_reg_CK , n11288 );
buf ( DFF_B_reg_D , n11902 );
buf ( n803 , n11903 );
buf ( n804 , n11904 );
buf ( n805 , n11905 );
buf ( n806 , n11938 );
buf ( n807 , n11939 );
buf ( n808 , n11940 );
buf ( n809 , n11941 );
buf ( n810 , n11972 );
buf ( n811 , n11973 );
buf ( n812 , n11974 );
buf ( n813 , n11975 );
buf ( n814 , n12006 );
buf ( n815 , n12007 );
buf ( n816 , n12008 );
buf ( n817 , n12009 );
buf ( n818 , n12040 );
buf ( n819 , n12041 );
buf ( n820 , n12042 );
buf ( n821 , n12043 );
buf ( n822 , n12074 );
buf ( n823 , n12075 );
buf ( n824 , n12076 );
buf ( n825 , n12077 );
buf ( n826 , n12108 );
buf ( n827 , n12109 );
buf ( n828 , n12110 );
buf ( n829 , n12111 );
buf ( n830 , n12142 );
buf ( n831 , n12143 );
buf ( n832 , n12144 );
buf ( n833 , n12145 );
buf ( n834 , n12176 );
buf ( n835 , n12177 );
buf ( n836 , n12178 );
buf ( n837 , n12179 );
buf ( n838 , n12210 );
buf ( n839 , n12211 );
buf ( n840 , n12212 );
buf ( n841 , n12213 );
buf ( n842 , n12244 );
buf ( n843 , n12245 );
buf ( n844 , n12246 );
buf ( n845 , n12247 );
buf ( n846 , n12278 );
buf ( n847 , n12279 );
buf ( n848 , n12280 );
buf ( n849 , n12281 );
buf ( n850 , n12312 );
buf ( n851 , n12313 );
buf ( n852 , n12314 );
buf ( n853 , n12315 );
buf ( n854 , n12346 );
buf ( n855 , n12347 );
buf ( n856 , n12348 );
buf ( n857 , n12349 );
buf ( n858 , n12380 );
buf ( n859 , n12381 );
buf ( n860 , n12382 );
buf ( n861 , n12383 );
buf ( n862 , n12414 );
buf ( n863 , n12415 );
buf ( n864 , n12416 );
buf ( n865 , n12417 );
buf ( n866 , n12448 );
buf ( n867 , n12449 );
buf ( n868 , n12450 );
buf ( n869 , n12451 );
buf ( n870 , n12482 );
buf ( n871 , n12483 );
buf ( n872 , n12484 );
buf ( n873 , n12485 );
buf ( n874 , n12516 );
buf ( n875 , n12517 );
buf ( n876 , n12518 );
buf ( n877 , n12519 );
buf ( n878 , n12550 );
buf ( n879 , n12551 );
buf ( n880 , n12552 );
buf ( n881 , n12553 );
buf ( n882 , n12584 );
buf ( n883 , n12585 );
buf ( n884 , n12586 );
buf ( n885 , n12587 );
buf ( n886 , n12618 );
buf ( n887 , n12619 );
buf ( n888 , n12620 );
buf ( n889 , n12621 );
buf ( n890 , n12652 );
buf ( n891 , n12653 );
buf ( n892 , n12654 );
buf ( n893 , n12655 );
buf ( n894 , n12686 );
buf ( n895 , n12687 );
buf ( n896 , n12688 );
buf ( n897 , n12689 );
buf ( n898 , n12720 );
buf ( n899 , n12721 );
buf ( n900 , n12722 );
buf ( n901 , n12723 );
buf ( n902 , n12754 );
buf ( n903 , n12755 );
buf ( n904 , n12756 );
buf ( n905 , n12757 );
buf ( n906 , n12788 );
buf ( n907 , n12789 );
buf ( n908 , n12790 );
buf ( n909 , n12791 );
buf ( n910 , n12822 );
buf ( n911 , n12823 );
buf ( n912 , n12824 );
buf ( n913 , n12825 );
buf ( n914 , n12856 );
buf ( n915 , n12857 );
buf ( n916 , n12858 );
buf ( n917 , n12859 );
buf ( n918 , n12890 );
buf ( n919 , n12891 );
buf ( n920 , n12892 );
buf ( n921 , n12893 );
buf ( n922 , n12924 );
buf ( n923 , n12925 );
buf ( n924 , n12926 );
buf ( n925 , n12927 );
buf ( n926 , n12957 );
buf ( n927 , n12958 );
buf ( n928 , n12959 );
buf ( n929 , n12960 );
buf ( n930 , n12986 );
buf ( n931 , n12987 );
buf ( n932 , n12988 );
buf ( n933 , n12989 );
buf ( n934 , n13678 );
buf ( n935 , n13679 );
buf ( n936 , n13680 );
buf ( n937 , n13681 );
buf ( n938 , n13719 );
buf ( n939 , n13720 );
buf ( n940 , n13721 );
buf ( n941 , n13722 );
buf ( n942 , n14170 );
buf ( n943 , n14171 );
buf ( n944 , n14172 );
buf ( n945 , n14173 );
buf ( n946 , n14211 );
buf ( n947 , n14212 );
buf ( n948 , n14213 );
buf ( n949 , n14214 );
buf ( n950 , n14253 );
buf ( n951 , n14254 );
buf ( n952 , n14255 );
buf ( n953 , n14256 );
buf ( n954 , n14294 );
buf ( n955 , n14295 );
buf ( n956 , n14296 );
buf ( n957 , n14297 );
buf ( n958 , n14335 );
buf ( n959 , n14336 );
buf ( n960 , n14337 );
buf ( n961 , n14338 );
buf ( n962 , n14376 );
buf ( n963 , n14377 );
buf ( n964 , n14378 );
buf ( n965 , n14379 );
buf ( n966 , n14417 );
buf ( n967 , n14418 );
buf ( n968 , n14419 );
buf ( n969 , n14420 );
buf ( n970 , n14458 );
buf ( n971 , n14459 );
buf ( n972 , n14460 );
buf ( n973 , n14461 );
buf ( n974 , n14499 );
buf ( n975 , n14500 );
buf ( n976 , n14501 );
buf ( n977 , n14502 );
buf ( n978 , n14540 );
buf ( n979 , n14541 );
buf ( n980 , n14542 );
buf ( n981 , n14543 );
buf ( n982 , n14581 );
buf ( n983 , n14582 );
buf ( n984 , n14583 );
buf ( n985 , n14584 );
buf ( n986 , n14622 );
buf ( n987 , n14623 );
buf ( n988 , n14624 );
buf ( n989 , n14625 );
buf ( n990 , n14663 );
buf ( n991 , n14664 );
buf ( n992 , n14665 );
buf ( n993 , n14666 );
buf ( n994 , n14704 );
buf ( n995 , n14705 );
buf ( n996 , n14706 );
buf ( n997 , n14707 );
buf ( n998 , n14745 );
buf ( n999 , n14746 );
buf ( n1000 , n14747 );
buf ( n1001 , n14748 );
buf ( n1002 , n14786 );
buf ( n1003 , n14787 );
buf ( n1004 , n14788 );
buf ( n1005 , n14789 );
buf ( n1006 , n14827 );
buf ( n1007 , n14828 );
buf ( n1008 , n14829 );
buf ( n1009 , n14830 );
buf ( n1010 , n14868 );
buf ( n1011 , n14869 );
buf ( n1012 , n14870 );
buf ( n1013 , n14871 );
buf ( n1014 , n14881 );
buf ( n1015 , n14882 );
buf ( n1016 , n14883 );
buf ( n1017 , n14884 );
buf ( n1018 , n14892 );
buf ( n1019 , n14893 );
buf ( n1020 , n14894 );
buf ( n1021 , n14895 );
buf ( n1022 , n14903 );
buf ( n1023 , n14904 );
buf ( n1024 , n14905 );
buf ( n1025 , n14906 );
buf ( n1026 , n14914 );
buf ( n1027 , n14915 );
buf ( n1028 , n14916 );
buf ( n1029 , n14917 );
buf ( n1030 , n14925 );
buf ( n1031 , n14926 );
buf ( n1032 , n14927 );
buf ( n1033 , n14928 );
buf ( n1034 , n14936 );
buf ( n1035 , n14937 );
buf ( n1036 , n14938 );
buf ( n1037 , n14939 );
buf ( n1038 , n14947 );
buf ( n1039 , n14948 );
buf ( n1040 , n14949 );
buf ( n1041 , n14950 );
buf ( n1042 , n14958 );
buf ( n1043 , n14959 );
buf ( n1044 , n14960 );
buf ( n1045 , n14961 );
buf ( n1046 , n14969 );
buf ( n1047 , n14970 );
buf ( n1048 , n14971 );
buf ( n1049 , n14972 );
buf ( n1050 , n14980 );
buf ( n1051 , n14981 );
buf ( n1052 , n14982 );
buf ( n1053 , n14983 );
buf ( n1054 , n14991 );
buf ( n1055 , n14992 );
buf ( n1056 , n14993 );
buf ( n1057 , n14994 );
buf ( n1058 , n15002 );
buf ( n1059 , n15003 );
buf ( n1060 , n15004 );
buf ( n1061 , n15005 );
buf ( n1062 , n15013 );
buf ( n1063 , n15014 );
buf ( n1064 , n15015 );
buf ( n1065 , n15016 );
buf ( n1066 , n15024 );
buf ( n1067 , n15025 );
buf ( n1068 , n15026 );
buf ( n1069 , n15027 );
buf ( n1070 , n15035 );
buf ( n1071 , n15036 );
buf ( n1072 , n15037 );
buf ( n1073 , n15038 );
buf ( n1074 , n15046 );
buf ( n1075 , n15047 );
buf ( n1076 , n15048 );
buf ( n1077 , n15049 );
buf ( n1078 , n15057 );
buf ( n1079 , n15058 );
buf ( n1080 , n15059 );
buf ( n1081 , n15060 );
buf ( n1082 , n15068 );
buf ( n1083 , n15069 );
buf ( n1084 , n15070 );
buf ( n1085 , n15071 );
buf ( n1086 , n15079 );
buf ( n1087 , n15080 );
buf ( n1088 , n15081 );
buf ( n1089 , n15082 );
buf ( n1090 , n15090 );
buf ( n1091 , n15091 );
buf ( n1092 , n15092 );
buf ( n1093 , n15093 );
buf ( n1094 , n15101 );
buf ( n1095 , n15102 );
buf ( n1096 , n15103 );
buf ( n1097 , n15104 );
buf ( n1098 , n15112 );
buf ( n1099 , n15113 );
buf ( n1100 , n15114 );
buf ( n1101 , n15115 );
buf ( n1102 , n15123 );
buf ( n1103 , n15124 );
buf ( n1104 , n15125 );
buf ( n1105 , n15126 );
buf ( n1106 , n15134 );
buf ( n1107 , n15135 );
buf ( n1108 , n15136 );
buf ( n1109 , n15137 );
buf ( n1110 , n15145 );
buf ( n1111 , n15146 );
buf ( n1112 , n15147 );
buf ( n1113 , n15148 );
buf ( n1114 , n15156 );
buf ( n1115 , n15157 );
buf ( n1116 , n15158 );
buf ( n1117 , n15159 );
buf ( n1118 , n15167 );
buf ( n1119 , n15168 );
buf ( n1120 , n15169 );
buf ( n1121 , n15170 );
buf ( n1122 , n15178 );
buf ( n1123 , n15179 );
buf ( n1124 , n15180 );
buf ( n1125 , n15181 );
buf ( n1126 , n15189 );
buf ( n1127 , n15190 );
buf ( n1128 , n15191 );
buf ( n1129 , n15192 );
buf ( n1130 , n15200 );
buf ( n1131 , n15201 );
buf ( n1132 , n15202 );
buf ( n1133 , n15203 );
buf ( n1134 , n15211 );
buf ( n1135 , n15212 );
buf ( n1136 , n15213 );
buf ( n1137 , n15214 );
buf ( n1138 , n15222 );
buf ( DFF_rd_reg_S , n15223 );
buf ( DFF_rd_reg_R , n15224 );
buf ( DFF_rd_reg_CK , n15225 );
buf ( DFF_rd_reg_D , n15235 );
buf ( DFF_wr_reg_S , n15236 );
buf ( DFF_wr_reg_R , n15237 );
buf ( DFF_wr_reg_CK , n15238 );
buf ( DFF_wr_reg_D , n15242 );
buf ( n2280 , PI_clock);
buf ( n2281 , PI_reset);
buf ( n2282 , n0 );
buf ( n2283 , n1 );
buf ( n2284 , n2 );
buf ( n2285 , n3 );
buf ( n2286 , n4 );
buf ( n2287 , n5 );
buf ( n2288 , n6 );
buf ( n2289 , n7 );
buf ( n2290 , n8 );
buf ( n2291 , n9 );
buf ( n2292 , n10 );
buf ( n2293 , n11 );
buf ( n2294 , n12 );
buf ( n2295 , n13 );
buf ( n2296 , n14 );
buf ( n2297 , n15 );
buf ( n2298 , n16 );
buf ( n2299 , n17 );
buf ( n2300 , n18 );
buf ( n2301 , n19 );
buf ( n2302 , n20 );
buf ( n2303 , n21 );
buf ( n2304 , n22 );
buf ( n2305 , n23 );
buf ( n2306 , n24 );
buf ( n2307 , n25 );
buf ( n2308 , n26 );
buf ( n2309 , n27 );
buf ( n2310 , n28 );
buf ( n2311 , n29 );
buf ( n2312 , n30 );
buf ( n2313 , n31 );
buf ( n2314 , n210 );
buf ( n2315 , n2314 );
buf ( n2316 , n209 );
buf ( n2317 , n2316 );
buf ( n2318 , n208 );
buf ( n2319 , n2318 );
buf ( n2320 , n207 );
buf ( n2321 , n2320 );
buf ( n2322 , n206 );
buf ( n2323 , n2322 );
buf ( n2324 , n205 );
buf ( n2325 , n2324 );
buf ( n2326 , n204 );
buf ( n2327 , n2326 );
buf ( n2328 , n203 );
buf ( n2329 , n2328 );
buf ( n2330 , n202 );
buf ( n2331 , n2330 );
buf ( n2332 , n201 );
buf ( n2333 , n2332 );
buf ( n2334 , n200 );
buf ( n2335 , n2334 );
buf ( n2336 , n199 );
buf ( n2337 , n2336 );
buf ( n2338 , n198 );
buf ( n2339 , n2338 );
buf ( n2340 , n197 );
buf ( n2341 , n2340 );
buf ( n2342 , n196 );
buf ( n2343 , n2342 );
buf ( n2344 , n195 );
buf ( n2345 , n2344 );
buf ( n2346 , n194 );
buf ( n2347 , n2346 );
buf ( n2348 , n193 );
buf ( n2349 , n2348 );
buf ( n2350 , n192 );
buf ( n2351 , n2350 );
buf ( n2352 , n191 );
buf ( n2353 , n2352 );
buf ( n2354 , n242 );
buf ( n2355 , n2354 );
buf ( n2356 , n241 );
buf ( n2357 , n2356 );
buf ( n2358 , n240 );
buf ( n2359 , n2358 );
buf ( n2360 , n239 );
buf ( n2361 , n2360 );
buf ( n2362 , n238 );
buf ( n2363 , n2362 );
buf ( n2364 , n237 );
buf ( n2365 , n2364 );
buf ( n2366 , n236 );
buf ( n2367 , n2366 );
buf ( n2368 , n235 );
buf ( n2369 , n2368 );
buf ( n2370 , n234 );
buf ( n2371 , n2370 );
buf ( n2372 , n233 );
buf ( n2373 , n2372 );
buf ( n2374 , n232 );
buf ( n2375 , n2374 );
buf ( n2376 , n231 );
buf ( n2377 , n2376 );
buf ( n2378 , n230 );
buf ( n2379 , n2378 );
buf ( n2380 , n229 );
buf ( n2381 , n2380 );
buf ( n2382 , n228 );
buf ( n2383 , n2382 );
buf ( n2384 , n227 );
buf ( n2385 , n2384 );
buf ( n2386 , n226 );
buf ( n2387 , n2386 );
buf ( n2388 , n225 );
buf ( n2389 , n2388 );
buf ( n2390 , n224 );
buf ( n2391 , n2390 );
buf ( n2392 , n223 );
buf ( n2393 , n2392 );
buf ( n2394 , n222 );
buf ( n2395 , n2394 );
buf ( n2396 , n221 );
buf ( n2397 , n2396 );
buf ( n2398 , n220 );
buf ( n2399 , n2398 );
buf ( n2400 , n219 );
buf ( n2401 , n2400 );
buf ( n2402 , n218 );
buf ( n2403 , n2402 );
buf ( n2404 , n217 );
buf ( n2405 , n2404 );
buf ( n2406 , n216 );
buf ( n2407 , n2406 );
buf ( n2408 , n215 );
buf ( n2409 , n2408 );
buf ( n2410 , n214 );
buf ( n2411 , n2410 );
buf ( n2412 , n213 );
buf ( n2413 , n2412 );
buf ( n2414 , n212 );
buf ( n2415 , n2414 );
buf ( n2416 , n211 );
buf ( n2417 , n2416 );
buf ( n2418 , DFF_rd_reg_Q);
buf ( n2419 , n2418 );
buf ( n2420 , DFF_wr_reg_Q);
buf ( n2421 , n2420 );
buf ( n2422 , DFF_state_reg_Q);
not ( n2423 , n2282 );
and ( n2424 , n2282 , n2423 );
buf ( n2425 , n2424 );
buf ( n2426 , n2281 );
buf ( n2427 , n2280 );
not ( n2428 , n2422 );
buf ( n2429 , n2428 );
buf ( n2430 , n32 );
buf ( n2431 , n2424 );
buf ( n2432 , n2281 );
buf ( n2433 , n2280 );
and ( n2434 , n2430 , n2422 );
and ( n2435 , n2313 , n2428 );
or ( n2436 , n2434 , n2435 );
buf ( n2437 , n2436 );
buf ( n2438 , n33 );
buf ( n2439 , n2424 );
buf ( n2440 , n2281 );
buf ( n2441 , n2280 );
buf ( n2442 , n63 );
not ( n2443 , n2442 );
and ( n2444 , n2443 , n2438 );
not ( n2445 , n2438 );
not ( n2446 , n2430 );
xor ( n2447 , n2445 , n2446 );
and ( n2448 , n2447 , n2442 );
or ( n2449 , n2444 , n2448 );
and ( n2450 , n2449 , n2422 );
and ( n2451 , n2312 , n2428 );
or ( n2452 , n2450 , n2451 );
buf ( n2453 , n2452 );
buf ( n2454 , n34 );
buf ( n2455 , n2424 );
buf ( n2456 , n2281 );
buf ( n2457 , n2280 );
not ( n2458 , n2442 );
and ( n2459 , n2458 , n2454 );
not ( n2460 , n2454 );
and ( n2461 , n2445 , n2446 );
xor ( n2462 , n2460 , n2461 );
and ( n2463 , n2462 , n2442 );
or ( n2464 , n2459 , n2463 );
and ( n2465 , n2464 , n2422 );
and ( n2466 , n2311 , n2428 );
or ( n2467 , n2465 , n2466 );
buf ( n2468 , n2467 );
buf ( n2469 , n35 );
buf ( n2470 , n2424 );
buf ( n2471 , n2281 );
buf ( n2472 , n2280 );
not ( n2473 , n2442 );
and ( n2474 , n2473 , n2469 );
not ( n2475 , n2469 );
and ( n2476 , n2460 , n2461 );
xor ( n2477 , n2475 , n2476 );
and ( n2478 , n2477 , n2442 );
or ( n2479 , n2474 , n2478 );
and ( n2480 , n2479 , n2422 );
and ( n2481 , n2310 , n2428 );
or ( n2482 , n2480 , n2481 );
buf ( n2483 , n2482 );
buf ( n2484 , n36 );
buf ( n2485 , n2424 );
buf ( n2486 , n2281 );
buf ( n2487 , n2280 );
not ( n2488 , n2442 );
and ( n2489 , n2488 , n2484 );
not ( n2490 , n2484 );
and ( n2491 , n2475 , n2476 );
xor ( n2492 , n2490 , n2491 );
and ( n2493 , n2492 , n2442 );
or ( n2494 , n2489 , n2493 );
and ( n2495 , n2494 , n2422 );
and ( n2496 , n2309 , n2428 );
or ( n2497 , n2495 , n2496 );
buf ( n2498 , n2497 );
buf ( n2499 , n37 );
buf ( n2500 , n2424 );
buf ( n2501 , n2281 );
buf ( n2502 , n2280 );
not ( n2503 , n2442 );
and ( n2504 , n2503 , n2499 );
not ( n2505 , n2499 );
and ( n2506 , n2490 , n2491 );
xor ( n2507 , n2505 , n2506 );
and ( n2508 , n2507 , n2442 );
or ( n2509 , n2504 , n2508 );
and ( n2510 , n2509 , n2422 );
and ( n2511 , n2308 , n2428 );
or ( n2512 , n2510 , n2511 );
buf ( n2513 , n2512 );
buf ( n2514 , n38 );
buf ( n2515 , n2424 );
buf ( n2516 , n2281 );
buf ( n2517 , n2280 );
not ( n2518 , n2442 );
and ( n2519 , n2518 , n2514 );
not ( n2520 , n2514 );
and ( n2521 , n2505 , n2506 );
xor ( n2522 , n2520 , n2521 );
and ( n2523 , n2522 , n2442 );
or ( n2524 , n2519 , n2523 );
and ( n2525 , n2524 , n2422 );
and ( n2526 , n2307 , n2428 );
or ( n2527 , n2525 , n2526 );
buf ( n2528 , n2527 );
buf ( n2529 , n39 );
buf ( n2530 , n2424 );
buf ( n2531 , n2281 );
buf ( n2532 , n2280 );
not ( n2533 , n2442 );
and ( n2534 , n2533 , n2529 );
not ( n2535 , n2529 );
and ( n2536 , n2520 , n2521 );
xor ( n2537 , n2535 , n2536 );
and ( n2538 , n2537 , n2442 );
or ( n2539 , n2534 , n2538 );
and ( n2540 , n2539 , n2422 );
and ( n2541 , n2306 , n2428 );
or ( n2542 , n2540 , n2541 );
buf ( n2543 , n2542 );
buf ( n2544 , n40 );
buf ( n2545 , n2424 );
buf ( n2546 , n2281 );
buf ( n2547 , n2280 );
not ( n2548 , n2442 );
and ( n2549 , n2548 , n2544 );
not ( n2550 , n2544 );
and ( n2551 , n2535 , n2536 );
xor ( n2552 , n2550 , n2551 );
and ( n2553 , n2552 , n2442 );
or ( n2554 , n2549 , n2553 );
and ( n2555 , n2554 , n2422 );
and ( n2556 , n2305 , n2428 );
or ( n2557 , n2555 , n2556 );
buf ( n2558 , n2557 );
buf ( n2559 , n41 );
buf ( n2560 , n2424 );
buf ( n2561 , n2281 );
buf ( n2562 , n2280 );
not ( n2563 , n2442 );
and ( n2564 , n2563 , n2559 );
not ( n2565 , n2559 );
and ( n2566 , n2550 , n2551 );
xor ( n2567 , n2565 , n2566 );
and ( n2568 , n2567 , n2442 );
or ( n2569 , n2564 , n2568 );
and ( n2570 , n2569 , n2422 );
and ( n2571 , n2304 , n2428 );
or ( n2572 , n2570 , n2571 );
buf ( n2573 , n2572 );
buf ( n2574 , n42 );
buf ( n2575 , n2424 );
buf ( n2576 , n2281 );
buf ( n2577 , n2280 );
not ( n2578 , n2442 );
and ( n2579 , n2578 , n2574 );
not ( n2580 , n2574 );
and ( n2581 , n2565 , n2566 );
xor ( n2582 , n2580 , n2581 );
and ( n2583 , n2582 , n2442 );
or ( n2584 , n2579 , n2583 );
and ( n2585 , n2584 , n2422 );
and ( n2586 , n2303 , n2428 );
or ( n2587 , n2585 , n2586 );
buf ( n2588 , n2587 );
buf ( n2589 , n43 );
buf ( n2590 , n2424 );
buf ( n2591 , n2281 );
buf ( n2592 , n2280 );
not ( n2593 , n2442 );
and ( n2594 , n2593 , n2589 );
not ( n2595 , n2589 );
and ( n2596 , n2580 , n2581 );
xor ( n2597 , n2595 , n2596 );
and ( n2598 , n2597 , n2442 );
or ( n2599 , n2594 , n2598 );
and ( n2600 , n2599 , n2422 );
and ( n2601 , n2302 , n2428 );
or ( n2602 , n2600 , n2601 );
buf ( n2603 , n2602 );
buf ( n2604 , n44 );
buf ( n2605 , n2424 );
buf ( n2606 , n2281 );
buf ( n2607 , n2280 );
not ( n2608 , n2442 );
and ( n2609 , n2608 , n2604 );
not ( n2610 , n2604 );
and ( n2611 , n2595 , n2596 );
xor ( n2612 , n2610 , n2611 );
and ( n2613 , n2612 , n2442 );
or ( n2614 , n2609 , n2613 );
and ( n2615 , n2614 , n2422 );
and ( n2616 , n2301 , n2428 );
or ( n2617 , n2615 , n2616 );
buf ( n2618 , n2617 );
buf ( n2619 , n45 );
buf ( n2620 , n2424 );
buf ( n2621 , n2281 );
buf ( n2622 , n2280 );
not ( n2623 , n2442 );
and ( n2624 , n2623 , n2619 );
not ( n2625 , n2619 );
and ( n2626 , n2610 , n2611 );
xor ( n2627 , n2625 , n2626 );
and ( n2628 , n2627 , n2442 );
or ( n2629 , n2624 , n2628 );
and ( n2630 , n2629 , n2422 );
and ( n2631 , n2300 , n2428 );
or ( n2632 , n2630 , n2631 );
buf ( n2633 , n2632 );
buf ( n2634 , n46 );
buf ( n2635 , n2424 );
buf ( n2636 , n2281 );
buf ( n2637 , n2280 );
not ( n2638 , n2442 );
and ( n2639 , n2638 , n2634 );
not ( n2640 , n2634 );
and ( n2641 , n2625 , n2626 );
xor ( n2642 , n2640 , n2641 );
and ( n2643 , n2642 , n2442 );
or ( n2644 , n2639 , n2643 );
and ( n2645 , n2644 , n2422 );
and ( n2646 , n2299 , n2428 );
or ( n2647 , n2645 , n2646 );
buf ( n2648 , n2647 );
buf ( n2649 , n47 );
buf ( n2650 , n2424 );
buf ( n2651 , n2281 );
buf ( n2652 , n2280 );
not ( n2653 , n2442 );
and ( n2654 , n2653 , n2649 );
not ( n2655 , n2649 );
and ( n2656 , n2640 , n2641 );
xor ( n2657 , n2655 , n2656 );
and ( n2658 , n2657 , n2442 );
or ( n2659 , n2654 , n2658 );
and ( n2660 , n2659 , n2422 );
and ( n2661 , n2298 , n2428 );
or ( n2662 , n2660 , n2661 );
buf ( n2663 , n2662 );
buf ( n2664 , n48 );
buf ( n2665 , n2424 );
buf ( n2666 , n2281 );
buf ( n2667 , n2280 );
not ( n2668 , n2442 );
and ( n2669 , n2668 , n2664 );
not ( n2670 , n2664 );
and ( n2671 , n2655 , n2656 );
xor ( n2672 , n2670 , n2671 );
and ( n2673 , n2672 , n2442 );
or ( n2674 , n2669 , n2673 );
and ( n2675 , n2674 , n2422 );
and ( n2676 , n2297 , n2428 );
or ( n2677 , n2675 , n2676 );
buf ( n2678 , n2677 );
buf ( n2679 , n49 );
buf ( n2680 , n2424 );
buf ( n2681 , n2281 );
buf ( n2682 , n2280 );
not ( n2683 , n2442 );
and ( n2684 , n2683 , n2679 );
not ( n2685 , n2679 );
and ( n2686 , n2670 , n2671 );
xor ( n2687 , n2685 , n2686 );
and ( n2688 , n2687 , n2442 );
or ( n2689 , n2684 , n2688 );
and ( n2690 , n2689 , n2422 );
and ( n2691 , n2296 , n2428 );
or ( n2692 , n2690 , n2691 );
buf ( n2693 , n2692 );
buf ( n2694 , n50 );
buf ( n2695 , n2424 );
buf ( n2696 , n2281 );
buf ( n2697 , n2280 );
not ( n2698 , n2442 );
and ( n2699 , n2698 , n2694 );
not ( n2700 , n2694 );
and ( n2701 , n2685 , n2686 );
xor ( n2702 , n2700 , n2701 );
and ( n2703 , n2702 , n2442 );
or ( n2704 , n2699 , n2703 );
and ( n2705 , n2704 , n2422 );
and ( n2706 , n2295 , n2428 );
or ( n2707 , n2705 , n2706 );
buf ( n2708 , n2707 );
buf ( n2709 , n51 );
buf ( n2710 , n2424 );
buf ( n2711 , n2281 );
buf ( n2712 , n2280 );
not ( n2713 , n2442 );
and ( n2714 , n2713 , n2709 );
not ( n2715 , n2709 );
and ( n2716 , n2700 , n2701 );
xor ( n2717 , n2715 , n2716 );
and ( n2718 , n2717 , n2442 );
or ( n2719 , n2714 , n2718 );
and ( n2720 , n2719 , n2422 );
and ( n2721 , n2294 , n2428 );
or ( n2722 , n2720 , n2721 );
buf ( n2723 , n2722 );
buf ( n2724 , n52 );
buf ( n2725 , n2424 );
buf ( n2726 , n2281 );
buf ( n2727 , n2280 );
not ( n2728 , n2442 );
and ( n2729 , n2728 , n2724 );
not ( n2730 , n2724 );
and ( n2731 , n2715 , n2716 );
xor ( n2732 , n2730 , n2731 );
and ( n2733 , n2732 , n2442 );
or ( n2734 , n2729 , n2733 );
and ( n2735 , n2734 , n2422 );
and ( n2736 , n2293 , n2428 );
or ( n2737 , n2735 , n2736 );
buf ( n2738 , n2737 );
buf ( n2739 , n53 );
buf ( n2740 , n2424 );
buf ( n2741 , n2281 );
buf ( n2742 , n2280 );
not ( n2743 , n2442 );
and ( n2744 , n2743 , n2739 );
not ( n2745 , n2739 );
and ( n2746 , n2730 , n2731 );
xor ( n2747 , n2745 , n2746 );
and ( n2748 , n2747 , n2442 );
or ( n2749 , n2744 , n2748 );
and ( n2750 , n2749 , n2422 );
and ( n2751 , n2292 , n2428 );
or ( n2752 , n2750 , n2751 );
buf ( n2753 , n2752 );
buf ( n2754 , n54 );
buf ( n2755 , n2424 );
buf ( n2756 , n2281 );
buf ( n2757 , n2280 );
not ( n2758 , n2442 );
and ( n2759 , n2758 , n2754 );
not ( n2760 , n2754 );
and ( n2761 , n2745 , n2746 );
xor ( n2762 , n2760 , n2761 );
and ( n2763 , n2762 , n2442 );
or ( n2764 , n2759 , n2763 );
and ( n2765 , n2764 , n2422 );
and ( n2766 , n2291 , n2428 );
or ( n2767 , n2765 , n2766 );
buf ( n2768 , n2767 );
buf ( n2769 , n55 );
buf ( n2770 , n2424 );
buf ( n2771 , n2281 );
buf ( n2772 , n2280 );
not ( n2773 , n2442 );
and ( n2774 , n2773 , n2769 );
not ( n2775 , n2769 );
and ( n2776 , n2760 , n2761 );
xor ( n2777 , n2775 , n2776 );
and ( n2778 , n2777 , n2442 );
or ( n2779 , n2774 , n2778 );
and ( n2780 , n2779 , n2422 );
and ( n2781 , n2290 , n2428 );
or ( n2782 , n2780 , n2781 );
buf ( n2783 , n2782 );
buf ( n2784 , n56 );
buf ( n2785 , n2424 );
buf ( n2786 , n2281 );
buf ( n2787 , n2280 );
not ( n2788 , n2442 );
and ( n2789 , n2788 , n2784 );
not ( n2790 , n2784 );
and ( n2791 , n2775 , n2776 );
xor ( n2792 , n2790 , n2791 );
and ( n2793 , n2792 , n2442 );
or ( n2794 , n2789 , n2793 );
and ( n2795 , n2794 , n2422 );
and ( n2796 , n2289 , n2428 );
or ( n2797 , n2795 , n2796 );
buf ( n2798 , n2797 );
buf ( n2799 , n57 );
buf ( n2800 , n2424 );
buf ( n2801 , n2281 );
buf ( n2802 , n2280 );
not ( n2803 , n2442 );
and ( n2804 , n2803 , n2799 );
not ( n2805 , n2799 );
and ( n2806 , n2790 , n2791 );
xor ( n2807 , n2805 , n2806 );
and ( n2808 , n2807 , n2442 );
or ( n2809 , n2804 , n2808 );
and ( n2810 , n2809 , n2422 );
and ( n2811 , n2288 , n2428 );
or ( n2812 , n2810 , n2811 );
buf ( n2813 , n2812 );
buf ( n2814 , n58 );
buf ( n2815 , n2424 );
buf ( n2816 , n2281 );
buf ( n2817 , n2280 );
not ( n2818 , n2442 );
and ( n2819 , n2818 , n2814 );
not ( n2820 , n2814 );
and ( n2821 , n2805 , n2806 );
xor ( n2822 , n2820 , n2821 );
and ( n2823 , n2822 , n2442 );
or ( n2824 , n2819 , n2823 );
and ( n2825 , n2824 , n2422 );
and ( n2826 , n2287 , n2428 );
or ( n2827 , n2825 , n2826 );
buf ( n2828 , n2827 );
buf ( n2829 , n59 );
buf ( n2830 , n2424 );
buf ( n2831 , n2281 );
buf ( n2832 , n2280 );
not ( n2833 , n2442 );
and ( n2834 , n2833 , n2829 );
not ( n2835 , n2829 );
and ( n2836 , n2820 , n2821 );
xor ( n2837 , n2835 , n2836 );
and ( n2838 , n2837 , n2442 );
or ( n2839 , n2834 , n2838 );
and ( n2840 , n2839 , n2422 );
and ( n2841 , n2286 , n2428 );
or ( n2842 , n2840 , n2841 );
buf ( n2843 , n2842 );
buf ( n2844 , n60 );
buf ( n2845 , n2424 );
buf ( n2846 , n2281 );
buf ( n2847 , n2280 );
not ( n2848 , n2442 );
and ( n2849 , n2848 , n2844 );
not ( n2850 , n2844 );
and ( n2851 , n2835 , n2836 );
xor ( n2852 , n2850 , n2851 );
and ( n2853 , n2852 , n2442 );
or ( n2854 , n2849 , n2853 );
and ( n2855 , n2854 , n2422 );
and ( n2856 , n2285 , n2428 );
or ( n2857 , n2855 , n2856 );
buf ( n2858 , n2857 );
buf ( n2859 , n61 );
buf ( n2860 , n2424 );
buf ( n2861 , n2281 );
buf ( n2862 , n2280 );
not ( n2863 , n2442 );
and ( n2864 , n2863 , n2859 );
not ( n2865 , n2859 );
and ( n2866 , n2850 , n2851 );
xor ( n2867 , n2865 , n2866 );
and ( n2868 , n2867 , n2442 );
or ( n2869 , n2864 , n2868 );
and ( n2870 , n2869 , n2422 );
and ( n2871 , n2284 , n2428 );
or ( n2872 , n2870 , n2871 );
buf ( n2873 , n2872 );
buf ( n2874 , n62 );
buf ( n2875 , n2424 );
buf ( n2876 , n2281 );
buf ( n2877 , n2280 );
not ( n2878 , n2442 );
and ( n2879 , n2878 , n2874 );
not ( n2880 , n2874 );
and ( n2881 , n2865 , n2866 );
xor ( n2882 , n2880 , n2881 );
and ( n2883 , n2882 , n2442 );
or ( n2884 , n2879 , n2883 );
and ( n2885 , n2884 , n2422 );
and ( n2886 , n2283 , n2428 );
or ( n2887 , n2885 , n2886 );
buf ( n2888 , n2887 );
buf ( n2889 , n2424 );
buf ( n2890 , n2281 );
buf ( n2891 , n2280 );
buf ( n2892 , n2442 );
not ( n2893 , n2892 );
and ( n2894 , n2893 , n2442 );
not ( n2895 , n2442 );
and ( n2896 , n2880 , n2881 );
xor ( n2897 , n2895 , n2896 );
and ( n2898 , n2897 , n2892 );
or ( n2899 , n2894 , n2898 );
and ( n2900 , n2899 , n2422 );
and ( n2901 , n2282 , n2428 );
or ( n2902 , n2900 , n2901 );
buf ( n2903 , n2902 );
buf ( n2904 , n64 );
buf ( n2905 , n2424 );
buf ( n2906 , n2281 );
buf ( n2907 , n2280 );
not ( n2908 , n2899 );
and ( n2909 , n2908 , n2779 );
not ( n2910 , n2779 );
not ( n2911 , n2764 );
not ( n2912 , n2749 );
not ( n2913 , n2734 );
not ( n2914 , n2719 );
not ( n2915 , n2704 );
not ( n2916 , n2689 );
not ( n2917 , n2674 );
not ( n2918 , n2659 );
not ( n2919 , n2644 );
not ( n2920 , n2629 );
not ( n2921 , n2614 );
not ( n2922 , n2599 );
not ( n2923 , n2584 );
not ( n2924 , n2569 );
not ( n2925 , n2554 );
not ( n2926 , n2539 );
not ( n2927 , n2524 );
not ( n2928 , n2509 );
not ( n2929 , n2494 );
not ( n2930 , n2479 );
not ( n2931 , n2464 );
not ( n2932 , n2449 );
not ( n2933 , n2430 );
and ( n2934 , n2932 , n2933 );
and ( n2935 , n2931 , n2934 );
and ( n2936 , n2930 , n2935 );
and ( n2937 , n2929 , n2936 );
and ( n2938 , n2928 , n2937 );
and ( n2939 , n2927 , n2938 );
and ( n2940 , n2926 , n2939 );
and ( n2941 , n2925 , n2940 );
and ( n2942 , n2924 , n2941 );
and ( n2943 , n2923 , n2942 );
and ( n2944 , n2922 , n2943 );
and ( n2945 , n2921 , n2944 );
and ( n2946 , n2920 , n2945 );
and ( n2947 , n2919 , n2946 );
and ( n2948 , n2918 , n2947 );
and ( n2949 , n2917 , n2948 );
and ( n2950 , n2916 , n2949 );
and ( n2951 , n2915 , n2950 );
and ( n2952 , n2914 , n2951 );
and ( n2953 , n2913 , n2952 );
and ( n2954 , n2912 , n2953 );
and ( n2955 , n2911 , n2954 );
xor ( n2956 , n2910 , n2955 );
and ( n2957 , n2956 , n2899 );
or ( n2958 , n2909 , n2957 );
not ( n2959 , n2958 );
not ( n2960 , n2959 );
not ( n2961 , n2960 );
not ( n2962 , n2961 );
buf ( n2963 , n2962 );
buf ( n2964 , n2963 );
not ( n2965 , n2899 );
and ( n2966 , n2965 , n2424 );
buf ( n2967 , n2899 );
not ( n2968 , n2967 );
and ( n2969 , n2968 , n2899 );
not ( n2970 , n2899 );
not ( n2971 , n2884 );
not ( n2972 , n2869 );
not ( n2973 , n2854 );
not ( n2974 , n2839 );
not ( n2975 , n2824 );
not ( n2976 , n2809 );
not ( n2977 , n2794 );
and ( n2978 , n2910 , n2955 );
and ( n2979 , n2977 , n2978 );
and ( n2980 , n2976 , n2979 );
and ( n2981 , n2975 , n2980 );
and ( n2982 , n2974 , n2981 );
and ( n2983 , n2973 , n2982 );
and ( n2984 , n2972 , n2983 );
and ( n2985 , n2971 , n2984 );
xor ( n2986 , n2970 , n2985 );
and ( n2987 , n2986 , n2967 );
or ( n2988 , n2969 , n2987 );
not ( n2989 , n2988 );
not ( n2990 , n2989 );
not ( n2991 , n2990 );
not ( n2992 , n2899 );
and ( n2993 , n2992 , n2884 );
xor ( n2994 , n2971 , n2984 );
and ( n2995 , n2994 , n2899 );
or ( n2996 , n2993 , n2995 );
not ( n2997 , n2996 );
not ( n2998 , n2997 );
not ( n2999 , n2998 );
not ( n3000 , n2899 );
and ( n3001 , n3000 , n2869 );
xor ( n3002 , n2972 , n2983 );
and ( n3003 , n3002 , n2899 );
or ( n3004 , n3001 , n3003 );
not ( n3005 , n3004 );
not ( n3006 , n3005 );
not ( n3007 , n3006 );
not ( n3008 , n2899 );
and ( n3009 , n3008 , n2854 );
xor ( n3010 , n2973 , n2982 );
and ( n3011 , n3010 , n2899 );
or ( n3012 , n3009 , n3011 );
not ( n3013 , n3012 );
not ( n3014 , n3013 );
not ( n3015 , n3014 );
not ( n3016 , n2899 );
and ( n3017 , n3016 , n2839 );
xor ( n3018 , n2974 , n2981 );
and ( n3019 , n3018 , n2899 );
or ( n3020 , n3017 , n3019 );
not ( n3021 , n3020 );
not ( n3022 , n3021 );
not ( n3023 , n3022 );
not ( n3024 , n2899 );
and ( n3025 , n3024 , n2824 );
xor ( n3026 , n2975 , n2980 );
and ( n3027 , n3026 , n2899 );
or ( n3028 , n3025 , n3027 );
not ( n3029 , n3028 );
not ( n3030 , n3029 );
not ( n3031 , n3030 );
not ( n3032 , n2899 );
and ( n3033 , n3032 , n2809 );
xor ( n3034 , n2976 , n2979 );
and ( n3035 , n3034 , n2899 );
or ( n3036 , n3033 , n3035 );
not ( n3037 , n3036 );
not ( n3038 , n3037 );
not ( n3039 , n3038 );
not ( n3040 , n2899 );
and ( n3041 , n3040 , n2794 );
xor ( n3042 , n2977 , n2978 );
and ( n3043 , n3042 , n2899 );
or ( n3044 , n3041 , n3043 );
not ( n3045 , n3044 );
not ( n3046 , n3045 );
not ( n3047 , n3046 );
not ( n3048 , n2960 );
and ( n3049 , n3047 , n3048 );
and ( n3050 , n3039 , n3049 );
and ( n3051 , n3031 , n3050 );
and ( n3052 , n3023 , n3051 );
and ( n3053 , n3015 , n3052 );
and ( n3054 , n3007 , n3053 );
and ( n3055 , n2999 , n3054 );
and ( n3056 , n2991 , n3055 );
not ( n3057 , n3056 );
and ( n3058 , n3057 , n2899 );
or ( n3059 , n2966 , n3058 );
and ( n3060 , n2964 , n3059 );
not ( n3061 , n3060 );
and ( n3062 , n3061 , n2962 );
xor ( n3063 , n2962 , n3059 );
xor ( n3064 , n3063 , n3059 );
and ( n3065 , n3064 , n3060 );
or ( n3066 , n3062 , n3065 );
not ( n3067 , n2899 );
and ( n3068 , n3067 , n2794 );
not ( n3069 , n2794 );
not ( n3070 , n2779 );
not ( n3071 , n2764 );
not ( n3072 , n2749 );
not ( n3073 , n2734 );
not ( n3074 , n2719 );
not ( n3075 , n2704 );
not ( n3076 , n2689 );
not ( n3077 , n2674 );
not ( n3078 , n2659 );
not ( n3079 , n2644 );
not ( n3080 , n2629 );
not ( n3081 , n2614 );
not ( n3082 , n2599 );
not ( n3083 , n2584 );
not ( n3084 , n2569 );
not ( n3085 , n2554 );
not ( n3086 , n2539 );
not ( n3087 , n2524 );
not ( n3088 , n2509 );
not ( n3089 , n2494 );
not ( n3090 , n2479 );
not ( n3091 , n2464 );
not ( n3092 , n2449 );
not ( n3093 , n2430 );
and ( n3094 , n3092 , n3093 );
and ( n3095 , n3091 , n3094 );
and ( n3096 , n3090 , n3095 );
and ( n3097 , n3089 , n3096 );
and ( n3098 , n3088 , n3097 );
and ( n3099 , n3087 , n3098 );
and ( n3100 , n3086 , n3099 );
and ( n3101 , n3085 , n3100 );
and ( n3102 , n3084 , n3101 );
and ( n3103 , n3083 , n3102 );
and ( n3104 , n3082 , n3103 );
and ( n3105 , n3081 , n3104 );
and ( n3106 , n3080 , n3105 );
and ( n3107 , n3079 , n3106 );
and ( n3108 , n3078 , n3107 );
and ( n3109 , n3077 , n3108 );
and ( n3110 , n3076 , n3109 );
and ( n3111 , n3075 , n3110 );
and ( n3112 , n3074 , n3111 );
and ( n3113 , n3073 , n3112 );
and ( n3114 , n3072 , n3113 );
and ( n3115 , n3071 , n3114 );
and ( n3116 , n3070 , n3115 );
xor ( n3117 , n3069 , n3116 );
and ( n3118 , n3117 , n2899 );
or ( n3119 , n3068 , n3118 );
not ( n3120 , n3119 );
not ( n3121 , n3120 );
not ( n3122 , n3121 );
not ( n3123 , n3122 );
not ( n3124 , n2899 );
and ( n3125 , n3124 , n2424 );
buf ( n3126 , n2899 );
not ( n3127 , n3126 );
and ( n3128 , n3127 , n2899 );
not ( n3129 , n2899 );
not ( n3130 , n2884 );
not ( n3131 , n2869 );
not ( n3132 , n2854 );
not ( n3133 , n2839 );
not ( n3134 , n2824 );
not ( n3135 , n2809 );
and ( n3136 , n3069 , n3116 );
and ( n3137 , n3135 , n3136 );
and ( n3138 , n3134 , n3137 );
and ( n3139 , n3133 , n3138 );
and ( n3140 , n3132 , n3139 );
and ( n3141 , n3131 , n3140 );
and ( n3142 , n3130 , n3141 );
xor ( n3143 , n3129 , n3142 );
and ( n3144 , n3143 , n3126 );
or ( n3145 , n3128 , n3144 );
not ( n3146 , n3145 );
not ( n3147 , n3146 );
not ( n3148 , n3147 );
not ( n3149 , n2899 );
and ( n3150 , n3149 , n2884 );
xor ( n3151 , n3130 , n3141 );
and ( n3152 , n3151 , n2899 );
or ( n3153 , n3150 , n3152 );
not ( n3154 , n3153 );
not ( n3155 , n3154 );
not ( n3156 , n3155 );
not ( n3157 , n2899 );
and ( n3158 , n3157 , n2869 );
xor ( n3159 , n3131 , n3140 );
and ( n3160 , n3159 , n2899 );
or ( n3161 , n3158 , n3160 );
not ( n3162 , n3161 );
not ( n3163 , n3162 );
not ( n3164 , n3163 );
not ( n3165 , n2899 );
and ( n3166 , n3165 , n2854 );
xor ( n3167 , n3132 , n3139 );
and ( n3168 , n3167 , n2899 );
or ( n3169 , n3166 , n3168 );
not ( n3170 , n3169 );
not ( n3171 , n3170 );
not ( n3172 , n3171 );
not ( n3173 , n2899 );
and ( n3174 , n3173 , n2839 );
xor ( n3175 , n3133 , n3138 );
and ( n3176 , n3175 , n2899 );
or ( n3177 , n3174 , n3176 );
not ( n3178 , n3177 );
not ( n3179 , n3178 );
not ( n3180 , n3179 );
not ( n3181 , n2899 );
and ( n3182 , n3181 , n2824 );
xor ( n3183 , n3134 , n3137 );
and ( n3184 , n3183 , n2899 );
or ( n3185 , n3182 , n3184 );
not ( n3186 , n3185 );
not ( n3187 , n3186 );
not ( n3188 , n3187 );
not ( n3189 , n2899 );
and ( n3190 , n3189 , n2809 );
xor ( n3191 , n3135 , n3136 );
and ( n3192 , n3191 , n2899 );
or ( n3193 , n3190 , n3192 );
not ( n3194 , n3193 );
not ( n3195 , n3194 );
not ( n3196 , n3195 );
not ( n3197 , n3121 );
and ( n3198 , n3196 , n3197 );
and ( n3199 , n3188 , n3198 );
and ( n3200 , n3180 , n3199 );
and ( n3201 , n3172 , n3200 );
and ( n3202 , n3164 , n3201 );
and ( n3203 , n3156 , n3202 );
and ( n3204 , n3148 , n3203 );
not ( n3205 , n3204 );
and ( n3206 , n3205 , n2899 );
or ( n3207 , n3125 , n3206 );
not ( n3208 , n3207 );
not ( n3209 , n2899 );
and ( n3210 , n3209 , n3195 );
xor ( n3211 , n3196 , n3197 );
and ( n3212 , n3211 , n2899 );
or ( n3213 , n3210 , n3212 );
and ( n3214 , n3208 , n3213 );
not ( n3215 , n3213 );
not ( n3216 , n3121 );
xor ( n3217 , n3215 , n3216 );
and ( n3218 , n3217 , n3207 );
or ( n3219 , n3214 , n3218 );
not ( n3220 , n3219 );
not ( n3221 , n3220 );
or ( n3222 , n3123 , n3221 );
not ( n3223 , n3207 );
not ( n3224 , n2899 );
and ( n3225 , n3224 , n3187 );
xor ( n3226 , n3188 , n3198 );
and ( n3227 , n3226 , n2899 );
or ( n3228 , n3225 , n3227 );
and ( n3229 , n3223 , n3228 );
not ( n3230 , n3228 );
and ( n3231 , n3215 , n3216 );
xor ( n3232 , n3230 , n3231 );
and ( n3233 , n3232 , n3207 );
or ( n3234 , n3229 , n3233 );
not ( n3235 , n3234 );
not ( n3236 , n3235 );
or ( n3237 , n3222 , n3236 );
and ( n3238 , n3237 , n3207 );
not ( n3239 , n3238 );
and ( n3240 , n3239 , n3123 );
xor ( n3241 , n3123 , n3207 );
xor ( n3242 , n3241 , n3207 );
and ( n3243 , n3242 , n3238 );
or ( n3244 , n3240 , n3243 );
not ( n3245 , n3238 );
and ( n3246 , n3245 , n3221 );
xor ( n3247 , n3221 , n3207 );
and ( n3248 , n3241 , n3207 );
xor ( n3249 , n3247 , n3248 );
and ( n3250 , n3249 , n3238 );
or ( n3251 , n3246 , n3250 );
not ( n3252 , n3238 );
and ( n3253 , n3252 , n3236 );
xor ( n3254 , n3236 , n3207 );
and ( n3255 , n3247 , n3248 );
xor ( n3256 , n3254 , n3255 );
and ( n3257 , n3256 , n3238 );
or ( n3258 , n3253 , n3257 );
and ( n3259 , n3244 , n3251 , n3258 );
or ( n3260 , n3066 , n3259 );
not ( n3261 , n3260 );
not ( n3262 , n3244 );
not ( n3263 , n3258 );
nor ( n3264 , n3262 , n3251 , n3263 );
not ( n3265 , n3264 );
nor ( n3266 , n3244 , n3251 , n3263 );
not ( n3267 , n3266 );
and ( n3268 , n3244 , n3251 , n3263 );
not ( n3269 , n3268 );
and ( n3270 , n3262 , n3251 , n3263 );
not ( n3271 , n3270 );
nor ( n3272 , n3262 , n3251 , n3258 );
not ( n3273 , n3272 );
nor ( n3274 , n3244 , n3251 , n3258 );
not ( n3275 , n3274 );
and ( n3276 , n3275 , n2904 );
and ( n3277 , n2424 , n3274 );
or ( n3278 , n3276 , n3277 );
and ( n3279 , n3273 , n3278 );
or ( n3280 , n2282 , n2423 );
and ( n3281 , n3280 , n3272 );
or ( n3282 , n3279 , n3281 );
and ( n3283 , n3271 , n3282 );
and ( n3284 , n2424 , n3270 );
or ( n3285 , n3283 , n3284 );
and ( n3286 , n3269 , n3285 );
and ( n3287 , n3280 , n3268 );
or ( n3288 , n3286 , n3287 );
and ( n3289 , n3267 , n3288 );
buf ( n3290 , DFF_B_reg_Q);
not ( n3291 , n3290 );
and ( n3292 , n3291 , n2904 );
and ( n3293 , n3280 , n3290 );
or ( n3294 , n3292 , n3293 );
and ( n3295 , n3294 , n3266 );
or ( n3296 , n3289 , n3295 );
and ( n3297 , n3265 , n3296 );
not ( n3298 , n3290 );
not ( n3299 , n3298 );
and ( n3300 , n3299 , n2904 );
and ( n3301 , n3280 , n3298 );
or ( n3302 , n3300 , n3301 );
and ( n3303 , n3302 , n3264 );
or ( n3304 , n3297 , n3303 );
and ( n3305 , n3261 , n3304 );
and ( n3306 , n2904 , n3260 );
or ( n3307 , n3305 , n3306 );
and ( n3308 , n3307 , n2422 );
and ( n3309 , n2904 , n2428 );
or ( n3310 , n3308 , n3309 );
buf ( n3311 , n3310 );
buf ( n3312 , n65 );
buf ( n3313 , n2424 );
buf ( n3314 , n2281 );
buf ( n3315 , n2280 );
not ( n3316 , n3260 );
not ( n3317 , n3264 );
not ( n3318 , n3266 );
not ( n3319 , n3268 );
not ( n3320 , n3270 );
not ( n3321 , n3272 );
not ( n3322 , n3274 );
and ( n3323 , n3322 , n3312 );
and ( n3324 , n2424 , n3274 );
or ( n3325 , n3323 , n3324 );
and ( n3326 , n3321 , n3325 );
and ( n3327 , n2424 , n3272 );
or ( n3328 , n3326 , n3327 );
and ( n3329 , n3320 , n3328 );
and ( n3330 , n3280 , n3270 );
or ( n3331 , n3329 , n3330 );
and ( n3332 , n3319 , n3331 );
and ( n3333 , n3280 , n3268 );
or ( n3334 , n3332 , n3333 );
and ( n3335 , n3318 , n3334 );
not ( n3336 , n3290 );
and ( n3337 , n3336 , n3312 );
and ( n3338 , n3280 , n3290 );
or ( n3339 , n3337 , n3338 );
and ( n3340 , n3339 , n3266 );
or ( n3341 , n3335 , n3340 );
and ( n3342 , n3317 , n3341 );
not ( n3343 , n3298 );
and ( n3344 , n3343 , n3312 );
and ( n3345 , n3280 , n3298 );
or ( n3346 , n3344 , n3345 );
and ( n3347 , n3346 , n3264 );
or ( n3348 , n3342 , n3347 );
and ( n3349 , n3316 , n3348 );
and ( n3350 , n3312 , n3260 );
or ( n3351 , n3349 , n3350 );
and ( n3352 , n3351 , n2422 );
and ( n3353 , n3312 , n2428 );
or ( n3354 , n3352 , n3353 );
buf ( n3355 , n3354 );
buf ( n3356 , n66 );
buf ( n3357 , n2424 );
buf ( n3358 , n2281 );
buf ( n3359 , n2280 );
not ( n3360 , n3260 );
not ( n3361 , n3356 );
not ( n3362 , n3361 );
buf ( n3363 , n3362 );
not ( n3364 , n2899 );
and ( n3365 , n3364 , n2719 );
not ( n3366 , n2719 );
not ( n3367 , n2704 );
not ( n3368 , n2689 );
not ( n3369 , n2674 );
not ( n3370 , n2659 );
not ( n3371 , n2644 );
not ( n3372 , n2629 );
not ( n3373 , n2614 );
not ( n3374 , n2599 );
not ( n3375 , n2584 );
not ( n3376 , n2569 );
not ( n3377 , n2554 );
not ( n3378 , n2539 );
not ( n3379 , n2524 );
not ( n3380 , n2509 );
not ( n3381 , n2494 );
not ( n3382 , n2479 );
not ( n3383 , n2464 );
not ( n3384 , n2449 );
not ( n3385 , n2430 );
and ( n3386 , n3384 , n3385 );
and ( n3387 , n3383 , n3386 );
and ( n3388 , n3382 , n3387 );
and ( n3389 , n3381 , n3388 );
and ( n3390 , n3380 , n3389 );
and ( n3391 , n3379 , n3390 );
and ( n3392 , n3378 , n3391 );
and ( n3393 , n3377 , n3392 );
and ( n3394 , n3376 , n3393 );
and ( n3395 , n3375 , n3394 );
and ( n3396 , n3374 , n3395 );
and ( n3397 , n3373 , n3396 );
and ( n3398 , n3372 , n3397 );
and ( n3399 , n3371 , n3398 );
and ( n3400 , n3370 , n3399 );
and ( n3401 , n3369 , n3400 );
and ( n3402 , n3368 , n3401 );
and ( n3403 , n3367 , n3402 );
xor ( n3404 , n3366 , n3403 );
and ( n3405 , n3404 , n2899 );
or ( n3406 , n3365 , n3405 );
not ( n3407 , n3406 );
not ( n3408 , n3407 );
not ( n3409 , n3408 );
not ( n3410 , n3409 );
not ( n3411 , n2899 );
and ( n3412 , n3411 , n2424 );
buf ( n3413 , n2899 );
not ( n3414 , n3413 );
and ( n3415 , n3414 , n2899 );
not ( n3416 , n2899 );
not ( n3417 , n2884 );
not ( n3418 , n2869 );
not ( n3419 , n2854 );
not ( n3420 , n2839 );
not ( n3421 , n2824 );
not ( n3422 , n2809 );
not ( n3423 , n2794 );
not ( n3424 , n2779 );
not ( n3425 , n2764 );
not ( n3426 , n2749 );
not ( n3427 , n2734 );
and ( n3428 , n3366 , n3403 );
and ( n3429 , n3427 , n3428 );
and ( n3430 , n3426 , n3429 );
and ( n3431 , n3425 , n3430 );
and ( n3432 , n3424 , n3431 );
and ( n3433 , n3423 , n3432 );
and ( n3434 , n3422 , n3433 );
and ( n3435 , n3421 , n3434 );
and ( n3436 , n3420 , n3435 );
and ( n3437 , n3419 , n3436 );
and ( n3438 , n3418 , n3437 );
and ( n3439 , n3417 , n3438 );
xor ( n3440 , n3416 , n3439 );
and ( n3441 , n3440 , n3413 );
or ( n3442 , n3415 , n3441 );
not ( n3443 , n3442 );
not ( n3444 , n3443 );
not ( n3445 , n3444 );
not ( n3446 , n2899 );
and ( n3447 , n3446 , n2884 );
xor ( n3448 , n3417 , n3438 );
and ( n3449 , n3448 , n2899 );
or ( n3450 , n3447 , n3449 );
not ( n3451 , n3450 );
not ( n3452 , n3451 );
not ( n3453 , n3452 );
not ( n3454 , n2899 );
and ( n3455 , n3454 , n2869 );
xor ( n3456 , n3418 , n3437 );
and ( n3457 , n3456 , n2899 );
or ( n3458 , n3455 , n3457 );
not ( n3459 , n3458 );
not ( n3460 , n3459 );
not ( n3461 , n3460 );
not ( n3462 , n2899 );
and ( n3463 , n3462 , n2854 );
xor ( n3464 , n3419 , n3436 );
and ( n3465 , n3464 , n2899 );
or ( n3466 , n3463 , n3465 );
not ( n3467 , n3466 );
not ( n3468 , n3467 );
not ( n3469 , n3468 );
not ( n3470 , n2899 );
and ( n3471 , n3470 , n2839 );
xor ( n3472 , n3420 , n3435 );
and ( n3473 , n3472 , n2899 );
or ( n3474 , n3471 , n3473 );
not ( n3475 , n3474 );
not ( n3476 , n3475 );
not ( n3477 , n3476 );
not ( n3478 , n2899 );
and ( n3479 , n3478 , n2824 );
xor ( n3480 , n3421 , n3434 );
and ( n3481 , n3480 , n2899 );
or ( n3482 , n3479 , n3481 );
not ( n3483 , n3482 );
not ( n3484 , n3483 );
not ( n3485 , n3484 );
not ( n3486 , n2899 );
and ( n3487 , n3486 , n2809 );
xor ( n3488 , n3422 , n3433 );
and ( n3489 , n3488 , n2899 );
or ( n3490 , n3487 , n3489 );
not ( n3491 , n3490 );
not ( n3492 , n3491 );
not ( n3493 , n3492 );
not ( n3494 , n2899 );
and ( n3495 , n3494 , n2794 );
xor ( n3496 , n3423 , n3432 );
and ( n3497 , n3496 , n2899 );
or ( n3498 , n3495 , n3497 );
not ( n3499 , n3498 );
not ( n3500 , n3499 );
not ( n3501 , n3500 );
not ( n3502 , n2899 );
and ( n3503 , n3502 , n2779 );
xor ( n3504 , n3424 , n3431 );
and ( n3505 , n3504 , n2899 );
or ( n3506 , n3503 , n3505 );
not ( n3507 , n3506 );
not ( n3508 , n3507 );
not ( n3509 , n3508 );
not ( n3510 , n2899 );
and ( n3511 , n3510 , n2764 );
xor ( n3512 , n3425 , n3430 );
and ( n3513 , n3512 , n2899 );
or ( n3514 , n3511 , n3513 );
not ( n3515 , n3514 );
not ( n3516 , n3515 );
not ( n3517 , n3516 );
not ( n3518 , n2899 );
and ( n3519 , n3518 , n2749 );
xor ( n3520 , n3426 , n3429 );
and ( n3521 , n3520 , n2899 );
or ( n3522 , n3519 , n3521 );
not ( n3523 , n3522 );
not ( n3524 , n3523 );
not ( n3525 , n3524 );
not ( n3526 , n2899 );
and ( n3527 , n3526 , n2734 );
xor ( n3528 , n3427 , n3428 );
and ( n3529 , n3528 , n2899 );
or ( n3530 , n3527 , n3529 );
not ( n3531 , n3530 );
not ( n3532 , n3531 );
not ( n3533 , n3532 );
not ( n3534 , n3408 );
and ( n3535 , n3533 , n3534 );
and ( n3536 , n3525 , n3535 );
and ( n3537 , n3517 , n3536 );
and ( n3538 , n3509 , n3537 );
and ( n3539 , n3501 , n3538 );
and ( n3540 , n3493 , n3539 );
and ( n3541 , n3485 , n3540 );
and ( n3542 , n3477 , n3541 );
and ( n3543 , n3469 , n3542 );
and ( n3544 , n3461 , n3543 );
and ( n3545 , n3453 , n3544 );
and ( n3546 , n3445 , n3545 );
not ( n3547 , n3546 );
and ( n3548 , n3547 , n2899 );
or ( n3549 , n3412 , n3548 );
not ( n3550 , n3549 );
not ( n3551 , n2899 );
and ( n3552 , n3551 , n3532 );
xor ( n3553 , n3533 , n3534 );
and ( n3554 , n3553 , n2899 );
or ( n3555 , n3552 , n3554 );
and ( n3556 , n3550 , n3555 );
not ( n3557 , n3555 );
not ( n3558 , n3408 );
xor ( n3559 , n3557 , n3558 );
and ( n3560 , n3559 , n3549 );
or ( n3561 , n3556 , n3560 );
not ( n3562 , n3561 );
not ( n3563 , n3562 );
or ( n3564 , n3410 , n3563 );
not ( n3565 , n3549 );
not ( n3566 , n2899 );
and ( n3567 , n3566 , n3524 );
xor ( n3568 , n3525 , n3535 );
and ( n3569 , n3568 , n2899 );
or ( n3570 , n3567 , n3569 );
and ( n3571 , n3565 , n3570 );
not ( n3572 , n3570 );
and ( n3573 , n3557 , n3558 );
xor ( n3574 , n3572 , n3573 );
and ( n3575 , n3574 , n3549 );
or ( n3576 , n3571 , n3575 );
not ( n3577 , n3576 );
not ( n3578 , n3577 );
or ( n3579 , n3564 , n3578 );
not ( n3580 , n3549 );
not ( n3581 , n2899 );
and ( n3582 , n3581 , n3516 );
xor ( n3583 , n3517 , n3536 );
and ( n3584 , n3583 , n2899 );
or ( n3585 , n3582 , n3584 );
and ( n3586 , n3580 , n3585 );
not ( n3587 , n3585 );
and ( n3588 , n3572 , n3573 );
xor ( n3589 , n3587 , n3588 );
and ( n3590 , n3589 , n3549 );
or ( n3591 , n3586 , n3590 );
not ( n3592 , n3591 );
not ( n3593 , n3592 );
or ( n3594 , n3579 , n3593 );
buf ( n3595 , n3594 );
buf ( n3596 , n3595 );
and ( n3597 , n3596 , n3549 );
not ( n3598 , n3597 );
and ( n3599 , n3598 , n3410 );
xor ( n3600 , n3410 , n3549 );
xor ( n3601 , n3600 , n3549 );
and ( n3602 , n3601 , n3597 );
or ( n3603 , n3599 , n3602 );
not ( n3604 , n3597 );
and ( n3605 , n3604 , n3563 );
xor ( n3606 , n3563 , n3549 );
and ( n3607 , n3600 , n3549 );
xor ( n3608 , n3606 , n3607 );
and ( n3609 , n3608 , n3597 );
or ( n3610 , n3605 , n3609 );
not ( n3611 , n3610 );
not ( n3612 , n3597 );
and ( n3613 , n3612 , n3578 );
xor ( n3614 , n3578 , n3549 );
and ( n3615 , n3606 , n3607 );
xor ( n3616 , n3614 , n3615 );
and ( n3617 , n3616 , n3597 );
or ( n3618 , n3613 , n3617 );
not ( n3619 , n3597 );
and ( n3620 , n3619 , n3593 );
xor ( n3621 , n3593 , n3549 );
and ( n3622 , n3614 , n3615 );
xor ( n3623 , n3621 , n3622 );
and ( n3624 , n3623 , n3597 );
or ( n3625 , n3620 , n3624 );
and ( n3626 , n3603 , n3611 , n3618 , n3625 );
not ( n3627 , n3603 );
and ( n3628 , n3627 , n3610 , n3618 , n3625 );
or ( n3629 , n3626 , n3628 );
and ( n3630 , n3603 , n3610 , n3618 , n3625 );
or ( n3631 , n3629 , n3630 );
and ( n3632 , n3363 , n3631 );
buf ( n3633 , n2424 );
not ( n3634 , n3290 );
buf ( n3635 , n190 );
not ( n3636 , n2899 );
and ( n3637 , n3636 , n2869 );
not ( n3638 , n2869 );
not ( n3639 , n2854 );
not ( n3640 , n2839 );
not ( n3641 , n2824 );
not ( n3642 , n2809 );
not ( n3643 , n2794 );
not ( n3644 , n2779 );
not ( n3645 , n2764 );
not ( n3646 , n2749 );
not ( n3647 , n2734 );
not ( n3648 , n2719 );
not ( n3649 , n2704 );
not ( n3650 , n2689 );
not ( n3651 , n2674 );
not ( n3652 , n2659 );
not ( n3653 , n2644 );
not ( n3654 , n2629 );
not ( n3655 , n2614 );
not ( n3656 , n2599 );
not ( n3657 , n2584 );
not ( n3658 , n2569 );
not ( n3659 , n2554 );
not ( n3660 , n2539 );
not ( n3661 , n2524 );
not ( n3662 , n2509 );
not ( n3663 , n2494 );
not ( n3664 , n2479 );
not ( n3665 , n2464 );
not ( n3666 , n2449 );
not ( n3667 , n2430 );
and ( n3668 , n3666 , n3667 );
and ( n3669 , n3665 , n3668 );
and ( n3670 , n3664 , n3669 );
and ( n3671 , n3663 , n3670 );
and ( n3672 , n3662 , n3671 );
and ( n3673 , n3661 , n3672 );
and ( n3674 , n3660 , n3673 );
and ( n3675 , n3659 , n3674 );
and ( n3676 , n3658 , n3675 );
and ( n3677 , n3657 , n3676 );
and ( n3678 , n3656 , n3677 );
and ( n3679 , n3655 , n3678 );
and ( n3680 , n3654 , n3679 );
and ( n3681 , n3653 , n3680 );
and ( n3682 , n3652 , n3681 );
and ( n3683 , n3651 , n3682 );
and ( n3684 , n3650 , n3683 );
and ( n3685 , n3649 , n3684 );
and ( n3686 , n3648 , n3685 );
and ( n3687 , n3647 , n3686 );
and ( n3688 , n3646 , n3687 );
and ( n3689 , n3645 , n3688 );
and ( n3690 , n3644 , n3689 );
and ( n3691 , n3643 , n3690 );
and ( n3692 , n3642 , n3691 );
and ( n3693 , n3641 , n3692 );
and ( n3694 , n3640 , n3693 );
and ( n3695 , n3639 , n3694 );
xor ( n3696 , n3638 , n3695 );
and ( n3697 , n3696 , n2899 );
or ( n3698 , n3637 , n3697 );
not ( n3699 , n3698 );
not ( n3700 , n3699 );
not ( n3701 , n3700 );
not ( n3702 , n3701 );
not ( n3703 , n2899 );
and ( n3704 , n3703 , n2424 );
buf ( n3705 , n2899 );
not ( n3706 , n3705 );
and ( n3707 , n3706 , n2899 );
not ( n3708 , n2899 );
not ( n3709 , n2884 );
and ( n3710 , n3638 , n3695 );
and ( n3711 , n3709 , n3710 );
xor ( n3712 , n3708 , n3711 );
and ( n3713 , n3712 , n3705 );
or ( n3714 , n3707 , n3713 );
not ( n3715 , n3714 );
not ( n3716 , n3715 );
not ( n3717 , n3716 );
not ( n3718 , n2899 );
and ( n3719 , n3718 , n2884 );
xor ( n3720 , n3709 , n3710 );
and ( n3721 , n3720 , n2899 );
or ( n3722 , n3719 , n3721 );
not ( n3723 , n3722 );
not ( n3724 , n3723 );
not ( n3725 , n3724 );
not ( n3726 , n3700 );
and ( n3727 , n3725 , n3726 );
and ( n3728 , n3717 , n3727 );
not ( n3729 , n3728 );
and ( n3730 , n3729 , n2899 );
or ( n3731 , n3704 , n3730 );
not ( n3732 , n3731 );
not ( n3733 , n2899 );
and ( n3734 , n3733 , n3724 );
xor ( n3735 , n3725 , n3726 );
and ( n3736 , n3735 , n2899 );
or ( n3737 , n3734 , n3736 );
and ( n3738 , n3732 , n3737 );
not ( n3739 , n3737 );
not ( n3740 , n3700 );
xor ( n3741 , n3739 , n3740 );
and ( n3742 , n3741 , n3731 );
or ( n3743 , n3738 , n3742 );
not ( n3744 , n3743 );
not ( n3745 , n3744 );
or ( n3746 , n3702 , n3745 );
and ( n3747 , n3746 , n3731 );
not ( n3748 , n3747 );
and ( n3749 , n3748 , n3702 );
xor ( n3750 , n3702 , n3731 );
xor ( n3751 , n3750 , n3731 );
and ( n3752 , n3751 , n3747 );
or ( n3753 , n3749 , n3752 );
not ( n3754 , n3753 );
not ( n3755 , n3747 );
and ( n3756 , n3755 , n3745 );
xor ( n3757 , n3745 , n3731 );
and ( n3758 , n3750 , n3731 );
xor ( n3759 , n3757 , n3758 );
and ( n3760 , n3759 , n3747 );
or ( n3761 , n3756 , n3760 );
and ( n3762 , n3754 , n3761 );
and ( n3763 , n3635 , n3762 );
buf ( n3764 , n126 );
nor ( n3765 , n3754 , n3761 );
and ( n3766 , n3764 , n3765 );
buf ( n3767 , n158 );
nor ( n3768 , n3753 , n3761 );
and ( n3769 , n3767 , n3768 );
or ( n3770 , n2424 , n3763 , n3766 , n3769 );
not ( n3771 , n3770 );
buf ( n3772 , n67 );
buf ( n3773 , n3772 );
not ( n3774 , n3773 );
not ( n3775 , n3774 );
buf ( n3776 , n3775 );
and ( n3777 , n3753 , n3761 );
and ( n3778 , n3776 , n3777 );
buf ( n3779 , n160 );
and ( n3780 , n3779 , n3762 );
buf ( n3781 , n96 );
and ( n3782 , n3781 , n3765 );
buf ( n3783 , n128 );
and ( n3784 , n3783 , n3768 );
or ( n3785 , n3778 , n3780 , n3782 , n3784 );
and ( n3786 , n3771 , n3785 );
not ( n3787 , n3785 );
and ( n3788 , n3363 , n3777 );
buf ( n3789 , n159 );
and ( n3790 , n3789 , n3762 );
buf ( n3791 , n95 );
and ( n3792 , n3791 , n3765 );
buf ( n3793 , n127 );
and ( n3794 , n3793 , n3768 );
or ( n3795 , n3788 , n3790 , n3792 , n3794 );
not ( n3796 , n3795 );
xor ( n3797 , n3787 , n3796 );
and ( n3798 , n3797 , n3770 );
or ( n3799 , n3786 , n3798 );
not ( n3800 , n3799 );
buf ( n3801 , n3800 );
buf ( n3802 , n3801 );
not ( n3803 , n3802 );
and ( n3804 , n3634 , n3803 );
not ( n3805 , n3803 );
not ( n3806 , n3805 );
not ( n3807 , n3770 );
and ( n3808 , n3807 , n2424 );
buf ( n3809 , n3770 );
not ( n3810 , n3809 );
and ( n3811 , n3810 , n3770 );
not ( n3812 , n3770 );
buf ( n3813 , n189 );
and ( n3814 , n3813 , n3762 );
buf ( n3815 , n125 );
and ( n3816 , n3815 , n3765 );
buf ( n3817 , n157 );
and ( n3818 , n3817 , n3768 );
or ( n3819 , n2424 , n3814 , n3816 , n3818 );
not ( n3820 , n3819 );
buf ( n3821 , n94 );
buf ( n3822 , n3821 );
not ( n3823 , n3822 );
not ( n3824 , n3823 );
buf ( n3825 , n3824 );
buf ( n3826 , n93 );
buf ( n3827 , n3826 );
not ( n3828 , n3827 );
not ( n3829 , n3828 );
buf ( n3830 , n3829 );
buf ( n3831 , n92 );
buf ( n3832 , n3831 );
not ( n3833 , n3832 );
not ( n3834 , n3833 );
buf ( n3835 , n3834 );
buf ( n3836 , n91 );
buf ( n3837 , n3836 );
not ( n3838 , n3837 );
not ( n3839 , n3838 );
buf ( n3840 , n3839 );
buf ( n3841 , n90 );
buf ( n3842 , n3841 );
not ( n3843 , n3842 );
not ( n3844 , n3843 );
buf ( n3845 , n3844 );
buf ( n3846 , n89 );
buf ( n3847 , n3846 );
not ( n3848 , n3847 );
not ( n3849 , n3848 );
buf ( n3850 , n3849 );
buf ( n3851 , n88 );
buf ( n3852 , n3851 );
not ( n3853 , n3852 );
not ( n3854 , n3853 );
buf ( n3855 , n3854 );
buf ( n3856 , n87 );
buf ( n3857 , n3856 );
not ( n3858 , n3857 );
not ( n3859 , n3858 );
buf ( n3860 , n3859 );
buf ( n3861 , n86 );
buf ( n3862 , n3861 );
not ( n3863 , n3862 );
not ( n3864 , n3863 );
buf ( n3865 , n3864 );
buf ( n3866 , n85 );
buf ( n3867 , n3866 );
not ( n3868 , n3867 );
not ( n3869 , n3868 );
buf ( n3870 , n3869 );
buf ( n3871 , n84 );
buf ( n3872 , n3871 );
not ( n3873 , n3872 );
not ( n3874 , n3873 );
buf ( n3875 , n3874 );
buf ( n3876 , n83 );
buf ( n3877 , n3876 );
not ( n3878 , n3877 );
not ( n3879 , n3878 );
buf ( n3880 , n3879 );
buf ( n3881 , n82 );
buf ( n3882 , n3881 );
not ( n3883 , n3882 );
not ( n3884 , n3883 );
buf ( n3885 , n3884 );
buf ( n3886 , n81 );
buf ( n3887 , n3886 );
not ( n3888 , n3887 );
not ( n3889 , n3888 );
buf ( n3890 , n3889 );
buf ( n3891 , n80 );
buf ( n3892 , n3891 );
not ( n3893 , n3892 );
not ( n3894 , n3893 );
buf ( n3895 , n3894 );
buf ( n3896 , n79 );
buf ( n3897 , n3896 );
not ( n3898 , n3897 );
not ( n3899 , n3898 );
buf ( n3900 , n3899 );
buf ( n3901 , n78 );
buf ( n3902 , n3901 );
not ( n3903 , n3902 );
not ( n3904 , n3903 );
buf ( n3905 , n3904 );
buf ( n3906 , n77 );
buf ( n3907 , n3906 );
not ( n3908 , n3907 );
not ( n3909 , n3908 );
buf ( n3910 , n3909 );
buf ( n3911 , n76 );
buf ( n3912 , n3911 );
not ( n3913 , n3912 );
not ( n3914 , n3913 );
buf ( n3915 , n3914 );
buf ( n3916 , n75 );
buf ( n3917 , n3916 );
not ( n3918 , n3917 );
not ( n3919 , n3918 );
buf ( n3920 , n3919 );
buf ( n3921 , n74 );
buf ( n3922 , n3921 );
not ( n3923 , n3922 );
not ( n3924 , n3923 );
buf ( n3925 , n3924 );
buf ( n3926 , n73 );
buf ( n3927 , n3926 );
not ( n3928 , n3927 );
not ( n3929 , n3928 );
buf ( n3930 , n3929 );
buf ( n3931 , n72 );
buf ( n3932 , n3931 );
not ( n3933 , n3932 );
not ( n3934 , n3933 );
buf ( n3935 , n3934 );
buf ( n3936 , n71 );
buf ( n3937 , n3936 );
not ( n3938 , n3937 );
not ( n3939 , n3938 );
buf ( n3940 , n3939 );
buf ( n3941 , n70 );
buf ( n3942 , n3941 );
not ( n3943 , n3942 );
not ( n3944 , n3943 );
buf ( n3945 , n3944 );
buf ( n3946 , n69 );
buf ( n3947 , n3946 );
not ( n3948 , n3947 );
not ( n3949 , n3948 );
buf ( n3950 , n3949 );
and ( n3951 , n3945 , n3950 );
and ( n3952 , n3940 , n3951 );
and ( n3953 , n3935 , n3952 );
and ( n3954 , n3930 , n3953 );
and ( n3955 , n3925 , n3954 );
and ( n3956 , n3920 , n3955 );
and ( n3957 , n3915 , n3956 );
and ( n3958 , n3910 , n3957 );
and ( n3959 , n3905 , n3958 );
and ( n3960 , n3900 , n3959 );
and ( n3961 , n3895 , n3960 );
and ( n3962 , n3890 , n3961 );
and ( n3963 , n3885 , n3962 );
and ( n3964 , n3880 , n3963 );
and ( n3965 , n3875 , n3964 );
and ( n3966 , n3870 , n3965 );
and ( n3967 , n3865 , n3966 );
and ( n3968 , n3860 , n3967 );
and ( n3969 , n3855 , n3968 );
and ( n3970 , n3850 , n3969 );
and ( n3971 , n3845 , n3970 );
and ( n3972 , n3840 , n3971 );
and ( n3973 , n3835 , n3972 );
and ( n3974 , n3830 , n3973 );
and ( n3975 , n3825 , n3974 );
buf ( n3976 , n3975 );
and ( n3977 , n3976 , n3777 );
buf ( n3978 , n188 );
and ( n3979 , n3978 , n3762 );
buf ( n3980 , n124 );
and ( n3981 , n3980 , n3765 );
buf ( n3982 , n156 );
and ( n3983 , n3982 , n3768 );
or ( n3984 , n3977 , n3979 , n3981 , n3983 );
not ( n3985 , n3984 );
xor ( n3986 , n3825 , n3974 );
and ( n3987 , n3986 , n3777 );
buf ( n3988 , n187 );
and ( n3989 , n3988 , n3762 );
buf ( n3990 , n123 );
and ( n3991 , n3990 , n3765 );
buf ( n3992 , n155 );
and ( n3993 , n3992 , n3768 );
or ( n3994 , n3987 , n3989 , n3991 , n3993 );
not ( n3995 , n3994 );
xor ( n3996 , n3830 , n3973 );
and ( n3997 , n3996 , n3777 );
buf ( n3998 , n186 );
and ( n3999 , n3998 , n3762 );
buf ( n4000 , n122 );
and ( n4001 , n4000 , n3765 );
buf ( n4002 , n154 );
and ( n4003 , n4002 , n3768 );
or ( n4004 , n3997 , n3999 , n4001 , n4003 );
not ( n4005 , n4004 );
xor ( n4006 , n3835 , n3972 );
and ( n4007 , n4006 , n3777 );
buf ( n4008 , n185 );
and ( n4009 , n4008 , n3762 );
buf ( n4010 , n121 );
and ( n4011 , n4010 , n3765 );
buf ( n4012 , n153 );
and ( n4013 , n4012 , n3768 );
or ( n4014 , n4007 , n4009 , n4011 , n4013 );
not ( n4015 , n4014 );
xor ( n4016 , n3840 , n3971 );
and ( n4017 , n4016 , n3777 );
buf ( n4018 , n184 );
and ( n4019 , n4018 , n3762 );
buf ( n4020 , n120 );
and ( n4021 , n4020 , n3765 );
buf ( n4022 , n152 );
and ( n4023 , n4022 , n3768 );
or ( n4024 , n4017 , n4019 , n4021 , n4023 );
not ( n4025 , n4024 );
xor ( n4026 , n3845 , n3970 );
and ( n4027 , n4026 , n3777 );
buf ( n4028 , n183 );
and ( n4029 , n4028 , n3762 );
buf ( n4030 , n119 );
and ( n4031 , n4030 , n3765 );
buf ( n4032 , n151 );
and ( n4033 , n4032 , n3768 );
or ( n4034 , n4027 , n4029 , n4031 , n4033 );
not ( n4035 , n4034 );
xor ( n4036 , n3850 , n3969 );
and ( n4037 , n4036 , n3777 );
buf ( n4038 , n182 );
and ( n4039 , n4038 , n3762 );
buf ( n4040 , n118 );
and ( n4041 , n4040 , n3765 );
buf ( n4042 , n150 );
and ( n4043 , n4042 , n3768 );
or ( n4044 , n4037 , n4039 , n4041 , n4043 );
not ( n4045 , n4044 );
xor ( n4046 , n3855 , n3968 );
and ( n4047 , n4046 , n3777 );
buf ( n4048 , n181 );
and ( n4049 , n4048 , n3762 );
buf ( n4050 , n117 );
and ( n4051 , n4050 , n3765 );
buf ( n4052 , n149 );
and ( n4053 , n4052 , n3768 );
or ( n4054 , n4047 , n4049 , n4051 , n4053 );
not ( n4055 , n4054 );
xor ( n4056 , n3860 , n3967 );
and ( n4057 , n4056 , n3777 );
buf ( n4058 , n180 );
and ( n4059 , n4058 , n3762 );
buf ( n4060 , n116 );
and ( n4061 , n4060 , n3765 );
buf ( n4062 , n148 );
and ( n4063 , n4062 , n3768 );
or ( n4064 , n4057 , n4059 , n4061 , n4063 );
not ( n4065 , n4064 );
xor ( n4066 , n3865 , n3966 );
and ( n4067 , n4066 , n3777 );
buf ( n4068 , n179 );
and ( n4069 , n4068 , n3762 );
buf ( n4070 , n115 );
and ( n4071 , n4070 , n3765 );
buf ( n4072 , n147 );
and ( n4073 , n4072 , n3768 );
or ( n4074 , n4067 , n4069 , n4071 , n4073 );
not ( n4075 , n4074 );
xor ( n4076 , n3870 , n3965 );
and ( n4077 , n4076 , n3777 );
buf ( n4078 , n178 );
and ( n4079 , n4078 , n3762 );
buf ( n4080 , n114 );
and ( n4081 , n4080 , n3765 );
buf ( n4082 , n146 );
and ( n4083 , n4082 , n3768 );
or ( n4084 , n4077 , n4079 , n4081 , n4083 );
not ( n4085 , n4084 );
xor ( n4086 , n3875 , n3964 );
and ( n4087 , n4086 , n3777 );
buf ( n4088 , n177 );
and ( n4089 , n4088 , n3762 );
buf ( n4090 , n113 );
and ( n4091 , n4090 , n3765 );
buf ( n4092 , n145 );
and ( n4093 , n4092 , n3768 );
or ( n4094 , n4087 , n4089 , n4091 , n4093 );
not ( n4095 , n4094 );
xor ( n4096 , n3880 , n3963 );
and ( n4097 , n4096 , n3777 );
buf ( n4098 , n176 );
and ( n4099 , n4098 , n3762 );
buf ( n4100 , n112 );
and ( n4101 , n4100 , n3765 );
buf ( n4102 , n144 );
and ( n4103 , n4102 , n3768 );
or ( n4104 , n4097 , n4099 , n4101 , n4103 );
not ( n4105 , n4104 );
xor ( n4106 , n3885 , n3962 );
and ( n4107 , n4106 , n3777 );
buf ( n4108 , n175 );
and ( n4109 , n4108 , n3762 );
buf ( n4110 , n111 );
and ( n4111 , n4110 , n3765 );
buf ( n4112 , n143 );
and ( n4113 , n4112 , n3768 );
or ( n4114 , n4107 , n4109 , n4111 , n4113 );
not ( n4115 , n4114 );
xor ( n4116 , n3890 , n3961 );
and ( n4117 , n4116 , n3777 );
buf ( n4118 , n174 );
and ( n4119 , n4118 , n3762 );
buf ( n4120 , n110 );
and ( n4121 , n4120 , n3765 );
buf ( n4122 , n142 );
and ( n4123 , n4122 , n3768 );
or ( n4124 , n4117 , n4119 , n4121 , n4123 );
not ( n4125 , n4124 );
xor ( n4126 , n3895 , n3960 );
and ( n4127 , n4126 , n3777 );
buf ( n4128 , n173 );
and ( n4129 , n4128 , n3762 );
buf ( n4130 , n109 );
and ( n4131 , n4130 , n3765 );
buf ( n4132 , n141 );
and ( n4133 , n4132 , n3768 );
or ( n4134 , n4127 , n4129 , n4131 , n4133 );
not ( n4135 , n4134 );
xor ( n4136 , n3900 , n3959 );
and ( n4137 , n4136 , n3777 );
buf ( n4138 , n172 );
and ( n4139 , n4138 , n3762 );
buf ( n4140 , n108 );
and ( n4141 , n4140 , n3765 );
buf ( n4142 , n140 );
and ( n4143 , n4142 , n3768 );
or ( n4144 , n4137 , n4139 , n4141 , n4143 );
not ( n4145 , n4144 );
xor ( n4146 , n3905 , n3958 );
and ( n4147 , n4146 , n3777 );
buf ( n4148 , n171 );
and ( n4149 , n4148 , n3762 );
buf ( n4150 , n107 );
and ( n4151 , n4150 , n3765 );
buf ( n4152 , n139 );
and ( n4153 , n4152 , n3768 );
or ( n4154 , n4147 , n4149 , n4151 , n4153 );
not ( n4155 , n4154 );
xor ( n4156 , n3910 , n3957 );
and ( n4157 , n4156 , n3777 );
buf ( n4158 , n170 );
and ( n4159 , n4158 , n3762 );
buf ( n4160 , n106 );
and ( n4161 , n4160 , n3765 );
buf ( n4162 , n138 );
and ( n4163 , n4162 , n3768 );
or ( n4164 , n4157 , n4159 , n4161 , n4163 );
not ( n4165 , n4164 );
xor ( n4166 , n3915 , n3956 );
and ( n4167 , n4166 , n3777 );
buf ( n4168 , n169 );
and ( n4169 , n4168 , n3762 );
buf ( n4170 , n105 );
and ( n4171 , n4170 , n3765 );
buf ( n4172 , n137 );
and ( n4173 , n4172 , n3768 );
or ( n4174 , n4167 , n4169 , n4171 , n4173 );
not ( n4175 , n4174 );
xor ( n4176 , n3920 , n3955 );
and ( n4177 , n4176 , n3777 );
buf ( n4178 , n168 );
and ( n4179 , n4178 , n3762 );
buf ( n4180 , n104 );
and ( n4181 , n4180 , n3765 );
buf ( n4182 , n136 );
and ( n4183 , n4182 , n3768 );
or ( n4184 , n4177 , n4179 , n4181 , n4183 );
not ( n4185 , n4184 );
xor ( n4186 , n3925 , n3954 );
and ( n4187 , n4186 , n3777 );
buf ( n4188 , n167 );
and ( n4189 , n4188 , n3762 );
buf ( n4190 , n103 );
and ( n4191 , n4190 , n3765 );
buf ( n4192 , n135 );
and ( n4193 , n4192 , n3768 );
or ( n4194 , n4187 , n4189 , n4191 , n4193 );
not ( n4195 , n4194 );
xor ( n4196 , n3930 , n3953 );
and ( n4197 , n4196 , n3777 );
buf ( n4198 , n166 );
and ( n4199 , n4198 , n3762 );
buf ( n4200 , n102 );
and ( n4201 , n4200 , n3765 );
buf ( n4202 , n134 );
and ( n4203 , n4202 , n3768 );
or ( n4204 , n4197 , n4199 , n4201 , n4203 );
not ( n4205 , n4204 );
xor ( n4206 , n3935 , n3952 );
and ( n4207 , n4206 , n3777 );
buf ( n4208 , n165 );
and ( n4209 , n4208 , n3762 );
buf ( n4210 , n101 );
and ( n4211 , n4210 , n3765 );
buf ( n4212 , n133 );
and ( n4213 , n4212 , n3768 );
or ( n4214 , n4207 , n4209 , n4211 , n4213 );
not ( n4215 , n4214 );
xor ( n4216 , n3940 , n3951 );
and ( n4217 , n4216 , n3777 );
buf ( n4218 , n164 );
and ( n4219 , n4218 , n3762 );
buf ( n4220 , n100 );
and ( n4221 , n4220 , n3765 );
buf ( n4222 , n132 );
and ( n4223 , n4222 , n3768 );
or ( n4224 , n4217 , n4219 , n4221 , n4223 );
not ( n4225 , n4224 );
xor ( n4226 , n3945 , n3950 );
and ( n4227 , n4226 , n3777 );
buf ( n4228 , n163 );
and ( n4229 , n4228 , n3762 );
buf ( n4230 , n99 );
and ( n4231 , n4230 , n3765 );
buf ( n4232 , n131 );
and ( n4233 , n4232 , n3768 );
or ( n4234 , n4227 , n4229 , n4231 , n4233 );
not ( n4235 , n4234 );
not ( n4236 , n3950 );
and ( n4237 , n4236 , n3777 );
buf ( n4238 , n162 );
and ( n4239 , n4238 , n3762 );
buf ( n4240 , n98 );
and ( n4241 , n4240 , n3765 );
buf ( n4242 , n130 );
and ( n4243 , n4242 , n3768 );
or ( n4244 , n4237 , n4239 , n4241 , n4243 );
not ( n4245 , n4244 );
buf ( n4246 , n68 );
buf ( n4247 , n4246 );
not ( n4248 , n4247 );
not ( n4249 , n4248 );
buf ( n4250 , n4249 );
and ( n4251 , n4250 , n3777 );
buf ( n4252 , n161 );
and ( n4253 , n4252 , n3762 );
buf ( n4254 , n97 );
and ( n4255 , n4254 , n3765 );
buf ( n4256 , n129 );
and ( n4257 , n4256 , n3768 );
or ( n4258 , n4251 , n4253 , n4255 , n4257 );
not ( n4259 , n4258 );
and ( n4260 , n3787 , n3796 );
and ( n4261 , n4259 , n4260 );
and ( n4262 , n4245 , n4261 );
and ( n4263 , n4235 , n4262 );
and ( n4264 , n4225 , n4263 );
and ( n4265 , n4215 , n4264 );
and ( n4266 , n4205 , n4265 );
and ( n4267 , n4195 , n4266 );
and ( n4268 , n4185 , n4267 );
and ( n4269 , n4175 , n4268 );
and ( n4270 , n4165 , n4269 );
and ( n4271 , n4155 , n4270 );
and ( n4272 , n4145 , n4271 );
and ( n4273 , n4135 , n4272 );
and ( n4274 , n4125 , n4273 );
and ( n4275 , n4115 , n4274 );
and ( n4276 , n4105 , n4275 );
and ( n4277 , n4095 , n4276 );
and ( n4278 , n4085 , n4277 );
and ( n4279 , n4075 , n4278 );
and ( n4280 , n4065 , n4279 );
and ( n4281 , n4055 , n4280 );
and ( n4282 , n4045 , n4281 );
and ( n4283 , n4035 , n4282 );
and ( n4284 , n4025 , n4283 );
and ( n4285 , n4015 , n4284 );
and ( n4286 , n4005 , n4285 );
and ( n4287 , n3995 , n4286 );
and ( n4288 , n3985 , n4287 );
and ( n4289 , n3820 , n4288 );
xor ( n4290 , n3812 , n4289 );
and ( n4291 , n4290 , n3809 );
or ( n4292 , n3811 , n4291 );
not ( n4293 , n4292 );
not ( n4294 , n4293 );
not ( n4295 , n4294 );
not ( n4296 , n3770 );
and ( n4297 , n4296 , n3819 );
xor ( n4298 , n3820 , n4288 );
and ( n4299 , n4298 , n3770 );
or ( n4300 , n4297 , n4299 );
not ( n4301 , n4300 );
not ( n4302 , n4301 );
not ( n4303 , n4302 );
not ( n4304 , n3770 );
and ( n4305 , n4304 , n3984 );
xor ( n4306 , n3985 , n4287 );
and ( n4307 , n4306 , n3770 );
or ( n4308 , n4305 , n4307 );
not ( n4309 , n4308 );
not ( n4310 , n4309 );
not ( n4311 , n4310 );
not ( n4312 , n3770 );
and ( n4313 , n4312 , n3994 );
xor ( n4314 , n3995 , n4286 );
and ( n4315 , n4314 , n3770 );
or ( n4316 , n4313 , n4315 );
not ( n4317 , n4316 );
not ( n4318 , n4317 );
not ( n4319 , n4318 );
not ( n4320 , n3770 );
and ( n4321 , n4320 , n4004 );
xor ( n4322 , n4005 , n4285 );
and ( n4323 , n4322 , n3770 );
or ( n4324 , n4321 , n4323 );
not ( n4325 , n4324 );
not ( n4326 , n4325 );
not ( n4327 , n4326 );
not ( n4328 , n3770 );
and ( n4329 , n4328 , n4014 );
xor ( n4330 , n4015 , n4284 );
and ( n4331 , n4330 , n3770 );
or ( n4332 , n4329 , n4331 );
not ( n4333 , n4332 );
not ( n4334 , n4333 );
not ( n4335 , n4334 );
not ( n4336 , n3770 );
and ( n4337 , n4336 , n4024 );
xor ( n4338 , n4025 , n4283 );
and ( n4339 , n4338 , n3770 );
or ( n4340 , n4337 , n4339 );
not ( n4341 , n4340 );
not ( n4342 , n4341 );
not ( n4343 , n4342 );
not ( n4344 , n3770 );
and ( n4345 , n4344 , n4034 );
xor ( n4346 , n4035 , n4282 );
and ( n4347 , n4346 , n3770 );
or ( n4348 , n4345 , n4347 );
not ( n4349 , n4348 );
not ( n4350 , n4349 );
not ( n4351 , n4350 );
not ( n4352 , n3770 );
and ( n4353 , n4352 , n4044 );
xor ( n4354 , n4045 , n4281 );
and ( n4355 , n4354 , n3770 );
or ( n4356 , n4353 , n4355 );
not ( n4357 , n4356 );
not ( n4358 , n4357 );
not ( n4359 , n4358 );
not ( n4360 , n3770 );
and ( n4361 , n4360 , n4054 );
xor ( n4362 , n4055 , n4280 );
and ( n4363 , n4362 , n3770 );
or ( n4364 , n4361 , n4363 );
not ( n4365 , n4364 );
not ( n4366 , n4365 );
not ( n4367 , n4366 );
not ( n4368 , n3770 );
and ( n4369 , n4368 , n4064 );
xor ( n4370 , n4065 , n4279 );
and ( n4371 , n4370 , n3770 );
or ( n4372 , n4369 , n4371 );
not ( n4373 , n4372 );
not ( n4374 , n4373 );
not ( n4375 , n4374 );
not ( n4376 , n3770 );
and ( n4377 , n4376 , n4074 );
xor ( n4378 , n4075 , n4278 );
and ( n4379 , n4378 , n3770 );
or ( n4380 , n4377 , n4379 );
not ( n4381 , n4380 );
not ( n4382 , n4381 );
not ( n4383 , n4382 );
not ( n4384 , n3770 );
and ( n4385 , n4384 , n4084 );
xor ( n4386 , n4085 , n4277 );
and ( n4387 , n4386 , n3770 );
or ( n4388 , n4385 , n4387 );
not ( n4389 , n4388 );
not ( n4390 , n4389 );
not ( n4391 , n4390 );
not ( n4392 , n3770 );
and ( n4393 , n4392 , n4094 );
xor ( n4394 , n4095 , n4276 );
and ( n4395 , n4394 , n3770 );
or ( n4396 , n4393 , n4395 );
not ( n4397 , n4396 );
not ( n4398 , n4397 );
not ( n4399 , n4398 );
not ( n4400 , n3770 );
and ( n4401 , n4400 , n4104 );
xor ( n4402 , n4105 , n4275 );
and ( n4403 , n4402 , n3770 );
or ( n4404 , n4401 , n4403 );
not ( n4405 , n4404 );
not ( n4406 , n4405 );
not ( n4407 , n4406 );
not ( n4408 , n3770 );
and ( n4409 , n4408 , n4114 );
xor ( n4410 , n4115 , n4274 );
and ( n4411 , n4410 , n3770 );
or ( n4412 , n4409 , n4411 );
not ( n4413 , n4412 );
not ( n4414 , n4413 );
not ( n4415 , n4414 );
not ( n4416 , n3770 );
and ( n4417 , n4416 , n4124 );
xor ( n4418 , n4125 , n4273 );
and ( n4419 , n4418 , n3770 );
or ( n4420 , n4417 , n4419 );
not ( n4421 , n4420 );
not ( n4422 , n4421 );
not ( n4423 , n4422 );
not ( n4424 , n3770 );
and ( n4425 , n4424 , n4134 );
xor ( n4426 , n4135 , n4272 );
and ( n4427 , n4426 , n3770 );
or ( n4428 , n4425 , n4427 );
not ( n4429 , n4428 );
not ( n4430 , n4429 );
not ( n4431 , n4430 );
not ( n4432 , n3770 );
and ( n4433 , n4432 , n4144 );
xor ( n4434 , n4145 , n4271 );
and ( n4435 , n4434 , n3770 );
or ( n4436 , n4433 , n4435 );
not ( n4437 , n4436 );
not ( n4438 , n4437 );
not ( n4439 , n4438 );
not ( n4440 , n3770 );
and ( n4441 , n4440 , n4154 );
xor ( n4442 , n4155 , n4270 );
and ( n4443 , n4442 , n3770 );
or ( n4444 , n4441 , n4443 );
not ( n4445 , n4444 );
not ( n4446 , n4445 );
not ( n4447 , n4446 );
not ( n4448 , n3770 );
and ( n4449 , n4448 , n4164 );
xor ( n4450 , n4165 , n4269 );
and ( n4451 , n4450 , n3770 );
or ( n4452 , n4449 , n4451 );
not ( n4453 , n4452 );
not ( n4454 , n4453 );
not ( n4455 , n4454 );
not ( n4456 , n3770 );
and ( n4457 , n4456 , n4174 );
xor ( n4458 , n4175 , n4268 );
and ( n4459 , n4458 , n3770 );
or ( n4460 , n4457 , n4459 );
not ( n4461 , n4460 );
buf ( n4462 , n4461 );
buf ( n4463 , n4462 );
not ( n4464 , n4463 );
not ( n4465 , n4464 );
not ( n4466 , n3770 );
and ( n4467 , n4466 , n4184 );
xor ( n4468 , n4185 , n4267 );
and ( n4469 , n4468 , n3770 );
or ( n4470 , n4467 , n4469 );
not ( n4471 , n4470 );
buf ( n4472 , n4471 );
buf ( n4473 , n4472 );
not ( n4474 , n4473 );
not ( n4475 , n4474 );
not ( n4476 , n3770 );
and ( n4477 , n4476 , n4194 );
xor ( n4478 , n4195 , n4266 );
and ( n4479 , n4478 , n3770 );
or ( n4480 , n4477 , n4479 );
not ( n4481 , n4480 );
buf ( n4482 , n4481 );
buf ( n4483 , n4482 );
not ( n4484 , n4483 );
not ( n4485 , n4484 );
not ( n4486 , n3770 );
and ( n4487 , n4486 , n4204 );
xor ( n4488 , n4205 , n4265 );
and ( n4489 , n4488 , n3770 );
or ( n4490 , n4487 , n4489 );
not ( n4491 , n4490 );
buf ( n4492 , n4491 );
buf ( n4493 , n4492 );
not ( n4494 , n4493 );
not ( n4495 , n4494 );
not ( n4496 , n3770 );
and ( n4497 , n4496 , n4214 );
xor ( n4498 , n4215 , n4264 );
and ( n4499 , n4498 , n3770 );
or ( n4500 , n4497 , n4499 );
not ( n4501 , n4500 );
buf ( n4502 , n4501 );
buf ( n4503 , n4502 );
not ( n4504 , n4503 );
not ( n4505 , n4504 );
not ( n4506 , n3770 );
and ( n4507 , n4506 , n4224 );
xor ( n4508 , n4225 , n4263 );
and ( n4509 , n4508 , n3770 );
or ( n4510 , n4507 , n4509 );
not ( n4511 , n4510 );
buf ( n4512 , n4511 );
buf ( n4513 , n4512 );
not ( n4514 , n4513 );
not ( n4515 , n4514 );
not ( n4516 , n3770 );
and ( n4517 , n4516 , n4234 );
xor ( n4518 , n4235 , n4262 );
and ( n4519 , n4518 , n3770 );
or ( n4520 , n4517 , n4519 );
not ( n4521 , n4520 );
buf ( n4522 , n4521 );
buf ( n4523 , n4522 );
not ( n4524 , n4523 );
not ( n4525 , n4524 );
not ( n4526 , n3770 );
and ( n4527 , n4526 , n4244 );
xor ( n4528 , n4245 , n4261 );
and ( n4529 , n4528 , n3770 );
or ( n4530 , n4527 , n4529 );
not ( n4531 , n4530 );
buf ( n4532 , n4531 );
buf ( n4533 , n4532 );
not ( n4534 , n4533 );
not ( n4535 , n4534 );
not ( n4536 , n3770 );
and ( n4537 , n4536 , n4258 );
xor ( n4538 , n4259 , n4260 );
and ( n4539 , n4538 , n3770 );
or ( n4540 , n4537 , n4539 );
not ( n4541 , n4540 );
buf ( n4542 , n4541 );
buf ( n4543 , n4542 );
not ( n4544 , n4543 );
not ( n4545 , n4544 );
not ( n4546 , n3803 );
and ( n4547 , n4545 , n4546 );
and ( n4548 , n4535 , n4547 );
and ( n4549 , n4525 , n4548 );
and ( n4550 , n4515 , n4549 );
and ( n4551 , n4505 , n4550 );
and ( n4552 , n4495 , n4551 );
and ( n4553 , n4485 , n4552 );
and ( n4554 , n4475 , n4553 );
and ( n4555 , n4465 , n4554 );
and ( n4556 , n4455 , n4555 );
and ( n4557 , n4447 , n4556 );
and ( n4558 , n4439 , n4557 );
and ( n4559 , n4431 , n4558 );
and ( n4560 , n4423 , n4559 );
and ( n4561 , n4415 , n4560 );
and ( n4562 , n4407 , n4561 );
and ( n4563 , n4399 , n4562 );
and ( n4564 , n4391 , n4563 );
and ( n4565 , n4383 , n4564 );
and ( n4566 , n4375 , n4565 );
and ( n4567 , n4367 , n4566 );
and ( n4568 , n4359 , n4567 );
and ( n4569 , n4351 , n4568 );
and ( n4570 , n4343 , n4569 );
and ( n4571 , n4335 , n4570 );
and ( n4572 , n4327 , n4571 );
and ( n4573 , n4319 , n4572 );
and ( n4574 , n4311 , n4573 );
and ( n4575 , n4303 , n4574 );
and ( n4576 , n4295 , n4575 );
not ( n4577 , n4576 );
and ( n4578 , n4577 , n3770 );
or ( n4579 , n3808 , n4578 );
not ( n4580 , n4579 );
not ( n4581 , n3770 );
and ( n4582 , n4581 , n4544 );
xor ( n4583 , n4545 , n4546 );
and ( n4584 , n4583 , n3770 );
or ( n4585 , n4582 , n4584 );
and ( n4586 , n4580 , n4585 );
not ( n4587 , n4585 );
not ( n4588 , n3803 );
xor ( n4589 , n4587 , n4588 );
and ( n4590 , n4589 , n4579 );
or ( n4591 , n4586 , n4590 );
not ( n4592 , n4591 );
not ( n4593 , n4592 );
or ( n4594 , n3806 , n4593 );
not ( n4595 , n4579 );
not ( n4596 , n3770 );
and ( n4597 , n4596 , n4534 );
xor ( n4598 , n4535 , n4547 );
and ( n4599 , n4598 , n3770 );
or ( n4600 , n4597 , n4599 );
and ( n4601 , n4595 , n4600 );
not ( n4602 , n4600 );
and ( n4603 , n4587 , n4588 );
xor ( n4604 , n4602 , n4603 );
and ( n4605 , n4604 , n4579 );
or ( n4606 , n4601 , n4605 );
not ( n4607 , n4606 );
not ( n4608 , n4607 );
or ( n4609 , n4594 , n4608 );
not ( n4610 , n4579 );
not ( n4611 , n3770 );
and ( n4612 , n4611 , n4524 );
xor ( n4613 , n4525 , n4548 );
and ( n4614 , n4613 , n3770 );
or ( n4615 , n4612 , n4614 );
and ( n4616 , n4610 , n4615 );
not ( n4617 , n4615 );
and ( n4618 , n4602 , n4603 );
xor ( n4619 , n4617 , n4618 );
and ( n4620 , n4619 , n4579 );
or ( n4621 , n4616 , n4620 );
not ( n4622 , n4621 );
not ( n4623 , n4622 );
or ( n4624 , n4609 , n4623 );
not ( n4625 , n4579 );
not ( n4626 , n3770 );
and ( n4627 , n4626 , n4514 );
xor ( n4628 , n4515 , n4549 );
and ( n4629 , n4628 , n3770 );
or ( n4630 , n4627 , n4629 );
and ( n4631 , n4625 , n4630 );
not ( n4632 , n4630 );
and ( n4633 , n4617 , n4618 );
xor ( n4634 , n4632 , n4633 );
and ( n4635 , n4634 , n4579 );
or ( n4636 , n4631 , n4635 );
not ( n4637 , n4636 );
not ( n4638 , n4637 );
or ( n4639 , n4624 , n4638 );
not ( n4640 , n4579 );
not ( n4641 , n3770 );
and ( n4642 , n4641 , n4504 );
xor ( n4643 , n4505 , n4550 );
and ( n4644 , n4643 , n3770 );
or ( n4645 , n4642 , n4644 );
and ( n4646 , n4640 , n4645 );
not ( n4647 , n4645 );
and ( n4648 , n4632 , n4633 );
xor ( n4649 , n4647 , n4648 );
and ( n4650 , n4649 , n4579 );
or ( n4651 , n4646 , n4650 );
not ( n4652 , n4651 );
not ( n4653 , n4652 );
or ( n4654 , n4639 , n4653 );
not ( n4655 , n4579 );
not ( n4656 , n3770 );
and ( n4657 , n4656 , n4494 );
xor ( n4658 , n4495 , n4551 );
and ( n4659 , n4658 , n3770 );
or ( n4660 , n4657 , n4659 );
and ( n4661 , n4655 , n4660 );
not ( n4662 , n4660 );
and ( n4663 , n4647 , n4648 );
xor ( n4664 , n4662 , n4663 );
and ( n4665 , n4664 , n4579 );
or ( n4666 , n4661 , n4665 );
not ( n4667 , n4666 );
not ( n4668 , n4667 );
or ( n4669 , n4654 , n4668 );
not ( n4670 , n4579 );
not ( n4671 , n3770 );
and ( n4672 , n4671 , n4484 );
xor ( n4673 , n4485 , n4552 );
and ( n4674 , n4673 , n3770 );
or ( n4675 , n4672 , n4674 );
and ( n4676 , n4670 , n4675 );
not ( n4677 , n4675 );
and ( n4678 , n4662 , n4663 );
xor ( n4679 , n4677 , n4678 );
and ( n4680 , n4679 , n4579 );
or ( n4681 , n4676 , n4680 );
not ( n4682 , n4681 );
not ( n4683 , n4682 );
or ( n4684 , n4669 , n4683 );
not ( n4685 , n4579 );
not ( n4686 , n3770 );
and ( n4687 , n4686 , n4474 );
xor ( n4688 , n4475 , n4553 );
and ( n4689 , n4688 , n3770 );
or ( n4690 , n4687 , n4689 );
and ( n4691 , n4685 , n4690 );
not ( n4692 , n4690 );
and ( n4693 , n4677 , n4678 );
xor ( n4694 , n4692 , n4693 );
and ( n4695 , n4694 , n4579 );
or ( n4696 , n4691 , n4695 );
not ( n4697 , n4696 );
not ( n4698 , n4697 );
or ( n4699 , n4684 , n4698 );
not ( n4700 , n4579 );
not ( n4701 , n3770 );
and ( n4702 , n4701 , n4464 );
xor ( n4703 , n4465 , n4554 );
and ( n4704 , n4703 , n3770 );
or ( n4705 , n4702 , n4704 );
and ( n4706 , n4700 , n4705 );
not ( n4707 , n4705 );
and ( n4708 , n4692 , n4693 );
xor ( n4709 , n4707 , n4708 );
and ( n4710 , n4709 , n4579 );
or ( n4711 , n4706 , n4710 );
not ( n4712 , n4711 );
not ( n4713 , n4712 );
or ( n4714 , n4699 , n4713 );
not ( n4715 , n4579 );
not ( n4716 , n3770 );
and ( n4717 , n4716 , n4454 );
xor ( n4718 , n4455 , n4555 );
and ( n4719 , n4718 , n3770 );
or ( n4720 , n4717 , n4719 );
and ( n4721 , n4715 , n4720 );
not ( n4722 , n4720 );
and ( n4723 , n4707 , n4708 );
xor ( n4724 , n4722 , n4723 );
and ( n4725 , n4724 , n4579 );
or ( n4726 , n4721 , n4725 );
not ( n4727 , n4726 );
not ( n4728 , n4727 );
or ( n4729 , n4714 , n4728 );
not ( n4730 , n4579 );
not ( n4731 , n3770 );
and ( n4732 , n4731 , n4446 );
xor ( n4733 , n4447 , n4556 );
and ( n4734 , n4733 , n3770 );
or ( n4735 , n4732 , n4734 );
and ( n4736 , n4730 , n4735 );
not ( n4737 , n4735 );
and ( n4738 , n4722 , n4723 );
xor ( n4739 , n4737 , n4738 );
and ( n4740 , n4739 , n4579 );
or ( n4741 , n4736 , n4740 );
not ( n4742 , n4741 );
not ( n4743 , n4742 );
or ( n4744 , n4729 , n4743 );
not ( n4745 , n4579 );
not ( n4746 , n3770 );
and ( n4747 , n4746 , n4438 );
xor ( n4748 , n4439 , n4557 );
and ( n4749 , n4748 , n3770 );
or ( n4750 , n4747 , n4749 );
and ( n4751 , n4745 , n4750 );
not ( n4752 , n4750 );
and ( n4753 , n4737 , n4738 );
xor ( n4754 , n4752 , n4753 );
and ( n4755 , n4754 , n4579 );
or ( n4756 , n4751 , n4755 );
not ( n4757 , n4756 );
not ( n4758 , n4757 );
or ( n4759 , n4744 , n4758 );
not ( n4760 , n4579 );
not ( n4761 , n3770 );
and ( n4762 , n4761 , n4430 );
xor ( n4763 , n4431 , n4558 );
and ( n4764 , n4763 , n3770 );
or ( n4765 , n4762 , n4764 );
and ( n4766 , n4760 , n4765 );
not ( n4767 , n4765 );
and ( n4768 , n4752 , n4753 );
xor ( n4769 , n4767 , n4768 );
and ( n4770 , n4769 , n4579 );
or ( n4771 , n4766 , n4770 );
not ( n4772 , n4771 );
not ( n4773 , n4772 );
or ( n4774 , n4759 , n4773 );
not ( n4775 , n4579 );
not ( n4776 , n3770 );
and ( n4777 , n4776 , n4422 );
xor ( n4778 , n4423 , n4559 );
and ( n4779 , n4778 , n3770 );
or ( n4780 , n4777 , n4779 );
and ( n4781 , n4775 , n4780 );
not ( n4782 , n4780 );
and ( n4783 , n4767 , n4768 );
xor ( n4784 , n4782 , n4783 );
and ( n4785 , n4784 , n4579 );
or ( n4786 , n4781 , n4785 );
not ( n4787 , n4786 );
not ( n4788 , n4787 );
or ( n4789 , n4774 , n4788 );
not ( n4790 , n4579 );
not ( n4791 , n3770 );
and ( n4792 , n4791 , n4414 );
xor ( n4793 , n4415 , n4560 );
and ( n4794 , n4793 , n3770 );
or ( n4795 , n4792 , n4794 );
and ( n4796 , n4790 , n4795 );
not ( n4797 , n4795 );
and ( n4798 , n4782 , n4783 );
xor ( n4799 , n4797 , n4798 );
and ( n4800 , n4799 , n4579 );
or ( n4801 , n4796 , n4800 );
not ( n4802 , n4801 );
not ( n4803 , n4802 );
or ( n4804 , n4789 , n4803 );
not ( n4805 , n4579 );
not ( n4806 , n3770 );
and ( n4807 , n4806 , n4406 );
xor ( n4808 , n4407 , n4561 );
and ( n4809 , n4808 , n3770 );
or ( n4810 , n4807 , n4809 );
and ( n4811 , n4805 , n4810 );
not ( n4812 , n4810 );
and ( n4813 , n4797 , n4798 );
xor ( n4814 , n4812 , n4813 );
and ( n4815 , n4814 , n4579 );
or ( n4816 , n4811 , n4815 );
not ( n4817 , n4816 );
not ( n4818 , n4817 );
or ( n4819 , n4804 , n4818 );
not ( n4820 , n4579 );
not ( n4821 , n3770 );
and ( n4822 , n4821 , n4398 );
xor ( n4823 , n4399 , n4562 );
and ( n4824 , n4823 , n3770 );
or ( n4825 , n4822 , n4824 );
and ( n4826 , n4820 , n4825 );
not ( n4827 , n4825 );
and ( n4828 , n4812 , n4813 );
xor ( n4829 , n4827 , n4828 );
and ( n4830 , n4829 , n4579 );
or ( n4831 , n4826 , n4830 );
not ( n4832 , n4831 );
not ( n4833 , n4832 );
or ( n4834 , n4819 , n4833 );
not ( n4835 , n4579 );
not ( n4836 , n3770 );
and ( n4837 , n4836 , n4390 );
xor ( n4838 , n4391 , n4563 );
and ( n4839 , n4838 , n3770 );
or ( n4840 , n4837 , n4839 );
and ( n4841 , n4835 , n4840 );
not ( n4842 , n4840 );
and ( n4843 , n4827 , n4828 );
xor ( n4844 , n4842 , n4843 );
and ( n4845 , n4844 , n4579 );
or ( n4846 , n4841 , n4845 );
not ( n4847 , n4846 );
not ( n4848 , n4847 );
or ( n4849 , n4834 , n4848 );
not ( n4850 , n4579 );
not ( n4851 , n3770 );
and ( n4852 , n4851 , n4382 );
xor ( n4853 , n4383 , n4564 );
and ( n4854 , n4853 , n3770 );
or ( n4855 , n4852 , n4854 );
and ( n4856 , n4850 , n4855 );
not ( n4857 , n4855 );
and ( n4858 , n4842 , n4843 );
xor ( n4859 , n4857 , n4858 );
and ( n4860 , n4859 , n4579 );
or ( n4861 , n4856 , n4860 );
not ( n4862 , n4861 );
not ( n4863 , n4862 );
or ( n4864 , n4849 , n4863 );
not ( n4865 , n4579 );
not ( n4866 , n3770 );
and ( n4867 , n4866 , n4374 );
xor ( n4868 , n4375 , n4565 );
and ( n4869 , n4868 , n3770 );
or ( n4870 , n4867 , n4869 );
and ( n4871 , n4865 , n4870 );
not ( n4872 , n4870 );
and ( n4873 , n4857 , n4858 );
xor ( n4874 , n4872 , n4873 );
and ( n4875 , n4874 , n4579 );
or ( n4876 , n4871 , n4875 );
not ( n4877 , n4876 );
not ( n4878 , n4877 );
or ( n4879 , n4864 , n4878 );
not ( n4880 , n4579 );
not ( n4881 , n3770 );
and ( n4882 , n4881 , n4366 );
xor ( n4883 , n4367 , n4566 );
and ( n4884 , n4883 , n3770 );
or ( n4885 , n4882 , n4884 );
and ( n4886 , n4880 , n4885 );
not ( n4887 , n4885 );
and ( n4888 , n4872 , n4873 );
xor ( n4889 , n4887 , n4888 );
and ( n4890 , n4889 , n4579 );
or ( n4891 , n4886 , n4890 );
not ( n4892 , n4891 );
not ( n4893 , n4892 );
or ( n4894 , n4879 , n4893 );
not ( n4895 , n4579 );
not ( n4896 , n3770 );
and ( n4897 , n4896 , n4358 );
xor ( n4898 , n4359 , n4567 );
and ( n4899 , n4898 , n3770 );
or ( n4900 , n4897 , n4899 );
and ( n4901 , n4895 , n4900 );
not ( n4902 , n4900 );
and ( n4903 , n4887 , n4888 );
xor ( n4904 , n4902 , n4903 );
and ( n4905 , n4904 , n4579 );
or ( n4906 , n4901 , n4905 );
not ( n4907 , n4906 );
not ( n4908 , n4907 );
or ( n4909 , n4894 , n4908 );
not ( n4910 , n4579 );
not ( n4911 , n3770 );
and ( n4912 , n4911 , n4350 );
xor ( n4913 , n4351 , n4568 );
and ( n4914 , n4913 , n3770 );
or ( n4915 , n4912 , n4914 );
and ( n4916 , n4910 , n4915 );
not ( n4917 , n4915 );
and ( n4918 , n4902 , n4903 );
xor ( n4919 , n4917 , n4918 );
and ( n4920 , n4919 , n4579 );
or ( n4921 , n4916 , n4920 );
not ( n4922 , n4921 );
not ( n4923 , n4922 );
or ( n4924 , n4909 , n4923 );
not ( n4925 , n4579 );
not ( n4926 , n3770 );
and ( n4927 , n4926 , n4342 );
xor ( n4928 , n4343 , n4569 );
and ( n4929 , n4928 , n3770 );
or ( n4930 , n4927 , n4929 );
and ( n4931 , n4925 , n4930 );
not ( n4932 , n4930 );
and ( n4933 , n4917 , n4918 );
xor ( n4934 , n4932 , n4933 );
and ( n4935 , n4934 , n4579 );
or ( n4936 , n4931 , n4935 );
not ( n4937 , n4936 );
not ( n4938 , n4937 );
or ( n4939 , n4924 , n4938 );
not ( n4940 , n4579 );
not ( n4941 , n3770 );
and ( n4942 , n4941 , n4334 );
xor ( n4943 , n4335 , n4570 );
and ( n4944 , n4943 , n3770 );
or ( n4945 , n4942 , n4944 );
and ( n4946 , n4940 , n4945 );
not ( n4947 , n4945 );
and ( n4948 , n4932 , n4933 );
xor ( n4949 , n4947 , n4948 );
and ( n4950 , n4949 , n4579 );
or ( n4951 , n4946 , n4950 );
not ( n4952 , n4951 );
not ( n4953 , n4952 );
or ( n4954 , n4939 , n4953 );
not ( n4955 , n4579 );
not ( n4956 , n3770 );
and ( n4957 , n4956 , n4326 );
xor ( n4958 , n4327 , n4571 );
and ( n4959 , n4958 , n3770 );
or ( n4960 , n4957 , n4959 );
and ( n4961 , n4955 , n4960 );
not ( n4962 , n4960 );
and ( n4963 , n4947 , n4948 );
xor ( n4964 , n4962 , n4963 );
and ( n4965 , n4964 , n4579 );
or ( n4966 , n4961 , n4965 );
not ( n4967 , n4966 );
not ( n4968 , n4967 );
or ( n4969 , n4954 , n4968 );
not ( n4970 , n4579 );
not ( n4971 , n3770 );
and ( n4972 , n4971 , n4318 );
xor ( n4973 , n4319 , n4572 );
and ( n4974 , n4973 , n3770 );
or ( n4975 , n4972 , n4974 );
and ( n4976 , n4970 , n4975 );
not ( n4977 , n4975 );
and ( n4978 , n4962 , n4963 );
xor ( n4979 , n4977 , n4978 );
and ( n4980 , n4979 , n4579 );
or ( n4981 , n4976 , n4980 );
not ( n4982 , n4981 );
not ( n4983 , n4982 );
or ( n4984 , n4969 , n4983 );
not ( n4985 , n4579 );
not ( n4986 , n3770 );
and ( n4987 , n4986 , n4310 );
xor ( n4988 , n4311 , n4573 );
and ( n4989 , n4988 , n3770 );
or ( n4990 , n4987 , n4989 );
and ( n4991 , n4985 , n4990 );
not ( n4992 , n4990 );
and ( n4993 , n4977 , n4978 );
xor ( n4994 , n4992 , n4993 );
and ( n4995 , n4994 , n4579 );
or ( n4996 , n4991 , n4995 );
not ( n4997 , n4996 );
not ( n4998 , n4997 );
or ( n4999 , n4984 , n4998 );
and ( n5000 , n4999 , n4579 );
not ( n5001 , n5000 );
and ( n5002 , n5001 , n3806 );
xor ( n5003 , n3806 , n4579 );
xor ( n5004 , n5003 , n4579 );
and ( n5005 , n5004 , n5000 );
or ( n5006 , n5002 , n5005 );
and ( n5007 , n5006 , n3290 );
or ( n5008 , n3804 , n5007 );
not ( n5009 , n2899 );
and ( n5010 , n5009 , n2839 );
not ( n5011 , n2839 );
not ( n5012 , n2824 );
not ( n5013 , n2809 );
not ( n5014 , n2794 );
not ( n5015 , n2779 );
not ( n5016 , n2764 );
not ( n5017 , n2749 );
not ( n5018 , n2734 );
not ( n5019 , n2719 );
not ( n5020 , n2704 );
not ( n5021 , n2689 );
not ( n5022 , n2674 );
not ( n5023 , n2659 );
not ( n5024 , n2644 );
not ( n5025 , n2629 );
not ( n5026 , n2614 );
not ( n5027 , n2599 );
not ( n5028 , n2584 );
not ( n5029 , n2569 );
not ( n5030 , n2554 );
not ( n5031 , n2539 );
not ( n5032 , n2524 );
not ( n5033 , n2509 );
not ( n5034 , n2494 );
not ( n5035 , n2479 );
not ( n5036 , n2464 );
not ( n5037 , n2449 );
not ( n5038 , n2430 );
and ( n5039 , n5037 , n5038 );
and ( n5040 , n5036 , n5039 );
and ( n5041 , n5035 , n5040 );
and ( n5042 , n5034 , n5041 );
and ( n5043 , n5033 , n5042 );
and ( n5044 , n5032 , n5043 );
and ( n5045 , n5031 , n5044 );
and ( n5046 , n5030 , n5045 );
and ( n5047 , n5029 , n5046 );
and ( n5048 , n5028 , n5047 );
and ( n5049 , n5027 , n5048 );
and ( n5050 , n5026 , n5049 );
and ( n5051 , n5025 , n5050 );
and ( n5052 , n5024 , n5051 );
and ( n5053 , n5023 , n5052 );
and ( n5054 , n5022 , n5053 );
and ( n5055 , n5021 , n5054 );
and ( n5056 , n5020 , n5055 );
and ( n5057 , n5019 , n5056 );
and ( n5058 , n5018 , n5057 );
and ( n5059 , n5017 , n5058 );
and ( n5060 , n5016 , n5059 );
and ( n5061 , n5015 , n5060 );
and ( n5062 , n5014 , n5061 );
and ( n5063 , n5013 , n5062 );
and ( n5064 , n5012 , n5063 );
xor ( n5065 , n5011 , n5064 );
and ( n5066 , n5065 , n2899 );
or ( n5067 , n5010 , n5066 );
not ( n5068 , n5067 );
not ( n5069 , n5068 );
not ( n5070 , n5069 );
not ( n5071 , n5070 );
not ( n5072 , n2899 );
and ( n5073 , n5072 , n2424 );
buf ( n5074 , n2899 );
not ( n5075 , n5074 );
and ( n5076 , n5075 , n2899 );
not ( n5077 , n2899 );
not ( n5078 , n2884 );
not ( n5079 , n2869 );
not ( n5080 , n2854 );
and ( n5081 , n5011 , n5064 );
and ( n5082 , n5080 , n5081 );
and ( n5083 , n5079 , n5082 );
and ( n5084 , n5078 , n5083 );
xor ( n5085 , n5077 , n5084 );
and ( n5086 , n5085 , n5074 );
or ( n5087 , n5076 , n5086 );
not ( n5088 , n5087 );
not ( n5089 , n5088 );
not ( n5090 , n5089 );
not ( n5091 , n2899 );
and ( n5092 , n5091 , n2884 );
xor ( n5093 , n5078 , n5083 );
and ( n5094 , n5093 , n2899 );
or ( n5095 , n5092 , n5094 );
not ( n5096 , n5095 );
not ( n5097 , n5096 );
not ( n5098 , n5097 );
not ( n5099 , n2899 );
and ( n5100 , n5099 , n2869 );
xor ( n5101 , n5079 , n5082 );
and ( n5102 , n5101 , n2899 );
or ( n5103 , n5100 , n5102 );
not ( n5104 , n5103 );
not ( n5105 , n5104 );
not ( n5106 , n5105 );
not ( n5107 , n2899 );
and ( n5108 , n5107 , n2854 );
xor ( n5109 , n5080 , n5081 );
and ( n5110 , n5109 , n2899 );
or ( n5111 , n5108 , n5110 );
not ( n5112 , n5111 );
not ( n5113 , n5112 );
not ( n5114 , n5113 );
not ( n5115 , n5069 );
and ( n5116 , n5114 , n5115 );
and ( n5117 , n5106 , n5116 );
and ( n5118 , n5098 , n5117 );
and ( n5119 , n5090 , n5118 );
not ( n5120 , n5119 );
and ( n5121 , n5120 , n2899 );
or ( n5122 , n5073 , n5121 );
not ( n5123 , n5122 );
not ( n5124 , n2899 );
and ( n5125 , n5124 , n5113 );
xor ( n5126 , n5114 , n5115 );
and ( n5127 , n5126 , n2899 );
or ( n5128 , n5125 , n5127 );
and ( n5129 , n5123 , n5128 );
not ( n5130 , n5128 );
not ( n5131 , n5069 );
xor ( n5132 , n5130 , n5131 );
and ( n5133 , n5132 , n5122 );
or ( n5134 , n5129 , n5133 );
not ( n5135 , n5134 );
not ( n5136 , n5135 );
or ( n5137 , n5071 , n5136 );
and ( n5138 , n5137 , n5122 );
not ( n5139 , n5138 );
and ( n5140 , n5139 , n5071 );
xor ( n5141 , n5071 , n5122 );
xor ( n5142 , n5141 , n5122 );
and ( n5143 , n5142 , n5138 );
or ( n5144 , n5140 , n5143 );
not ( n5145 , n5144 );
not ( n5146 , n5138 );
and ( n5147 , n5146 , n5136 );
xor ( n5148 , n5136 , n5122 );
and ( n5149 , n5141 , n5122 );
xor ( n5150 , n5148 , n5149 );
and ( n5151 , n5150 , n5138 );
or ( n5152 , n5147 , n5151 );
nor ( n5153 , n5145 , n5152 );
and ( n5154 , n5008 , n5153 );
nor ( n5155 , n5144 , n5152 );
and ( n5156 , n3803 , n5155 );
or ( n5157 , n2424 , n3633 , n5154 , n5156 );
not ( n5158 , n3304 );
not ( n5159 , n3348 );
buf ( n5160 , n2424 );
buf ( n5161 , n2424 );
buf ( n5162 , n2424 );
buf ( n5163 , n2424 );
buf ( n5164 , n2424 );
buf ( n5165 , n2424 );
buf ( n5166 , n2424 );
buf ( n5167 , n2424 );
buf ( n5168 , n2424 );
buf ( n5169 , n2424 );
buf ( n5170 , n2424 );
buf ( n5171 , n2424 );
buf ( n5172 , n2424 );
buf ( n5173 , n2424 );
buf ( n5174 , n2424 );
buf ( n5175 , n2424 );
buf ( n5176 , n2424 );
buf ( n5177 , n2424 );
buf ( n5178 , n2424 );
buf ( n5179 , n2424 );
buf ( n5180 , n2424 );
buf ( n5181 , n2424 );
buf ( n5182 , n2424 );
buf ( n5183 , n2424 );
buf ( n5184 , n2424 );
buf ( n5185 , n2424 );
buf ( n5186 , n2424 );
buf ( n5187 , n2424 );
buf ( n5188 , n2424 );
nor ( n5189 , n5158 , n5159 , n2424 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 );
and ( n5190 , n5157 , n5189 );
buf ( n5191 , n2424 );
buf ( n5192 , n2424 );
buf ( n5193 , n2424 );
buf ( n5194 , n2424 );
buf ( n5195 , n2424 );
buf ( n5196 , n2424 );
buf ( n5197 , n2424 );
buf ( n5198 , n2424 );
buf ( n5199 , n2424 );
buf ( n5200 , n2424 );
buf ( n5201 , n2424 );
buf ( n5202 , n2424 );
buf ( n5203 , n2424 );
buf ( n5204 , n2424 );
buf ( n5205 , n2424 );
buf ( n5206 , n2424 );
buf ( n5207 , n2424 );
buf ( n5208 , n2424 );
buf ( n5209 , n2424 );
buf ( n5210 , n2424 );
buf ( n5211 , n2424 );
buf ( n5212 , n2424 );
buf ( n5213 , n2424 );
buf ( n5214 , n2424 );
buf ( n5215 , n2424 );
buf ( n5216 , n2424 );
buf ( n5217 , n2424 );
buf ( n5218 , n2424 );
buf ( n5219 , n2424 );
nor ( n5220 , n5158 , n3348 , n2424 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 );
buf ( n5221 , n2424 );
buf ( n5222 , n2424 );
buf ( n5223 , n2424 );
buf ( n5224 , n2424 );
buf ( n5225 , n2424 );
buf ( n5226 , n2424 );
buf ( n5227 , n2424 );
buf ( n5228 , n2424 );
buf ( n5229 , n2424 );
buf ( n5230 , n2424 );
buf ( n5231 , n2424 );
buf ( n5232 , n2424 );
buf ( n5233 , n2424 );
buf ( n5234 , n2424 );
buf ( n5235 , n2424 );
buf ( n5236 , n2424 );
buf ( n5237 , n2424 );
buf ( n5238 , n2424 );
buf ( n5239 , n2424 );
buf ( n5240 , n2424 );
buf ( n5241 , n2424 );
buf ( n5242 , n2424 );
buf ( n5243 , n2424 );
buf ( n5244 , n2424 );
buf ( n5245 , n2424 );
buf ( n5246 , n2424 );
buf ( n5247 , n2424 );
buf ( n5248 , n2424 );
buf ( n5249 , n2424 );
nor ( n5250 , n3304 , n3348 , n2424 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 );
or ( n5251 , n5220 , n5250 );
buf ( n5252 , n2424 );
buf ( n5253 , n2424 );
buf ( n5254 , n2424 );
buf ( n5255 , n2424 );
buf ( n5256 , n2424 );
buf ( n5257 , n2424 );
buf ( n5258 , n2424 );
buf ( n5259 , n2424 );
buf ( n5260 , n2424 );
buf ( n5261 , n2424 );
buf ( n5262 , n2424 );
buf ( n5263 , n2424 );
buf ( n5264 , n2424 );
buf ( n5265 , n2424 );
buf ( n5266 , n2424 );
buf ( n5267 , n2424 );
buf ( n5268 , n2424 );
buf ( n5269 , n2424 );
buf ( n5270 , n2424 );
buf ( n5271 , n2424 );
buf ( n5272 , n2424 );
buf ( n5273 , n2424 );
buf ( n5274 , n2424 );
buf ( n5275 , n2424 );
buf ( n5276 , n2424 );
buf ( n5277 , n2424 );
buf ( n5278 , n2424 );
buf ( n5279 , n2424 );
buf ( n5280 , n2424 );
nor ( n5281 , n3304 , n5159 , n2424 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 );
or ( n5282 , n5251 , n5281 );
buf ( n5283 , n5282 );
and ( n5284 , n3363 , n5283 );
or ( n5285 , n5190 , n5284 );
and ( n5286 , n3627 , n3611 , n3618 , n3625 );
and ( n5287 , n5285 , n5286 );
and ( n5288 , n5145 , n5152 );
or ( n5289 , n5153 , n5288 );
and ( n5290 , n5144 , n5152 );
or ( n5291 , n5289 , n5290 );
and ( n5292 , n2313 , n5291 );
not ( n5293 , n2430 );
not ( n5294 , n5293 );
not ( n5295 , n2899 );
and ( n5296 , n5295 , n2449 );
not ( n5297 , n2449 );
not ( n5298 , n2430 );
xor ( n5299 , n5297 , n5298 );
and ( n5300 , n5299 , n2899 );
or ( n5301 , n5296 , n5300 );
not ( n5302 , n5301 );
not ( n5303 , n5302 );
or ( n5304 , n5294 , n5303 );
not ( n5305 , n2899 );
and ( n5306 , n5305 , n2464 );
not ( n5307 , n2464 );
and ( n5308 , n5297 , n5298 );
xor ( n5309 , n5307 , n5308 );
and ( n5310 , n5309 , n2899 );
or ( n5311 , n5306 , n5310 );
not ( n5312 , n5311 );
not ( n5313 , n5312 );
or ( n5314 , n5304 , n5313 );
not ( n5315 , n2899 );
and ( n5316 , n5315 , n2479 );
not ( n5317 , n2479 );
and ( n5318 , n5307 , n5308 );
xor ( n5319 , n5317 , n5318 );
and ( n5320 , n5319 , n2899 );
or ( n5321 , n5316 , n5320 );
not ( n5322 , n5321 );
not ( n5323 , n5322 );
or ( n5324 , n5314 , n5323 );
not ( n5325 , n2899 );
and ( n5326 , n5325 , n2494 );
not ( n5327 , n2494 );
and ( n5328 , n5317 , n5318 );
xor ( n5329 , n5327 , n5328 );
and ( n5330 , n5329 , n2899 );
or ( n5331 , n5326 , n5330 );
not ( n5332 , n5331 );
not ( n5333 , n5332 );
or ( n5334 , n5324 , n5333 );
not ( n5335 , n2899 );
and ( n5336 , n5335 , n2509 );
not ( n5337 , n2509 );
and ( n5338 , n5327 , n5328 );
xor ( n5339 , n5337 , n5338 );
and ( n5340 , n5339 , n2899 );
or ( n5341 , n5336 , n5340 );
not ( n5342 , n5341 );
not ( n5343 , n5342 );
or ( n5344 , n5334 , n5343 );
not ( n5345 , n2899 );
and ( n5346 , n5345 , n2524 );
not ( n5347 , n2524 );
and ( n5348 , n5337 , n5338 );
xor ( n5349 , n5347 , n5348 );
and ( n5350 , n5349 , n2899 );
or ( n5351 , n5346 , n5350 );
not ( n5352 , n5351 );
not ( n5353 , n5352 );
or ( n5354 , n5344 , n5353 );
not ( n5355 , n2899 );
and ( n5356 , n5355 , n2539 );
not ( n5357 , n2539 );
and ( n5358 , n5347 , n5348 );
xor ( n5359 , n5357 , n5358 );
and ( n5360 , n5359 , n2899 );
or ( n5361 , n5356 , n5360 );
not ( n5362 , n5361 );
not ( n5363 , n5362 );
or ( n5364 , n5354 , n5363 );
not ( n5365 , n2899 );
and ( n5366 , n5365 , n2554 );
not ( n5367 , n2554 );
and ( n5368 , n5357 , n5358 );
xor ( n5369 , n5367 , n5368 );
and ( n5370 , n5369 , n2899 );
or ( n5371 , n5366 , n5370 );
not ( n5372 , n5371 );
not ( n5373 , n5372 );
or ( n5374 , n5364 , n5373 );
not ( n5375 , n2899 );
and ( n5376 , n5375 , n2569 );
not ( n5377 , n2569 );
and ( n5378 , n5367 , n5368 );
xor ( n5379 , n5377 , n5378 );
and ( n5380 , n5379 , n2899 );
or ( n5381 , n5376 , n5380 );
not ( n5382 , n5381 );
not ( n5383 , n5382 );
or ( n5384 , n5374 , n5383 );
not ( n5385 , n2899 );
and ( n5386 , n5385 , n2584 );
not ( n5387 , n2584 );
and ( n5388 , n5377 , n5378 );
xor ( n5389 , n5387 , n5388 );
and ( n5390 , n5389 , n2899 );
or ( n5391 , n5386 , n5390 );
not ( n5392 , n5391 );
not ( n5393 , n5392 );
or ( n5394 , n5384 , n5393 );
not ( n5395 , n2899 );
and ( n5396 , n5395 , n2599 );
not ( n5397 , n2599 );
and ( n5398 , n5387 , n5388 );
xor ( n5399 , n5397 , n5398 );
and ( n5400 , n5399 , n2899 );
or ( n5401 , n5396 , n5400 );
not ( n5402 , n5401 );
not ( n5403 , n5402 );
or ( n5404 , n5394 , n5403 );
not ( n5405 , n2899 );
and ( n5406 , n5405 , n2614 );
not ( n5407 , n2614 );
and ( n5408 , n5397 , n5398 );
xor ( n5409 , n5407 , n5408 );
and ( n5410 , n5409 , n2899 );
or ( n5411 , n5406 , n5410 );
not ( n5412 , n5411 );
not ( n5413 , n5412 );
or ( n5414 , n5404 , n5413 );
not ( n5415 , n2899 );
and ( n5416 , n5415 , n2629 );
not ( n5417 , n2629 );
and ( n5418 , n5407 , n5408 );
xor ( n5419 , n5417 , n5418 );
and ( n5420 , n5419 , n2899 );
or ( n5421 , n5416 , n5420 );
not ( n5422 , n5421 );
not ( n5423 , n5422 );
or ( n5424 , n5414 , n5423 );
not ( n5425 , n2899 );
and ( n5426 , n5425 , n2644 );
not ( n5427 , n2644 );
and ( n5428 , n5417 , n5418 );
xor ( n5429 , n5427 , n5428 );
and ( n5430 , n5429 , n2899 );
or ( n5431 , n5426 , n5430 );
not ( n5432 , n5431 );
not ( n5433 , n5432 );
or ( n5434 , n5424 , n5433 );
not ( n5435 , n2899 );
and ( n5436 , n5435 , n2659 );
not ( n5437 , n2659 );
and ( n5438 , n5427 , n5428 );
xor ( n5439 , n5437 , n5438 );
and ( n5440 , n5439 , n2899 );
or ( n5441 , n5436 , n5440 );
not ( n5442 , n5441 );
not ( n5443 , n5442 );
or ( n5444 , n5434 , n5443 );
not ( n5445 , n2899 );
and ( n5446 , n5445 , n2674 );
not ( n5447 , n2674 );
and ( n5448 , n5437 , n5438 );
xor ( n5449 , n5447 , n5448 );
and ( n5450 , n5449 , n2899 );
or ( n5451 , n5446 , n5450 );
not ( n5452 , n5451 );
not ( n5453 , n5452 );
or ( n5454 , n5444 , n5453 );
not ( n5455 , n2899 );
and ( n5456 , n5455 , n2689 );
not ( n5457 , n2689 );
and ( n5458 , n5447 , n5448 );
xor ( n5459 , n5457 , n5458 );
and ( n5460 , n5459 , n2899 );
or ( n5461 , n5456 , n5460 );
not ( n5462 , n5461 );
not ( n5463 , n5462 );
or ( n5464 , n5454 , n5463 );
not ( n5465 , n2899 );
and ( n5466 , n5465 , n2704 );
not ( n5467 , n2704 );
and ( n5468 , n5457 , n5458 );
xor ( n5469 , n5467 , n5468 );
and ( n5470 , n5469 , n2899 );
or ( n5471 , n5466 , n5470 );
not ( n5472 , n5471 );
not ( n5473 , n5472 );
or ( n5474 , n5464 , n5473 );
not ( n5475 , n2899 );
and ( n5476 , n5475 , n2719 );
not ( n5477 , n2719 );
and ( n5478 , n5467 , n5468 );
xor ( n5479 , n5477 , n5478 );
and ( n5480 , n5479 , n2899 );
or ( n5481 , n5476 , n5480 );
not ( n5482 , n5481 );
not ( n5483 , n5482 );
or ( n5484 , n5474 , n5483 );
and ( n5485 , n5484 , n2899 );
not ( n5486 , n5485 );
and ( n5487 , n5486 , n5294 );
xor ( n5488 , n5294 , n2899 );
xor ( n5489 , n5488 , n2899 );
and ( n5490 , n5489 , n5485 );
or ( n5491 , n5487 , n5490 );
and ( n5492 , n5491 , n5155 );
or ( n5493 , n5292 , n5492 );
xor ( n5494 , n3795 , n5493 );
not ( n5495 , n5494 );
not ( n5496 , n5495 );
and ( n5497 , n2282 , n5291 );
not ( n5498 , n5497 );
xor ( n5499 , n3770 , n5498 );
and ( n5500 , n2283 , n5291 );
not ( n5501 , n5500 );
and ( n5502 , n3819 , n5501 );
and ( n5503 , n2284 , n5291 );
not ( n5504 , n5503 );
and ( n5505 , n3984 , n5504 );
and ( n5506 , n2285 , n5291 );
not ( n5507 , n5506 );
and ( n5508 , n3994 , n5507 );
and ( n5509 , n2286 , n5291 );
not ( n5510 , n5509 );
and ( n5511 , n4004 , n5510 );
and ( n5512 , n2287 , n5291 );
not ( n5513 , n5512 );
and ( n5514 , n4014 , n5513 );
and ( n5515 , n2288 , n5291 );
not ( n5516 , n5515 );
and ( n5517 , n4024 , n5516 );
and ( n5518 , n2289 , n5291 );
not ( n5519 , n5518 );
and ( n5520 , n4034 , n5519 );
and ( n5521 , n2290 , n5291 );
not ( n5522 , n5521 );
and ( n5523 , n4044 , n5522 );
and ( n5524 , n2291 , n5291 );
not ( n5525 , n5524 );
and ( n5526 , n4054 , n5525 );
and ( n5527 , n2292 , n5291 );
not ( n5528 , n5527 );
and ( n5529 , n4064 , n5528 );
and ( n5530 , n2293 , n5291 );
not ( n5531 , n5530 );
and ( n5532 , n4074 , n5531 );
and ( n5533 , n2294 , n5291 );
not ( n5534 , n5485 );
and ( n5535 , n5534 , n5483 );
xor ( n5536 , n5483 , n2899 );
xor ( n5537 , n5473 , n2899 );
xor ( n5538 , n5463 , n2899 );
xor ( n5539 , n5453 , n2899 );
xor ( n5540 , n5443 , n2899 );
xor ( n5541 , n5433 , n2899 );
xor ( n5542 , n5423 , n2899 );
xor ( n5543 , n5413 , n2899 );
xor ( n5544 , n5403 , n2899 );
xor ( n5545 , n5393 , n2899 );
xor ( n5546 , n5383 , n2899 );
xor ( n5547 , n5373 , n2899 );
xor ( n5548 , n5363 , n2899 );
xor ( n5549 , n5353 , n2899 );
xor ( n5550 , n5343 , n2899 );
xor ( n5551 , n5333 , n2899 );
xor ( n5552 , n5323 , n2899 );
xor ( n5553 , n5313 , n2899 );
xor ( n5554 , n5303 , n2899 );
and ( n5555 , n5488 , n2899 );
and ( n5556 , n5554 , n5555 );
and ( n5557 , n5553 , n5556 );
and ( n5558 , n5552 , n5557 );
and ( n5559 , n5551 , n5558 );
and ( n5560 , n5550 , n5559 );
and ( n5561 , n5549 , n5560 );
and ( n5562 , n5548 , n5561 );
and ( n5563 , n5547 , n5562 );
and ( n5564 , n5546 , n5563 );
and ( n5565 , n5545 , n5564 );
and ( n5566 , n5544 , n5565 );
and ( n5567 , n5543 , n5566 );
and ( n5568 , n5542 , n5567 );
and ( n5569 , n5541 , n5568 );
and ( n5570 , n5540 , n5569 );
and ( n5571 , n5539 , n5570 );
and ( n5572 , n5538 , n5571 );
and ( n5573 , n5537 , n5572 );
xor ( n5574 , n5536 , n5573 );
and ( n5575 , n5574 , n5485 );
or ( n5576 , n5535 , n5575 );
and ( n5577 , n5576 , n5155 );
or ( n5578 , n5533 , n5577 );
not ( n5579 , n5578 );
and ( n5580 , n4084 , n5579 );
and ( n5581 , n2295 , n5291 );
not ( n5582 , n5485 );
and ( n5583 , n5582 , n5473 );
xor ( n5584 , n5537 , n5572 );
and ( n5585 , n5584 , n5485 );
or ( n5586 , n5583 , n5585 );
and ( n5587 , n5586 , n5155 );
or ( n5588 , n5581 , n5587 );
not ( n5589 , n5588 );
and ( n5590 , n4094 , n5589 );
and ( n5591 , n2296 , n5291 );
not ( n5592 , n5485 );
and ( n5593 , n5592 , n5463 );
xor ( n5594 , n5538 , n5571 );
and ( n5595 , n5594 , n5485 );
or ( n5596 , n5593 , n5595 );
and ( n5597 , n5596 , n5155 );
or ( n5598 , n5591 , n5597 );
not ( n5599 , n5598 );
and ( n5600 , n4104 , n5599 );
and ( n5601 , n2297 , n5291 );
not ( n5602 , n5485 );
and ( n5603 , n5602 , n5453 );
xor ( n5604 , n5539 , n5570 );
and ( n5605 , n5604 , n5485 );
or ( n5606 , n5603 , n5605 );
and ( n5607 , n5606 , n5155 );
or ( n5608 , n5601 , n5607 );
not ( n5609 , n5608 );
and ( n5610 , n4114 , n5609 );
and ( n5611 , n2298 , n5291 );
not ( n5612 , n5485 );
and ( n5613 , n5612 , n5443 );
xor ( n5614 , n5540 , n5569 );
and ( n5615 , n5614 , n5485 );
or ( n5616 , n5613 , n5615 );
and ( n5617 , n5616 , n5155 );
or ( n5618 , n5611 , n5617 );
not ( n5619 , n5618 );
and ( n5620 , n4124 , n5619 );
and ( n5621 , n2299 , n5291 );
not ( n5622 , n5485 );
and ( n5623 , n5622 , n5433 );
xor ( n5624 , n5541 , n5568 );
and ( n5625 , n5624 , n5485 );
or ( n5626 , n5623 , n5625 );
and ( n5627 , n5626 , n5155 );
or ( n5628 , n5621 , n5627 );
not ( n5629 , n5628 );
and ( n5630 , n4134 , n5629 );
and ( n5631 , n2300 , n5291 );
not ( n5632 , n5485 );
and ( n5633 , n5632 , n5423 );
xor ( n5634 , n5542 , n5567 );
and ( n5635 , n5634 , n5485 );
or ( n5636 , n5633 , n5635 );
and ( n5637 , n5636 , n5155 );
or ( n5638 , n5631 , n5637 );
not ( n5639 , n5638 );
and ( n5640 , n4144 , n5639 );
and ( n5641 , n2301 , n5291 );
not ( n5642 , n5485 );
and ( n5643 , n5642 , n5413 );
xor ( n5644 , n5543 , n5566 );
and ( n5645 , n5644 , n5485 );
or ( n5646 , n5643 , n5645 );
and ( n5647 , n5646 , n5155 );
or ( n5648 , n5641 , n5647 );
not ( n5649 , n5648 );
and ( n5650 , n4154 , n5649 );
and ( n5651 , n2302 , n5291 );
not ( n5652 , n5485 );
and ( n5653 , n5652 , n5403 );
xor ( n5654 , n5544 , n5565 );
and ( n5655 , n5654 , n5485 );
or ( n5656 , n5653 , n5655 );
and ( n5657 , n5656 , n5155 );
or ( n5658 , n5651 , n5657 );
not ( n5659 , n5658 );
and ( n5660 , n4164 , n5659 );
and ( n5661 , n2303 , n5291 );
not ( n5662 , n5485 );
and ( n5663 , n5662 , n5393 );
xor ( n5664 , n5545 , n5564 );
and ( n5665 , n5664 , n5485 );
or ( n5666 , n5663 , n5665 );
and ( n5667 , n5666 , n5155 );
or ( n5668 , n5661 , n5667 );
not ( n5669 , n5668 );
and ( n5670 , n4174 , n5669 );
and ( n5671 , n2304 , n5291 );
not ( n5672 , n5485 );
and ( n5673 , n5672 , n5383 );
xor ( n5674 , n5546 , n5563 );
and ( n5675 , n5674 , n5485 );
or ( n5676 , n5673 , n5675 );
and ( n5677 , n5676 , n5155 );
or ( n5678 , n5671 , n5677 );
not ( n5679 , n5678 );
and ( n5680 , n4184 , n5679 );
and ( n5681 , n2305 , n5291 );
not ( n5682 , n5485 );
and ( n5683 , n5682 , n5373 );
xor ( n5684 , n5547 , n5562 );
and ( n5685 , n5684 , n5485 );
or ( n5686 , n5683 , n5685 );
and ( n5687 , n5686 , n5155 );
or ( n5688 , n5681 , n5687 );
not ( n5689 , n5688 );
and ( n5690 , n4194 , n5689 );
and ( n5691 , n2306 , n5291 );
not ( n5692 , n5485 );
and ( n5693 , n5692 , n5363 );
xor ( n5694 , n5548 , n5561 );
and ( n5695 , n5694 , n5485 );
or ( n5696 , n5693 , n5695 );
and ( n5697 , n5696 , n5155 );
or ( n5698 , n5691 , n5697 );
not ( n5699 , n5698 );
and ( n5700 , n4204 , n5699 );
and ( n5701 , n2307 , n5291 );
not ( n5702 , n5485 );
and ( n5703 , n5702 , n5353 );
xor ( n5704 , n5549 , n5560 );
and ( n5705 , n5704 , n5485 );
or ( n5706 , n5703 , n5705 );
and ( n5707 , n5706 , n5155 );
or ( n5708 , n5701 , n5707 );
not ( n5709 , n5708 );
and ( n5710 , n4214 , n5709 );
and ( n5711 , n2308 , n5291 );
not ( n5712 , n5485 );
and ( n5713 , n5712 , n5343 );
xor ( n5714 , n5550 , n5559 );
and ( n5715 , n5714 , n5485 );
or ( n5716 , n5713 , n5715 );
and ( n5717 , n5716 , n5155 );
or ( n5718 , n5711 , n5717 );
not ( n5719 , n5718 );
and ( n5720 , n4224 , n5719 );
and ( n5721 , n2309 , n5291 );
not ( n5722 , n5485 );
and ( n5723 , n5722 , n5333 );
xor ( n5724 , n5551 , n5558 );
and ( n5725 , n5724 , n5485 );
or ( n5726 , n5723 , n5725 );
and ( n5727 , n5726 , n5155 );
or ( n5728 , n5721 , n5727 );
not ( n5729 , n5728 );
and ( n5730 , n4234 , n5729 );
and ( n5731 , n2310 , n5291 );
not ( n5732 , n5485 );
and ( n5733 , n5732 , n5323 );
xor ( n5734 , n5552 , n5557 );
and ( n5735 , n5734 , n5485 );
or ( n5736 , n5733 , n5735 );
and ( n5737 , n5736 , n5155 );
or ( n5738 , n5731 , n5737 );
not ( n5739 , n5738 );
and ( n5740 , n4244 , n5739 );
and ( n5741 , n2311 , n5291 );
not ( n5742 , n5485 );
and ( n5743 , n5742 , n5313 );
xor ( n5744 , n5553 , n5556 );
and ( n5745 , n5744 , n5485 );
or ( n5746 , n5743 , n5745 );
and ( n5747 , n5746 , n5155 );
or ( n5748 , n5741 , n5747 );
not ( n5749 , n5748 );
and ( n5750 , n4258 , n5749 );
and ( n5751 , n2312 , n5291 );
not ( n5752 , n5485 );
and ( n5753 , n5752 , n5303 );
xor ( n5754 , n5554 , n5555 );
and ( n5755 , n5754 , n5485 );
or ( n5756 , n5753 , n5755 );
and ( n5757 , n5756 , n5155 );
or ( n5758 , n5751 , n5757 );
not ( n5759 , n5758 );
and ( n5760 , n3785 , n5759 );
not ( n5761 , n5493 );
or ( n5762 , n3795 , n5761 );
and ( n5763 , n5759 , n5762 );
and ( n5764 , n3785 , n5762 );
or ( n5765 , n5760 , n5763 , n5764 );
and ( n5766 , n5749 , n5765 );
and ( n5767 , n4258 , n5765 );
or ( n5768 , n5750 , n5766 , n5767 );
and ( n5769 , n5739 , n5768 );
and ( n5770 , n4244 , n5768 );
or ( n5771 , n5740 , n5769 , n5770 );
and ( n5772 , n5729 , n5771 );
and ( n5773 , n4234 , n5771 );
or ( n5774 , n5730 , n5772 , n5773 );
and ( n5775 , n5719 , n5774 );
and ( n5776 , n4224 , n5774 );
or ( n5777 , n5720 , n5775 , n5776 );
and ( n5778 , n5709 , n5777 );
and ( n5779 , n4214 , n5777 );
or ( n5780 , n5710 , n5778 , n5779 );
and ( n5781 , n5699 , n5780 );
and ( n5782 , n4204 , n5780 );
or ( n5783 , n5700 , n5781 , n5782 );
and ( n5784 , n5689 , n5783 );
and ( n5785 , n4194 , n5783 );
or ( n5786 , n5690 , n5784 , n5785 );
and ( n5787 , n5679 , n5786 );
and ( n5788 , n4184 , n5786 );
or ( n5789 , n5680 , n5787 , n5788 );
and ( n5790 , n5669 , n5789 );
and ( n5791 , n4174 , n5789 );
or ( n5792 , n5670 , n5790 , n5791 );
and ( n5793 , n5659 , n5792 );
and ( n5794 , n4164 , n5792 );
or ( n5795 , n5660 , n5793 , n5794 );
and ( n5796 , n5649 , n5795 );
and ( n5797 , n4154 , n5795 );
or ( n5798 , n5650 , n5796 , n5797 );
and ( n5799 , n5639 , n5798 );
and ( n5800 , n4144 , n5798 );
or ( n5801 , n5640 , n5799 , n5800 );
and ( n5802 , n5629 , n5801 );
and ( n5803 , n4134 , n5801 );
or ( n5804 , n5630 , n5802 , n5803 );
and ( n5805 , n5619 , n5804 );
and ( n5806 , n4124 , n5804 );
or ( n5807 , n5620 , n5805 , n5806 );
and ( n5808 , n5609 , n5807 );
and ( n5809 , n4114 , n5807 );
or ( n5810 , n5610 , n5808 , n5809 );
and ( n5811 , n5599 , n5810 );
and ( n5812 , n4104 , n5810 );
or ( n5813 , n5600 , n5811 , n5812 );
and ( n5814 , n5589 , n5813 );
and ( n5815 , n4094 , n5813 );
or ( n5816 , n5590 , n5814 , n5815 );
and ( n5817 , n5579 , n5816 );
and ( n5818 , n4084 , n5816 );
or ( n5819 , n5580 , n5817 , n5818 );
and ( n5820 , n5531 , n5819 );
and ( n5821 , n4074 , n5819 );
or ( n5822 , n5532 , n5820 , n5821 );
and ( n5823 , n5528 , n5822 );
and ( n5824 , n4064 , n5822 );
or ( n5825 , n5529 , n5823 , n5824 );
and ( n5826 , n5525 , n5825 );
and ( n5827 , n4054 , n5825 );
or ( n5828 , n5526 , n5826 , n5827 );
and ( n5829 , n5522 , n5828 );
and ( n5830 , n4044 , n5828 );
or ( n5831 , n5523 , n5829 , n5830 );
and ( n5832 , n5519 , n5831 );
and ( n5833 , n4034 , n5831 );
or ( n5834 , n5520 , n5832 , n5833 );
and ( n5835 , n5516 , n5834 );
and ( n5836 , n4024 , n5834 );
or ( n5837 , n5517 , n5835 , n5836 );
and ( n5838 , n5513 , n5837 );
and ( n5839 , n4014 , n5837 );
or ( n5840 , n5514 , n5838 , n5839 );
and ( n5841 , n5510 , n5840 );
and ( n5842 , n4004 , n5840 );
or ( n5843 , n5511 , n5841 , n5842 );
and ( n5844 , n5507 , n5843 );
and ( n5845 , n3994 , n5843 );
or ( n5846 , n5508 , n5844 , n5845 );
and ( n5847 , n5504 , n5846 );
and ( n5848 , n3984 , n5846 );
or ( n5849 , n5505 , n5847 , n5848 );
and ( n5850 , n5501 , n5849 );
and ( n5851 , n3819 , n5849 );
or ( n5852 , n5502 , n5850 , n5851 );
xor ( n5853 , n5499 , n5852 );
not ( n5854 , n5853 );
xor ( n5855 , n3785 , n5759 );
xor ( n5856 , n5855 , n5762 );
and ( n5857 , n5854 , n5856 );
not ( n5858 , n5856 );
not ( n5859 , n5494 );
xor ( n5860 , n5858 , n5859 );
and ( n5861 , n5860 , n5853 );
or ( n5862 , n5857 , n5861 );
not ( n5863 , n5862 );
not ( n5864 , n5863 );
or ( n5865 , n5496 , n5864 );
not ( n5866 , n5853 );
xor ( n5867 , n4258 , n5749 );
xor ( n5868 , n5867 , n5765 );
and ( n5869 , n5866 , n5868 );
not ( n5870 , n5868 );
and ( n5871 , n5858 , n5859 );
xor ( n5872 , n5870 , n5871 );
and ( n5873 , n5872 , n5853 );
or ( n5874 , n5869 , n5873 );
not ( n5875 , n5874 );
not ( n5876 , n5875 );
or ( n5877 , n5865 , n5876 );
not ( n5878 , n5853 );
xor ( n5879 , n4244 , n5739 );
xor ( n5880 , n5879 , n5768 );
and ( n5881 , n5878 , n5880 );
not ( n5882 , n5880 );
and ( n5883 , n5870 , n5871 );
xor ( n5884 , n5882 , n5883 );
and ( n5885 , n5884 , n5853 );
or ( n5886 , n5881 , n5885 );
not ( n5887 , n5886 );
not ( n5888 , n5887 );
or ( n5889 , n5877 , n5888 );
not ( n5890 , n5853 );
xor ( n5891 , n4234 , n5729 );
xor ( n5892 , n5891 , n5771 );
and ( n5893 , n5890 , n5892 );
not ( n5894 , n5892 );
and ( n5895 , n5882 , n5883 );
xor ( n5896 , n5894 , n5895 );
and ( n5897 , n5896 , n5853 );
or ( n5898 , n5893 , n5897 );
not ( n5899 , n5898 );
not ( n5900 , n5899 );
or ( n5901 , n5889 , n5900 );
not ( n5902 , n5853 );
xor ( n5903 , n4224 , n5719 );
xor ( n5904 , n5903 , n5774 );
and ( n5905 , n5902 , n5904 );
not ( n5906 , n5904 );
and ( n5907 , n5894 , n5895 );
xor ( n5908 , n5906 , n5907 );
and ( n5909 , n5908 , n5853 );
or ( n5910 , n5905 , n5909 );
not ( n5911 , n5910 );
not ( n5912 , n5911 );
or ( n5913 , n5901 , n5912 );
not ( n5914 , n5853 );
xor ( n5915 , n4214 , n5709 );
xor ( n5916 , n5915 , n5777 );
and ( n5917 , n5914 , n5916 );
not ( n5918 , n5916 );
and ( n5919 , n5906 , n5907 );
xor ( n5920 , n5918 , n5919 );
and ( n5921 , n5920 , n5853 );
or ( n5922 , n5917 , n5921 );
not ( n5923 , n5922 );
not ( n5924 , n5923 );
or ( n5925 , n5913 , n5924 );
not ( n5926 , n5853 );
xor ( n5927 , n4204 , n5699 );
xor ( n5928 , n5927 , n5780 );
and ( n5929 , n5926 , n5928 );
not ( n5930 , n5928 );
and ( n5931 , n5918 , n5919 );
xor ( n5932 , n5930 , n5931 );
and ( n5933 , n5932 , n5853 );
or ( n5934 , n5929 , n5933 );
not ( n5935 , n5934 );
not ( n5936 , n5935 );
or ( n5937 , n5925 , n5936 );
not ( n5938 , n5853 );
xor ( n5939 , n4194 , n5689 );
xor ( n5940 , n5939 , n5783 );
and ( n5941 , n5938 , n5940 );
not ( n5942 , n5940 );
and ( n5943 , n5930 , n5931 );
xor ( n5944 , n5942 , n5943 );
and ( n5945 , n5944 , n5853 );
or ( n5946 , n5941 , n5945 );
not ( n5947 , n5946 );
not ( n5948 , n5947 );
or ( n5949 , n5937 , n5948 );
not ( n5950 , n5853 );
xor ( n5951 , n4184 , n5679 );
xor ( n5952 , n5951 , n5786 );
and ( n5953 , n5950 , n5952 );
not ( n5954 , n5952 );
and ( n5955 , n5942 , n5943 );
xor ( n5956 , n5954 , n5955 );
and ( n5957 , n5956 , n5853 );
or ( n5958 , n5953 , n5957 );
not ( n5959 , n5958 );
not ( n5960 , n5959 );
or ( n5961 , n5949 , n5960 );
not ( n5962 , n5853 );
xor ( n5963 , n4174 , n5669 );
xor ( n5964 , n5963 , n5789 );
and ( n5965 , n5962 , n5964 );
not ( n5966 , n5964 );
and ( n5967 , n5954 , n5955 );
xor ( n5968 , n5966 , n5967 );
and ( n5969 , n5968 , n5853 );
or ( n5970 , n5965 , n5969 );
not ( n5971 , n5970 );
not ( n5972 , n5971 );
or ( n5973 , n5961 , n5972 );
not ( n5974 , n5853 );
xor ( n5975 , n4164 , n5659 );
xor ( n5976 , n5975 , n5792 );
and ( n5977 , n5974 , n5976 );
not ( n5978 , n5976 );
and ( n5979 , n5966 , n5967 );
xor ( n5980 , n5978 , n5979 );
and ( n5981 , n5980 , n5853 );
or ( n5982 , n5977 , n5981 );
not ( n5983 , n5982 );
not ( n5984 , n5983 );
or ( n5985 , n5973 , n5984 );
not ( n5986 , n5853 );
xor ( n5987 , n4154 , n5649 );
xor ( n5988 , n5987 , n5795 );
and ( n5989 , n5986 , n5988 );
not ( n5990 , n5988 );
and ( n5991 , n5978 , n5979 );
xor ( n5992 , n5990 , n5991 );
and ( n5993 , n5992 , n5853 );
or ( n5994 , n5989 , n5993 );
not ( n5995 , n5994 );
not ( n5996 , n5995 );
or ( n5997 , n5985 , n5996 );
not ( n5998 , n5853 );
xor ( n5999 , n4144 , n5639 );
xor ( n6000 , n5999 , n5798 );
and ( n6001 , n5998 , n6000 );
not ( n6002 , n6000 );
and ( n6003 , n5990 , n5991 );
xor ( n6004 , n6002 , n6003 );
and ( n6005 , n6004 , n5853 );
or ( n6006 , n6001 , n6005 );
not ( n6007 , n6006 );
not ( n6008 , n6007 );
or ( n6009 , n5997 , n6008 );
not ( n6010 , n5853 );
xor ( n6011 , n4134 , n5629 );
xor ( n6012 , n6011 , n5801 );
and ( n6013 , n6010 , n6012 );
not ( n6014 , n6012 );
and ( n6015 , n6002 , n6003 );
xor ( n6016 , n6014 , n6015 );
and ( n6017 , n6016 , n5853 );
or ( n6018 , n6013 , n6017 );
not ( n6019 , n6018 );
not ( n6020 , n6019 );
or ( n6021 , n6009 , n6020 );
not ( n6022 , n5853 );
xor ( n6023 , n4124 , n5619 );
xor ( n6024 , n6023 , n5804 );
and ( n6025 , n6022 , n6024 );
not ( n6026 , n6024 );
and ( n6027 , n6014 , n6015 );
xor ( n6028 , n6026 , n6027 );
and ( n6029 , n6028 , n5853 );
or ( n6030 , n6025 , n6029 );
not ( n6031 , n6030 );
not ( n6032 , n6031 );
or ( n6033 , n6021 , n6032 );
not ( n6034 , n5853 );
xor ( n6035 , n4114 , n5609 );
xor ( n6036 , n6035 , n5807 );
and ( n6037 , n6034 , n6036 );
not ( n6038 , n6036 );
and ( n6039 , n6026 , n6027 );
xor ( n6040 , n6038 , n6039 );
and ( n6041 , n6040 , n5853 );
or ( n6042 , n6037 , n6041 );
not ( n6043 , n6042 );
not ( n6044 , n6043 );
or ( n6045 , n6033 , n6044 );
not ( n6046 , n5853 );
xor ( n6047 , n4104 , n5599 );
xor ( n6048 , n6047 , n5810 );
and ( n6049 , n6046 , n6048 );
not ( n6050 , n6048 );
and ( n6051 , n6038 , n6039 );
xor ( n6052 , n6050 , n6051 );
and ( n6053 , n6052 , n5853 );
or ( n6054 , n6049 , n6053 );
not ( n6055 , n6054 );
not ( n6056 , n6055 );
or ( n6057 , n6045 , n6056 );
not ( n6058 , n5853 );
xor ( n6059 , n4094 , n5589 );
xor ( n6060 , n6059 , n5813 );
and ( n6061 , n6058 , n6060 );
not ( n6062 , n6060 );
and ( n6063 , n6050 , n6051 );
xor ( n6064 , n6062 , n6063 );
and ( n6065 , n6064 , n5853 );
or ( n6066 , n6061 , n6065 );
not ( n6067 , n6066 );
not ( n6068 , n6067 );
or ( n6069 , n6057 , n6068 );
not ( n6070 , n5853 );
xor ( n6071 , n4084 , n5579 );
xor ( n6072 , n6071 , n5816 );
and ( n6073 , n6070 , n6072 );
not ( n6074 , n6072 );
and ( n6075 , n6062 , n6063 );
xor ( n6076 , n6074 , n6075 );
and ( n6077 , n6076 , n5853 );
or ( n6078 , n6073 , n6077 );
not ( n6079 , n6078 );
not ( n6080 , n6079 );
or ( n6081 , n6069 , n6080 );
not ( n6082 , n5853 );
xor ( n6083 , n4074 , n5531 );
xor ( n6084 , n6083 , n5819 );
and ( n6085 , n6082 , n6084 );
not ( n6086 , n6084 );
and ( n6087 , n6074 , n6075 );
xor ( n6088 , n6086 , n6087 );
and ( n6089 , n6088 , n5853 );
or ( n6090 , n6085 , n6089 );
not ( n6091 , n6090 );
not ( n6092 , n6091 );
or ( n6093 , n6081 , n6092 );
not ( n6094 , n5853 );
xor ( n6095 , n4064 , n5528 );
xor ( n6096 , n6095 , n5822 );
and ( n6097 , n6094 , n6096 );
not ( n6098 , n6096 );
and ( n6099 , n6086 , n6087 );
xor ( n6100 , n6098 , n6099 );
and ( n6101 , n6100 , n5853 );
or ( n6102 , n6097 , n6101 );
not ( n6103 , n6102 );
not ( n6104 , n6103 );
or ( n6105 , n6093 , n6104 );
not ( n6106 , n5853 );
xor ( n6107 , n4054 , n5525 );
xor ( n6108 , n6107 , n5825 );
and ( n6109 , n6106 , n6108 );
not ( n6110 , n6108 );
and ( n6111 , n6098 , n6099 );
xor ( n6112 , n6110 , n6111 );
and ( n6113 , n6112 , n5853 );
or ( n6114 , n6109 , n6113 );
not ( n6115 , n6114 );
not ( n6116 , n6115 );
or ( n6117 , n6105 , n6116 );
not ( n6118 , n5853 );
xor ( n6119 , n4044 , n5522 );
xor ( n6120 , n6119 , n5828 );
and ( n6121 , n6118 , n6120 );
not ( n6122 , n6120 );
and ( n6123 , n6110 , n6111 );
xor ( n6124 , n6122 , n6123 );
and ( n6125 , n6124 , n5853 );
or ( n6126 , n6121 , n6125 );
not ( n6127 , n6126 );
not ( n6128 , n6127 );
or ( n6129 , n6117 , n6128 );
not ( n6130 , n5853 );
xor ( n6131 , n4034 , n5519 );
xor ( n6132 , n6131 , n5831 );
and ( n6133 , n6130 , n6132 );
not ( n6134 , n6132 );
and ( n6135 , n6122 , n6123 );
xor ( n6136 , n6134 , n6135 );
and ( n6137 , n6136 , n5853 );
or ( n6138 , n6133 , n6137 );
not ( n6139 , n6138 );
not ( n6140 , n6139 );
or ( n6141 , n6129 , n6140 );
not ( n6142 , n5853 );
xor ( n6143 , n4024 , n5516 );
xor ( n6144 , n6143 , n5834 );
and ( n6145 , n6142 , n6144 );
not ( n6146 , n6144 );
and ( n6147 , n6134 , n6135 );
xor ( n6148 , n6146 , n6147 );
and ( n6149 , n6148 , n5853 );
or ( n6150 , n6145 , n6149 );
not ( n6151 , n6150 );
not ( n6152 , n6151 );
or ( n6153 , n6141 , n6152 );
not ( n6154 , n5853 );
xor ( n6155 , n4014 , n5513 );
xor ( n6156 , n6155 , n5837 );
and ( n6157 , n6154 , n6156 );
not ( n6158 , n6156 );
and ( n6159 , n6146 , n6147 );
xor ( n6160 , n6158 , n6159 );
and ( n6161 , n6160 , n5853 );
or ( n6162 , n6157 , n6161 );
not ( n6163 , n6162 );
not ( n6164 , n6163 );
or ( n6165 , n6153 , n6164 );
not ( n6166 , n5853 );
xor ( n6167 , n4004 , n5510 );
xor ( n6168 , n6167 , n5840 );
and ( n6169 , n6166 , n6168 );
not ( n6170 , n6168 );
and ( n6171 , n6158 , n6159 );
xor ( n6172 , n6170 , n6171 );
and ( n6173 , n6172 , n5853 );
or ( n6174 , n6169 , n6173 );
not ( n6175 , n6174 );
not ( n6176 , n6175 );
or ( n6177 , n6165 , n6176 );
not ( n6178 , n5853 );
xor ( n6179 , n3994 , n5507 );
xor ( n6180 , n6179 , n5843 );
and ( n6181 , n6178 , n6180 );
not ( n6182 , n6180 );
and ( n6183 , n6170 , n6171 );
xor ( n6184 , n6182 , n6183 );
and ( n6185 , n6184 , n5853 );
or ( n6186 , n6181 , n6185 );
not ( n6187 , n6186 );
not ( n6188 , n6187 );
or ( n6189 , n6177 , n6188 );
not ( n6190 , n5853 );
xor ( n6191 , n3984 , n5504 );
xor ( n6192 , n6191 , n5846 );
and ( n6193 , n6190 , n6192 );
not ( n6194 , n6192 );
and ( n6195 , n6182 , n6183 );
xor ( n6196 , n6194 , n6195 );
and ( n6197 , n6196 , n5853 );
or ( n6198 , n6193 , n6197 );
not ( n6199 , n6198 );
not ( n6200 , n6199 );
or ( n6201 , n6189 , n6200 );
and ( n6202 , n6201 , n5853 );
not ( n6203 , n6202 );
and ( n6204 , n6203 , n5496 );
xor ( n6205 , n5496 , n5853 );
xor ( n6206 , n6205 , n5853 );
and ( n6207 , n6206 , n6202 );
or ( n6208 , n6204 , n6207 );
and ( n6209 , n6208 , n5189 );
and ( n6210 , n3363 , n5283 );
or ( n6211 , n6209 , n6210 );
not ( n6212 , n3625 );
and ( n6213 , n3627 , n3610 , n3618 , n6212 );
and ( n6214 , n3603 , n3610 , n3618 , n6212 );
or ( n6215 , n6213 , n6214 );
nor ( n6216 , n3627 , n3610 , n3618 , n6212 );
or ( n6217 , n6215 , n6216 );
nor ( n6218 , n3627 , n3611 , n3618 , n6212 );
or ( n6219 , n6217 , n6218 );
and ( n6220 , n6211 , n6219 );
xor ( n6221 , n3795 , n5493 );
not ( n6222 , n6221 );
not ( n6223 , n6222 );
xor ( n6224 , n3770 , n5497 );
and ( n6225 , n3819 , n5500 );
and ( n6226 , n3984 , n5503 );
and ( n6227 , n3994 , n5506 );
and ( n6228 , n4004 , n5509 );
and ( n6229 , n4014 , n5512 );
and ( n6230 , n4024 , n5515 );
and ( n6231 , n4034 , n5518 );
and ( n6232 , n4044 , n5521 );
and ( n6233 , n4054 , n5524 );
and ( n6234 , n4064 , n5527 );
and ( n6235 , n4074 , n5530 );
and ( n6236 , n4084 , n5578 );
and ( n6237 , n4094 , n5588 );
and ( n6238 , n4104 , n5598 );
and ( n6239 , n4114 , n5608 );
and ( n6240 , n4124 , n5618 );
and ( n6241 , n4134 , n5628 );
and ( n6242 , n4144 , n5638 );
and ( n6243 , n4154 , n5648 );
and ( n6244 , n4164 , n5658 );
and ( n6245 , n4174 , n5668 );
and ( n6246 , n4184 , n5678 );
and ( n6247 , n4194 , n5688 );
and ( n6248 , n4204 , n5698 );
and ( n6249 , n4214 , n5708 );
and ( n6250 , n4224 , n5718 );
and ( n6251 , n4234 , n5728 );
and ( n6252 , n4244 , n5738 );
and ( n6253 , n4258 , n5748 );
and ( n6254 , n3785 , n5758 );
and ( n6255 , n3795 , n5493 );
and ( n6256 , n5758 , n6255 );
and ( n6257 , n3785 , n6255 );
or ( n6258 , n6254 , n6256 , n6257 );
and ( n6259 , n5748 , n6258 );
and ( n6260 , n4258 , n6258 );
or ( n6261 , n6253 , n6259 , n6260 );
and ( n6262 , n5738 , n6261 );
and ( n6263 , n4244 , n6261 );
or ( n6264 , n6252 , n6262 , n6263 );
and ( n6265 , n5728 , n6264 );
and ( n6266 , n4234 , n6264 );
or ( n6267 , n6251 , n6265 , n6266 );
and ( n6268 , n5718 , n6267 );
and ( n6269 , n4224 , n6267 );
or ( n6270 , n6250 , n6268 , n6269 );
and ( n6271 , n5708 , n6270 );
and ( n6272 , n4214 , n6270 );
or ( n6273 , n6249 , n6271 , n6272 );
and ( n6274 , n5698 , n6273 );
and ( n6275 , n4204 , n6273 );
or ( n6276 , n6248 , n6274 , n6275 );
and ( n6277 , n5688 , n6276 );
and ( n6278 , n4194 , n6276 );
or ( n6279 , n6247 , n6277 , n6278 );
and ( n6280 , n5678 , n6279 );
and ( n6281 , n4184 , n6279 );
or ( n6282 , n6246 , n6280 , n6281 );
and ( n6283 , n5668 , n6282 );
and ( n6284 , n4174 , n6282 );
or ( n6285 , n6245 , n6283 , n6284 );
and ( n6286 , n5658 , n6285 );
and ( n6287 , n4164 , n6285 );
or ( n6288 , n6244 , n6286 , n6287 );
and ( n6289 , n5648 , n6288 );
and ( n6290 , n4154 , n6288 );
or ( n6291 , n6243 , n6289 , n6290 );
and ( n6292 , n5638 , n6291 );
and ( n6293 , n4144 , n6291 );
or ( n6294 , n6242 , n6292 , n6293 );
and ( n6295 , n5628 , n6294 );
and ( n6296 , n4134 , n6294 );
or ( n6297 , n6241 , n6295 , n6296 );
and ( n6298 , n5618 , n6297 );
and ( n6299 , n4124 , n6297 );
or ( n6300 , n6240 , n6298 , n6299 );
and ( n6301 , n5608 , n6300 );
and ( n6302 , n4114 , n6300 );
or ( n6303 , n6239 , n6301 , n6302 );
and ( n6304 , n5598 , n6303 );
and ( n6305 , n4104 , n6303 );
or ( n6306 , n6238 , n6304 , n6305 );
and ( n6307 , n5588 , n6306 );
and ( n6308 , n4094 , n6306 );
or ( n6309 , n6237 , n6307 , n6308 );
and ( n6310 , n5578 , n6309 );
and ( n6311 , n4084 , n6309 );
or ( n6312 , n6236 , n6310 , n6311 );
and ( n6313 , n5530 , n6312 );
and ( n6314 , n4074 , n6312 );
or ( n6315 , n6235 , n6313 , n6314 );
and ( n6316 , n5527 , n6315 );
and ( n6317 , n4064 , n6315 );
or ( n6318 , n6234 , n6316 , n6317 );
and ( n6319 , n5524 , n6318 );
and ( n6320 , n4054 , n6318 );
or ( n6321 , n6233 , n6319 , n6320 );
and ( n6322 , n5521 , n6321 );
and ( n6323 , n4044 , n6321 );
or ( n6324 , n6232 , n6322 , n6323 );
and ( n6325 , n5518 , n6324 );
and ( n6326 , n4034 , n6324 );
or ( n6327 , n6231 , n6325 , n6326 );
and ( n6328 , n5515 , n6327 );
and ( n6329 , n4024 , n6327 );
or ( n6330 , n6230 , n6328 , n6329 );
and ( n6331 , n5512 , n6330 );
and ( n6332 , n4014 , n6330 );
or ( n6333 , n6229 , n6331 , n6332 );
and ( n6334 , n5509 , n6333 );
and ( n6335 , n4004 , n6333 );
or ( n6336 , n6228 , n6334 , n6335 );
and ( n6337 , n5506 , n6336 );
and ( n6338 , n3994 , n6336 );
or ( n6339 , n6227 , n6337 , n6338 );
and ( n6340 , n5503 , n6339 );
and ( n6341 , n3984 , n6339 );
or ( n6342 , n6226 , n6340 , n6341 );
and ( n6343 , n5500 , n6342 );
and ( n6344 , n3819 , n6342 );
or ( n6345 , n6225 , n6343 , n6344 );
xor ( n6346 , n6224 , n6345 );
not ( n6347 , n6346 );
xor ( n6348 , n3785 , n5758 );
xor ( n6349 , n6348 , n6255 );
and ( n6350 , n6347 , n6349 );
not ( n6351 , n6349 );
not ( n6352 , n6221 );
xor ( n6353 , n6351 , n6352 );
and ( n6354 , n6353 , n6346 );
or ( n6355 , n6350 , n6354 );
not ( n6356 , n6355 );
not ( n6357 , n6356 );
or ( n6358 , n6223 , n6357 );
not ( n6359 , n6346 );
xor ( n6360 , n4258 , n5748 );
xor ( n6361 , n6360 , n6258 );
and ( n6362 , n6359 , n6361 );
not ( n6363 , n6361 );
and ( n6364 , n6351 , n6352 );
xor ( n6365 , n6363 , n6364 );
and ( n6366 , n6365 , n6346 );
or ( n6367 , n6362 , n6366 );
not ( n6368 , n6367 );
not ( n6369 , n6368 );
or ( n6370 , n6358 , n6369 );
not ( n6371 , n6346 );
xor ( n6372 , n4244 , n5738 );
xor ( n6373 , n6372 , n6261 );
and ( n6374 , n6371 , n6373 );
not ( n6375 , n6373 );
and ( n6376 , n6363 , n6364 );
xor ( n6377 , n6375 , n6376 );
and ( n6378 , n6377 , n6346 );
or ( n6379 , n6374 , n6378 );
not ( n6380 , n6379 );
not ( n6381 , n6380 );
or ( n6382 , n6370 , n6381 );
not ( n6383 , n6346 );
xor ( n6384 , n4234 , n5728 );
xor ( n6385 , n6384 , n6264 );
and ( n6386 , n6383 , n6385 );
not ( n6387 , n6385 );
and ( n6388 , n6375 , n6376 );
xor ( n6389 , n6387 , n6388 );
and ( n6390 , n6389 , n6346 );
or ( n6391 , n6386 , n6390 );
not ( n6392 , n6391 );
not ( n6393 , n6392 );
or ( n6394 , n6382 , n6393 );
not ( n6395 , n6346 );
xor ( n6396 , n4224 , n5718 );
xor ( n6397 , n6396 , n6267 );
and ( n6398 , n6395 , n6397 );
not ( n6399 , n6397 );
and ( n6400 , n6387 , n6388 );
xor ( n6401 , n6399 , n6400 );
and ( n6402 , n6401 , n6346 );
or ( n6403 , n6398 , n6402 );
not ( n6404 , n6403 );
not ( n6405 , n6404 );
or ( n6406 , n6394 , n6405 );
not ( n6407 , n6346 );
xor ( n6408 , n4214 , n5708 );
xor ( n6409 , n6408 , n6270 );
and ( n6410 , n6407 , n6409 );
not ( n6411 , n6409 );
and ( n6412 , n6399 , n6400 );
xor ( n6413 , n6411 , n6412 );
and ( n6414 , n6413 , n6346 );
or ( n6415 , n6410 , n6414 );
not ( n6416 , n6415 );
not ( n6417 , n6416 );
or ( n6418 , n6406 , n6417 );
not ( n6419 , n6346 );
xor ( n6420 , n4204 , n5698 );
xor ( n6421 , n6420 , n6273 );
and ( n6422 , n6419 , n6421 );
not ( n6423 , n6421 );
and ( n6424 , n6411 , n6412 );
xor ( n6425 , n6423 , n6424 );
and ( n6426 , n6425 , n6346 );
or ( n6427 , n6422 , n6426 );
not ( n6428 , n6427 );
not ( n6429 , n6428 );
or ( n6430 , n6418 , n6429 );
not ( n6431 , n6346 );
xor ( n6432 , n4194 , n5688 );
xor ( n6433 , n6432 , n6276 );
and ( n6434 , n6431 , n6433 );
not ( n6435 , n6433 );
and ( n6436 , n6423 , n6424 );
xor ( n6437 , n6435 , n6436 );
and ( n6438 , n6437 , n6346 );
or ( n6439 , n6434 , n6438 );
not ( n6440 , n6439 );
not ( n6441 , n6440 );
or ( n6442 , n6430 , n6441 );
not ( n6443 , n6346 );
xor ( n6444 , n4184 , n5678 );
xor ( n6445 , n6444 , n6279 );
and ( n6446 , n6443 , n6445 );
not ( n6447 , n6445 );
and ( n6448 , n6435 , n6436 );
xor ( n6449 , n6447 , n6448 );
and ( n6450 , n6449 , n6346 );
or ( n6451 , n6446 , n6450 );
not ( n6452 , n6451 );
not ( n6453 , n6452 );
or ( n6454 , n6442 , n6453 );
not ( n6455 , n6346 );
xor ( n6456 , n4174 , n5668 );
xor ( n6457 , n6456 , n6282 );
and ( n6458 , n6455 , n6457 );
not ( n6459 , n6457 );
and ( n6460 , n6447 , n6448 );
xor ( n6461 , n6459 , n6460 );
and ( n6462 , n6461 , n6346 );
or ( n6463 , n6458 , n6462 );
not ( n6464 , n6463 );
not ( n6465 , n6464 );
or ( n6466 , n6454 , n6465 );
not ( n6467 , n6346 );
xor ( n6468 , n4164 , n5658 );
xor ( n6469 , n6468 , n6285 );
and ( n6470 , n6467 , n6469 );
not ( n6471 , n6469 );
and ( n6472 , n6459 , n6460 );
xor ( n6473 , n6471 , n6472 );
and ( n6474 , n6473 , n6346 );
or ( n6475 , n6470 , n6474 );
not ( n6476 , n6475 );
not ( n6477 , n6476 );
or ( n6478 , n6466 , n6477 );
not ( n6479 , n6346 );
xor ( n6480 , n4154 , n5648 );
xor ( n6481 , n6480 , n6288 );
and ( n6482 , n6479 , n6481 );
not ( n6483 , n6481 );
and ( n6484 , n6471 , n6472 );
xor ( n6485 , n6483 , n6484 );
and ( n6486 , n6485 , n6346 );
or ( n6487 , n6482 , n6486 );
not ( n6488 , n6487 );
not ( n6489 , n6488 );
or ( n6490 , n6478 , n6489 );
not ( n6491 , n6346 );
xor ( n6492 , n4144 , n5638 );
xor ( n6493 , n6492 , n6291 );
and ( n6494 , n6491 , n6493 );
not ( n6495 , n6493 );
and ( n6496 , n6483 , n6484 );
xor ( n6497 , n6495 , n6496 );
and ( n6498 , n6497 , n6346 );
or ( n6499 , n6494 , n6498 );
not ( n6500 , n6499 );
not ( n6501 , n6500 );
or ( n6502 , n6490 , n6501 );
not ( n6503 , n6346 );
xor ( n6504 , n4134 , n5628 );
xor ( n6505 , n6504 , n6294 );
and ( n6506 , n6503 , n6505 );
not ( n6507 , n6505 );
and ( n6508 , n6495 , n6496 );
xor ( n6509 , n6507 , n6508 );
and ( n6510 , n6509 , n6346 );
or ( n6511 , n6506 , n6510 );
not ( n6512 , n6511 );
not ( n6513 , n6512 );
or ( n6514 , n6502 , n6513 );
not ( n6515 , n6346 );
xor ( n6516 , n4124 , n5618 );
xor ( n6517 , n6516 , n6297 );
and ( n6518 , n6515 , n6517 );
not ( n6519 , n6517 );
and ( n6520 , n6507 , n6508 );
xor ( n6521 , n6519 , n6520 );
and ( n6522 , n6521 , n6346 );
or ( n6523 , n6518 , n6522 );
not ( n6524 , n6523 );
not ( n6525 , n6524 );
or ( n6526 , n6514 , n6525 );
not ( n6527 , n6346 );
xor ( n6528 , n4114 , n5608 );
xor ( n6529 , n6528 , n6300 );
and ( n6530 , n6527 , n6529 );
not ( n6531 , n6529 );
and ( n6532 , n6519 , n6520 );
xor ( n6533 , n6531 , n6532 );
and ( n6534 , n6533 , n6346 );
or ( n6535 , n6530 , n6534 );
not ( n6536 , n6535 );
not ( n6537 , n6536 );
or ( n6538 , n6526 , n6537 );
not ( n6539 , n6346 );
xor ( n6540 , n4104 , n5598 );
xor ( n6541 , n6540 , n6303 );
and ( n6542 , n6539 , n6541 );
not ( n6543 , n6541 );
and ( n6544 , n6531 , n6532 );
xor ( n6545 , n6543 , n6544 );
and ( n6546 , n6545 , n6346 );
or ( n6547 , n6542 , n6546 );
not ( n6548 , n6547 );
not ( n6549 , n6548 );
or ( n6550 , n6538 , n6549 );
not ( n6551 , n6346 );
xor ( n6552 , n4094 , n5588 );
xor ( n6553 , n6552 , n6306 );
and ( n6554 , n6551 , n6553 );
not ( n6555 , n6553 );
and ( n6556 , n6543 , n6544 );
xor ( n6557 , n6555 , n6556 );
and ( n6558 , n6557 , n6346 );
or ( n6559 , n6554 , n6558 );
not ( n6560 , n6559 );
not ( n6561 , n6560 );
or ( n6562 , n6550 , n6561 );
not ( n6563 , n6346 );
xor ( n6564 , n4084 , n5578 );
xor ( n6565 , n6564 , n6309 );
and ( n6566 , n6563 , n6565 );
not ( n6567 , n6565 );
and ( n6568 , n6555 , n6556 );
xor ( n6569 , n6567 , n6568 );
and ( n6570 , n6569 , n6346 );
or ( n6571 , n6566 , n6570 );
not ( n6572 , n6571 );
not ( n6573 , n6572 );
or ( n6574 , n6562 , n6573 );
not ( n6575 , n6346 );
xor ( n6576 , n4074 , n5530 );
xor ( n6577 , n6576 , n6312 );
and ( n6578 , n6575 , n6577 );
not ( n6579 , n6577 );
and ( n6580 , n6567 , n6568 );
xor ( n6581 , n6579 , n6580 );
and ( n6582 , n6581 , n6346 );
or ( n6583 , n6578 , n6582 );
not ( n6584 , n6583 );
not ( n6585 , n6584 );
or ( n6586 , n6574 , n6585 );
not ( n6587 , n6346 );
xor ( n6588 , n4064 , n5527 );
xor ( n6589 , n6588 , n6315 );
and ( n6590 , n6587 , n6589 );
not ( n6591 , n6589 );
and ( n6592 , n6579 , n6580 );
xor ( n6593 , n6591 , n6592 );
and ( n6594 , n6593 , n6346 );
or ( n6595 , n6590 , n6594 );
not ( n6596 , n6595 );
not ( n6597 , n6596 );
or ( n6598 , n6586 , n6597 );
not ( n6599 , n6346 );
xor ( n6600 , n4054 , n5524 );
xor ( n6601 , n6600 , n6318 );
and ( n6602 , n6599 , n6601 );
not ( n6603 , n6601 );
and ( n6604 , n6591 , n6592 );
xor ( n6605 , n6603 , n6604 );
and ( n6606 , n6605 , n6346 );
or ( n6607 , n6602 , n6606 );
not ( n6608 , n6607 );
not ( n6609 , n6608 );
or ( n6610 , n6598 , n6609 );
not ( n6611 , n6346 );
xor ( n6612 , n4044 , n5521 );
xor ( n6613 , n6612 , n6321 );
and ( n6614 , n6611 , n6613 );
not ( n6615 , n6613 );
and ( n6616 , n6603 , n6604 );
xor ( n6617 , n6615 , n6616 );
and ( n6618 , n6617 , n6346 );
or ( n6619 , n6614 , n6618 );
not ( n6620 , n6619 );
not ( n6621 , n6620 );
or ( n6622 , n6610 , n6621 );
not ( n6623 , n6346 );
xor ( n6624 , n4034 , n5518 );
xor ( n6625 , n6624 , n6324 );
and ( n6626 , n6623 , n6625 );
not ( n6627 , n6625 );
and ( n6628 , n6615 , n6616 );
xor ( n6629 , n6627 , n6628 );
and ( n6630 , n6629 , n6346 );
or ( n6631 , n6626 , n6630 );
not ( n6632 , n6631 );
not ( n6633 , n6632 );
or ( n6634 , n6622 , n6633 );
not ( n6635 , n6346 );
xor ( n6636 , n4024 , n5515 );
xor ( n6637 , n6636 , n6327 );
and ( n6638 , n6635 , n6637 );
not ( n6639 , n6637 );
and ( n6640 , n6627 , n6628 );
xor ( n6641 , n6639 , n6640 );
and ( n6642 , n6641 , n6346 );
or ( n6643 , n6638 , n6642 );
not ( n6644 , n6643 );
not ( n6645 , n6644 );
or ( n6646 , n6634 , n6645 );
not ( n6647 , n6346 );
xor ( n6648 , n4014 , n5512 );
xor ( n6649 , n6648 , n6330 );
and ( n6650 , n6647 , n6649 );
not ( n6651 , n6649 );
and ( n6652 , n6639 , n6640 );
xor ( n6653 , n6651 , n6652 );
and ( n6654 , n6653 , n6346 );
or ( n6655 , n6650 , n6654 );
not ( n6656 , n6655 );
not ( n6657 , n6656 );
or ( n6658 , n6646 , n6657 );
not ( n6659 , n6346 );
xor ( n6660 , n4004 , n5509 );
xor ( n6661 , n6660 , n6333 );
and ( n6662 , n6659 , n6661 );
not ( n6663 , n6661 );
and ( n6664 , n6651 , n6652 );
xor ( n6665 , n6663 , n6664 );
and ( n6666 , n6665 , n6346 );
or ( n6667 , n6662 , n6666 );
not ( n6668 , n6667 );
not ( n6669 , n6668 );
or ( n6670 , n6658 , n6669 );
not ( n6671 , n6346 );
xor ( n6672 , n3994 , n5506 );
xor ( n6673 , n6672 , n6336 );
and ( n6674 , n6671 , n6673 );
not ( n6675 , n6673 );
and ( n6676 , n6663 , n6664 );
xor ( n6677 , n6675 , n6676 );
and ( n6678 , n6677 , n6346 );
or ( n6679 , n6674 , n6678 );
not ( n6680 , n6679 );
not ( n6681 , n6680 );
or ( n6682 , n6670 , n6681 );
not ( n6683 , n6346 );
xor ( n6684 , n3984 , n5503 );
xor ( n6685 , n6684 , n6339 );
and ( n6686 , n6683 , n6685 );
not ( n6687 , n6685 );
and ( n6688 , n6675 , n6676 );
xor ( n6689 , n6687 , n6688 );
and ( n6690 , n6689 , n6346 );
or ( n6691 , n6686 , n6690 );
not ( n6692 , n6691 );
not ( n6693 , n6692 );
or ( n6694 , n6682 , n6693 );
and ( n6695 , n6694 , n6346 );
not ( n6696 , n6695 );
and ( n6697 , n6696 , n6223 );
xor ( n6698 , n6223 , n6346 );
xor ( n6699 , n6698 , n6346 );
and ( n6700 , n6699 , n6695 );
or ( n6701 , n6697 , n6700 );
and ( n6702 , n6701 , n5189 );
and ( n6703 , n3363 , n5283 );
or ( n6704 , n6702 , n6703 );
and ( n6705 , n3627 , n3611 , n3618 , n6212 );
and ( n6706 , n3603 , n3611 , n3618 , n6212 );
or ( n6707 , n6705 , n6706 );
nor ( n6708 , n3603 , n3610 , n3618 , n6212 );
or ( n6709 , n6707 , n6708 );
nor ( n6710 , n3603 , n3611 , n3618 , n6212 );
or ( n6711 , n6709 , n6710 );
and ( n6712 , n6704 , n6711 );
and ( n6713 , n5493 , n5189 );
and ( n6714 , n3363 , n5283 );
or ( n6715 , n6713 , n6714 );
nor ( n6716 , n3603 , n3611 , n3618 , n3625 );
nor ( n6717 , n3627 , n3611 , n3618 , n3625 );
or ( n6718 , n6716 , n6717 );
and ( n6719 , n6715 , n6718 );
nor ( n6720 , n3627 , n3610 , n3618 , n3625 );
and ( n6721 , n5493 , n6720 );
and ( n6722 , n5493 , n5189 );
and ( n6723 , n3363 , n5283 );
or ( n6724 , n6722 , n6723 );
nor ( n6725 , n3603 , n3610 , n3618 , n3625 );
and ( n6726 , n6724 , n6725 );
or ( n6727 , n3632 , n5287 , n6220 , n6712 , n6719 , n6721 , n6726 );
and ( n6728 , n3360 , n6727 );
and ( n6729 , n3363 , n3260 );
or ( n6730 , n6728 , n6729 );
and ( n6731 , n6730 , n2422 );
and ( n6732 , n3356 , n2428 );
or ( n6733 , n6731 , n6732 );
buf ( n6734 , n6733 );
buf ( n6735 , n2424 );
buf ( n6736 , n2281 );
buf ( n6737 , n2280 );
not ( n6738 , n3260 );
and ( n6739 , n3776 , n3631 );
not ( n6740 , n3795 );
not ( n6741 , n6740 );
not ( n6742 , n3770 );
and ( n6743 , n6742 , n3785 );
not ( n6744 , n3785 );
not ( n6745 , n3795 );
xor ( n6746 , n6744 , n6745 );
and ( n6747 , n6746 , n3770 );
or ( n6748 , n6743 , n6747 );
not ( n6749 , n6748 );
not ( n6750 , n6749 );
or ( n6751 , n6741 , n6750 );
not ( n6752 , n3770 );
and ( n6753 , n6752 , n4258 );
not ( n6754 , n4258 );
and ( n6755 , n6744 , n6745 );
xor ( n6756 , n6754 , n6755 );
and ( n6757 , n6756 , n3770 );
or ( n6758 , n6753 , n6757 );
not ( n6759 , n6758 );
not ( n6760 , n6759 );
or ( n6761 , n6751 , n6760 );
not ( n6762 , n3770 );
and ( n6763 , n6762 , n4244 );
not ( n6764 , n4244 );
and ( n6765 , n6754 , n6755 );
xor ( n6766 , n6764 , n6765 );
and ( n6767 , n6766 , n3770 );
or ( n6768 , n6763 , n6767 );
not ( n6769 , n6768 );
not ( n6770 , n6769 );
or ( n6771 , n6761 , n6770 );
not ( n6772 , n3770 );
and ( n6773 , n6772 , n4234 );
not ( n6774 , n4234 );
and ( n6775 , n6764 , n6765 );
xor ( n6776 , n6774 , n6775 );
and ( n6777 , n6776 , n3770 );
or ( n6778 , n6773 , n6777 );
not ( n6779 , n6778 );
not ( n6780 , n6779 );
or ( n6781 , n6771 , n6780 );
not ( n6782 , n3770 );
and ( n6783 , n6782 , n4224 );
not ( n6784 , n4224 );
and ( n6785 , n6774 , n6775 );
xor ( n6786 , n6784 , n6785 );
and ( n6787 , n6786 , n3770 );
or ( n6788 , n6783 , n6787 );
not ( n6789 , n6788 );
not ( n6790 , n6789 );
or ( n6791 , n6781 , n6790 );
not ( n6792 , n3770 );
and ( n6793 , n6792 , n4214 );
not ( n6794 , n4214 );
and ( n6795 , n6784 , n6785 );
xor ( n6796 , n6794 , n6795 );
and ( n6797 , n6796 , n3770 );
or ( n6798 , n6793 , n6797 );
not ( n6799 , n6798 );
not ( n6800 , n6799 );
or ( n6801 , n6791 , n6800 );
not ( n6802 , n3770 );
and ( n6803 , n6802 , n4204 );
not ( n6804 , n4204 );
and ( n6805 , n6794 , n6795 );
xor ( n6806 , n6804 , n6805 );
and ( n6807 , n6806 , n3770 );
or ( n6808 , n6803 , n6807 );
not ( n6809 , n6808 );
not ( n6810 , n6809 );
or ( n6811 , n6801 , n6810 );
not ( n6812 , n3770 );
and ( n6813 , n6812 , n4194 );
not ( n6814 , n4194 );
and ( n6815 , n6804 , n6805 );
xor ( n6816 , n6814 , n6815 );
and ( n6817 , n6816 , n3770 );
or ( n6818 , n6813 , n6817 );
not ( n6819 , n6818 );
not ( n6820 , n6819 );
or ( n6821 , n6811 , n6820 );
not ( n6822 , n3770 );
and ( n6823 , n6822 , n4184 );
not ( n6824 , n4184 );
and ( n6825 , n6814 , n6815 );
xor ( n6826 , n6824 , n6825 );
and ( n6827 , n6826 , n3770 );
or ( n6828 , n6823 , n6827 );
not ( n6829 , n6828 );
not ( n6830 , n6829 );
or ( n6831 , n6821 , n6830 );
not ( n6832 , n3770 );
and ( n6833 , n6832 , n4174 );
not ( n6834 , n4174 );
and ( n6835 , n6824 , n6825 );
xor ( n6836 , n6834 , n6835 );
and ( n6837 , n6836 , n3770 );
or ( n6838 , n6833 , n6837 );
not ( n6839 , n6838 );
not ( n6840 , n6839 );
or ( n6841 , n6831 , n6840 );
not ( n6842 , n3770 );
and ( n6843 , n6842 , n4164 );
not ( n6844 , n4164 );
and ( n6845 , n6834 , n6835 );
xor ( n6846 , n6844 , n6845 );
and ( n6847 , n6846 , n3770 );
or ( n6848 , n6843 , n6847 );
not ( n6849 , n6848 );
not ( n6850 , n6849 );
or ( n6851 , n6841 , n6850 );
not ( n6852 , n3770 );
and ( n6853 , n6852 , n4154 );
not ( n6854 , n4154 );
and ( n6855 , n6844 , n6845 );
xor ( n6856 , n6854 , n6855 );
and ( n6857 , n6856 , n3770 );
or ( n6858 , n6853 , n6857 );
not ( n6859 , n6858 );
not ( n6860 , n6859 );
or ( n6861 , n6851 , n6860 );
not ( n6862 , n3770 );
and ( n6863 , n6862 , n4144 );
not ( n6864 , n4144 );
and ( n6865 , n6854 , n6855 );
xor ( n6866 , n6864 , n6865 );
and ( n6867 , n6866 , n3770 );
or ( n6868 , n6863 , n6867 );
not ( n6869 , n6868 );
not ( n6870 , n6869 );
or ( n6871 , n6861 , n6870 );
not ( n6872 , n3770 );
and ( n6873 , n6872 , n4134 );
not ( n6874 , n4134 );
and ( n6875 , n6864 , n6865 );
xor ( n6876 , n6874 , n6875 );
and ( n6877 , n6876 , n3770 );
or ( n6878 , n6873 , n6877 );
not ( n6879 , n6878 );
not ( n6880 , n6879 );
or ( n6881 , n6871 , n6880 );
not ( n6882 , n3770 );
and ( n6883 , n6882 , n4124 );
not ( n6884 , n4124 );
and ( n6885 , n6874 , n6875 );
xor ( n6886 , n6884 , n6885 );
and ( n6887 , n6886 , n3770 );
or ( n6888 , n6883 , n6887 );
not ( n6889 , n6888 );
not ( n6890 , n6889 );
or ( n6891 , n6881 , n6890 );
not ( n6892 , n3770 );
and ( n6893 , n6892 , n4114 );
not ( n6894 , n4114 );
and ( n6895 , n6884 , n6885 );
xor ( n6896 , n6894 , n6895 );
and ( n6897 , n6896 , n3770 );
or ( n6898 , n6893 , n6897 );
not ( n6899 , n6898 );
not ( n6900 , n6899 );
or ( n6901 , n6891 , n6900 );
not ( n6902 , n3770 );
and ( n6903 , n6902 , n4104 );
not ( n6904 , n4104 );
and ( n6905 , n6894 , n6895 );
xor ( n6906 , n6904 , n6905 );
and ( n6907 , n6906 , n3770 );
or ( n6908 , n6903 , n6907 );
not ( n6909 , n6908 );
not ( n6910 , n6909 );
or ( n6911 , n6901 , n6910 );
not ( n6912 , n3770 );
and ( n6913 , n6912 , n4094 );
not ( n6914 , n4094 );
and ( n6915 , n6904 , n6905 );
xor ( n6916 , n6914 , n6915 );
and ( n6917 , n6916 , n3770 );
or ( n6918 , n6913 , n6917 );
not ( n6919 , n6918 );
not ( n6920 , n6919 );
or ( n6921 , n6911 , n6920 );
not ( n6922 , n3770 );
and ( n6923 , n6922 , n4084 );
not ( n6924 , n4084 );
and ( n6925 , n6914 , n6915 );
xor ( n6926 , n6924 , n6925 );
and ( n6927 , n6926 , n3770 );
or ( n6928 , n6923 , n6927 );
not ( n6929 , n6928 );
not ( n6930 , n6929 );
or ( n6931 , n6921 , n6930 );
not ( n6932 , n3770 );
and ( n6933 , n6932 , n4074 );
not ( n6934 , n4074 );
and ( n6935 , n6924 , n6925 );
xor ( n6936 , n6934 , n6935 );
and ( n6937 , n6936 , n3770 );
or ( n6938 , n6933 , n6937 );
not ( n6939 , n6938 );
not ( n6940 , n6939 );
or ( n6941 , n6931 , n6940 );
not ( n6942 , n3770 );
and ( n6943 , n6942 , n4064 );
not ( n6944 , n4064 );
and ( n6945 , n6934 , n6935 );
xor ( n6946 , n6944 , n6945 );
and ( n6947 , n6946 , n3770 );
or ( n6948 , n6943 , n6947 );
not ( n6949 , n6948 );
not ( n6950 , n6949 );
or ( n6951 , n6941 , n6950 );
not ( n6952 , n3770 );
and ( n6953 , n6952 , n4054 );
not ( n6954 , n4054 );
and ( n6955 , n6944 , n6945 );
xor ( n6956 , n6954 , n6955 );
and ( n6957 , n6956 , n3770 );
or ( n6958 , n6953 , n6957 );
not ( n6959 , n6958 );
not ( n6960 , n6959 );
or ( n6961 , n6951 , n6960 );
not ( n6962 , n3770 );
and ( n6963 , n6962 , n4044 );
not ( n6964 , n4044 );
and ( n6965 , n6954 , n6955 );
xor ( n6966 , n6964 , n6965 );
and ( n6967 , n6966 , n3770 );
or ( n6968 , n6963 , n6967 );
not ( n6969 , n6968 );
not ( n6970 , n6969 );
or ( n6971 , n6961 , n6970 );
not ( n6972 , n3770 );
and ( n6973 , n6972 , n4034 );
not ( n6974 , n4034 );
and ( n6975 , n6964 , n6965 );
xor ( n6976 , n6974 , n6975 );
and ( n6977 , n6976 , n3770 );
or ( n6978 , n6973 , n6977 );
not ( n6979 , n6978 );
not ( n6980 , n6979 );
or ( n6981 , n6971 , n6980 );
not ( n6982 , n3770 );
and ( n6983 , n6982 , n4024 );
not ( n6984 , n4024 );
and ( n6985 , n6974 , n6975 );
xor ( n6986 , n6984 , n6985 );
and ( n6987 , n6986 , n3770 );
or ( n6988 , n6983 , n6987 );
not ( n6989 , n6988 );
not ( n6990 , n6989 );
or ( n6991 , n6981 , n6990 );
not ( n6992 , n3770 );
and ( n6993 , n6992 , n4014 );
not ( n6994 , n4014 );
and ( n6995 , n6984 , n6985 );
xor ( n6996 , n6994 , n6995 );
and ( n6997 , n6996 , n3770 );
or ( n6998 , n6993 , n6997 );
not ( n6999 , n6998 );
not ( n7000 , n6999 );
or ( n7001 , n6991 , n7000 );
not ( n7002 , n3770 );
and ( n7003 , n7002 , n4004 );
not ( n7004 , n4004 );
and ( n7005 , n6994 , n6995 );
xor ( n7006 , n7004 , n7005 );
and ( n7007 , n7006 , n3770 );
or ( n7008 , n7003 , n7007 );
not ( n7009 , n7008 );
not ( n7010 , n7009 );
or ( n7011 , n7001 , n7010 );
not ( n7012 , n3770 );
and ( n7013 , n7012 , n3994 );
not ( n7014 , n3994 );
and ( n7015 , n7004 , n7005 );
xor ( n7016 , n7014 , n7015 );
and ( n7017 , n7016 , n3770 );
or ( n7018 , n7013 , n7017 );
not ( n7019 , n7018 );
not ( n7020 , n7019 );
or ( n7021 , n7011 , n7020 );
and ( n7022 , n7021 , n3770 );
not ( n7023 , n7022 );
and ( n7024 , n7023 , n6741 );
xor ( n7025 , n6741 , n3770 );
xor ( n7026 , n7025 , n3770 );
and ( n7027 , n7026 , n7022 );
or ( n7028 , n7024 , n7027 );
and ( n7029 , n7028 , n5290 );
and ( n7030 , n7028 , n5288 );
not ( n7031 , n3290 );
and ( n7032 , n7031 , n4585 );
not ( n7033 , n5000 );
and ( n7034 , n7033 , n4593 );
xor ( n7035 , n4593 , n4579 );
and ( n7036 , n5003 , n4579 );
xor ( n7037 , n7035 , n7036 );
and ( n7038 , n7037 , n5000 );
or ( n7039 , n7034 , n7038 );
and ( n7040 , n7039 , n3290 );
or ( n7041 , n7032 , n7040 );
and ( n7042 , n7041 , n5153 );
and ( n7043 , n4585 , n5155 );
or ( n7044 , n7029 , n7030 , n7042 , n7043 );
and ( n7045 , n7044 , n5189 );
and ( n7046 , n3776 , n5283 );
or ( n7047 , n7045 , n7046 );
and ( n7048 , n7047 , n5286 );
not ( n7049 , n6202 );
and ( n7050 , n7049 , n5864 );
xor ( n7051 , n5864 , n5853 );
and ( n7052 , n6205 , n5853 );
xor ( n7053 , n7051 , n7052 );
and ( n7054 , n7053 , n6202 );
or ( n7055 , n7050 , n7054 );
and ( n7056 , n7055 , n5189 );
and ( n7057 , n3776 , n5283 );
or ( n7058 , n7056 , n7057 );
and ( n7059 , n7058 , n6219 );
not ( n7060 , n6695 );
and ( n7061 , n7060 , n6357 );
xor ( n7062 , n6357 , n6346 );
and ( n7063 , n6698 , n6346 );
xor ( n7064 , n7062 , n7063 );
and ( n7065 , n7064 , n6695 );
or ( n7066 , n7061 , n7065 );
and ( n7067 , n7066 , n5189 );
and ( n7068 , n3776 , n5283 );
or ( n7069 , n7067 , n7068 );
and ( n7070 , n7069 , n6711 );
and ( n7071 , n5758 , n5189 );
and ( n7072 , n3776 , n5283 );
or ( n7073 , n7071 , n7072 );
and ( n7074 , n7073 , n6718 );
and ( n7075 , n5758 , n6720 );
not ( n7076 , n5758 );
not ( n7077 , n5493 );
xor ( n7078 , n7076 , n7077 );
and ( n7079 , n7078 , n5189 );
and ( n7080 , n3776 , n5283 );
or ( n7081 , n7079 , n7080 );
and ( n7082 , n7081 , n6725 );
or ( n7083 , n6739 , n7048 , n7059 , n7070 , n7074 , n7075 , n7082 );
and ( n7084 , n6738 , n7083 );
and ( n7085 , n3776 , n3260 );
or ( n7086 , n7084 , n7085 );
and ( n7087 , n7086 , n2422 );
and ( n7088 , n3772 , n2428 );
or ( n7089 , n7087 , n7088 );
buf ( n7090 , n7089 );
buf ( n7091 , n2424 );
buf ( n7092 , n2281 );
buf ( n7093 , n2280 );
not ( n7094 , n3260 );
and ( n7095 , n4250 , n3631 );
not ( n7096 , n7022 );
and ( n7097 , n7096 , n6750 );
xor ( n7098 , n6750 , n3770 );
and ( n7099 , n7025 , n3770 );
xor ( n7100 , n7098 , n7099 );
and ( n7101 , n7100 , n7022 );
or ( n7102 , n7097 , n7101 );
and ( n7103 , n7102 , n5290 );
and ( n7104 , n7102 , n5288 );
not ( n7105 , n3290 );
and ( n7106 , n7105 , n4600 );
not ( n7107 , n5000 );
and ( n7108 , n7107 , n4608 );
xor ( n7109 , n4608 , n4579 );
and ( n7110 , n7035 , n7036 );
xor ( n7111 , n7109 , n7110 );
and ( n7112 , n7111 , n5000 );
or ( n7113 , n7108 , n7112 );
and ( n7114 , n7113 , n3290 );
or ( n7115 , n7106 , n7114 );
and ( n7116 , n7115 , n5153 );
and ( n7117 , n4600 , n5155 );
or ( n7118 , n7103 , n7104 , n7116 , n7117 );
and ( n7119 , n7118 , n5189 );
and ( n7120 , n4250 , n5283 );
or ( n7121 , n7119 , n7120 );
and ( n7122 , n7121 , n5286 );
not ( n7123 , n6202 );
and ( n7124 , n7123 , n5876 );
xor ( n7125 , n5876 , n5853 );
and ( n7126 , n7051 , n7052 );
xor ( n7127 , n7125 , n7126 );
and ( n7128 , n7127 , n6202 );
or ( n7129 , n7124 , n7128 );
and ( n7130 , n7129 , n5189 );
and ( n7131 , n4250 , n5283 );
or ( n7132 , n7130 , n7131 );
and ( n7133 , n7132 , n6219 );
not ( n7134 , n6695 );
and ( n7135 , n7134 , n6369 );
xor ( n7136 , n6369 , n6346 );
and ( n7137 , n7062 , n7063 );
xor ( n7138 , n7136 , n7137 );
and ( n7139 , n7138 , n6695 );
or ( n7140 , n7135 , n7139 );
and ( n7141 , n7140 , n5189 );
and ( n7142 , n4250 , n5283 );
or ( n7143 , n7141 , n7142 );
and ( n7144 , n7143 , n6711 );
and ( n7145 , n5748 , n5189 );
and ( n7146 , n4250 , n5283 );
or ( n7147 , n7145 , n7146 );
and ( n7148 , n7147 , n6718 );
and ( n7149 , n5748 , n6720 );
not ( n7150 , n5748 );
and ( n7151 , n7076 , n7077 );
xor ( n7152 , n7150 , n7151 );
and ( n7153 , n7152 , n5189 );
and ( n7154 , n4250 , n5283 );
or ( n7155 , n7153 , n7154 );
and ( n7156 , n7155 , n6725 );
or ( n7157 , n7095 , n7122 , n7133 , n7144 , n7148 , n7149 , n7156 );
and ( n7158 , n7094 , n7157 );
and ( n7159 , n4250 , n3260 );
or ( n7160 , n7158 , n7159 );
and ( n7161 , n7160 , n2422 );
and ( n7162 , n4246 , n2428 );
or ( n7163 , n7161 , n7162 );
buf ( n7164 , n7163 );
buf ( n7165 , n2424 );
buf ( n7166 , n2281 );
buf ( n7167 , n2280 );
not ( n7168 , n3260 );
and ( n7169 , n4236 , n3631 );
not ( n7170 , n7022 );
and ( n7171 , n7170 , n6760 );
xor ( n7172 , n6760 , n3770 );
and ( n7173 , n7098 , n7099 );
xor ( n7174 , n7172 , n7173 );
and ( n7175 , n7174 , n7022 );
or ( n7176 , n7171 , n7175 );
and ( n7177 , n7176 , n5290 );
and ( n7178 , n7176 , n5288 );
not ( n7179 , n3290 );
and ( n7180 , n7179 , n4615 );
not ( n7181 , n5000 );
and ( n7182 , n7181 , n4623 );
xor ( n7183 , n4623 , n4579 );
and ( n7184 , n7109 , n7110 );
xor ( n7185 , n7183 , n7184 );
and ( n7186 , n7185 , n5000 );
or ( n7187 , n7182 , n7186 );
and ( n7188 , n7187 , n3290 );
or ( n7189 , n7180 , n7188 );
and ( n7190 , n7189 , n5153 );
and ( n7191 , n4615 , n5155 );
or ( n7192 , n7177 , n7178 , n7190 , n7191 );
and ( n7193 , n7192 , n5189 );
and ( n7194 , n4236 , n5283 );
or ( n7195 , n7193 , n7194 );
and ( n7196 , n7195 , n5286 );
not ( n7197 , n6202 );
and ( n7198 , n7197 , n5888 );
xor ( n7199 , n5888 , n5853 );
and ( n7200 , n7125 , n7126 );
xor ( n7201 , n7199 , n7200 );
and ( n7202 , n7201 , n6202 );
or ( n7203 , n7198 , n7202 );
and ( n7204 , n7203 , n5189 );
and ( n7205 , n4236 , n5283 );
or ( n7206 , n7204 , n7205 );
and ( n7207 , n7206 , n6219 );
not ( n7208 , n6695 );
and ( n7209 , n7208 , n6381 );
xor ( n7210 , n6381 , n6346 );
and ( n7211 , n7136 , n7137 );
xor ( n7212 , n7210 , n7211 );
and ( n7213 , n7212 , n6695 );
or ( n7214 , n7209 , n7213 );
and ( n7215 , n7214 , n5189 );
and ( n7216 , n4236 , n5283 );
or ( n7217 , n7215 , n7216 );
and ( n7218 , n7217 , n6711 );
and ( n7219 , n5738 , n5189 );
and ( n7220 , n4236 , n5283 );
or ( n7221 , n7219 , n7220 );
and ( n7222 , n7221 , n6718 );
and ( n7223 , n5738 , n6720 );
not ( n7224 , n5738 );
and ( n7225 , n7150 , n7151 );
xor ( n7226 , n7224 , n7225 );
and ( n7227 , n7226 , n5189 );
and ( n7228 , n4236 , n5283 );
or ( n7229 , n7227 , n7228 );
and ( n7230 , n7229 , n6725 );
or ( n7231 , n7169 , n7196 , n7207 , n7218 , n7222 , n7223 , n7230 );
and ( n7232 , n7168 , n7231 );
and ( n7233 , n4236 , n3260 );
or ( n7234 , n7232 , n7233 );
and ( n7235 , n7234 , n2422 );
and ( n7236 , n3946 , n2428 );
or ( n7237 , n7235 , n7236 );
buf ( n7238 , n7237 );
buf ( n7239 , n2424 );
buf ( n7240 , n2281 );
buf ( n7241 , n2280 );
not ( n7242 , n3260 );
and ( n7243 , n4226 , n3631 );
not ( n7244 , n7022 );
and ( n7245 , n7244 , n6770 );
xor ( n7246 , n6770 , n3770 );
and ( n7247 , n7172 , n7173 );
xor ( n7248 , n7246 , n7247 );
and ( n7249 , n7248 , n7022 );
or ( n7250 , n7245 , n7249 );
and ( n7251 , n7250 , n5290 );
and ( n7252 , n7250 , n5288 );
not ( n7253 , n3290 );
and ( n7254 , n7253 , n4630 );
not ( n7255 , n5000 );
and ( n7256 , n7255 , n4638 );
xor ( n7257 , n4638 , n4579 );
and ( n7258 , n7183 , n7184 );
xor ( n7259 , n7257 , n7258 );
and ( n7260 , n7259 , n5000 );
or ( n7261 , n7256 , n7260 );
and ( n7262 , n7261 , n3290 );
or ( n7263 , n7254 , n7262 );
and ( n7264 , n7263 , n5153 );
and ( n7265 , n4630 , n5155 );
or ( n7266 , n7251 , n7252 , n7264 , n7265 );
and ( n7267 , n7266 , n5189 );
and ( n7268 , n4226 , n5283 );
or ( n7269 , n7267 , n7268 );
and ( n7270 , n7269 , n5286 );
not ( n7271 , n6202 );
and ( n7272 , n7271 , n5900 );
xor ( n7273 , n5900 , n5853 );
and ( n7274 , n7199 , n7200 );
xor ( n7275 , n7273 , n7274 );
and ( n7276 , n7275 , n6202 );
or ( n7277 , n7272 , n7276 );
and ( n7278 , n7277 , n5189 );
and ( n7279 , n4226 , n5283 );
or ( n7280 , n7278 , n7279 );
and ( n7281 , n7280 , n6219 );
not ( n7282 , n6695 );
and ( n7283 , n7282 , n6393 );
xor ( n7284 , n6393 , n6346 );
and ( n7285 , n7210 , n7211 );
xor ( n7286 , n7284 , n7285 );
and ( n7287 , n7286 , n6695 );
or ( n7288 , n7283 , n7287 );
and ( n7289 , n7288 , n5189 );
and ( n7290 , n4226 , n5283 );
or ( n7291 , n7289 , n7290 );
and ( n7292 , n7291 , n6711 );
and ( n7293 , n5728 , n5189 );
and ( n7294 , n4226 , n5283 );
or ( n7295 , n7293 , n7294 );
and ( n7296 , n7295 , n6718 );
and ( n7297 , n5728 , n6720 );
not ( n7298 , n5728 );
and ( n7299 , n7224 , n7225 );
xor ( n7300 , n7298 , n7299 );
and ( n7301 , n7300 , n5189 );
and ( n7302 , n4226 , n5283 );
or ( n7303 , n7301 , n7302 );
and ( n7304 , n7303 , n6725 );
or ( n7305 , n7243 , n7270 , n7281 , n7292 , n7296 , n7297 , n7304 );
and ( n7306 , n7242 , n7305 );
and ( n7307 , n4226 , n3260 );
or ( n7308 , n7306 , n7307 );
and ( n7309 , n7308 , n2422 );
and ( n7310 , n3941 , n2428 );
or ( n7311 , n7309 , n7310 );
buf ( n7312 , n7311 );
buf ( n7313 , n2424 );
buf ( n7314 , n2281 );
buf ( n7315 , n2280 );
not ( n7316 , n3260 );
and ( n7317 , n4216 , n3631 );
not ( n7318 , n7022 );
and ( n7319 , n7318 , n6780 );
xor ( n7320 , n6780 , n3770 );
and ( n7321 , n7246 , n7247 );
xor ( n7322 , n7320 , n7321 );
and ( n7323 , n7322 , n7022 );
or ( n7324 , n7319 , n7323 );
and ( n7325 , n7324 , n5290 );
and ( n7326 , n7324 , n5288 );
not ( n7327 , n3290 );
and ( n7328 , n7327 , n4645 );
not ( n7329 , n5000 );
and ( n7330 , n7329 , n4653 );
xor ( n7331 , n4653 , n4579 );
and ( n7332 , n7257 , n7258 );
xor ( n7333 , n7331 , n7332 );
and ( n7334 , n7333 , n5000 );
or ( n7335 , n7330 , n7334 );
and ( n7336 , n7335 , n3290 );
or ( n7337 , n7328 , n7336 );
and ( n7338 , n7337 , n5153 );
and ( n7339 , n4645 , n5155 );
or ( n7340 , n7325 , n7326 , n7338 , n7339 );
and ( n7341 , n7340 , n5189 );
and ( n7342 , n4216 , n5283 );
or ( n7343 , n7341 , n7342 );
and ( n7344 , n7343 , n5286 );
not ( n7345 , n6202 );
and ( n7346 , n7345 , n5912 );
xor ( n7347 , n5912 , n5853 );
and ( n7348 , n7273 , n7274 );
xor ( n7349 , n7347 , n7348 );
and ( n7350 , n7349 , n6202 );
or ( n7351 , n7346 , n7350 );
and ( n7352 , n7351 , n5189 );
and ( n7353 , n4216 , n5283 );
or ( n7354 , n7352 , n7353 );
and ( n7355 , n7354 , n6219 );
not ( n7356 , n6695 );
and ( n7357 , n7356 , n6405 );
xor ( n7358 , n6405 , n6346 );
and ( n7359 , n7284 , n7285 );
xor ( n7360 , n7358 , n7359 );
and ( n7361 , n7360 , n6695 );
or ( n7362 , n7357 , n7361 );
and ( n7363 , n7362 , n5189 );
and ( n7364 , n4216 , n5283 );
or ( n7365 , n7363 , n7364 );
and ( n7366 , n7365 , n6711 );
and ( n7367 , n5718 , n5189 );
and ( n7368 , n4216 , n5283 );
or ( n7369 , n7367 , n7368 );
and ( n7370 , n7369 , n6718 );
and ( n7371 , n5718 , n6720 );
not ( n7372 , n5718 );
and ( n7373 , n7298 , n7299 );
xor ( n7374 , n7372 , n7373 );
and ( n7375 , n7374 , n5189 );
and ( n7376 , n4216 , n5283 );
or ( n7377 , n7375 , n7376 );
and ( n7378 , n7377 , n6725 );
or ( n7379 , n7317 , n7344 , n7355 , n7366 , n7370 , n7371 , n7378 );
and ( n7380 , n7316 , n7379 );
and ( n7381 , n4216 , n3260 );
or ( n7382 , n7380 , n7381 );
and ( n7383 , n7382 , n2422 );
and ( n7384 , n3936 , n2428 );
or ( n7385 , n7383 , n7384 );
buf ( n7386 , n7385 );
buf ( n7387 , n2424 );
buf ( n7388 , n2281 );
buf ( n7389 , n2280 );
not ( n7390 , n3260 );
and ( n7391 , n4206 , n3631 );
not ( n7392 , n7022 );
and ( n7393 , n7392 , n6790 );
xor ( n7394 , n6790 , n3770 );
and ( n7395 , n7320 , n7321 );
xor ( n7396 , n7394 , n7395 );
and ( n7397 , n7396 , n7022 );
or ( n7398 , n7393 , n7397 );
and ( n7399 , n7398 , n5290 );
and ( n7400 , n7398 , n5288 );
not ( n7401 , n3290 );
and ( n7402 , n7401 , n4660 );
not ( n7403 , n5000 );
and ( n7404 , n7403 , n4668 );
xor ( n7405 , n4668 , n4579 );
and ( n7406 , n7331 , n7332 );
xor ( n7407 , n7405 , n7406 );
and ( n7408 , n7407 , n5000 );
or ( n7409 , n7404 , n7408 );
and ( n7410 , n7409 , n3290 );
or ( n7411 , n7402 , n7410 );
and ( n7412 , n7411 , n5153 );
and ( n7413 , n4660 , n5155 );
or ( n7414 , n7399 , n7400 , n7412 , n7413 );
and ( n7415 , n7414 , n5189 );
and ( n7416 , n4206 , n5283 );
or ( n7417 , n7415 , n7416 );
and ( n7418 , n7417 , n5286 );
not ( n7419 , n6202 );
and ( n7420 , n7419 , n5924 );
xor ( n7421 , n5924 , n5853 );
and ( n7422 , n7347 , n7348 );
xor ( n7423 , n7421 , n7422 );
and ( n7424 , n7423 , n6202 );
or ( n7425 , n7420 , n7424 );
and ( n7426 , n7425 , n5189 );
and ( n7427 , n4206 , n5283 );
or ( n7428 , n7426 , n7427 );
and ( n7429 , n7428 , n6219 );
not ( n7430 , n6695 );
and ( n7431 , n7430 , n6417 );
xor ( n7432 , n6417 , n6346 );
and ( n7433 , n7358 , n7359 );
xor ( n7434 , n7432 , n7433 );
and ( n7435 , n7434 , n6695 );
or ( n7436 , n7431 , n7435 );
and ( n7437 , n7436 , n5189 );
and ( n7438 , n4206 , n5283 );
or ( n7439 , n7437 , n7438 );
and ( n7440 , n7439 , n6711 );
and ( n7441 , n5708 , n5189 );
and ( n7442 , n4206 , n5283 );
or ( n7443 , n7441 , n7442 );
and ( n7444 , n7443 , n6718 );
and ( n7445 , n5708 , n6720 );
not ( n7446 , n5708 );
and ( n7447 , n7372 , n7373 );
xor ( n7448 , n7446 , n7447 );
and ( n7449 , n7448 , n5189 );
and ( n7450 , n4206 , n5283 );
or ( n7451 , n7449 , n7450 );
and ( n7452 , n7451 , n6725 );
or ( n7453 , n7391 , n7418 , n7429 , n7440 , n7444 , n7445 , n7452 );
and ( n7454 , n7390 , n7453 );
and ( n7455 , n4206 , n3260 );
or ( n7456 , n7454 , n7455 );
and ( n7457 , n7456 , n2422 );
and ( n7458 , n3931 , n2428 );
or ( n7459 , n7457 , n7458 );
buf ( n7460 , n7459 );
buf ( n7461 , n2424 );
buf ( n7462 , n2281 );
buf ( n7463 , n2280 );
not ( n7464 , n3260 );
and ( n7465 , n4196 , n3631 );
not ( n7466 , n7022 );
and ( n7467 , n7466 , n6800 );
xor ( n7468 , n6800 , n3770 );
and ( n7469 , n7394 , n7395 );
xor ( n7470 , n7468 , n7469 );
and ( n7471 , n7470 , n7022 );
or ( n7472 , n7467 , n7471 );
and ( n7473 , n7472 , n5290 );
and ( n7474 , n7472 , n5288 );
not ( n7475 , n3290 );
and ( n7476 , n7475 , n4675 );
not ( n7477 , n5000 );
and ( n7478 , n7477 , n4683 );
xor ( n7479 , n4683 , n4579 );
and ( n7480 , n7405 , n7406 );
xor ( n7481 , n7479 , n7480 );
and ( n7482 , n7481 , n5000 );
or ( n7483 , n7478 , n7482 );
and ( n7484 , n7483 , n3290 );
or ( n7485 , n7476 , n7484 );
and ( n7486 , n7485 , n5153 );
and ( n7487 , n4675 , n5155 );
or ( n7488 , n7473 , n7474 , n7486 , n7487 );
and ( n7489 , n7488 , n5189 );
and ( n7490 , n4196 , n5283 );
or ( n7491 , n7489 , n7490 );
and ( n7492 , n7491 , n5286 );
not ( n7493 , n6202 );
and ( n7494 , n7493 , n5936 );
xor ( n7495 , n5936 , n5853 );
and ( n7496 , n7421 , n7422 );
xor ( n7497 , n7495 , n7496 );
and ( n7498 , n7497 , n6202 );
or ( n7499 , n7494 , n7498 );
and ( n7500 , n7499 , n5189 );
and ( n7501 , n4196 , n5283 );
or ( n7502 , n7500 , n7501 );
and ( n7503 , n7502 , n6219 );
not ( n7504 , n6695 );
and ( n7505 , n7504 , n6429 );
xor ( n7506 , n6429 , n6346 );
and ( n7507 , n7432 , n7433 );
xor ( n7508 , n7506 , n7507 );
and ( n7509 , n7508 , n6695 );
or ( n7510 , n7505 , n7509 );
and ( n7511 , n7510 , n5189 );
and ( n7512 , n4196 , n5283 );
or ( n7513 , n7511 , n7512 );
and ( n7514 , n7513 , n6711 );
and ( n7515 , n5698 , n5189 );
and ( n7516 , n4196 , n5283 );
or ( n7517 , n7515 , n7516 );
and ( n7518 , n7517 , n6718 );
and ( n7519 , n5698 , n6720 );
not ( n7520 , n5698 );
and ( n7521 , n7446 , n7447 );
xor ( n7522 , n7520 , n7521 );
and ( n7523 , n7522 , n5189 );
and ( n7524 , n4196 , n5283 );
or ( n7525 , n7523 , n7524 );
and ( n7526 , n7525 , n6725 );
or ( n7527 , n7465 , n7492 , n7503 , n7514 , n7518 , n7519 , n7526 );
and ( n7528 , n7464 , n7527 );
and ( n7529 , n4196 , n3260 );
or ( n7530 , n7528 , n7529 );
and ( n7531 , n7530 , n2422 );
and ( n7532 , n3926 , n2428 );
or ( n7533 , n7531 , n7532 );
buf ( n7534 , n7533 );
buf ( n7535 , n2424 );
buf ( n7536 , n2281 );
buf ( n7537 , n2280 );
not ( n7538 , n3260 );
and ( n7539 , n4186 , n3631 );
not ( n7540 , n7022 );
and ( n7541 , n7540 , n6810 );
xor ( n7542 , n6810 , n3770 );
and ( n7543 , n7468 , n7469 );
xor ( n7544 , n7542 , n7543 );
and ( n7545 , n7544 , n7022 );
or ( n7546 , n7541 , n7545 );
and ( n7547 , n7546 , n5290 );
and ( n7548 , n7546 , n5288 );
not ( n7549 , n3290 );
and ( n7550 , n7549 , n4690 );
not ( n7551 , n5000 );
and ( n7552 , n7551 , n4698 );
xor ( n7553 , n4698 , n4579 );
and ( n7554 , n7479 , n7480 );
xor ( n7555 , n7553 , n7554 );
and ( n7556 , n7555 , n5000 );
or ( n7557 , n7552 , n7556 );
and ( n7558 , n7557 , n3290 );
or ( n7559 , n7550 , n7558 );
and ( n7560 , n7559 , n5153 );
and ( n7561 , n4690 , n5155 );
or ( n7562 , n7547 , n7548 , n7560 , n7561 );
and ( n7563 , n7562 , n5189 );
and ( n7564 , n4186 , n5283 );
or ( n7565 , n7563 , n7564 );
and ( n7566 , n7565 , n5286 );
not ( n7567 , n6202 );
and ( n7568 , n7567 , n5948 );
xor ( n7569 , n5948 , n5853 );
and ( n7570 , n7495 , n7496 );
xor ( n7571 , n7569 , n7570 );
and ( n7572 , n7571 , n6202 );
or ( n7573 , n7568 , n7572 );
and ( n7574 , n7573 , n5189 );
and ( n7575 , n4186 , n5283 );
or ( n7576 , n7574 , n7575 );
and ( n7577 , n7576 , n6219 );
not ( n7578 , n6695 );
and ( n7579 , n7578 , n6441 );
xor ( n7580 , n6441 , n6346 );
and ( n7581 , n7506 , n7507 );
xor ( n7582 , n7580 , n7581 );
and ( n7583 , n7582 , n6695 );
or ( n7584 , n7579 , n7583 );
and ( n7585 , n7584 , n5189 );
and ( n7586 , n4186 , n5283 );
or ( n7587 , n7585 , n7586 );
and ( n7588 , n7587 , n6711 );
and ( n7589 , n5688 , n5189 );
and ( n7590 , n4186 , n5283 );
or ( n7591 , n7589 , n7590 );
and ( n7592 , n7591 , n6718 );
and ( n7593 , n5688 , n6720 );
not ( n7594 , n5688 );
and ( n7595 , n7520 , n7521 );
xor ( n7596 , n7594 , n7595 );
and ( n7597 , n7596 , n5189 );
and ( n7598 , n4186 , n5283 );
or ( n7599 , n7597 , n7598 );
and ( n7600 , n7599 , n6725 );
or ( n7601 , n7539 , n7566 , n7577 , n7588 , n7592 , n7593 , n7600 );
and ( n7602 , n7538 , n7601 );
and ( n7603 , n4186 , n3260 );
or ( n7604 , n7602 , n7603 );
and ( n7605 , n7604 , n2422 );
and ( n7606 , n3921 , n2428 );
or ( n7607 , n7605 , n7606 );
buf ( n7608 , n7607 );
buf ( n7609 , n2424 );
buf ( n7610 , n2281 );
buf ( n7611 , n2280 );
not ( n7612 , n3260 );
and ( n7613 , n4176 , n3631 );
not ( n7614 , n7022 );
and ( n7615 , n7614 , n6820 );
xor ( n7616 , n6820 , n3770 );
and ( n7617 , n7542 , n7543 );
xor ( n7618 , n7616 , n7617 );
and ( n7619 , n7618 , n7022 );
or ( n7620 , n7615 , n7619 );
and ( n7621 , n7620 , n5290 );
and ( n7622 , n7620 , n5288 );
not ( n7623 , n3290 );
and ( n7624 , n7623 , n4705 );
not ( n7625 , n5000 );
and ( n7626 , n7625 , n4713 );
xor ( n7627 , n4713 , n4579 );
and ( n7628 , n7553 , n7554 );
xor ( n7629 , n7627 , n7628 );
and ( n7630 , n7629 , n5000 );
or ( n7631 , n7626 , n7630 );
and ( n7632 , n7631 , n3290 );
or ( n7633 , n7624 , n7632 );
and ( n7634 , n7633 , n5153 );
and ( n7635 , n4705 , n5155 );
or ( n7636 , n7621 , n7622 , n7634 , n7635 );
and ( n7637 , n7636 , n5189 );
and ( n7638 , n4176 , n5283 );
or ( n7639 , n7637 , n7638 );
and ( n7640 , n7639 , n5286 );
not ( n7641 , n6202 );
and ( n7642 , n7641 , n5960 );
xor ( n7643 , n5960 , n5853 );
and ( n7644 , n7569 , n7570 );
xor ( n7645 , n7643 , n7644 );
and ( n7646 , n7645 , n6202 );
or ( n7647 , n7642 , n7646 );
and ( n7648 , n7647 , n5189 );
and ( n7649 , n4176 , n5283 );
or ( n7650 , n7648 , n7649 );
and ( n7651 , n7650 , n6219 );
not ( n7652 , n6695 );
and ( n7653 , n7652 , n6453 );
xor ( n7654 , n6453 , n6346 );
and ( n7655 , n7580 , n7581 );
xor ( n7656 , n7654 , n7655 );
and ( n7657 , n7656 , n6695 );
or ( n7658 , n7653 , n7657 );
and ( n7659 , n7658 , n5189 );
and ( n7660 , n4176 , n5283 );
or ( n7661 , n7659 , n7660 );
and ( n7662 , n7661 , n6711 );
and ( n7663 , n5678 , n5189 );
and ( n7664 , n4176 , n5283 );
or ( n7665 , n7663 , n7664 );
and ( n7666 , n7665 , n6718 );
and ( n7667 , n5678 , n6720 );
not ( n7668 , n5678 );
and ( n7669 , n7594 , n7595 );
xor ( n7670 , n7668 , n7669 );
and ( n7671 , n7670 , n5189 );
and ( n7672 , n4176 , n5283 );
or ( n7673 , n7671 , n7672 );
and ( n7674 , n7673 , n6725 );
or ( n7675 , n7613 , n7640 , n7651 , n7662 , n7666 , n7667 , n7674 );
and ( n7676 , n7612 , n7675 );
and ( n7677 , n4176 , n3260 );
or ( n7678 , n7676 , n7677 );
and ( n7679 , n7678 , n2422 );
and ( n7680 , n3916 , n2428 );
or ( n7681 , n7679 , n7680 );
buf ( n7682 , n7681 );
buf ( n7683 , n2424 );
buf ( n7684 , n2281 );
buf ( n7685 , n2280 );
not ( n7686 , n3260 );
and ( n7687 , n4166 , n3631 );
not ( n7688 , n7022 );
and ( n7689 , n7688 , n6830 );
xor ( n7690 , n6830 , n3770 );
and ( n7691 , n7616 , n7617 );
xor ( n7692 , n7690 , n7691 );
and ( n7693 , n7692 , n7022 );
or ( n7694 , n7689 , n7693 );
and ( n7695 , n7694 , n5290 );
and ( n7696 , n7694 , n5288 );
not ( n7697 , n3290 );
and ( n7698 , n7697 , n4720 );
not ( n7699 , n5000 );
and ( n7700 , n7699 , n4728 );
xor ( n7701 , n4728 , n4579 );
and ( n7702 , n7627 , n7628 );
xor ( n7703 , n7701 , n7702 );
and ( n7704 , n7703 , n5000 );
or ( n7705 , n7700 , n7704 );
and ( n7706 , n7705 , n3290 );
or ( n7707 , n7698 , n7706 );
and ( n7708 , n7707 , n5153 );
and ( n7709 , n4720 , n5155 );
or ( n7710 , n7695 , n7696 , n7708 , n7709 );
and ( n7711 , n7710 , n5189 );
and ( n7712 , n4166 , n5283 );
or ( n7713 , n7711 , n7712 );
and ( n7714 , n7713 , n5286 );
not ( n7715 , n6202 );
and ( n7716 , n7715 , n5972 );
xor ( n7717 , n5972 , n5853 );
and ( n7718 , n7643 , n7644 );
xor ( n7719 , n7717 , n7718 );
and ( n7720 , n7719 , n6202 );
or ( n7721 , n7716 , n7720 );
and ( n7722 , n7721 , n5189 );
and ( n7723 , n4166 , n5283 );
or ( n7724 , n7722 , n7723 );
and ( n7725 , n7724 , n6219 );
not ( n7726 , n6695 );
and ( n7727 , n7726 , n6465 );
xor ( n7728 , n6465 , n6346 );
and ( n7729 , n7654 , n7655 );
xor ( n7730 , n7728 , n7729 );
and ( n7731 , n7730 , n6695 );
or ( n7732 , n7727 , n7731 );
and ( n7733 , n7732 , n5189 );
and ( n7734 , n4166 , n5283 );
or ( n7735 , n7733 , n7734 );
and ( n7736 , n7735 , n6711 );
and ( n7737 , n5668 , n5189 );
and ( n7738 , n4166 , n5283 );
or ( n7739 , n7737 , n7738 );
and ( n7740 , n7739 , n6718 );
and ( n7741 , n5668 , n6720 );
not ( n7742 , n5668 );
and ( n7743 , n7668 , n7669 );
xor ( n7744 , n7742 , n7743 );
and ( n7745 , n7744 , n5189 );
and ( n7746 , n4166 , n5283 );
or ( n7747 , n7745 , n7746 );
and ( n7748 , n7747 , n6725 );
or ( n7749 , n7687 , n7714 , n7725 , n7736 , n7740 , n7741 , n7748 );
and ( n7750 , n7686 , n7749 );
and ( n7751 , n4166 , n3260 );
or ( n7752 , n7750 , n7751 );
and ( n7753 , n7752 , n2422 );
and ( n7754 , n3911 , n2428 );
or ( n7755 , n7753 , n7754 );
buf ( n7756 , n7755 );
buf ( n7757 , n2424 );
buf ( n7758 , n2281 );
buf ( n7759 , n2280 );
not ( n7760 , n3260 );
and ( n7761 , n4156 , n3631 );
not ( n7762 , n7022 );
and ( n7763 , n7762 , n6840 );
xor ( n7764 , n6840 , n3770 );
and ( n7765 , n7690 , n7691 );
xor ( n7766 , n7764 , n7765 );
and ( n7767 , n7766 , n7022 );
or ( n7768 , n7763 , n7767 );
and ( n7769 , n7768 , n5290 );
and ( n7770 , n7768 , n5288 );
not ( n7771 , n3290 );
and ( n7772 , n7771 , n4735 );
not ( n7773 , n5000 );
and ( n7774 , n7773 , n4743 );
xor ( n7775 , n4743 , n4579 );
and ( n7776 , n7701 , n7702 );
xor ( n7777 , n7775 , n7776 );
and ( n7778 , n7777 , n5000 );
or ( n7779 , n7774 , n7778 );
and ( n7780 , n7779 , n3290 );
or ( n7781 , n7772 , n7780 );
and ( n7782 , n7781 , n5153 );
and ( n7783 , n4735 , n5155 );
or ( n7784 , n7769 , n7770 , n7782 , n7783 );
and ( n7785 , n7784 , n5189 );
and ( n7786 , n4156 , n5283 );
or ( n7787 , n7785 , n7786 );
and ( n7788 , n7787 , n5286 );
not ( n7789 , n6202 );
and ( n7790 , n7789 , n5984 );
xor ( n7791 , n5984 , n5853 );
and ( n7792 , n7717 , n7718 );
xor ( n7793 , n7791 , n7792 );
and ( n7794 , n7793 , n6202 );
or ( n7795 , n7790 , n7794 );
and ( n7796 , n7795 , n5189 );
and ( n7797 , n4156 , n5283 );
or ( n7798 , n7796 , n7797 );
and ( n7799 , n7798 , n6219 );
not ( n7800 , n6695 );
and ( n7801 , n7800 , n6477 );
xor ( n7802 , n6477 , n6346 );
and ( n7803 , n7728 , n7729 );
xor ( n7804 , n7802 , n7803 );
and ( n7805 , n7804 , n6695 );
or ( n7806 , n7801 , n7805 );
and ( n7807 , n7806 , n5189 );
and ( n7808 , n4156 , n5283 );
or ( n7809 , n7807 , n7808 );
and ( n7810 , n7809 , n6711 );
and ( n7811 , n5658 , n5189 );
and ( n7812 , n4156 , n5283 );
or ( n7813 , n7811 , n7812 );
and ( n7814 , n7813 , n6718 );
and ( n7815 , n5658 , n6720 );
not ( n7816 , n5658 );
and ( n7817 , n7742 , n7743 );
xor ( n7818 , n7816 , n7817 );
and ( n7819 , n7818 , n5189 );
and ( n7820 , n4156 , n5283 );
or ( n7821 , n7819 , n7820 );
and ( n7822 , n7821 , n6725 );
or ( n7823 , n7761 , n7788 , n7799 , n7810 , n7814 , n7815 , n7822 );
and ( n7824 , n7760 , n7823 );
and ( n7825 , n4156 , n3260 );
or ( n7826 , n7824 , n7825 );
and ( n7827 , n7826 , n2422 );
and ( n7828 , n3906 , n2428 );
or ( n7829 , n7827 , n7828 );
buf ( n7830 , n7829 );
buf ( n7831 , n2424 );
buf ( n7832 , n2281 );
buf ( n7833 , n2280 );
not ( n7834 , n3260 );
and ( n7835 , n4146 , n3631 );
not ( n7836 , n7022 );
and ( n7837 , n7836 , n6850 );
xor ( n7838 , n6850 , n3770 );
and ( n7839 , n7764 , n7765 );
xor ( n7840 , n7838 , n7839 );
and ( n7841 , n7840 , n7022 );
or ( n7842 , n7837 , n7841 );
and ( n7843 , n7842 , n5290 );
and ( n7844 , n7842 , n5288 );
not ( n7845 , n3290 );
and ( n7846 , n7845 , n4750 );
not ( n7847 , n5000 );
and ( n7848 , n7847 , n4758 );
xor ( n7849 , n4758 , n4579 );
and ( n7850 , n7775 , n7776 );
xor ( n7851 , n7849 , n7850 );
and ( n7852 , n7851 , n5000 );
or ( n7853 , n7848 , n7852 );
and ( n7854 , n7853 , n3290 );
or ( n7855 , n7846 , n7854 );
and ( n7856 , n7855 , n5153 );
and ( n7857 , n4750 , n5155 );
or ( n7858 , n7843 , n7844 , n7856 , n7857 );
and ( n7859 , n7858 , n5189 );
and ( n7860 , n4146 , n5283 );
or ( n7861 , n7859 , n7860 );
and ( n7862 , n7861 , n5286 );
not ( n7863 , n6202 );
and ( n7864 , n7863 , n5996 );
xor ( n7865 , n5996 , n5853 );
and ( n7866 , n7791 , n7792 );
xor ( n7867 , n7865 , n7866 );
and ( n7868 , n7867 , n6202 );
or ( n7869 , n7864 , n7868 );
and ( n7870 , n7869 , n5189 );
and ( n7871 , n4146 , n5283 );
or ( n7872 , n7870 , n7871 );
and ( n7873 , n7872 , n6219 );
not ( n7874 , n6695 );
and ( n7875 , n7874 , n6489 );
xor ( n7876 , n6489 , n6346 );
and ( n7877 , n7802 , n7803 );
xor ( n7878 , n7876 , n7877 );
and ( n7879 , n7878 , n6695 );
or ( n7880 , n7875 , n7879 );
and ( n7881 , n7880 , n5189 );
and ( n7882 , n4146 , n5283 );
or ( n7883 , n7881 , n7882 );
and ( n7884 , n7883 , n6711 );
and ( n7885 , n5648 , n5189 );
and ( n7886 , n4146 , n5283 );
or ( n7887 , n7885 , n7886 );
and ( n7888 , n7887 , n6718 );
and ( n7889 , n5648 , n6720 );
not ( n7890 , n5648 );
and ( n7891 , n7816 , n7817 );
xor ( n7892 , n7890 , n7891 );
and ( n7893 , n7892 , n5189 );
and ( n7894 , n4146 , n5283 );
or ( n7895 , n7893 , n7894 );
and ( n7896 , n7895 , n6725 );
or ( n7897 , n7835 , n7862 , n7873 , n7884 , n7888 , n7889 , n7896 );
and ( n7898 , n7834 , n7897 );
and ( n7899 , n4146 , n3260 );
or ( n7900 , n7898 , n7899 );
and ( n7901 , n7900 , n2422 );
and ( n7902 , n3901 , n2428 );
or ( n7903 , n7901 , n7902 );
buf ( n7904 , n7903 );
buf ( n7905 , n2424 );
buf ( n7906 , n2281 );
buf ( n7907 , n2280 );
not ( n7908 , n3260 );
and ( n7909 , n4136 , n3631 );
not ( n7910 , n7022 );
and ( n7911 , n7910 , n6860 );
xor ( n7912 , n6860 , n3770 );
and ( n7913 , n7838 , n7839 );
xor ( n7914 , n7912 , n7913 );
and ( n7915 , n7914 , n7022 );
or ( n7916 , n7911 , n7915 );
and ( n7917 , n7916 , n5290 );
and ( n7918 , n7916 , n5288 );
not ( n7919 , n3290 );
and ( n7920 , n7919 , n4765 );
not ( n7921 , n5000 );
and ( n7922 , n7921 , n4773 );
xor ( n7923 , n4773 , n4579 );
and ( n7924 , n7849 , n7850 );
xor ( n7925 , n7923 , n7924 );
and ( n7926 , n7925 , n5000 );
or ( n7927 , n7922 , n7926 );
and ( n7928 , n7927 , n3290 );
or ( n7929 , n7920 , n7928 );
and ( n7930 , n7929 , n5153 );
and ( n7931 , n4765 , n5155 );
or ( n7932 , n7917 , n7918 , n7930 , n7931 );
and ( n7933 , n7932 , n5189 );
and ( n7934 , n4136 , n5283 );
or ( n7935 , n7933 , n7934 );
and ( n7936 , n7935 , n5286 );
not ( n7937 , n6202 );
and ( n7938 , n7937 , n6008 );
xor ( n7939 , n6008 , n5853 );
and ( n7940 , n7865 , n7866 );
xor ( n7941 , n7939 , n7940 );
and ( n7942 , n7941 , n6202 );
or ( n7943 , n7938 , n7942 );
and ( n7944 , n7943 , n5189 );
and ( n7945 , n4136 , n5283 );
or ( n7946 , n7944 , n7945 );
and ( n7947 , n7946 , n6219 );
not ( n7948 , n6695 );
and ( n7949 , n7948 , n6501 );
xor ( n7950 , n6501 , n6346 );
and ( n7951 , n7876 , n7877 );
xor ( n7952 , n7950 , n7951 );
and ( n7953 , n7952 , n6695 );
or ( n7954 , n7949 , n7953 );
and ( n7955 , n7954 , n5189 );
and ( n7956 , n4136 , n5283 );
or ( n7957 , n7955 , n7956 );
and ( n7958 , n7957 , n6711 );
and ( n7959 , n5638 , n5189 );
and ( n7960 , n4136 , n5283 );
or ( n7961 , n7959 , n7960 );
and ( n7962 , n7961 , n6718 );
and ( n7963 , n5638 , n6720 );
not ( n7964 , n5638 );
and ( n7965 , n7890 , n7891 );
xor ( n7966 , n7964 , n7965 );
and ( n7967 , n7966 , n5189 );
and ( n7968 , n4136 , n5283 );
or ( n7969 , n7967 , n7968 );
and ( n7970 , n7969 , n6725 );
or ( n7971 , n7909 , n7936 , n7947 , n7958 , n7962 , n7963 , n7970 );
and ( n7972 , n7908 , n7971 );
and ( n7973 , n4136 , n3260 );
or ( n7974 , n7972 , n7973 );
and ( n7975 , n7974 , n2422 );
and ( n7976 , n3896 , n2428 );
or ( n7977 , n7975 , n7976 );
buf ( n7978 , n7977 );
buf ( n7979 , n2424 );
buf ( n7980 , n2281 );
buf ( n7981 , n2280 );
not ( n7982 , n3260 );
and ( n7983 , n4126 , n3631 );
not ( n7984 , n7022 );
and ( n7985 , n7984 , n6870 );
xor ( n7986 , n6870 , n3770 );
and ( n7987 , n7912 , n7913 );
xor ( n7988 , n7986 , n7987 );
and ( n7989 , n7988 , n7022 );
or ( n7990 , n7985 , n7989 );
and ( n7991 , n7990 , n5290 );
and ( n7992 , n7990 , n5288 );
not ( n7993 , n3290 );
and ( n7994 , n7993 , n4780 );
not ( n7995 , n5000 );
and ( n7996 , n7995 , n4788 );
xor ( n7997 , n4788 , n4579 );
and ( n7998 , n7923 , n7924 );
xor ( n7999 , n7997 , n7998 );
and ( n8000 , n7999 , n5000 );
or ( n8001 , n7996 , n8000 );
and ( n8002 , n8001 , n3290 );
or ( n8003 , n7994 , n8002 );
and ( n8004 , n8003 , n5153 );
and ( n8005 , n4780 , n5155 );
or ( n8006 , n7991 , n7992 , n8004 , n8005 );
and ( n8007 , n8006 , n5189 );
and ( n8008 , n4126 , n5283 );
or ( n8009 , n8007 , n8008 );
and ( n8010 , n8009 , n5286 );
not ( n8011 , n6202 );
and ( n8012 , n8011 , n6020 );
xor ( n8013 , n6020 , n5853 );
and ( n8014 , n7939 , n7940 );
xor ( n8015 , n8013 , n8014 );
and ( n8016 , n8015 , n6202 );
or ( n8017 , n8012 , n8016 );
and ( n8018 , n8017 , n5189 );
and ( n8019 , n4126 , n5283 );
or ( n8020 , n8018 , n8019 );
and ( n8021 , n8020 , n6219 );
not ( n8022 , n6695 );
and ( n8023 , n8022 , n6513 );
xor ( n8024 , n6513 , n6346 );
and ( n8025 , n7950 , n7951 );
xor ( n8026 , n8024 , n8025 );
and ( n8027 , n8026 , n6695 );
or ( n8028 , n8023 , n8027 );
and ( n8029 , n8028 , n5189 );
and ( n8030 , n4126 , n5283 );
or ( n8031 , n8029 , n8030 );
and ( n8032 , n8031 , n6711 );
and ( n8033 , n5628 , n5189 );
and ( n8034 , n4126 , n5283 );
or ( n8035 , n8033 , n8034 );
and ( n8036 , n8035 , n6718 );
and ( n8037 , n5628 , n6720 );
not ( n8038 , n5628 );
and ( n8039 , n7964 , n7965 );
xor ( n8040 , n8038 , n8039 );
and ( n8041 , n8040 , n5189 );
and ( n8042 , n4126 , n5283 );
or ( n8043 , n8041 , n8042 );
and ( n8044 , n8043 , n6725 );
or ( n8045 , n7983 , n8010 , n8021 , n8032 , n8036 , n8037 , n8044 );
and ( n8046 , n7982 , n8045 );
and ( n8047 , n4126 , n3260 );
or ( n8048 , n8046 , n8047 );
and ( n8049 , n8048 , n2422 );
and ( n8050 , n3891 , n2428 );
or ( n8051 , n8049 , n8050 );
buf ( n8052 , n8051 );
buf ( n8053 , n2424 );
buf ( n8054 , n2281 );
buf ( n8055 , n2280 );
not ( n8056 , n3260 );
and ( n8057 , n4116 , n3631 );
not ( n8058 , n7022 );
and ( n8059 , n8058 , n6880 );
xor ( n8060 , n6880 , n3770 );
and ( n8061 , n7986 , n7987 );
xor ( n8062 , n8060 , n8061 );
and ( n8063 , n8062 , n7022 );
or ( n8064 , n8059 , n8063 );
and ( n8065 , n8064 , n5290 );
and ( n8066 , n8064 , n5288 );
not ( n8067 , n3290 );
and ( n8068 , n8067 , n4795 );
not ( n8069 , n5000 );
and ( n8070 , n8069 , n4803 );
xor ( n8071 , n4803 , n4579 );
and ( n8072 , n7997 , n7998 );
xor ( n8073 , n8071 , n8072 );
and ( n8074 , n8073 , n5000 );
or ( n8075 , n8070 , n8074 );
and ( n8076 , n8075 , n3290 );
or ( n8077 , n8068 , n8076 );
and ( n8078 , n8077 , n5153 );
and ( n8079 , n4795 , n5155 );
or ( n8080 , n8065 , n8066 , n8078 , n8079 );
and ( n8081 , n8080 , n5189 );
and ( n8082 , n4116 , n5283 );
or ( n8083 , n8081 , n8082 );
and ( n8084 , n8083 , n5286 );
not ( n8085 , n6202 );
and ( n8086 , n8085 , n6032 );
xor ( n8087 , n6032 , n5853 );
and ( n8088 , n8013 , n8014 );
xor ( n8089 , n8087 , n8088 );
and ( n8090 , n8089 , n6202 );
or ( n8091 , n8086 , n8090 );
and ( n8092 , n8091 , n5189 );
and ( n8093 , n4116 , n5283 );
or ( n8094 , n8092 , n8093 );
and ( n8095 , n8094 , n6219 );
not ( n8096 , n6695 );
and ( n8097 , n8096 , n6525 );
xor ( n8098 , n6525 , n6346 );
and ( n8099 , n8024 , n8025 );
xor ( n8100 , n8098 , n8099 );
and ( n8101 , n8100 , n6695 );
or ( n8102 , n8097 , n8101 );
and ( n8103 , n8102 , n5189 );
and ( n8104 , n4116 , n5283 );
or ( n8105 , n8103 , n8104 );
and ( n8106 , n8105 , n6711 );
and ( n8107 , n5618 , n5189 );
and ( n8108 , n4116 , n5283 );
or ( n8109 , n8107 , n8108 );
and ( n8110 , n8109 , n6718 );
and ( n8111 , n5618 , n6720 );
not ( n8112 , n5618 );
and ( n8113 , n8038 , n8039 );
xor ( n8114 , n8112 , n8113 );
and ( n8115 , n8114 , n5189 );
and ( n8116 , n4116 , n5283 );
or ( n8117 , n8115 , n8116 );
and ( n8118 , n8117 , n6725 );
or ( n8119 , n8057 , n8084 , n8095 , n8106 , n8110 , n8111 , n8118 );
and ( n8120 , n8056 , n8119 );
and ( n8121 , n4116 , n3260 );
or ( n8122 , n8120 , n8121 );
and ( n8123 , n8122 , n2422 );
and ( n8124 , n3886 , n2428 );
or ( n8125 , n8123 , n8124 );
buf ( n8126 , n8125 );
buf ( n8127 , n2424 );
buf ( n8128 , n2281 );
buf ( n8129 , n2280 );
not ( n8130 , n3260 );
and ( n8131 , n4106 , n3631 );
not ( n8132 , n7022 );
and ( n8133 , n8132 , n6890 );
xor ( n8134 , n6890 , n3770 );
and ( n8135 , n8060 , n8061 );
xor ( n8136 , n8134 , n8135 );
and ( n8137 , n8136 , n7022 );
or ( n8138 , n8133 , n8137 );
and ( n8139 , n8138 , n5290 );
and ( n8140 , n8138 , n5288 );
not ( n8141 , n3290 );
and ( n8142 , n8141 , n4810 );
not ( n8143 , n5000 );
and ( n8144 , n8143 , n4818 );
xor ( n8145 , n4818 , n4579 );
and ( n8146 , n8071 , n8072 );
xor ( n8147 , n8145 , n8146 );
and ( n8148 , n8147 , n5000 );
or ( n8149 , n8144 , n8148 );
and ( n8150 , n8149 , n3290 );
or ( n8151 , n8142 , n8150 );
and ( n8152 , n8151 , n5153 );
and ( n8153 , n4810 , n5155 );
or ( n8154 , n8139 , n8140 , n8152 , n8153 );
and ( n8155 , n8154 , n5189 );
and ( n8156 , n4106 , n5283 );
or ( n8157 , n8155 , n8156 );
and ( n8158 , n8157 , n5286 );
not ( n8159 , n6202 );
and ( n8160 , n8159 , n6044 );
xor ( n8161 , n6044 , n5853 );
and ( n8162 , n8087 , n8088 );
xor ( n8163 , n8161 , n8162 );
and ( n8164 , n8163 , n6202 );
or ( n8165 , n8160 , n8164 );
and ( n8166 , n8165 , n5189 );
and ( n8167 , n4106 , n5283 );
or ( n8168 , n8166 , n8167 );
and ( n8169 , n8168 , n6219 );
not ( n8170 , n6695 );
and ( n8171 , n8170 , n6537 );
xor ( n8172 , n6537 , n6346 );
and ( n8173 , n8098 , n8099 );
xor ( n8174 , n8172 , n8173 );
and ( n8175 , n8174 , n6695 );
or ( n8176 , n8171 , n8175 );
and ( n8177 , n8176 , n5189 );
and ( n8178 , n4106 , n5283 );
or ( n8179 , n8177 , n8178 );
and ( n8180 , n8179 , n6711 );
and ( n8181 , n5608 , n5189 );
and ( n8182 , n4106 , n5283 );
or ( n8183 , n8181 , n8182 );
and ( n8184 , n8183 , n6718 );
and ( n8185 , n5608 , n6720 );
not ( n8186 , n5608 );
and ( n8187 , n8112 , n8113 );
xor ( n8188 , n8186 , n8187 );
and ( n8189 , n8188 , n5189 );
and ( n8190 , n4106 , n5283 );
or ( n8191 , n8189 , n8190 );
and ( n8192 , n8191 , n6725 );
or ( n8193 , n8131 , n8158 , n8169 , n8180 , n8184 , n8185 , n8192 );
and ( n8194 , n8130 , n8193 );
and ( n8195 , n4106 , n3260 );
or ( n8196 , n8194 , n8195 );
and ( n8197 , n8196 , n2422 );
and ( n8198 , n3881 , n2428 );
or ( n8199 , n8197 , n8198 );
buf ( n8200 , n8199 );
buf ( n8201 , n2424 );
buf ( n8202 , n2281 );
buf ( n8203 , n2280 );
not ( n8204 , n3260 );
and ( n8205 , n4096 , n3631 );
not ( n8206 , n7022 );
and ( n8207 , n8206 , n6900 );
xor ( n8208 , n6900 , n3770 );
and ( n8209 , n8134 , n8135 );
xor ( n8210 , n8208 , n8209 );
and ( n8211 , n8210 , n7022 );
or ( n8212 , n8207 , n8211 );
and ( n8213 , n8212 , n5290 );
and ( n8214 , n8212 , n5288 );
not ( n8215 , n3290 );
and ( n8216 , n8215 , n4825 );
not ( n8217 , n5000 );
and ( n8218 , n8217 , n4833 );
xor ( n8219 , n4833 , n4579 );
and ( n8220 , n8145 , n8146 );
xor ( n8221 , n8219 , n8220 );
and ( n8222 , n8221 , n5000 );
or ( n8223 , n8218 , n8222 );
and ( n8224 , n8223 , n3290 );
or ( n8225 , n8216 , n8224 );
and ( n8226 , n8225 , n5153 );
and ( n8227 , n4825 , n5155 );
or ( n8228 , n8213 , n8214 , n8226 , n8227 );
and ( n8229 , n8228 , n5189 );
and ( n8230 , n4096 , n5283 );
or ( n8231 , n8229 , n8230 );
and ( n8232 , n8231 , n5286 );
not ( n8233 , n6202 );
and ( n8234 , n8233 , n6056 );
xor ( n8235 , n6056 , n5853 );
and ( n8236 , n8161 , n8162 );
xor ( n8237 , n8235 , n8236 );
and ( n8238 , n8237 , n6202 );
or ( n8239 , n8234 , n8238 );
and ( n8240 , n8239 , n5189 );
and ( n8241 , n4096 , n5283 );
or ( n8242 , n8240 , n8241 );
and ( n8243 , n8242 , n6219 );
not ( n8244 , n6695 );
and ( n8245 , n8244 , n6549 );
xor ( n8246 , n6549 , n6346 );
and ( n8247 , n8172 , n8173 );
xor ( n8248 , n8246 , n8247 );
and ( n8249 , n8248 , n6695 );
or ( n8250 , n8245 , n8249 );
and ( n8251 , n8250 , n5189 );
and ( n8252 , n4096 , n5283 );
or ( n8253 , n8251 , n8252 );
and ( n8254 , n8253 , n6711 );
and ( n8255 , n5598 , n5189 );
and ( n8256 , n4096 , n5283 );
or ( n8257 , n8255 , n8256 );
and ( n8258 , n8257 , n6718 );
and ( n8259 , n5598 , n6720 );
not ( n8260 , n5598 );
and ( n8261 , n8186 , n8187 );
xor ( n8262 , n8260 , n8261 );
and ( n8263 , n8262 , n5189 );
and ( n8264 , n4096 , n5283 );
or ( n8265 , n8263 , n8264 );
and ( n8266 , n8265 , n6725 );
or ( n8267 , n8205 , n8232 , n8243 , n8254 , n8258 , n8259 , n8266 );
and ( n8268 , n8204 , n8267 );
and ( n8269 , n4096 , n3260 );
or ( n8270 , n8268 , n8269 );
and ( n8271 , n8270 , n2422 );
and ( n8272 , n3876 , n2428 );
or ( n8273 , n8271 , n8272 );
buf ( n8274 , n8273 );
buf ( n8275 , n2424 );
buf ( n8276 , n2281 );
buf ( n8277 , n2280 );
not ( n8278 , n3260 );
and ( n8279 , n4086 , n3631 );
not ( n8280 , n7022 );
and ( n8281 , n8280 , n6910 );
xor ( n8282 , n6910 , n3770 );
and ( n8283 , n8208 , n8209 );
xor ( n8284 , n8282 , n8283 );
and ( n8285 , n8284 , n7022 );
or ( n8286 , n8281 , n8285 );
and ( n8287 , n8286 , n5290 );
and ( n8288 , n8286 , n5288 );
not ( n8289 , n3290 );
and ( n8290 , n8289 , n4840 );
not ( n8291 , n5000 );
and ( n8292 , n8291 , n4848 );
xor ( n8293 , n4848 , n4579 );
and ( n8294 , n8219 , n8220 );
xor ( n8295 , n8293 , n8294 );
and ( n8296 , n8295 , n5000 );
or ( n8297 , n8292 , n8296 );
and ( n8298 , n8297 , n3290 );
or ( n8299 , n8290 , n8298 );
and ( n8300 , n8299 , n5153 );
and ( n8301 , n4840 , n5155 );
or ( n8302 , n8287 , n8288 , n8300 , n8301 );
and ( n8303 , n8302 , n5189 );
and ( n8304 , n4086 , n5283 );
or ( n8305 , n8303 , n8304 );
and ( n8306 , n8305 , n5286 );
not ( n8307 , n6202 );
and ( n8308 , n8307 , n6068 );
xor ( n8309 , n6068 , n5853 );
and ( n8310 , n8235 , n8236 );
xor ( n8311 , n8309 , n8310 );
and ( n8312 , n8311 , n6202 );
or ( n8313 , n8308 , n8312 );
and ( n8314 , n8313 , n5189 );
and ( n8315 , n4086 , n5283 );
or ( n8316 , n8314 , n8315 );
and ( n8317 , n8316 , n6219 );
not ( n8318 , n6695 );
and ( n8319 , n8318 , n6561 );
xor ( n8320 , n6561 , n6346 );
and ( n8321 , n8246 , n8247 );
xor ( n8322 , n8320 , n8321 );
and ( n8323 , n8322 , n6695 );
or ( n8324 , n8319 , n8323 );
and ( n8325 , n8324 , n5189 );
and ( n8326 , n4086 , n5283 );
or ( n8327 , n8325 , n8326 );
and ( n8328 , n8327 , n6711 );
and ( n8329 , n5588 , n5189 );
and ( n8330 , n4086 , n5283 );
or ( n8331 , n8329 , n8330 );
and ( n8332 , n8331 , n6718 );
and ( n8333 , n5588 , n6720 );
not ( n8334 , n5588 );
and ( n8335 , n8260 , n8261 );
xor ( n8336 , n8334 , n8335 );
and ( n8337 , n8336 , n5189 );
and ( n8338 , n4086 , n5283 );
or ( n8339 , n8337 , n8338 );
and ( n8340 , n8339 , n6725 );
or ( n8341 , n8279 , n8306 , n8317 , n8328 , n8332 , n8333 , n8340 );
and ( n8342 , n8278 , n8341 );
and ( n8343 , n4086 , n3260 );
or ( n8344 , n8342 , n8343 );
and ( n8345 , n8344 , n2422 );
and ( n8346 , n3871 , n2428 );
or ( n8347 , n8345 , n8346 );
buf ( n8348 , n8347 );
buf ( n8349 , n2424 );
buf ( n8350 , n2281 );
buf ( n8351 , n2280 );
not ( n8352 , n3260 );
and ( n8353 , n4076 , n3631 );
not ( n8354 , n7022 );
and ( n8355 , n8354 , n6920 );
xor ( n8356 , n6920 , n3770 );
and ( n8357 , n8282 , n8283 );
xor ( n8358 , n8356 , n8357 );
and ( n8359 , n8358 , n7022 );
or ( n8360 , n8355 , n8359 );
and ( n8361 , n8360 , n5290 );
and ( n8362 , n8360 , n5288 );
not ( n8363 , n3290 );
and ( n8364 , n8363 , n4855 );
not ( n8365 , n5000 );
and ( n8366 , n8365 , n4863 );
xor ( n8367 , n4863 , n4579 );
and ( n8368 , n8293 , n8294 );
xor ( n8369 , n8367 , n8368 );
and ( n8370 , n8369 , n5000 );
or ( n8371 , n8366 , n8370 );
and ( n8372 , n8371 , n3290 );
or ( n8373 , n8364 , n8372 );
and ( n8374 , n8373 , n5153 );
and ( n8375 , n4855 , n5155 );
or ( n8376 , n8361 , n8362 , n8374 , n8375 );
and ( n8377 , n8376 , n5189 );
and ( n8378 , n4076 , n5283 );
or ( n8379 , n8377 , n8378 );
and ( n8380 , n8379 , n5286 );
not ( n8381 , n6202 );
and ( n8382 , n8381 , n6080 );
xor ( n8383 , n6080 , n5853 );
and ( n8384 , n8309 , n8310 );
xor ( n8385 , n8383 , n8384 );
and ( n8386 , n8385 , n6202 );
or ( n8387 , n8382 , n8386 );
and ( n8388 , n8387 , n5189 );
and ( n8389 , n4076 , n5283 );
or ( n8390 , n8388 , n8389 );
and ( n8391 , n8390 , n6219 );
not ( n8392 , n6695 );
and ( n8393 , n8392 , n6573 );
xor ( n8394 , n6573 , n6346 );
and ( n8395 , n8320 , n8321 );
xor ( n8396 , n8394 , n8395 );
and ( n8397 , n8396 , n6695 );
or ( n8398 , n8393 , n8397 );
and ( n8399 , n8398 , n5189 );
and ( n8400 , n4076 , n5283 );
or ( n8401 , n8399 , n8400 );
and ( n8402 , n8401 , n6711 );
and ( n8403 , n5578 , n5189 );
and ( n8404 , n4076 , n5283 );
or ( n8405 , n8403 , n8404 );
and ( n8406 , n8405 , n6718 );
and ( n8407 , n5578 , n6720 );
not ( n8408 , n5578 );
and ( n8409 , n8334 , n8335 );
xor ( n8410 , n8408 , n8409 );
and ( n8411 , n8410 , n5189 );
and ( n8412 , n4076 , n5283 );
or ( n8413 , n8411 , n8412 );
and ( n8414 , n8413 , n6725 );
or ( n8415 , n8353 , n8380 , n8391 , n8402 , n8406 , n8407 , n8414 );
and ( n8416 , n8352 , n8415 );
and ( n8417 , n4076 , n3260 );
or ( n8418 , n8416 , n8417 );
and ( n8419 , n8418 , n2422 );
and ( n8420 , n3866 , n2428 );
or ( n8421 , n8419 , n8420 );
buf ( n8422 , n8421 );
buf ( n8423 , n2424 );
buf ( n8424 , n2281 );
buf ( n8425 , n2280 );
not ( n8426 , n3260 );
and ( n8427 , n4066 , n3631 );
not ( n8428 , n7022 );
and ( n8429 , n8428 , n6930 );
xor ( n8430 , n6930 , n3770 );
and ( n8431 , n8356 , n8357 );
xor ( n8432 , n8430 , n8431 );
and ( n8433 , n8432 , n7022 );
or ( n8434 , n8429 , n8433 );
and ( n8435 , n8434 , n5290 );
and ( n8436 , n8434 , n5288 );
not ( n8437 , n3290 );
and ( n8438 , n8437 , n4870 );
not ( n8439 , n5000 );
and ( n8440 , n8439 , n4878 );
xor ( n8441 , n4878 , n4579 );
and ( n8442 , n8367 , n8368 );
xor ( n8443 , n8441 , n8442 );
and ( n8444 , n8443 , n5000 );
or ( n8445 , n8440 , n8444 );
and ( n8446 , n8445 , n3290 );
or ( n8447 , n8438 , n8446 );
and ( n8448 , n8447 , n5153 );
and ( n8449 , n4870 , n5155 );
or ( n8450 , n8435 , n8436 , n8448 , n8449 );
and ( n8451 , n8450 , n5189 );
and ( n8452 , n4066 , n5283 );
or ( n8453 , n8451 , n8452 );
and ( n8454 , n8453 , n5286 );
not ( n8455 , n6202 );
and ( n8456 , n8455 , n6092 );
xor ( n8457 , n6092 , n5853 );
and ( n8458 , n8383 , n8384 );
xor ( n8459 , n8457 , n8458 );
and ( n8460 , n8459 , n6202 );
or ( n8461 , n8456 , n8460 );
and ( n8462 , n8461 , n5189 );
and ( n8463 , n4066 , n5283 );
or ( n8464 , n8462 , n8463 );
and ( n8465 , n8464 , n6219 );
not ( n8466 , n6695 );
and ( n8467 , n8466 , n6585 );
xor ( n8468 , n6585 , n6346 );
and ( n8469 , n8394 , n8395 );
xor ( n8470 , n8468 , n8469 );
and ( n8471 , n8470 , n6695 );
or ( n8472 , n8467 , n8471 );
and ( n8473 , n8472 , n5189 );
and ( n8474 , n4066 , n5283 );
or ( n8475 , n8473 , n8474 );
and ( n8476 , n8475 , n6711 );
and ( n8477 , n5530 , n5189 );
and ( n8478 , n4066 , n5283 );
or ( n8479 , n8477 , n8478 );
and ( n8480 , n8479 , n6718 );
and ( n8481 , n5530 , n6720 );
not ( n8482 , n5530 );
and ( n8483 , n8408 , n8409 );
xor ( n8484 , n8482 , n8483 );
and ( n8485 , n8484 , n5189 );
and ( n8486 , n4066 , n5283 );
or ( n8487 , n8485 , n8486 );
and ( n8488 , n8487 , n6725 );
or ( n8489 , n8427 , n8454 , n8465 , n8476 , n8480 , n8481 , n8488 );
and ( n8490 , n8426 , n8489 );
and ( n8491 , n4066 , n3260 );
or ( n8492 , n8490 , n8491 );
and ( n8493 , n8492 , n2422 );
and ( n8494 , n3861 , n2428 );
or ( n8495 , n8493 , n8494 );
buf ( n8496 , n8495 );
buf ( n8497 , n2424 );
buf ( n8498 , n2281 );
buf ( n8499 , n2280 );
not ( n8500 , n3260 );
and ( n8501 , n4056 , n3631 );
not ( n8502 , n7022 );
and ( n8503 , n8502 , n6940 );
xor ( n8504 , n6940 , n3770 );
and ( n8505 , n8430 , n8431 );
xor ( n8506 , n8504 , n8505 );
and ( n8507 , n8506 , n7022 );
or ( n8508 , n8503 , n8507 );
and ( n8509 , n8508 , n5290 );
and ( n8510 , n8508 , n5288 );
not ( n8511 , n3290 );
and ( n8512 , n8511 , n4885 );
not ( n8513 , n5000 );
and ( n8514 , n8513 , n4893 );
xor ( n8515 , n4893 , n4579 );
and ( n8516 , n8441 , n8442 );
xor ( n8517 , n8515 , n8516 );
and ( n8518 , n8517 , n5000 );
or ( n8519 , n8514 , n8518 );
and ( n8520 , n8519 , n3290 );
or ( n8521 , n8512 , n8520 );
and ( n8522 , n8521 , n5153 );
and ( n8523 , n4885 , n5155 );
or ( n8524 , n8509 , n8510 , n8522 , n8523 );
and ( n8525 , n8524 , n5189 );
and ( n8526 , n4056 , n5283 );
or ( n8527 , n8525 , n8526 );
and ( n8528 , n8527 , n5286 );
not ( n8529 , n6202 );
and ( n8530 , n8529 , n6104 );
xor ( n8531 , n6104 , n5853 );
and ( n8532 , n8457 , n8458 );
xor ( n8533 , n8531 , n8532 );
and ( n8534 , n8533 , n6202 );
or ( n8535 , n8530 , n8534 );
and ( n8536 , n8535 , n5189 );
and ( n8537 , n4056 , n5283 );
or ( n8538 , n8536 , n8537 );
and ( n8539 , n8538 , n6219 );
not ( n8540 , n6695 );
and ( n8541 , n8540 , n6597 );
xor ( n8542 , n6597 , n6346 );
and ( n8543 , n8468 , n8469 );
xor ( n8544 , n8542 , n8543 );
and ( n8545 , n8544 , n6695 );
or ( n8546 , n8541 , n8545 );
and ( n8547 , n8546 , n5189 );
and ( n8548 , n4056 , n5283 );
or ( n8549 , n8547 , n8548 );
and ( n8550 , n8549 , n6711 );
and ( n8551 , n5527 , n5189 );
and ( n8552 , n4056 , n5283 );
or ( n8553 , n8551 , n8552 );
and ( n8554 , n8553 , n6718 );
and ( n8555 , n5527 , n6720 );
not ( n8556 , n5527 );
and ( n8557 , n8482 , n8483 );
xor ( n8558 , n8556 , n8557 );
and ( n8559 , n8558 , n5189 );
and ( n8560 , n4056 , n5283 );
or ( n8561 , n8559 , n8560 );
and ( n8562 , n8561 , n6725 );
or ( n8563 , n8501 , n8528 , n8539 , n8550 , n8554 , n8555 , n8562 );
and ( n8564 , n8500 , n8563 );
and ( n8565 , n4056 , n3260 );
or ( n8566 , n8564 , n8565 );
and ( n8567 , n8566 , n2422 );
and ( n8568 , n3856 , n2428 );
or ( n8569 , n8567 , n8568 );
buf ( n8570 , n8569 );
buf ( n8571 , n2424 );
buf ( n8572 , n2281 );
buf ( n8573 , n2280 );
not ( n8574 , n3260 );
and ( n8575 , n4046 , n3631 );
not ( n8576 , n7022 );
and ( n8577 , n8576 , n6950 );
xor ( n8578 , n6950 , n3770 );
and ( n8579 , n8504 , n8505 );
xor ( n8580 , n8578 , n8579 );
and ( n8581 , n8580 , n7022 );
or ( n8582 , n8577 , n8581 );
and ( n8583 , n8582 , n5290 );
and ( n8584 , n8582 , n5288 );
not ( n8585 , n3290 );
and ( n8586 , n8585 , n4900 );
not ( n8587 , n5000 );
and ( n8588 , n8587 , n4908 );
xor ( n8589 , n4908 , n4579 );
and ( n8590 , n8515 , n8516 );
xor ( n8591 , n8589 , n8590 );
and ( n8592 , n8591 , n5000 );
or ( n8593 , n8588 , n8592 );
and ( n8594 , n8593 , n3290 );
or ( n8595 , n8586 , n8594 );
and ( n8596 , n8595 , n5153 );
and ( n8597 , n4900 , n5155 );
or ( n8598 , n8583 , n8584 , n8596 , n8597 );
and ( n8599 , n8598 , n5189 );
and ( n8600 , n4046 , n5283 );
or ( n8601 , n8599 , n8600 );
and ( n8602 , n8601 , n5286 );
not ( n8603 , n6202 );
and ( n8604 , n8603 , n6116 );
xor ( n8605 , n6116 , n5853 );
and ( n8606 , n8531 , n8532 );
xor ( n8607 , n8605 , n8606 );
and ( n8608 , n8607 , n6202 );
or ( n8609 , n8604 , n8608 );
and ( n8610 , n8609 , n5189 );
and ( n8611 , n4046 , n5283 );
or ( n8612 , n8610 , n8611 );
and ( n8613 , n8612 , n6219 );
not ( n8614 , n6695 );
and ( n8615 , n8614 , n6609 );
xor ( n8616 , n6609 , n6346 );
and ( n8617 , n8542 , n8543 );
xor ( n8618 , n8616 , n8617 );
and ( n8619 , n8618 , n6695 );
or ( n8620 , n8615 , n8619 );
and ( n8621 , n8620 , n5189 );
and ( n8622 , n4046 , n5283 );
or ( n8623 , n8621 , n8622 );
and ( n8624 , n8623 , n6711 );
and ( n8625 , n5524 , n5189 );
and ( n8626 , n4046 , n5283 );
or ( n8627 , n8625 , n8626 );
and ( n8628 , n8627 , n6718 );
and ( n8629 , n5524 , n6720 );
not ( n8630 , n5524 );
and ( n8631 , n8556 , n8557 );
xor ( n8632 , n8630 , n8631 );
and ( n8633 , n8632 , n5189 );
and ( n8634 , n4046 , n5283 );
or ( n8635 , n8633 , n8634 );
and ( n8636 , n8635 , n6725 );
or ( n8637 , n8575 , n8602 , n8613 , n8624 , n8628 , n8629 , n8636 );
and ( n8638 , n8574 , n8637 );
and ( n8639 , n4046 , n3260 );
or ( n8640 , n8638 , n8639 );
and ( n8641 , n8640 , n2422 );
and ( n8642 , n3851 , n2428 );
or ( n8643 , n8641 , n8642 );
buf ( n8644 , n8643 );
buf ( n8645 , n2424 );
buf ( n8646 , n2281 );
buf ( n8647 , n2280 );
not ( n8648 , n3260 );
and ( n8649 , n4036 , n3631 );
not ( n8650 , n7022 );
and ( n8651 , n8650 , n6960 );
xor ( n8652 , n6960 , n3770 );
and ( n8653 , n8578 , n8579 );
xor ( n8654 , n8652 , n8653 );
and ( n8655 , n8654 , n7022 );
or ( n8656 , n8651 , n8655 );
and ( n8657 , n8656 , n5290 );
and ( n8658 , n8656 , n5288 );
not ( n8659 , n3290 );
and ( n8660 , n8659 , n4915 );
not ( n8661 , n5000 );
and ( n8662 , n8661 , n4923 );
xor ( n8663 , n4923 , n4579 );
and ( n8664 , n8589 , n8590 );
xor ( n8665 , n8663 , n8664 );
and ( n8666 , n8665 , n5000 );
or ( n8667 , n8662 , n8666 );
and ( n8668 , n8667 , n3290 );
or ( n8669 , n8660 , n8668 );
and ( n8670 , n8669 , n5153 );
and ( n8671 , n4915 , n5155 );
or ( n8672 , n8657 , n8658 , n8670 , n8671 );
and ( n8673 , n8672 , n5189 );
and ( n8674 , n4036 , n5283 );
or ( n8675 , n8673 , n8674 );
and ( n8676 , n8675 , n5286 );
not ( n8677 , n6202 );
and ( n8678 , n8677 , n6128 );
xor ( n8679 , n6128 , n5853 );
and ( n8680 , n8605 , n8606 );
xor ( n8681 , n8679 , n8680 );
and ( n8682 , n8681 , n6202 );
or ( n8683 , n8678 , n8682 );
and ( n8684 , n8683 , n5189 );
and ( n8685 , n4036 , n5283 );
or ( n8686 , n8684 , n8685 );
and ( n8687 , n8686 , n6219 );
not ( n8688 , n6695 );
and ( n8689 , n8688 , n6621 );
xor ( n8690 , n6621 , n6346 );
and ( n8691 , n8616 , n8617 );
xor ( n8692 , n8690 , n8691 );
and ( n8693 , n8692 , n6695 );
or ( n8694 , n8689 , n8693 );
and ( n8695 , n8694 , n5189 );
and ( n8696 , n4036 , n5283 );
or ( n8697 , n8695 , n8696 );
and ( n8698 , n8697 , n6711 );
and ( n8699 , n5521 , n5189 );
and ( n8700 , n4036 , n5283 );
or ( n8701 , n8699 , n8700 );
and ( n8702 , n8701 , n6718 );
and ( n8703 , n5521 , n6720 );
not ( n8704 , n5521 );
and ( n8705 , n8630 , n8631 );
xor ( n8706 , n8704 , n8705 );
and ( n8707 , n8706 , n5189 );
and ( n8708 , n4036 , n5283 );
or ( n8709 , n8707 , n8708 );
and ( n8710 , n8709 , n6725 );
or ( n8711 , n8649 , n8676 , n8687 , n8698 , n8702 , n8703 , n8710 );
and ( n8712 , n8648 , n8711 );
and ( n8713 , n4036 , n3260 );
or ( n8714 , n8712 , n8713 );
and ( n8715 , n8714 , n2422 );
and ( n8716 , n3846 , n2428 );
or ( n8717 , n8715 , n8716 );
buf ( n8718 , n8717 );
buf ( n8719 , n2424 );
buf ( n8720 , n2281 );
buf ( n8721 , n2280 );
not ( n8722 , n3260 );
and ( n8723 , n4026 , n3631 );
not ( n8724 , n7022 );
and ( n8725 , n8724 , n6970 );
xor ( n8726 , n6970 , n3770 );
and ( n8727 , n8652 , n8653 );
xor ( n8728 , n8726 , n8727 );
and ( n8729 , n8728 , n7022 );
or ( n8730 , n8725 , n8729 );
and ( n8731 , n8730 , n5290 );
and ( n8732 , n8730 , n5288 );
not ( n8733 , n3290 );
and ( n8734 , n8733 , n4930 );
not ( n8735 , n5000 );
and ( n8736 , n8735 , n4938 );
xor ( n8737 , n4938 , n4579 );
and ( n8738 , n8663 , n8664 );
xor ( n8739 , n8737 , n8738 );
and ( n8740 , n8739 , n5000 );
or ( n8741 , n8736 , n8740 );
and ( n8742 , n8741 , n3290 );
or ( n8743 , n8734 , n8742 );
and ( n8744 , n8743 , n5153 );
and ( n8745 , n4930 , n5155 );
or ( n8746 , n8731 , n8732 , n8744 , n8745 );
and ( n8747 , n8746 , n5189 );
and ( n8748 , n4026 , n5283 );
or ( n8749 , n8747 , n8748 );
and ( n8750 , n8749 , n5286 );
not ( n8751 , n6202 );
and ( n8752 , n8751 , n6140 );
xor ( n8753 , n6140 , n5853 );
and ( n8754 , n8679 , n8680 );
xor ( n8755 , n8753 , n8754 );
and ( n8756 , n8755 , n6202 );
or ( n8757 , n8752 , n8756 );
and ( n8758 , n8757 , n5189 );
and ( n8759 , n4026 , n5283 );
or ( n8760 , n8758 , n8759 );
and ( n8761 , n8760 , n6219 );
not ( n8762 , n6695 );
and ( n8763 , n8762 , n6633 );
xor ( n8764 , n6633 , n6346 );
and ( n8765 , n8690 , n8691 );
xor ( n8766 , n8764 , n8765 );
and ( n8767 , n8766 , n6695 );
or ( n8768 , n8763 , n8767 );
and ( n8769 , n8768 , n5189 );
and ( n8770 , n4026 , n5283 );
or ( n8771 , n8769 , n8770 );
and ( n8772 , n8771 , n6711 );
and ( n8773 , n5518 , n5189 );
and ( n8774 , n4026 , n5283 );
or ( n8775 , n8773 , n8774 );
and ( n8776 , n8775 , n6718 );
and ( n8777 , n5518 , n6720 );
not ( n8778 , n5518 );
and ( n8779 , n8704 , n8705 );
xor ( n8780 , n8778 , n8779 );
and ( n8781 , n8780 , n5189 );
and ( n8782 , n4026 , n5283 );
or ( n8783 , n8781 , n8782 );
and ( n8784 , n8783 , n6725 );
or ( n8785 , n8723 , n8750 , n8761 , n8772 , n8776 , n8777 , n8784 );
and ( n8786 , n8722 , n8785 );
and ( n8787 , n4026 , n3260 );
or ( n8788 , n8786 , n8787 );
and ( n8789 , n8788 , n2422 );
and ( n8790 , n3841 , n2428 );
or ( n8791 , n8789 , n8790 );
buf ( n8792 , n8791 );
buf ( n8793 , n2424 );
buf ( n8794 , n2281 );
buf ( n8795 , n2280 );
not ( n8796 , n3260 );
and ( n8797 , n4016 , n3631 );
not ( n8798 , n7022 );
and ( n8799 , n8798 , n6980 );
xor ( n8800 , n6980 , n3770 );
and ( n8801 , n8726 , n8727 );
xor ( n8802 , n8800 , n8801 );
and ( n8803 , n8802 , n7022 );
or ( n8804 , n8799 , n8803 );
and ( n8805 , n8804 , n5290 );
and ( n8806 , n8804 , n5288 );
not ( n8807 , n3290 );
and ( n8808 , n8807 , n4945 );
not ( n8809 , n5000 );
and ( n8810 , n8809 , n4953 );
xor ( n8811 , n4953 , n4579 );
and ( n8812 , n8737 , n8738 );
xor ( n8813 , n8811 , n8812 );
and ( n8814 , n8813 , n5000 );
or ( n8815 , n8810 , n8814 );
and ( n8816 , n8815 , n3290 );
or ( n8817 , n8808 , n8816 );
and ( n8818 , n8817 , n5153 );
and ( n8819 , n4945 , n5155 );
or ( n8820 , n8805 , n8806 , n8818 , n8819 );
and ( n8821 , n8820 , n5189 );
and ( n8822 , n4016 , n5283 );
or ( n8823 , n8821 , n8822 );
and ( n8824 , n8823 , n5286 );
not ( n8825 , n6202 );
and ( n8826 , n8825 , n6152 );
xor ( n8827 , n6152 , n5853 );
and ( n8828 , n8753 , n8754 );
xor ( n8829 , n8827 , n8828 );
and ( n8830 , n8829 , n6202 );
or ( n8831 , n8826 , n8830 );
and ( n8832 , n8831 , n5189 );
and ( n8833 , n4016 , n5283 );
or ( n8834 , n8832 , n8833 );
and ( n8835 , n8834 , n6219 );
not ( n8836 , n6695 );
and ( n8837 , n8836 , n6645 );
xor ( n8838 , n6645 , n6346 );
and ( n8839 , n8764 , n8765 );
xor ( n8840 , n8838 , n8839 );
and ( n8841 , n8840 , n6695 );
or ( n8842 , n8837 , n8841 );
and ( n8843 , n8842 , n5189 );
and ( n8844 , n4016 , n5283 );
or ( n8845 , n8843 , n8844 );
and ( n8846 , n8845 , n6711 );
and ( n8847 , n5515 , n5189 );
and ( n8848 , n4016 , n5283 );
or ( n8849 , n8847 , n8848 );
and ( n8850 , n8849 , n6718 );
and ( n8851 , n5515 , n6720 );
not ( n8852 , n5515 );
and ( n8853 , n8778 , n8779 );
xor ( n8854 , n8852 , n8853 );
and ( n8855 , n8854 , n5189 );
and ( n8856 , n4016 , n5283 );
or ( n8857 , n8855 , n8856 );
and ( n8858 , n8857 , n6725 );
or ( n8859 , n8797 , n8824 , n8835 , n8846 , n8850 , n8851 , n8858 );
and ( n8860 , n8796 , n8859 );
and ( n8861 , n4016 , n3260 );
or ( n8862 , n8860 , n8861 );
and ( n8863 , n8862 , n2422 );
and ( n8864 , n3836 , n2428 );
or ( n8865 , n8863 , n8864 );
buf ( n8866 , n8865 );
buf ( n8867 , n2424 );
buf ( n8868 , n2281 );
buf ( n8869 , n2280 );
not ( n8870 , n3260 );
and ( n8871 , n4006 , n3631 );
not ( n8872 , n7022 );
and ( n8873 , n8872 , n6990 );
xor ( n8874 , n6990 , n3770 );
and ( n8875 , n8800 , n8801 );
xor ( n8876 , n8874 , n8875 );
and ( n8877 , n8876 , n7022 );
or ( n8878 , n8873 , n8877 );
and ( n8879 , n8878 , n5290 );
and ( n8880 , n8878 , n5288 );
not ( n8881 , n3290 );
and ( n8882 , n8881 , n4960 );
not ( n8883 , n5000 );
and ( n8884 , n8883 , n4968 );
xor ( n8885 , n4968 , n4579 );
and ( n8886 , n8811 , n8812 );
xor ( n8887 , n8885 , n8886 );
and ( n8888 , n8887 , n5000 );
or ( n8889 , n8884 , n8888 );
and ( n8890 , n8889 , n3290 );
or ( n8891 , n8882 , n8890 );
and ( n8892 , n8891 , n5153 );
and ( n8893 , n4960 , n5155 );
or ( n8894 , n8879 , n8880 , n8892 , n8893 );
and ( n8895 , n8894 , n5189 );
and ( n8896 , n4006 , n5283 );
or ( n8897 , n8895 , n8896 );
and ( n8898 , n8897 , n5286 );
not ( n8899 , n6202 );
and ( n8900 , n8899 , n6164 );
xor ( n8901 , n6164 , n5853 );
and ( n8902 , n8827 , n8828 );
xor ( n8903 , n8901 , n8902 );
and ( n8904 , n8903 , n6202 );
or ( n8905 , n8900 , n8904 );
and ( n8906 , n8905 , n5189 );
and ( n8907 , n4006 , n5283 );
or ( n8908 , n8906 , n8907 );
and ( n8909 , n8908 , n6219 );
not ( n8910 , n6695 );
and ( n8911 , n8910 , n6657 );
xor ( n8912 , n6657 , n6346 );
and ( n8913 , n8838 , n8839 );
xor ( n8914 , n8912 , n8913 );
and ( n8915 , n8914 , n6695 );
or ( n8916 , n8911 , n8915 );
and ( n8917 , n8916 , n5189 );
and ( n8918 , n4006 , n5283 );
or ( n8919 , n8917 , n8918 );
and ( n8920 , n8919 , n6711 );
and ( n8921 , n5512 , n5189 );
and ( n8922 , n4006 , n5283 );
or ( n8923 , n8921 , n8922 );
and ( n8924 , n8923 , n6718 );
and ( n8925 , n5512 , n6720 );
not ( n8926 , n5512 );
and ( n8927 , n8852 , n8853 );
xor ( n8928 , n8926 , n8927 );
and ( n8929 , n8928 , n5189 );
and ( n8930 , n4006 , n5283 );
or ( n8931 , n8929 , n8930 );
and ( n8932 , n8931 , n6725 );
or ( n8933 , n8871 , n8898 , n8909 , n8920 , n8924 , n8925 , n8932 );
and ( n8934 , n8870 , n8933 );
and ( n8935 , n4006 , n3260 );
or ( n8936 , n8934 , n8935 );
and ( n8937 , n8936 , n2422 );
and ( n8938 , n3831 , n2428 );
or ( n8939 , n8937 , n8938 );
buf ( n8940 , n8939 );
buf ( n8941 , n2424 );
buf ( n8942 , n2281 );
buf ( n8943 , n2280 );
not ( n8944 , n3260 );
and ( n8945 , n3996 , n3631 );
not ( n8946 , n7022 );
and ( n8947 , n8946 , n7000 );
xor ( n8948 , n7000 , n3770 );
and ( n8949 , n8874 , n8875 );
xor ( n8950 , n8948 , n8949 );
and ( n8951 , n8950 , n7022 );
or ( n8952 , n8947 , n8951 );
and ( n8953 , n8952 , n5290 );
and ( n8954 , n8952 , n5288 );
not ( n8955 , n3290 );
and ( n8956 , n8955 , n4975 );
not ( n8957 , n5000 );
and ( n8958 , n8957 , n4983 );
xor ( n8959 , n4983 , n4579 );
and ( n8960 , n8885 , n8886 );
xor ( n8961 , n8959 , n8960 );
and ( n8962 , n8961 , n5000 );
or ( n8963 , n8958 , n8962 );
and ( n8964 , n8963 , n3290 );
or ( n8965 , n8956 , n8964 );
and ( n8966 , n8965 , n5153 );
and ( n8967 , n4975 , n5155 );
or ( n8968 , n8953 , n8954 , n8966 , n8967 );
and ( n8969 , n8968 , n5189 );
and ( n8970 , n3996 , n5283 );
or ( n8971 , n8969 , n8970 );
and ( n8972 , n8971 , n5286 );
not ( n8973 , n6202 );
and ( n8974 , n8973 , n6176 );
xor ( n8975 , n6176 , n5853 );
and ( n8976 , n8901 , n8902 );
xor ( n8977 , n8975 , n8976 );
and ( n8978 , n8977 , n6202 );
or ( n8979 , n8974 , n8978 );
and ( n8980 , n8979 , n5189 );
and ( n8981 , n3996 , n5283 );
or ( n8982 , n8980 , n8981 );
and ( n8983 , n8982 , n6219 );
not ( n8984 , n6695 );
and ( n8985 , n8984 , n6669 );
xor ( n8986 , n6669 , n6346 );
and ( n8987 , n8912 , n8913 );
xor ( n8988 , n8986 , n8987 );
and ( n8989 , n8988 , n6695 );
or ( n8990 , n8985 , n8989 );
and ( n8991 , n8990 , n5189 );
and ( n8992 , n3996 , n5283 );
or ( n8993 , n8991 , n8992 );
and ( n8994 , n8993 , n6711 );
and ( n8995 , n5509 , n5189 );
and ( n8996 , n3996 , n5283 );
or ( n8997 , n8995 , n8996 );
and ( n8998 , n8997 , n6718 );
and ( n8999 , n5509 , n6720 );
not ( n9000 , n5509 );
and ( n9001 , n8926 , n8927 );
xor ( n9002 , n9000 , n9001 );
and ( n9003 , n9002 , n5189 );
and ( n9004 , n3996 , n5283 );
or ( n9005 , n9003 , n9004 );
and ( n9006 , n9005 , n6725 );
or ( n9007 , n8945 , n8972 , n8983 , n8994 , n8998 , n8999 , n9006 );
and ( n9008 , n8944 , n9007 );
and ( n9009 , n3996 , n3260 );
or ( n9010 , n9008 , n9009 );
and ( n9011 , n9010 , n2422 );
and ( n9012 , n3826 , n2428 );
or ( n9013 , n9011 , n9012 );
buf ( n9014 , n9013 );
buf ( n9015 , n2424 );
buf ( n9016 , n2281 );
buf ( n9017 , n2280 );
not ( n9018 , n3260 );
and ( n9019 , n3986 , n3631 );
not ( n9020 , n7022 );
and ( n9021 , n9020 , n7010 );
xor ( n9022 , n7010 , n3770 );
and ( n9023 , n8948 , n8949 );
xor ( n9024 , n9022 , n9023 );
and ( n9025 , n9024 , n7022 );
or ( n9026 , n9021 , n9025 );
and ( n9027 , n9026 , n5290 );
and ( n9028 , n9026 , n5288 );
not ( n9029 , n3290 );
and ( n9030 , n9029 , n4990 );
not ( n9031 , n5000 );
and ( n9032 , n9031 , n4998 );
xor ( n9033 , n4998 , n4579 );
and ( n9034 , n8959 , n8960 );
xor ( n9035 , n9033 , n9034 );
and ( n9036 , n9035 , n5000 );
or ( n9037 , n9032 , n9036 );
and ( n9038 , n9037 , n3290 );
or ( n9039 , n9030 , n9038 );
and ( n9040 , n9039 , n5153 );
and ( n9041 , n4990 , n5155 );
or ( n9042 , n9027 , n9028 , n9040 , n9041 );
and ( n9043 , n9042 , n5189 );
and ( n9044 , n3986 , n5283 );
or ( n9045 , n9043 , n9044 );
and ( n9046 , n9045 , n5286 );
not ( n9047 , n6202 );
and ( n9048 , n9047 , n6188 );
xor ( n9049 , n6188 , n5853 );
and ( n9050 , n8975 , n8976 );
xor ( n9051 , n9049 , n9050 );
and ( n9052 , n9051 , n6202 );
or ( n9053 , n9048 , n9052 );
and ( n9054 , n9053 , n5189 );
and ( n9055 , n3986 , n5283 );
or ( n9056 , n9054 , n9055 );
and ( n9057 , n9056 , n6219 );
not ( n9058 , n6695 );
and ( n9059 , n9058 , n6681 );
xor ( n9060 , n6681 , n6346 );
and ( n9061 , n8986 , n8987 );
xor ( n9062 , n9060 , n9061 );
and ( n9063 , n9062 , n6695 );
or ( n9064 , n9059 , n9063 );
and ( n9065 , n9064 , n5189 );
and ( n9066 , n3986 , n5283 );
or ( n9067 , n9065 , n9066 );
and ( n9068 , n9067 , n6711 );
and ( n9069 , n5506 , n5189 );
and ( n9070 , n3986 , n5283 );
or ( n9071 , n9069 , n9070 );
and ( n9072 , n9071 , n6718 );
and ( n9073 , n5506 , n6720 );
not ( n9074 , n5506 );
and ( n9075 , n9000 , n9001 );
xor ( n9076 , n9074 , n9075 );
and ( n9077 , n9076 , n5189 );
and ( n9078 , n3986 , n5283 );
or ( n9079 , n9077 , n9078 );
and ( n9080 , n9079 , n6725 );
or ( n9081 , n9019 , n9046 , n9057 , n9068 , n9072 , n9073 , n9080 );
and ( n9082 , n9018 , n9081 );
and ( n9083 , n3986 , n3260 );
or ( n9084 , n9082 , n9083 );
and ( n9085 , n9084 , n2422 );
and ( n9086 , n3821 , n2428 );
or ( n9087 , n9085 , n9086 );
buf ( n9088 , n9087 );
buf ( n9089 , n2424 );
buf ( n9090 , n2281 );
buf ( n9091 , n2280 );
not ( n9092 , n3260 );
and ( n9093 , n5157 , n5220 );
or ( n9094 , n5250 , n5281 );
or ( n9095 , n9094 , n5189 );
buf ( n9096 , n9095 );
and ( n9097 , n3791 , n9096 );
or ( n9098 , n9093 , n9097 );
and ( n9099 , n9098 , n5286 );
and ( n9100 , n6208 , n5220 );
and ( n9101 , n3791 , n9096 );
or ( n9102 , n9100 , n9101 );
and ( n9103 , n9102 , n6219 );
and ( n9104 , n6701 , n5220 );
and ( n9105 , n3791 , n9096 );
or ( n9106 , n9104 , n9105 );
and ( n9107 , n9106 , n6711 );
and ( n9108 , n5493 , n5220 );
and ( n9109 , n3791 , n9096 );
or ( n9110 , n9108 , n9109 );
and ( n9111 , n9110 , n6718 );
and ( n9112 , n5493 , n5220 );
and ( n9113 , n3791 , n9096 );
or ( n9114 , n9112 , n9113 );
and ( n9115 , n9114 , n6725 );
or ( n9116 , n6720 , n3631 );
and ( n9117 , n3791 , n9116 );
or ( n9118 , n9099 , n9103 , n9107 , n9111 , n9115 , n9117 );
and ( n9119 , n9092 , n9118 );
and ( n9120 , n3791 , n3260 );
or ( n9121 , n9119 , n9120 );
and ( n9122 , n9121 , n2422 );
and ( n9123 , n3791 , n2428 );
or ( n9124 , n9122 , n9123 );
buf ( n9125 , n9124 );
buf ( n9126 , n2424 );
buf ( n9127 , n2281 );
buf ( n9128 , n2280 );
not ( n9129 , n3260 );
and ( n9130 , n7044 , n5220 );
and ( n9131 , n3781 , n9096 );
or ( n9132 , n9130 , n9131 );
and ( n9133 , n9132 , n5286 );
and ( n9134 , n7055 , n5220 );
and ( n9135 , n3781 , n9096 );
or ( n9136 , n9134 , n9135 );
and ( n9137 , n9136 , n6219 );
and ( n9138 , n7066 , n5220 );
and ( n9139 , n3781 , n9096 );
or ( n9140 , n9138 , n9139 );
and ( n9141 , n9140 , n6711 );
and ( n9142 , n5758 , n5220 );
and ( n9143 , n3781 , n9096 );
or ( n9144 , n9142 , n9143 );
and ( n9145 , n9144 , n6718 );
and ( n9146 , n7078 , n5220 );
and ( n9147 , n3781 , n9096 );
or ( n9148 , n9146 , n9147 );
and ( n9149 , n9148 , n6725 );
and ( n9150 , n3781 , n9116 );
or ( n9151 , n9133 , n9137 , n9141 , n9145 , n9149 , n9150 );
and ( n9152 , n9129 , n9151 );
and ( n9153 , n3781 , n3260 );
or ( n9154 , n9152 , n9153 );
and ( n9155 , n9154 , n2422 );
and ( n9156 , n3781 , n2428 );
or ( n9157 , n9155 , n9156 );
buf ( n9158 , n9157 );
buf ( n9159 , n2424 );
buf ( n9160 , n2281 );
buf ( n9161 , n2280 );
not ( n9162 , n3260 );
and ( n9163 , n7118 , n5220 );
and ( n9164 , n4254 , n9096 );
or ( n9165 , n9163 , n9164 );
and ( n9166 , n9165 , n5286 );
and ( n9167 , n7129 , n5220 );
and ( n9168 , n4254 , n9096 );
or ( n9169 , n9167 , n9168 );
and ( n9170 , n9169 , n6219 );
and ( n9171 , n7140 , n5220 );
and ( n9172 , n4254 , n9096 );
or ( n9173 , n9171 , n9172 );
and ( n9174 , n9173 , n6711 );
and ( n9175 , n5748 , n5220 );
and ( n9176 , n4254 , n9096 );
or ( n9177 , n9175 , n9176 );
and ( n9178 , n9177 , n6718 );
and ( n9179 , n7152 , n5220 );
and ( n9180 , n4254 , n9096 );
or ( n9181 , n9179 , n9180 );
and ( n9182 , n9181 , n6725 );
and ( n9183 , n4254 , n9116 );
or ( n9184 , n9166 , n9170 , n9174 , n9178 , n9182 , n9183 );
and ( n9185 , n9162 , n9184 );
and ( n9186 , n4254 , n3260 );
or ( n9187 , n9185 , n9186 );
and ( n9188 , n9187 , n2422 );
and ( n9189 , n4254 , n2428 );
or ( n9190 , n9188 , n9189 );
buf ( n9191 , n9190 );
buf ( n9192 , n2424 );
buf ( n9193 , n2281 );
buf ( n9194 , n2280 );
not ( n9195 , n3260 );
and ( n9196 , n7192 , n5220 );
and ( n9197 , n4240 , n9096 );
or ( n9198 , n9196 , n9197 );
and ( n9199 , n9198 , n5286 );
and ( n9200 , n7203 , n5220 );
and ( n9201 , n4240 , n9096 );
or ( n9202 , n9200 , n9201 );
and ( n9203 , n9202 , n6219 );
and ( n9204 , n7214 , n5220 );
and ( n9205 , n4240 , n9096 );
or ( n9206 , n9204 , n9205 );
and ( n9207 , n9206 , n6711 );
and ( n9208 , n5738 , n5220 );
and ( n9209 , n4240 , n9096 );
or ( n9210 , n9208 , n9209 );
and ( n9211 , n9210 , n6718 );
and ( n9212 , n7226 , n5220 );
and ( n9213 , n4240 , n9096 );
or ( n9214 , n9212 , n9213 );
and ( n9215 , n9214 , n6725 );
and ( n9216 , n4240 , n9116 );
or ( n9217 , n9199 , n9203 , n9207 , n9211 , n9215 , n9216 );
and ( n9218 , n9195 , n9217 );
and ( n9219 , n4240 , n3260 );
or ( n9220 , n9218 , n9219 );
and ( n9221 , n9220 , n2422 );
and ( n9222 , n4240 , n2428 );
or ( n9223 , n9221 , n9222 );
buf ( n9224 , n9223 );
buf ( n9225 , n2424 );
buf ( n9226 , n2281 );
buf ( n9227 , n2280 );
not ( n9228 , n3260 );
and ( n9229 , n7266 , n5220 );
and ( n9230 , n4230 , n9096 );
or ( n9231 , n9229 , n9230 );
and ( n9232 , n9231 , n5286 );
and ( n9233 , n7277 , n5220 );
and ( n9234 , n4230 , n9096 );
or ( n9235 , n9233 , n9234 );
and ( n9236 , n9235 , n6219 );
and ( n9237 , n7288 , n5220 );
and ( n9238 , n4230 , n9096 );
or ( n9239 , n9237 , n9238 );
and ( n9240 , n9239 , n6711 );
and ( n9241 , n5728 , n5220 );
and ( n9242 , n4230 , n9096 );
or ( n9243 , n9241 , n9242 );
and ( n9244 , n9243 , n6718 );
and ( n9245 , n7300 , n5220 );
and ( n9246 , n4230 , n9096 );
or ( n9247 , n9245 , n9246 );
and ( n9248 , n9247 , n6725 );
and ( n9249 , n4230 , n9116 );
or ( n9250 , n9232 , n9236 , n9240 , n9244 , n9248 , n9249 );
and ( n9251 , n9228 , n9250 );
and ( n9252 , n4230 , n3260 );
or ( n9253 , n9251 , n9252 );
and ( n9254 , n9253 , n2422 );
and ( n9255 , n4230 , n2428 );
or ( n9256 , n9254 , n9255 );
buf ( n9257 , n9256 );
buf ( n9258 , n2424 );
buf ( n9259 , n2281 );
buf ( n9260 , n2280 );
not ( n9261 , n3260 );
and ( n9262 , n7340 , n5220 );
and ( n9263 , n4220 , n9096 );
or ( n9264 , n9262 , n9263 );
and ( n9265 , n9264 , n5286 );
and ( n9266 , n7351 , n5220 );
and ( n9267 , n4220 , n9096 );
or ( n9268 , n9266 , n9267 );
and ( n9269 , n9268 , n6219 );
and ( n9270 , n7362 , n5220 );
and ( n9271 , n4220 , n9096 );
or ( n9272 , n9270 , n9271 );
and ( n9273 , n9272 , n6711 );
and ( n9274 , n5718 , n5220 );
and ( n9275 , n4220 , n9096 );
or ( n9276 , n9274 , n9275 );
and ( n9277 , n9276 , n6718 );
and ( n9278 , n7374 , n5220 );
and ( n9279 , n4220 , n9096 );
or ( n9280 , n9278 , n9279 );
and ( n9281 , n9280 , n6725 );
and ( n9282 , n4220 , n9116 );
or ( n9283 , n9265 , n9269 , n9273 , n9277 , n9281 , n9282 );
and ( n9284 , n9261 , n9283 );
and ( n9285 , n4220 , n3260 );
or ( n9286 , n9284 , n9285 );
and ( n9287 , n9286 , n2422 );
and ( n9288 , n4220 , n2428 );
or ( n9289 , n9287 , n9288 );
buf ( n9290 , n9289 );
buf ( n9291 , n2424 );
buf ( n9292 , n2281 );
buf ( n9293 , n2280 );
not ( n9294 , n3260 );
and ( n9295 , n7414 , n5220 );
and ( n9296 , n4210 , n9096 );
or ( n9297 , n9295 , n9296 );
and ( n9298 , n9297 , n5286 );
and ( n9299 , n7425 , n5220 );
and ( n9300 , n4210 , n9096 );
or ( n9301 , n9299 , n9300 );
and ( n9302 , n9301 , n6219 );
and ( n9303 , n7436 , n5220 );
and ( n9304 , n4210 , n9096 );
or ( n9305 , n9303 , n9304 );
and ( n9306 , n9305 , n6711 );
and ( n9307 , n5708 , n5220 );
and ( n9308 , n4210 , n9096 );
or ( n9309 , n9307 , n9308 );
and ( n9310 , n9309 , n6718 );
and ( n9311 , n7448 , n5220 );
and ( n9312 , n4210 , n9096 );
or ( n9313 , n9311 , n9312 );
and ( n9314 , n9313 , n6725 );
and ( n9315 , n4210 , n9116 );
or ( n9316 , n9298 , n9302 , n9306 , n9310 , n9314 , n9315 );
and ( n9317 , n9294 , n9316 );
and ( n9318 , n4210 , n3260 );
or ( n9319 , n9317 , n9318 );
and ( n9320 , n9319 , n2422 );
and ( n9321 , n4210 , n2428 );
or ( n9322 , n9320 , n9321 );
buf ( n9323 , n9322 );
buf ( n9324 , n2424 );
buf ( n9325 , n2281 );
buf ( n9326 , n2280 );
not ( n9327 , n3260 );
and ( n9328 , n7488 , n5220 );
and ( n9329 , n4200 , n9096 );
or ( n9330 , n9328 , n9329 );
and ( n9331 , n9330 , n5286 );
and ( n9332 , n7499 , n5220 );
and ( n9333 , n4200 , n9096 );
or ( n9334 , n9332 , n9333 );
and ( n9335 , n9334 , n6219 );
and ( n9336 , n7510 , n5220 );
and ( n9337 , n4200 , n9096 );
or ( n9338 , n9336 , n9337 );
and ( n9339 , n9338 , n6711 );
and ( n9340 , n5698 , n5220 );
and ( n9341 , n4200 , n9096 );
or ( n9342 , n9340 , n9341 );
and ( n9343 , n9342 , n6718 );
and ( n9344 , n7522 , n5220 );
and ( n9345 , n4200 , n9096 );
or ( n9346 , n9344 , n9345 );
and ( n9347 , n9346 , n6725 );
and ( n9348 , n4200 , n9116 );
or ( n9349 , n9331 , n9335 , n9339 , n9343 , n9347 , n9348 );
and ( n9350 , n9327 , n9349 );
and ( n9351 , n4200 , n3260 );
or ( n9352 , n9350 , n9351 );
and ( n9353 , n9352 , n2422 );
and ( n9354 , n4200 , n2428 );
or ( n9355 , n9353 , n9354 );
buf ( n9356 , n9355 );
buf ( n9357 , n2424 );
buf ( n9358 , n2281 );
buf ( n9359 , n2280 );
not ( n9360 , n3260 );
and ( n9361 , n7562 , n5220 );
and ( n9362 , n4190 , n9096 );
or ( n9363 , n9361 , n9362 );
and ( n9364 , n9363 , n5286 );
and ( n9365 , n7573 , n5220 );
and ( n9366 , n4190 , n9096 );
or ( n9367 , n9365 , n9366 );
and ( n9368 , n9367 , n6219 );
and ( n9369 , n7584 , n5220 );
and ( n9370 , n4190 , n9096 );
or ( n9371 , n9369 , n9370 );
and ( n9372 , n9371 , n6711 );
and ( n9373 , n5688 , n5220 );
and ( n9374 , n4190 , n9096 );
or ( n9375 , n9373 , n9374 );
and ( n9376 , n9375 , n6718 );
and ( n9377 , n7596 , n5220 );
and ( n9378 , n4190 , n9096 );
or ( n9379 , n9377 , n9378 );
and ( n9380 , n9379 , n6725 );
and ( n9381 , n4190 , n9116 );
or ( n9382 , n9364 , n9368 , n9372 , n9376 , n9380 , n9381 );
and ( n9383 , n9360 , n9382 );
and ( n9384 , n4190 , n3260 );
or ( n9385 , n9383 , n9384 );
and ( n9386 , n9385 , n2422 );
and ( n9387 , n4190 , n2428 );
or ( n9388 , n9386 , n9387 );
buf ( n9389 , n9388 );
buf ( n9390 , n2424 );
buf ( n9391 , n2281 );
buf ( n9392 , n2280 );
not ( n9393 , n3260 );
and ( n9394 , n7636 , n5220 );
and ( n9395 , n4180 , n9096 );
or ( n9396 , n9394 , n9395 );
and ( n9397 , n9396 , n5286 );
and ( n9398 , n7647 , n5220 );
and ( n9399 , n4180 , n9096 );
or ( n9400 , n9398 , n9399 );
and ( n9401 , n9400 , n6219 );
and ( n9402 , n7658 , n5220 );
and ( n9403 , n4180 , n9096 );
or ( n9404 , n9402 , n9403 );
and ( n9405 , n9404 , n6711 );
and ( n9406 , n5678 , n5220 );
and ( n9407 , n4180 , n9096 );
or ( n9408 , n9406 , n9407 );
and ( n9409 , n9408 , n6718 );
and ( n9410 , n7670 , n5220 );
and ( n9411 , n4180 , n9096 );
or ( n9412 , n9410 , n9411 );
and ( n9413 , n9412 , n6725 );
and ( n9414 , n4180 , n9116 );
or ( n9415 , n9397 , n9401 , n9405 , n9409 , n9413 , n9414 );
and ( n9416 , n9393 , n9415 );
and ( n9417 , n4180 , n3260 );
or ( n9418 , n9416 , n9417 );
and ( n9419 , n9418 , n2422 );
and ( n9420 , n4180 , n2428 );
or ( n9421 , n9419 , n9420 );
buf ( n9422 , n9421 );
buf ( n9423 , n2424 );
buf ( n9424 , n2281 );
buf ( n9425 , n2280 );
not ( n9426 , n3260 );
and ( n9427 , n7710 , n5220 );
and ( n9428 , n4170 , n9096 );
or ( n9429 , n9427 , n9428 );
and ( n9430 , n9429 , n5286 );
and ( n9431 , n7721 , n5220 );
and ( n9432 , n4170 , n9096 );
or ( n9433 , n9431 , n9432 );
and ( n9434 , n9433 , n6219 );
and ( n9435 , n7732 , n5220 );
and ( n9436 , n4170 , n9096 );
or ( n9437 , n9435 , n9436 );
and ( n9438 , n9437 , n6711 );
and ( n9439 , n5668 , n5220 );
and ( n9440 , n4170 , n9096 );
or ( n9441 , n9439 , n9440 );
and ( n9442 , n9441 , n6718 );
and ( n9443 , n7744 , n5220 );
and ( n9444 , n4170 , n9096 );
or ( n9445 , n9443 , n9444 );
and ( n9446 , n9445 , n6725 );
and ( n9447 , n4170 , n9116 );
or ( n9448 , n9430 , n9434 , n9438 , n9442 , n9446 , n9447 );
and ( n9449 , n9426 , n9448 );
and ( n9450 , n4170 , n3260 );
or ( n9451 , n9449 , n9450 );
and ( n9452 , n9451 , n2422 );
and ( n9453 , n4170 , n2428 );
or ( n9454 , n9452 , n9453 );
buf ( n9455 , n9454 );
buf ( n9456 , n2424 );
buf ( n9457 , n2281 );
buf ( n9458 , n2280 );
not ( n9459 , n3260 );
and ( n9460 , n7784 , n5220 );
and ( n9461 , n4160 , n9096 );
or ( n9462 , n9460 , n9461 );
and ( n9463 , n9462 , n5286 );
and ( n9464 , n7795 , n5220 );
and ( n9465 , n4160 , n9096 );
or ( n9466 , n9464 , n9465 );
and ( n9467 , n9466 , n6219 );
and ( n9468 , n7806 , n5220 );
and ( n9469 , n4160 , n9096 );
or ( n9470 , n9468 , n9469 );
and ( n9471 , n9470 , n6711 );
and ( n9472 , n5658 , n5220 );
and ( n9473 , n4160 , n9096 );
or ( n9474 , n9472 , n9473 );
and ( n9475 , n9474 , n6718 );
and ( n9476 , n7818 , n5220 );
and ( n9477 , n4160 , n9096 );
or ( n9478 , n9476 , n9477 );
and ( n9479 , n9478 , n6725 );
and ( n9480 , n4160 , n9116 );
or ( n9481 , n9463 , n9467 , n9471 , n9475 , n9479 , n9480 );
and ( n9482 , n9459 , n9481 );
and ( n9483 , n4160 , n3260 );
or ( n9484 , n9482 , n9483 );
and ( n9485 , n9484 , n2422 );
and ( n9486 , n4160 , n2428 );
or ( n9487 , n9485 , n9486 );
buf ( n9488 , n9487 );
buf ( n9489 , n2424 );
buf ( n9490 , n2281 );
buf ( n9491 , n2280 );
not ( n9492 , n3260 );
and ( n9493 , n7858 , n5220 );
and ( n9494 , n4150 , n9096 );
or ( n9495 , n9493 , n9494 );
and ( n9496 , n9495 , n5286 );
and ( n9497 , n7869 , n5220 );
and ( n9498 , n4150 , n9096 );
or ( n9499 , n9497 , n9498 );
and ( n9500 , n9499 , n6219 );
and ( n9501 , n7880 , n5220 );
and ( n9502 , n4150 , n9096 );
or ( n9503 , n9501 , n9502 );
and ( n9504 , n9503 , n6711 );
and ( n9505 , n5648 , n5220 );
and ( n9506 , n4150 , n9096 );
or ( n9507 , n9505 , n9506 );
and ( n9508 , n9507 , n6718 );
and ( n9509 , n7892 , n5220 );
and ( n9510 , n4150 , n9096 );
or ( n9511 , n9509 , n9510 );
and ( n9512 , n9511 , n6725 );
and ( n9513 , n4150 , n9116 );
or ( n9514 , n9496 , n9500 , n9504 , n9508 , n9512 , n9513 );
and ( n9515 , n9492 , n9514 );
and ( n9516 , n4150 , n3260 );
or ( n9517 , n9515 , n9516 );
and ( n9518 , n9517 , n2422 );
and ( n9519 , n4150 , n2428 );
or ( n9520 , n9518 , n9519 );
buf ( n9521 , n9520 );
buf ( n9522 , n2424 );
buf ( n9523 , n2281 );
buf ( n9524 , n2280 );
not ( n9525 , n3260 );
and ( n9526 , n7932 , n5220 );
and ( n9527 , n4140 , n9096 );
or ( n9528 , n9526 , n9527 );
and ( n9529 , n9528 , n5286 );
and ( n9530 , n7943 , n5220 );
and ( n9531 , n4140 , n9096 );
or ( n9532 , n9530 , n9531 );
and ( n9533 , n9532 , n6219 );
and ( n9534 , n7954 , n5220 );
and ( n9535 , n4140 , n9096 );
or ( n9536 , n9534 , n9535 );
and ( n9537 , n9536 , n6711 );
and ( n9538 , n5638 , n5220 );
and ( n9539 , n4140 , n9096 );
or ( n9540 , n9538 , n9539 );
and ( n9541 , n9540 , n6718 );
and ( n9542 , n7966 , n5220 );
and ( n9543 , n4140 , n9096 );
or ( n9544 , n9542 , n9543 );
and ( n9545 , n9544 , n6725 );
and ( n9546 , n4140 , n9116 );
or ( n9547 , n9529 , n9533 , n9537 , n9541 , n9545 , n9546 );
and ( n9548 , n9525 , n9547 );
and ( n9549 , n4140 , n3260 );
or ( n9550 , n9548 , n9549 );
and ( n9551 , n9550 , n2422 );
and ( n9552 , n4140 , n2428 );
or ( n9553 , n9551 , n9552 );
buf ( n9554 , n9553 );
buf ( n9555 , n2424 );
buf ( n9556 , n2281 );
buf ( n9557 , n2280 );
not ( n9558 , n3260 );
and ( n9559 , n8006 , n5220 );
and ( n9560 , n4130 , n9096 );
or ( n9561 , n9559 , n9560 );
and ( n9562 , n9561 , n5286 );
and ( n9563 , n8017 , n5220 );
and ( n9564 , n4130 , n9096 );
or ( n9565 , n9563 , n9564 );
and ( n9566 , n9565 , n6219 );
and ( n9567 , n8028 , n5220 );
and ( n9568 , n4130 , n9096 );
or ( n9569 , n9567 , n9568 );
and ( n9570 , n9569 , n6711 );
and ( n9571 , n5628 , n5220 );
and ( n9572 , n4130 , n9096 );
or ( n9573 , n9571 , n9572 );
and ( n9574 , n9573 , n6718 );
and ( n9575 , n8040 , n5220 );
and ( n9576 , n4130 , n9096 );
or ( n9577 , n9575 , n9576 );
and ( n9578 , n9577 , n6725 );
and ( n9579 , n4130 , n9116 );
or ( n9580 , n9562 , n9566 , n9570 , n9574 , n9578 , n9579 );
and ( n9581 , n9558 , n9580 );
and ( n9582 , n4130 , n3260 );
or ( n9583 , n9581 , n9582 );
and ( n9584 , n9583 , n2422 );
and ( n9585 , n4130 , n2428 );
or ( n9586 , n9584 , n9585 );
buf ( n9587 , n9586 );
buf ( n9588 , n2424 );
buf ( n9589 , n2281 );
buf ( n9590 , n2280 );
not ( n9591 , n3260 );
and ( n9592 , n8080 , n5220 );
and ( n9593 , n4120 , n9096 );
or ( n9594 , n9592 , n9593 );
and ( n9595 , n9594 , n5286 );
and ( n9596 , n8091 , n5220 );
and ( n9597 , n4120 , n9096 );
or ( n9598 , n9596 , n9597 );
and ( n9599 , n9598 , n6219 );
and ( n9600 , n8102 , n5220 );
and ( n9601 , n4120 , n9096 );
or ( n9602 , n9600 , n9601 );
and ( n9603 , n9602 , n6711 );
and ( n9604 , n5618 , n5220 );
and ( n9605 , n4120 , n9096 );
or ( n9606 , n9604 , n9605 );
and ( n9607 , n9606 , n6718 );
and ( n9608 , n8114 , n5220 );
and ( n9609 , n4120 , n9096 );
or ( n9610 , n9608 , n9609 );
and ( n9611 , n9610 , n6725 );
and ( n9612 , n4120 , n9116 );
or ( n9613 , n9595 , n9599 , n9603 , n9607 , n9611 , n9612 );
and ( n9614 , n9591 , n9613 );
and ( n9615 , n4120 , n3260 );
or ( n9616 , n9614 , n9615 );
and ( n9617 , n9616 , n2422 );
and ( n9618 , n4120 , n2428 );
or ( n9619 , n9617 , n9618 );
buf ( n9620 , n9619 );
buf ( n9621 , n2424 );
buf ( n9622 , n2281 );
buf ( n9623 , n2280 );
not ( n9624 , n3260 );
and ( n9625 , n8154 , n5220 );
and ( n9626 , n4110 , n9096 );
or ( n9627 , n9625 , n9626 );
and ( n9628 , n9627 , n5286 );
and ( n9629 , n8165 , n5220 );
and ( n9630 , n4110 , n9096 );
or ( n9631 , n9629 , n9630 );
and ( n9632 , n9631 , n6219 );
and ( n9633 , n8176 , n5220 );
and ( n9634 , n4110 , n9096 );
or ( n9635 , n9633 , n9634 );
and ( n9636 , n9635 , n6711 );
and ( n9637 , n5608 , n5220 );
and ( n9638 , n4110 , n9096 );
or ( n9639 , n9637 , n9638 );
and ( n9640 , n9639 , n6718 );
and ( n9641 , n8188 , n5220 );
and ( n9642 , n4110 , n9096 );
or ( n9643 , n9641 , n9642 );
and ( n9644 , n9643 , n6725 );
and ( n9645 , n4110 , n9116 );
or ( n9646 , n9628 , n9632 , n9636 , n9640 , n9644 , n9645 );
and ( n9647 , n9624 , n9646 );
and ( n9648 , n4110 , n3260 );
or ( n9649 , n9647 , n9648 );
and ( n9650 , n9649 , n2422 );
and ( n9651 , n4110 , n2428 );
or ( n9652 , n9650 , n9651 );
buf ( n9653 , n9652 );
buf ( n9654 , n2424 );
buf ( n9655 , n2281 );
buf ( n9656 , n2280 );
not ( n9657 , n3260 );
and ( n9658 , n8228 , n5220 );
and ( n9659 , n4100 , n9096 );
or ( n9660 , n9658 , n9659 );
and ( n9661 , n9660 , n5286 );
and ( n9662 , n8239 , n5220 );
and ( n9663 , n4100 , n9096 );
or ( n9664 , n9662 , n9663 );
and ( n9665 , n9664 , n6219 );
and ( n9666 , n8250 , n5220 );
and ( n9667 , n4100 , n9096 );
or ( n9668 , n9666 , n9667 );
and ( n9669 , n9668 , n6711 );
and ( n9670 , n5598 , n5220 );
and ( n9671 , n4100 , n9096 );
or ( n9672 , n9670 , n9671 );
and ( n9673 , n9672 , n6718 );
and ( n9674 , n8262 , n5220 );
and ( n9675 , n4100 , n9096 );
or ( n9676 , n9674 , n9675 );
and ( n9677 , n9676 , n6725 );
and ( n9678 , n4100 , n9116 );
or ( n9679 , n9661 , n9665 , n9669 , n9673 , n9677 , n9678 );
and ( n9680 , n9657 , n9679 );
and ( n9681 , n4100 , n3260 );
or ( n9682 , n9680 , n9681 );
and ( n9683 , n9682 , n2422 );
and ( n9684 , n4100 , n2428 );
or ( n9685 , n9683 , n9684 );
buf ( n9686 , n9685 );
buf ( n9687 , n2424 );
buf ( n9688 , n2281 );
buf ( n9689 , n2280 );
not ( n9690 , n3260 );
and ( n9691 , n8302 , n5220 );
and ( n9692 , n4090 , n9096 );
or ( n9693 , n9691 , n9692 );
and ( n9694 , n9693 , n5286 );
and ( n9695 , n8313 , n5220 );
and ( n9696 , n4090 , n9096 );
or ( n9697 , n9695 , n9696 );
and ( n9698 , n9697 , n6219 );
and ( n9699 , n8324 , n5220 );
and ( n9700 , n4090 , n9096 );
or ( n9701 , n9699 , n9700 );
and ( n9702 , n9701 , n6711 );
and ( n9703 , n5588 , n5220 );
and ( n9704 , n4090 , n9096 );
or ( n9705 , n9703 , n9704 );
and ( n9706 , n9705 , n6718 );
and ( n9707 , n8336 , n5220 );
and ( n9708 , n4090 , n9096 );
or ( n9709 , n9707 , n9708 );
and ( n9710 , n9709 , n6725 );
and ( n9711 , n4090 , n9116 );
or ( n9712 , n9694 , n9698 , n9702 , n9706 , n9710 , n9711 );
and ( n9713 , n9690 , n9712 );
and ( n9714 , n4090 , n3260 );
or ( n9715 , n9713 , n9714 );
and ( n9716 , n9715 , n2422 );
and ( n9717 , n4090 , n2428 );
or ( n9718 , n9716 , n9717 );
buf ( n9719 , n9718 );
buf ( n9720 , n2424 );
buf ( n9721 , n2281 );
buf ( n9722 , n2280 );
not ( n9723 , n3260 );
and ( n9724 , n8376 , n5220 );
and ( n9725 , n4080 , n9096 );
or ( n9726 , n9724 , n9725 );
and ( n9727 , n9726 , n5286 );
and ( n9728 , n8387 , n5220 );
and ( n9729 , n4080 , n9096 );
or ( n9730 , n9728 , n9729 );
and ( n9731 , n9730 , n6219 );
and ( n9732 , n8398 , n5220 );
and ( n9733 , n4080 , n9096 );
or ( n9734 , n9732 , n9733 );
and ( n9735 , n9734 , n6711 );
and ( n9736 , n5578 , n5220 );
and ( n9737 , n4080 , n9096 );
or ( n9738 , n9736 , n9737 );
and ( n9739 , n9738 , n6718 );
and ( n9740 , n8410 , n5220 );
and ( n9741 , n4080 , n9096 );
or ( n9742 , n9740 , n9741 );
and ( n9743 , n9742 , n6725 );
and ( n9744 , n4080 , n9116 );
or ( n9745 , n9727 , n9731 , n9735 , n9739 , n9743 , n9744 );
and ( n9746 , n9723 , n9745 );
and ( n9747 , n4080 , n3260 );
or ( n9748 , n9746 , n9747 );
and ( n9749 , n9748 , n2422 );
and ( n9750 , n4080 , n2428 );
or ( n9751 , n9749 , n9750 );
buf ( n9752 , n9751 );
buf ( n9753 , n2424 );
buf ( n9754 , n2281 );
buf ( n9755 , n2280 );
not ( n9756 , n3260 );
and ( n9757 , n8450 , n5220 );
and ( n9758 , n4070 , n9096 );
or ( n9759 , n9757 , n9758 );
and ( n9760 , n9759 , n5286 );
and ( n9761 , n8461 , n5220 );
and ( n9762 , n4070 , n9096 );
or ( n9763 , n9761 , n9762 );
and ( n9764 , n9763 , n6219 );
and ( n9765 , n8472 , n5220 );
and ( n9766 , n4070 , n9096 );
or ( n9767 , n9765 , n9766 );
and ( n9768 , n9767 , n6711 );
and ( n9769 , n5530 , n5220 );
and ( n9770 , n4070 , n9096 );
or ( n9771 , n9769 , n9770 );
and ( n9772 , n9771 , n6718 );
and ( n9773 , n8484 , n5220 );
and ( n9774 , n4070 , n9096 );
or ( n9775 , n9773 , n9774 );
and ( n9776 , n9775 , n6725 );
and ( n9777 , n4070 , n9116 );
or ( n9778 , n9760 , n9764 , n9768 , n9772 , n9776 , n9777 );
and ( n9779 , n9756 , n9778 );
and ( n9780 , n4070 , n3260 );
or ( n9781 , n9779 , n9780 );
and ( n9782 , n9781 , n2422 );
and ( n9783 , n4070 , n2428 );
or ( n9784 , n9782 , n9783 );
buf ( n9785 , n9784 );
buf ( n9786 , n2424 );
buf ( n9787 , n2281 );
buf ( n9788 , n2280 );
not ( n9789 , n3260 );
and ( n9790 , n8524 , n5220 );
and ( n9791 , n4060 , n9096 );
or ( n9792 , n9790 , n9791 );
and ( n9793 , n9792 , n5286 );
and ( n9794 , n8535 , n5220 );
and ( n9795 , n4060 , n9096 );
or ( n9796 , n9794 , n9795 );
and ( n9797 , n9796 , n6219 );
and ( n9798 , n8546 , n5220 );
and ( n9799 , n4060 , n9096 );
or ( n9800 , n9798 , n9799 );
and ( n9801 , n9800 , n6711 );
and ( n9802 , n5527 , n5220 );
and ( n9803 , n4060 , n9096 );
or ( n9804 , n9802 , n9803 );
and ( n9805 , n9804 , n6718 );
and ( n9806 , n8558 , n5220 );
and ( n9807 , n4060 , n9096 );
or ( n9808 , n9806 , n9807 );
and ( n9809 , n9808 , n6725 );
and ( n9810 , n4060 , n9116 );
or ( n9811 , n9793 , n9797 , n9801 , n9805 , n9809 , n9810 );
and ( n9812 , n9789 , n9811 );
and ( n9813 , n4060 , n3260 );
or ( n9814 , n9812 , n9813 );
and ( n9815 , n9814 , n2422 );
and ( n9816 , n4060 , n2428 );
or ( n9817 , n9815 , n9816 );
buf ( n9818 , n9817 );
buf ( n9819 , n2424 );
buf ( n9820 , n2281 );
buf ( n9821 , n2280 );
not ( n9822 , n3260 );
and ( n9823 , n8598 , n5220 );
and ( n9824 , n4050 , n9096 );
or ( n9825 , n9823 , n9824 );
and ( n9826 , n9825 , n5286 );
and ( n9827 , n8609 , n5220 );
and ( n9828 , n4050 , n9096 );
or ( n9829 , n9827 , n9828 );
and ( n9830 , n9829 , n6219 );
and ( n9831 , n8620 , n5220 );
and ( n9832 , n4050 , n9096 );
or ( n9833 , n9831 , n9832 );
and ( n9834 , n9833 , n6711 );
and ( n9835 , n5524 , n5220 );
and ( n9836 , n4050 , n9096 );
or ( n9837 , n9835 , n9836 );
and ( n9838 , n9837 , n6718 );
and ( n9839 , n8632 , n5220 );
and ( n9840 , n4050 , n9096 );
or ( n9841 , n9839 , n9840 );
and ( n9842 , n9841 , n6725 );
and ( n9843 , n4050 , n9116 );
or ( n9844 , n9826 , n9830 , n9834 , n9838 , n9842 , n9843 );
and ( n9845 , n9822 , n9844 );
and ( n9846 , n4050 , n3260 );
or ( n9847 , n9845 , n9846 );
and ( n9848 , n9847 , n2422 );
and ( n9849 , n4050 , n2428 );
or ( n9850 , n9848 , n9849 );
buf ( n9851 , n9850 );
buf ( n9852 , n2424 );
buf ( n9853 , n2281 );
buf ( n9854 , n2280 );
not ( n9855 , n3260 );
and ( n9856 , n8672 , n5220 );
and ( n9857 , n4040 , n9096 );
or ( n9858 , n9856 , n9857 );
and ( n9859 , n9858 , n5286 );
and ( n9860 , n8683 , n5220 );
and ( n9861 , n4040 , n9096 );
or ( n9862 , n9860 , n9861 );
and ( n9863 , n9862 , n6219 );
and ( n9864 , n8694 , n5220 );
and ( n9865 , n4040 , n9096 );
or ( n9866 , n9864 , n9865 );
and ( n9867 , n9866 , n6711 );
and ( n9868 , n5521 , n5220 );
and ( n9869 , n4040 , n9096 );
or ( n9870 , n9868 , n9869 );
and ( n9871 , n9870 , n6718 );
and ( n9872 , n8706 , n5220 );
and ( n9873 , n4040 , n9096 );
or ( n9874 , n9872 , n9873 );
and ( n9875 , n9874 , n6725 );
and ( n9876 , n4040 , n9116 );
or ( n9877 , n9859 , n9863 , n9867 , n9871 , n9875 , n9876 );
and ( n9878 , n9855 , n9877 );
and ( n9879 , n4040 , n3260 );
or ( n9880 , n9878 , n9879 );
and ( n9881 , n9880 , n2422 );
and ( n9882 , n4040 , n2428 );
or ( n9883 , n9881 , n9882 );
buf ( n9884 , n9883 );
buf ( n9885 , n2424 );
buf ( n9886 , n2281 );
buf ( n9887 , n2280 );
not ( n9888 , n3260 );
and ( n9889 , n8746 , n5220 );
and ( n9890 , n4030 , n9096 );
or ( n9891 , n9889 , n9890 );
and ( n9892 , n9891 , n5286 );
and ( n9893 , n8757 , n5220 );
and ( n9894 , n4030 , n9096 );
or ( n9895 , n9893 , n9894 );
and ( n9896 , n9895 , n6219 );
and ( n9897 , n8768 , n5220 );
and ( n9898 , n4030 , n9096 );
or ( n9899 , n9897 , n9898 );
and ( n9900 , n9899 , n6711 );
and ( n9901 , n5518 , n5220 );
and ( n9902 , n4030 , n9096 );
or ( n9903 , n9901 , n9902 );
and ( n9904 , n9903 , n6718 );
and ( n9905 , n8780 , n5220 );
and ( n9906 , n4030 , n9096 );
or ( n9907 , n9905 , n9906 );
and ( n9908 , n9907 , n6725 );
and ( n9909 , n4030 , n9116 );
or ( n9910 , n9892 , n9896 , n9900 , n9904 , n9908 , n9909 );
and ( n9911 , n9888 , n9910 );
and ( n9912 , n4030 , n3260 );
or ( n9913 , n9911 , n9912 );
and ( n9914 , n9913 , n2422 );
and ( n9915 , n4030 , n2428 );
or ( n9916 , n9914 , n9915 );
buf ( n9917 , n9916 );
buf ( n9918 , n2424 );
buf ( n9919 , n2281 );
buf ( n9920 , n2280 );
not ( n9921 , n3260 );
and ( n9922 , n8820 , n5220 );
and ( n9923 , n4020 , n9096 );
or ( n9924 , n9922 , n9923 );
and ( n9925 , n9924 , n5286 );
and ( n9926 , n8831 , n5220 );
and ( n9927 , n4020 , n9096 );
or ( n9928 , n9926 , n9927 );
and ( n9929 , n9928 , n6219 );
and ( n9930 , n8842 , n5220 );
and ( n9931 , n4020 , n9096 );
or ( n9932 , n9930 , n9931 );
and ( n9933 , n9932 , n6711 );
and ( n9934 , n5515 , n5220 );
and ( n9935 , n4020 , n9096 );
or ( n9936 , n9934 , n9935 );
and ( n9937 , n9936 , n6718 );
and ( n9938 , n8854 , n5220 );
and ( n9939 , n4020 , n9096 );
or ( n9940 , n9938 , n9939 );
and ( n9941 , n9940 , n6725 );
and ( n9942 , n4020 , n9116 );
or ( n9943 , n9925 , n9929 , n9933 , n9937 , n9941 , n9942 );
and ( n9944 , n9921 , n9943 );
and ( n9945 , n4020 , n3260 );
or ( n9946 , n9944 , n9945 );
and ( n9947 , n9946 , n2422 );
and ( n9948 , n4020 , n2428 );
or ( n9949 , n9947 , n9948 );
buf ( n9950 , n9949 );
buf ( n9951 , n2424 );
buf ( n9952 , n2281 );
buf ( n9953 , n2280 );
not ( n9954 , n3260 );
and ( n9955 , n8894 , n5220 );
and ( n9956 , n4010 , n9096 );
or ( n9957 , n9955 , n9956 );
and ( n9958 , n9957 , n5286 );
and ( n9959 , n8905 , n5220 );
and ( n9960 , n4010 , n9096 );
or ( n9961 , n9959 , n9960 );
and ( n9962 , n9961 , n6219 );
and ( n9963 , n8916 , n5220 );
and ( n9964 , n4010 , n9096 );
or ( n9965 , n9963 , n9964 );
and ( n9966 , n9965 , n6711 );
and ( n9967 , n5512 , n5220 );
and ( n9968 , n4010 , n9096 );
or ( n9969 , n9967 , n9968 );
and ( n9970 , n9969 , n6718 );
and ( n9971 , n8928 , n5220 );
and ( n9972 , n4010 , n9096 );
or ( n9973 , n9971 , n9972 );
and ( n9974 , n9973 , n6725 );
and ( n9975 , n4010 , n9116 );
or ( n9976 , n9958 , n9962 , n9966 , n9970 , n9974 , n9975 );
and ( n9977 , n9954 , n9976 );
and ( n9978 , n4010 , n3260 );
or ( n9979 , n9977 , n9978 );
and ( n9980 , n9979 , n2422 );
and ( n9981 , n4010 , n2428 );
or ( n9982 , n9980 , n9981 );
buf ( n9983 , n9982 );
buf ( n9984 , n2424 );
buf ( n9985 , n2281 );
buf ( n9986 , n2280 );
not ( n9987 , n3260 );
and ( n9988 , n8968 , n5220 );
and ( n9989 , n4000 , n9096 );
or ( n9990 , n9988 , n9989 );
and ( n9991 , n9990 , n5286 );
and ( n9992 , n8979 , n5220 );
and ( n9993 , n4000 , n9096 );
or ( n9994 , n9992 , n9993 );
and ( n9995 , n9994 , n6219 );
and ( n9996 , n8990 , n5220 );
and ( n9997 , n4000 , n9096 );
or ( n9998 , n9996 , n9997 );
and ( n9999 , n9998 , n6711 );
and ( n10000 , n5509 , n5220 );
and ( n10001 , n4000 , n9096 );
or ( n10002 , n10000 , n10001 );
and ( n10003 , n10002 , n6718 );
and ( n10004 , n9002 , n5220 );
and ( n10005 , n4000 , n9096 );
or ( n10006 , n10004 , n10005 );
and ( n10007 , n10006 , n6725 );
and ( n10008 , n4000 , n9116 );
or ( n10009 , n9991 , n9995 , n9999 , n10003 , n10007 , n10008 );
and ( n10010 , n9987 , n10009 );
and ( n10011 , n4000 , n3260 );
or ( n10012 , n10010 , n10011 );
and ( n10013 , n10012 , n2422 );
and ( n10014 , n4000 , n2428 );
or ( n10015 , n10013 , n10014 );
buf ( n10016 , n10015 );
buf ( n10017 , n2424 );
buf ( n10018 , n2281 );
buf ( n10019 , n2280 );
not ( n10020 , n3260 );
and ( n10021 , n9042 , n5220 );
and ( n10022 , n3990 , n9096 );
or ( n10023 , n10021 , n10022 );
and ( n10024 , n10023 , n5286 );
and ( n10025 , n9053 , n5220 );
and ( n10026 , n3990 , n9096 );
or ( n10027 , n10025 , n10026 );
and ( n10028 , n10027 , n6219 );
and ( n10029 , n9064 , n5220 );
and ( n10030 , n3990 , n9096 );
or ( n10031 , n10029 , n10030 );
and ( n10032 , n10031 , n6711 );
and ( n10033 , n5506 , n5220 );
and ( n10034 , n3990 , n9096 );
or ( n10035 , n10033 , n10034 );
and ( n10036 , n10035 , n6718 );
and ( n10037 , n9076 , n5220 );
and ( n10038 , n3990 , n9096 );
or ( n10039 , n10037 , n10038 );
and ( n10040 , n10039 , n6725 );
and ( n10041 , n3990 , n9116 );
or ( n10042 , n10024 , n10028 , n10032 , n10036 , n10040 , n10041 );
and ( n10043 , n10020 , n10042 );
and ( n10044 , n3990 , n3260 );
or ( n10045 , n10043 , n10044 );
and ( n10046 , n10045 , n2422 );
and ( n10047 , n3990 , n2428 );
or ( n10048 , n10046 , n10047 );
buf ( n10049 , n10048 );
buf ( n10050 , n2424 );
buf ( n10051 , n2281 );
buf ( n10052 , n2280 );
not ( n10053 , n3260 );
not ( n10054 , n7022 );
and ( n10055 , n10054 , n7020 );
xor ( n10056 , n7020 , n3770 );
and ( n10057 , n9022 , n9023 );
xor ( n10058 , n10056 , n10057 );
and ( n10059 , n10058 , n7022 );
or ( n10060 , n10055 , n10059 );
and ( n10061 , n10060 , n5290 );
and ( n10062 , n10060 , n5288 );
not ( n10063 , n3290 );
not ( n10064 , n3770 );
and ( n10065 , n10064 , n4302 );
xor ( n10066 , n4303 , n4574 );
and ( n10067 , n10066 , n3770 );
or ( n10068 , n10065 , n10067 );
and ( n10069 , n10063 , n10068 );
not ( n10070 , n5000 );
and ( n10071 , n10070 , n2424 );
and ( n10072 , n9033 , n9034 );
and ( n10073 , n10072 , n5000 );
or ( n10074 , n10071 , n10073 );
and ( n10075 , n10074 , n3290 );
or ( n10076 , n10069 , n10075 );
and ( n10077 , n10076 , n5153 );
and ( n10078 , n10068 , n5155 );
or ( n10079 , n10061 , n10062 , n10077 , n10078 );
and ( n10080 , n10079 , n5220 );
and ( n10081 , n3980 , n9096 );
or ( n10082 , n10080 , n10081 );
and ( n10083 , n10082 , n5286 );
not ( n10084 , n6202 );
and ( n10085 , n10084 , n6200 );
xor ( n10086 , n6200 , n5853 );
and ( n10087 , n9049 , n9050 );
xor ( n10088 , n10086 , n10087 );
and ( n10089 , n10088 , n6202 );
or ( n10090 , n10085 , n10089 );
and ( n10091 , n10090 , n5220 );
and ( n10092 , n3980 , n9096 );
or ( n10093 , n10091 , n10092 );
and ( n10094 , n10093 , n6219 );
not ( n10095 , n6695 );
and ( n10096 , n10095 , n6693 );
xor ( n10097 , n6693 , n6346 );
and ( n10098 , n9060 , n9061 );
xor ( n10099 , n10097 , n10098 );
and ( n10100 , n10099 , n6695 );
or ( n10101 , n10096 , n10100 );
and ( n10102 , n10101 , n5220 );
and ( n10103 , n3980 , n9096 );
or ( n10104 , n10102 , n10103 );
and ( n10105 , n10104 , n6711 );
and ( n10106 , n5503 , n5220 );
and ( n10107 , n3980 , n9096 );
or ( n10108 , n10106 , n10107 );
and ( n10109 , n10108 , n6718 );
not ( n10110 , n5503 );
and ( n10111 , n9074 , n9075 );
xor ( n10112 , n10110 , n10111 );
and ( n10113 , n10112 , n5220 );
and ( n10114 , n3980 , n9096 );
or ( n10115 , n10113 , n10114 );
and ( n10116 , n10115 , n6725 );
and ( n10117 , n3980 , n9116 );
or ( n10118 , n10083 , n10094 , n10105 , n10109 , n10116 , n10117 );
and ( n10119 , n10053 , n10118 );
and ( n10120 , n3980 , n3260 );
or ( n10121 , n10119 , n10120 );
and ( n10122 , n10121 , n2422 );
and ( n10123 , n3980 , n2428 );
or ( n10124 , n10122 , n10123 );
buf ( n10125 , n10124 );
buf ( n10126 , n2424 );
buf ( n10127 , n2281 );
buf ( n10128 , n2280 );
not ( n10129 , n3260 );
not ( n10130 , n7022 );
and ( n10131 , n10130 , n2424 );
and ( n10132 , n10056 , n10057 );
and ( n10133 , n10132 , n7022 );
or ( n10134 , n10131 , n10133 );
and ( n10135 , n10134 , n5290 );
and ( n10136 , n10134 , n5288 );
not ( n10137 , n3290 );
not ( n10138 , n3770 );
and ( n10139 , n10138 , n4294 );
xor ( n10140 , n4295 , n4575 );
and ( n10141 , n10140 , n3770 );
or ( n10142 , n10139 , n10141 );
and ( n10143 , n10137 , n10142 );
and ( n10144 , n2424 , n3290 );
or ( n10145 , n10143 , n10144 );
and ( n10146 , n10145 , n5153 );
and ( n10147 , n10142 , n5155 );
or ( n10148 , n10135 , n10136 , n10146 , n10147 );
and ( n10149 , n10148 , n5220 );
and ( n10150 , n3815 , n9096 );
or ( n10151 , n10149 , n10150 );
and ( n10152 , n10151 , n5286 );
not ( n10153 , n6202 );
and ( n10154 , n10153 , n2424 );
and ( n10155 , n10086 , n10087 );
and ( n10156 , n10155 , n6202 );
or ( n10157 , n10154 , n10156 );
and ( n10158 , n10157 , n5220 );
and ( n10159 , n3815 , n9096 );
or ( n10160 , n10158 , n10159 );
and ( n10161 , n10160 , n6219 );
not ( n10162 , n6695 );
and ( n10163 , n10162 , n2424 );
and ( n10164 , n10097 , n10098 );
and ( n10165 , n10164 , n6695 );
or ( n10166 , n10163 , n10165 );
and ( n10167 , n10166 , n5220 );
and ( n10168 , n3815 , n9096 );
or ( n10169 , n10167 , n10168 );
and ( n10170 , n10169 , n6711 );
and ( n10171 , n5500 , n5220 );
and ( n10172 , n3815 , n9096 );
or ( n10173 , n10171 , n10172 );
and ( n10174 , n10173 , n6718 );
not ( n10175 , n5500 );
and ( n10176 , n10110 , n10111 );
xor ( n10177 , n10175 , n10176 );
and ( n10178 , n10177 , n5220 );
and ( n10179 , n3815 , n9096 );
or ( n10180 , n10178 , n10179 );
and ( n10181 , n10180 , n6725 );
and ( n10182 , n3815 , n9116 );
or ( n10183 , n10152 , n10161 , n10170 , n10174 , n10181 , n10182 );
and ( n10184 , n10129 , n10183 );
and ( n10185 , n3815 , n3260 );
or ( n10186 , n10184 , n10185 );
and ( n10187 , n10186 , n2422 );
and ( n10188 , n3815 , n2428 );
or ( n10189 , n10187 , n10188 );
buf ( n10190 , n10189 );
buf ( n10191 , n2424 );
buf ( n10192 , n2281 );
buf ( n10193 , n2280 );
not ( n10194 , n3260 );
buf ( n10195 , n2424 );
not ( n10196 , n3290 );
and ( n10197 , n10196 , n4579 );
and ( n10198 , n2424 , n3290 );
or ( n10199 , n10197 , n10198 );
and ( n10200 , n10199 , n5153 );
and ( n10201 , n4579 , n5155 );
or ( n10202 , n2424 , n10195 , n10200 , n10201 );
and ( n10203 , n10202 , n5220 );
and ( n10204 , n3764 , n9096 );
or ( n10205 , n10203 , n10204 );
and ( n10206 , n10205 , n5286 );
and ( n10207 , n3764 , n9096 );
and ( n10208 , n10207 , n6219 );
and ( n10209 , n3764 , n9096 );
and ( n10210 , n10209 , n6711 );
and ( n10211 , n5497 , n5220 );
and ( n10212 , n3764 , n9096 );
or ( n10213 , n10211 , n10212 );
and ( n10214 , n10213 , n6718 );
not ( n10215 , n5497 );
and ( n10216 , n10175 , n10176 );
xor ( n10217 , n10215 , n10216 );
and ( n10218 , n10217 , n5220 );
and ( n10219 , n3764 , n9096 );
or ( n10220 , n10218 , n10219 );
and ( n10221 , n10220 , n6725 );
and ( n10222 , n3764 , n9116 );
or ( n10223 , n10206 , n10208 , n10210 , n10214 , n10221 , n10222 );
and ( n10224 , n10194 , n10223 );
and ( n10225 , n3764 , n3260 );
or ( n10226 , n10224 , n10225 );
and ( n10227 , n10226 , n2422 );
and ( n10228 , n3764 , n2428 );
or ( n10229 , n10227 , n10228 );
buf ( n10230 , n10229 );
buf ( n10231 , n2424 );
buf ( n10232 , n2281 );
buf ( n10233 , n2280 );
not ( n10234 , n3260 );
and ( n10235 , n5157 , n5250 );
or ( n10236 , n5220 , n5281 );
or ( n10237 , n10236 , n5189 );
buf ( n10238 , n10237 );
and ( n10239 , n3793 , n10238 );
or ( n10240 , n10235 , n10239 );
and ( n10241 , n10240 , n5286 );
and ( n10242 , n6208 , n5250 );
and ( n10243 , n3793 , n10238 );
or ( n10244 , n10242 , n10243 );
and ( n10245 , n10244 , n6219 );
and ( n10246 , n6701 , n5250 );
and ( n10247 , n3793 , n10238 );
or ( n10248 , n10246 , n10247 );
and ( n10249 , n10248 , n6711 );
and ( n10250 , n5493 , n5250 );
and ( n10251 , n3793 , n10238 );
or ( n10252 , n10250 , n10251 );
and ( n10253 , n10252 , n6718 );
and ( n10254 , n5493 , n5250 );
and ( n10255 , n3793 , n10238 );
or ( n10256 , n10254 , n10255 );
and ( n10257 , n10256 , n6725 );
and ( n10258 , n3793 , n9116 );
or ( n10259 , n10241 , n10245 , n10249 , n10253 , n10257 , n10258 );
and ( n10260 , n10234 , n10259 );
and ( n10261 , n3793 , n3260 );
or ( n10262 , n10260 , n10261 );
and ( n10263 , n10262 , n2422 );
and ( n10264 , n3793 , n2428 );
or ( n10265 , n10263 , n10264 );
buf ( n10266 , n10265 );
buf ( n10267 , n2424 );
buf ( n10268 , n2281 );
buf ( n10269 , n2280 );
not ( n10270 , n3260 );
and ( n10271 , n7044 , n5250 );
and ( n10272 , n3783 , n10238 );
or ( n10273 , n10271 , n10272 );
and ( n10274 , n10273 , n5286 );
and ( n10275 , n7055 , n5250 );
and ( n10276 , n3783 , n10238 );
or ( n10277 , n10275 , n10276 );
and ( n10278 , n10277 , n6219 );
and ( n10279 , n7066 , n5250 );
and ( n10280 , n3783 , n10238 );
or ( n10281 , n10279 , n10280 );
and ( n10282 , n10281 , n6711 );
and ( n10283 , n5758 , n5250 );
and ( n10284 , n3783 , n10238 );
or ( n10285 , n10283 , n10284 );
and ( n10286 , n10285 , n6718 );
and ( n10287 , n7078 , n5250 );
and ( n10288 , n3783 , n10238 );
or ( n10289 , n10287 , n10288 );
and ( n10290 , n10289 , n6725 );
and ( n10291 , n3783 , n9116 );
or ( n10292 , n10274 , n10278 , n10282 , n10286 , n10290 , n10291 );
and ( n10293 , n10270 , n10292 );
and ( n10294 , n3783 , n3260 );
or ( n10295 , n10293 , n10294 );
and ( n10296 , n10295 , n2422 );
and ( n10297 , n3783 , n2428 );
or ( n10298 , n10296 , n10297 );
buf ( n10299 , n10298 );
buf ( n10300 , n2424 );
buf ( n10301 , n2281 );
buf ( n10302 , n2280 );
not ( n10303 , n3260 );
and ( n10304 , n7118 , n5250 );
and ( n10305 , n4256 , n10238 );
or ( n10306 , n10304 , n10305 );
and ( n10307 , n10306 , n5286 );
and ( n10308 , n7129 , n5250 );
and ( n10309 , n4256 , n10238 );
or ( n10310 , n10308 , n10309 );
and ( n10311 , n10310 , n6219 );
and ( n10312 , n7140 , n5250 );
and ( n10313 , n4256 , n10238 );
or ( n10314 , n10312 , n10313 );
and ( n10315 , n10314 , n6711 );
and ( n10316 , n5748 , n5250 );
and ( n10317 , n4256 , n10238 );
or ( n10318 , n10316 , n10317 );
and ( n10319 , n10318 , n6718 );
and ( n10320 , n7152 , n5250 );
and ( n10321 , n4256 , n10238 );
or ( n10322 , n10320 , n10321 );
and ( n10323 , n10322 , n6725 );
and ( n10324 , n4256 , n9116 );
or ( n10325 , n10307 , n10311 , n10315 , n10319 , n10323 , n10324 );
and ( n10326 , n10303 , n10325 );
and ( n10327 , n4256 , n3260 );
or ( n10328 , n10326 , n10327 );
and ( n10329 , n10328 , n2422 );
and ( n10330 , n4256 , n2428 );
or ( n10331 , n10329 , n10330 );
buf ( n10332 , n10331 );
buf ( n10333 , n2424 );
buf ( n10334 , n2281 );
buf ( n10335 , n2280 );
not ( n10336 , n3260 );
and ( n10337 , n7192 , n5250 );
and ( n10338 , n4242 , n10238 );
or ( n10339 , n10337 , n10338 );
and ( n10340 , n10339 , n5286 );
and ( n10341 , n7203 , n5250 );
and ( n10342 , n4242 , n10238 );
or ( n10343 , n10341 , n10342 );
and ( n10344 , n10343 , n6219 );
and ( n10345 , n7214 , n5250 );
and ( n10346 , n4242 , n10238 );
or ( n10347 , n10345 , n10346 );
and ( n10348 , n10347 , n6711 );
and ( n10349 , n5738 , n5250 );
and ( n10350 , n4242 , n10238 );
or ( n10351 , n10349 , n10350 );
and ( n10352 , n10351 , n6718 );
and ( n10353 , n7226 , n5250 );
and ( n10354 , n4242 , n10238 );
or ( n10355 , n10353 , n10354 );
and ( n10356 , n10355 , n6725 );
and ( n10357 , n4242 , n9116 );
or ( n10358 , n10340 , n10344 , n10348 , n10352 , n10356 , n10357 );
and ( n10359 , n10336 , n10358 );
and ( n10360 , n4242 , n3260 );
or ( n10361 , n10359 , n10360 );
and ( n10362 , n10361 , n2422 );
and ( n10363 , n4242 , n2428 );
or ( n10364 , n10362 , n10363 );
buf ( n10365 , n10364 );
buf ( n10366 , n2424 );
buf ( n10367 , n2281 );
buf ( n10368 , n2280 );
not ( n10369 , n3260 );
and ( n10370 , n7266 , n5250 );
and ( n10371 , n4232 , n10238 );
or ( n10372 , n10370 , n10371 );
and ( n10373 , n10372 , n5286 );
and ( n10374 , n7277 , n5250 );
and ( n10375 , n4232 , n10238 );
or ( n10376 , n10374 , n10375 );
and ( n10377 , n10376 , n6219 );
and ( n10378 , n7288 , n5250 );
and ( n10379 , n4232 , n10238 );
or ( n10380 , n10378 , n10379 );
and ( n10381 , n10380 , n6711 );
and ( n10382 , n5728 , n5250 );
and ( n10383 , n4232 , n10238 );
or ( n10384 , n10382 , n10383 );
and ( n10385 , n10384 , n6718 );
and ( n10386 , n7300 , n5250 );
and ( n10387 , n4232 , n10238 );
or ( n10388 , n10386 , n10387 );
and ( n10389 , n10388 , n6725 );
and ( n10390 , n4232 , n9116 );
or ( n10391 , n10373 , n10377 , n10381 , n10385 , n10389 , n10390 );
and ( n10392 , n10369 , n10391 );
and ( n10393 , n4232 , n3260 );
or ( n10394 , n10392 , n10393 );
and ( n10395 , n10394 , n2422 );
and ( n10396 , n4232 , n2428 );
or ( n10397 , n10395 , n10396 );
buf ( n10398 , n10397 );
buf ( n10399 , n2424 );
buf ( n10400 , n2281 );
buf ( n10401 , n2280 );
not ( n10402 , n3260 );
and ( n10403 , n7340 , n5250 );
and ( n10404 , n4222 , n10238 );
or ( n10405 , n10403 , n10404 );
and ( n10406 , n10405 , n5286 );
and ( n10407 , n7351 , n5250 );
and ( n10408 , n4222 , n10238 );
or ( n10409 , n10407 , n10408 );
and ( n10410 , n10409 , n6219 );
and ( n10411 , n7362 , n5250 );
and ( n10412 , n4222 , n10238 );
or ( n10413 , n10411 , n10412 );
and ( n10414 , n10413 , n6711 );
and ( n10415 , n5718 , n5250 );
and ( n10416 , n4222 , n10238 );
or ( n10417 , n10415 , n10416 );
and ( n10418 , n10417 , n6718 );
and ( n10419 , n7374 , n5250 );
and ( n10420 , n4222 , n10238 );
or ( n10421 , n10419 , n10420 );
and ( n10422 , n10421 , n6725 );
and ( n10423 , n4222 , n9116 );
or ( n10424 , n10406 , n10410 , n10414 , n10418 , n10422 , n10423 );
and ( n10425 , n10402 , n10424 );
and ( n10426 , n4222 , n3260 );
or ( n10427 , n10425 , n10426 );
and ( n10428 , n10427 , n2422 );
and ( n10429 , n4222 , n2428 );
or ( n10430 , n10428 , n10429 );
buf ( n10431 , n10430 );
buf ( n10432 , n2424 );
buf ( n10433 , n2281 );
buf ( n10434 , n2280 );
not ( n10435 , n3260 );
and ( n10436 , n7414 , n5250 );
and ( n10437 , n4212 , n10238 );
or ( n10438 , n10436 , n10437 );
and ( n10439 , n10438 , n5286 );
and ( n10440 , n7425 , n5250 );
and ( n10441 , n4212 , n10238 );
or ( n10442 , n10440 , n10441 );
and ( n10443 , n10442 , n6219 );
and ( n10444 , n7436 , n5250 );
and ( n10445 , n4212 , n10238 );
or ( n10446 , n10444 , n10445 );
and ( n10447 , n10446 , n6711 );
and ( n10448 , n5708 , n5250 );
and ( n10449 , n4212 , n10238 );
or ( n10450 , n10448 , n10449 );
and ( n10451 , n10450 , n6718 );
and ( n10452 , n7448 , n5250 );
and ( n10453 , n4212 , n10238 );
or ( n10454 , n10452 , n10453 );
and ( n10455 , n10454 , n6725 );
and ( n10456 , n4212 , n9116 );
or ( n10457 , n10439 , n10443 , n10447 , n10451 , n10455 , n10456 );
and ( n10458 , n10435 , n10457 );
and ( n10459 , n4212 , n3260 );
or ( n10460 , n10458 , n10459 );
and ( n10461 , n10460 , n2422 );
and ( n10462 , n4212 , n2428 );
or ( n10463 , n10461 , n10462 );
buf ( n10464 , n10463 );
buf ( n10465 , n2424 );
buf ( n10466 , n2281 );
buf ( n10467 , n2280 );
not ( n10468 , n3260 );
and ( n10469 , n7488 , n5250 );
and ( n10470 , n4202 , n10238 );
or ( n10471 , n10469 , n10470 );
and ( n10472 , n10471 , n5286 );
and ( n10473 , n7499 , n5250 );
and ( n10474 , n4202 , n10238 );
or ( n10475 , n10473 , n10474 );
and ( n10476 , n10475 , n6219 );
and ( n10477 , n7510 , n5250 );
and ( n10478 , n4202 , n10238 );
or ( n10479 , n10477 , n10478 );
and ( n10480 , n10479 , n6711 );
and ( n10481 , n5698 , n5250 );
and ( n10482 , n4202 , n10238 );
or ( n10483 , n10481 , n10482 );
and ( n10484 , n10483 , n6718 );
and ( n10485 , n7522 , n5250 );
and ( n10486 , n4202 , n10238 );
or ( n10487 , n10485 , n10486 );
and ( n10488 , n10487 , n6725 );
and ( n10489 , n4202 , n9116 );
or ( n10490 , n10472 , n10476 , n10480 , n10484 , n10488 , n10489 );
and ( n10491 , n10468 , n10490 );
and ( n10492 , n4202 , n3260 );
or ( n10493 , n10491 , n10492 );
and ( n10494 , n10493 , n2422 );
and ( n10495 , n4202 , n2428 );
or ( n10496 , n10494 , n10495 );
buf ( n10497 , n10496 );
buf ( n10498 , n2424 );
buf ( n10499 , n2281 );
buf ( n10500 , n2280 );
not ( n10501 , n3260 );
and ( n10502 , n7562 , n5250 );
and ( n10503 , n4192 , n10238 );
or ( n10504 , n10502 , n10503 );
and ( n10505 , n10504 , n5286 );
and ( n10506 , n7573 , n5250 );
and ( n10507 , n4192 , n10238 );
or ( n10508 , n10506 , n10507 );
and ( n10509 , n10508 , n6219 );
and ( n10510 , n7584 , n5250 );
and ( n10511 , n4192 , n10238 );
or ( n10512 , n10510 , n10511 );
and ( n10513 , n10512 , n6711 );
and ( n10514 , n5688 , n5250 );
and ( n10515 , n4192 , n10238 );
or ( n10516 , n10514 , n10515 );
and ( n10517 , n10516 , n6718 );
and ( n10518 , n7596 , n5250 );
and ( n10519 , n4192 , n10238 );
or ( n10520 , n10518 , n10519 );
and ( n10521 , n10520 , n6725 );
and ( n10522 , n4192 , n9116 );
or ( n10523 , n10505 , n10509 , n10513 , n10517 , n10521 , n10522 );
and ( n10524 , n10501 , n10523 );
and ( n10525 , n4192 , n3260 );
or ( n10526 , n10524 , n10525 );
and ( n10527 , n10526 , n2422 );
and ( n10528 , n4192 , n2428 );
or ( n10529 , n10527 , n10528 );
buf ( n10530 , n10529 );
buf ( n10531 , n2424 );
buf ( n10532 , n2281 );
buf ( n10533 , n2280 );
not ( n10534 , n3260 );
and ( n10535 , n7636 , n5250 );
and ( n10536 , n4182 , n10238 );
or ( n10537 , n10535 , n10536 );
and ( n10538 , n10537 , n5286 );
and ( n10539 , n7647 , n5250 );
and ( n10540 , n4182 , n10238 );
or ( n10541 , n10539 , n10540 );
and ( n10542 , n10541 , n6219 );
and ( n10543 , n7658 , n5250 );
and ( n10544 , n4182 , n10238 );
or ( n10545 , n10543 , n10544 );
and ( n10546 , n10545 , n6711 );
and ( n10547 , n5678 , n5250 );
and ( n10548 , n4182 , n10238 );
or ( n10549 , n10547 , n10548 );
and ( n10550 , n10549 , n6718 );
and ( n10551 , n7670 , n5250 );
and ( n10552 , n4182 , n10238 );
or ( n10553 , n10551 , n10552 );
and ( n10554 , n10553 , n6725 );
and ( n10555 , n4182 , n9116 );
or ( n10556 , n10538 , n10542 , n10546 , n10550 , n10554 , n10555 );
and ( n10557 , n10534 , n10556 );
and ( n10558 , n4182 , n3260 );
or ( n10559 , n10557 , n10558 );
and ( n10560 , n10559 , n2422 );
and ( n10561 , n4182 , n2428 );
or ( n10562 , n10560 , n10561 );
buf ( n10563 , n10562 );
buf ( n10564 , n2424 );
buf ( n10565 , n2281 );
buf ( n10566 , n2280 );
not ( n10567 , n3260 );
and ( n10568 , n7710 , n5250 );
and ( n10569 , n4172 , n10238 );
or ( n10570 , n10568 , n10569 );
and ( n10571 , n10570 , n5286 );
and ( n10572 , n7721 , n5250 );
and ( n10573 , n4172 , n10238 );
or ( n10574 , n10572 , n10573 );
and ( n10575 , n10574 , n6219 );
and ( n10576 , n7732 , n5250 );
and ( n10577 , n4172 , n10238 );
or ( n10578 , n10576 , n10577 );
and ( n10579 , n10578 , n6711 );
and ( n10580 , n5668 , n5250 );
and ( n10581 , n4172 , n10238 );
or ( n10582 , n10580 , n10581 );
and ( n10583 , n10582 , n6718 );
and ( n10584 , n7744 , n5250 );
and ( n10585 , n4172 , n10238 );
or ( n10586 , n10584 , n10585 );
and ( n10587 , n10586 , n6725 );
and ( n10588 , n4172 , n9116 );
or ( n10589 , n10571 , n10575 , n10579 , n10583 , n10587 , n10588 );
and ( n10590 , n10567 , n10589 );
and ( n10591 , n4172 , n3260 );
or ( n10592 , n10590 , n10591 );
and ( n10593 , n10592 , n2422 );
and ( n10594 , n4172 , n2428 );
or ( n10595 , n10593 , n10594 );
buf ( n10596 , n10595 );
buf ( n10597 , n2424 );
buf ( n10598 , n2281 );
buf ( n10599 , n2280 );
not ( n10600 , n3260 );
and ( n10601 , n7784 , n5250 );
and ( n10602 , n4162 , n10238 );
or ( n10603 , n10601 , n10602 );
and ( n10604 , n10603 , n5286 );
and ( n10605 , n7795 , n5250 );
and ( n10606 , n4162 , n10238 );
or ( n10607 , n10605 , n10606 );
and ( n10608 , n10607 , n6219 );
and ( n10609 , n7806 , n5250 );
and ( n10610 , n4162 , n10238 );
or ( n10611 , n10609 , n10610 );
and ( n10612 , n10611 , n6711 );
and ( n10613 , n5658 , n5250 );
and ( n10614 , n4162 , n10238 );
or ( n10615 , n10613 , n10614 );
and ( n10616 , n10615 , n6718 );
and ( n10617 , n7818 , n5250 );
and ( n10618 , n4162 , n10238 );
or ( n10619 , n10617 , n10618 );
and ( n10620 , n10619 , n6725 );
and ( n10621 , n4162 , n9116 );
or ( n10622 , n10604 , n10608 , n10612 , n10616 , n10620 , n10621 );
and ( n10623 , n10600 , n10622 );
and ( n10624 , n4162 , n3260 );
or ( n10625 , n10623 , n10624 );
and ( n10626 , n10625 , n2422 );
and ( n10627 , n4162 , n2428 );
or ( n10628 , n10626 , n10627 );
buf ( n10629 , n10628 );
buf ( n10630 , n2424 );
buf ( n10631 , n2281 );
buf ( n10632 , n2280 );
not ( n10633 , n3260 );
and ( n10634 , n7858 , n5250 );
and ( n10635 , n4152 , n10238 );
or ( n10636 , n10634 , n10635 );
and ( n10637 , n10636 , n5286 );
and ( n10638 , n7869 , n5250 );
and ( n10639 , n4152 , n10238 );
or ( n10640 , n10638 , n10639 );
and ( n10641 , n10640 , n6219 );
and ( n10642 , n7880 , n5250 );
and ( n10643 , n4152 , n10238 );
or ( n10644 , n10642 , n10643 );
and ( n10645 , n10644 , n6711 );
and ( n10646 , n5648 , n5250 );
and ( n10647 , n4152 , n10238 );
or ( n10648 , n10646 , n10647 );
and ( n10649 , n10648 , n6718 );
and ( n10650 , n7892 , n5250 );
and ( n10651 , n4152 , n10238 );
or ( n10652 , n10650 , n10651 );
and ( n10653 , n10652 , n6725 );
and ( n10654 , n4152 , n9116 );
or ( n10655 , n10637 , n10641 , n10645 , n10649 , n10653 , n10654 );
and ( n10656 , n10633 , n10655 );
and ( n10657 , n4152 , n3260 );
or ( n10658 , n10656 , n10657 );
and ( n10659 , n10658 , n2422 );
and ( n10660 , n4152 , n2428 );
or ( n10661 , n10659 , n10660 );
buf ( n10662 , n10661 );
buf ( n10663 , n2424 );
buf ( n10664 , n2281 );
buf ( n10665 , n2280 );
not ( n10666 , n3260 );
and ( n10667 , n7932 , n5250 );
and ( n10668 , n4142 , n10238 );
or ( n10669 , n10667 , n10668 );
and ( n10670 , n10669 , n5286 );
and ( n10671 , n7943 , n5250 );
and ( n10672 , n4142 , n10238 );
or ( n10673 , n10671 , n10672 );
and ( n10674 , n10673 , n6219 );
and ( n10675 , n7954 , n5250 );
and ( n10676 , n4142 , n10238 );
or ( n10677 , n10675 , n10676 );
and ( n10678 , n10677 , n6711 );
and ( n10679 , n5638 , n5250 );
and ( n10680 , n4142 , n10238 );
or ( n10681 , n10679 , n10680 );
and ( n10682 , n10681 , n6718 );
and ( n10683 , n7966 , n5250 );
and ( n10684 , n4142 , n10238 );
or ( n10685 , n10683 , n10684 );
and ( n10686 , n10685 , n6725 );
and ( n10687 , n4142 , n9116 );
or ( n10688 , n10670 , n10674 , n10678 , n10682 , n10686 , n10687 );
and ( n10689 , n10666 , n10688 );
and ( n10690 , n4142 , n3260 );
or ( n10691 , n10689 , n10690 );
and ( n10692 , n10691 , n2422 );
and ( n10693 , n4142 , n2428 );
or ( n10694 , n10692 , n10693 );
buf ( n10695 , n10694 );
buf ( n10696 , n2424 );
buf ( n10697 , n2281 );
buf ( n10698 , n2280 );
not ( n10699 , n3260 );
and ( n10700 , n8006 , n5250 );
and ( n10701 , n4132 , n10238 );
or ( n10702 , n10700 , n10701 );
and ( n10703 , n10702 , n5286 );
and ( n10704 , n8017 , n5250 );
and ( n10705 , n4132 , n10238 );
or ( n10706 , n10704 , n10705 );
and ( n10707 , n10706 , n6219 );
and ( n10708 , n8028 , n5250 );
and ( n10709 , n4132 , n10238 );
or ( n10710 , n10708 , n10709 );
and ( n10711 , n10710 , n6711 );
and ( n10712 , n5628 , n5250 );
and ( n10713 , n4132 , n10238 );
or ( n10714 , n10712 , n10713 );
and ( n10715 , n10714 , n6718 );
and ( n10716 , n8040 , n5250 );
and ( n10717 , n4132 , n10238 );
or ( n10718 , n10716 , n10717 );
and ( n10719 , n10718 , n6725 );
and ( n10720 , n4132 , n9116 );
or ( n10721 , n10703 , n10707 , n10711 , n10715 , n10719 , n10720 );
and ( n10722 , n10699 , n10721 );
and ( n10723 , n4132 , n3260 );
or ( n10724 , n10722 , n10723 );
and ( n10725 , n10724 , n2422 );
and ( n10726 , n4132 , n2428 );
or ( n10727 , n10725 , n10726 );
buf ( n10728 , n10727 );
buf ( n10729 , n2424 );
buf ( n10730 , n2281 );
buf ( n10731 , n2280 );
not ( n10732 , n3260 );
and ( n10733 , n8080 , n5250 );
and ( n10734 , n4122 , n10238 );
or ( n10735 , n10733 , n10734 );
and ( n10736 , n10735 , n5286 );
and ( n10737 , n8091 , n5250 );
and ( n10738 , n4122 , n10238 );
or ( n10739 , n10737 , n10738 );
and ( n10740 , n10739 , n6219 );
and ( n10741 , n8102 , n5250 );
and ( n10742 , n4122 , n10238 );
or ( n10743 , n10741 , n10742 );
and ( n10744 , n10743 , n6711 );
and ( n10745 , n5618 , n5250 );
and ( n10746 , n4122 , n10238 );
or ( n10747 , n10745 , n10746 );
and ( n10748 , n10747 , n6718 );
and ( n10749 , n8114 , n5250 );
and ( n10750 , n4122 , n10238 );
or ( n10751 , n10749 , n10750 );
and ( n10752 , n10751 , n6725 );
and ( n10753 , n4122 , n9116 );
or ( n10754 , n10736 , n10740 , n10744 , n10748 , n10752 , n10753 );
and ( n10755 , n10732 , n10754 );
and ( n10756 , n4122 , n3260 );
or ( n10757 , n10755 , n10756 );
and ( n10758 , n10757 , n2422 );
and ( n10759 , n4122 , n2428 );
or ( n10760 , n10758 , n10759 );
buf ( n10761 , n10760 );
buf ( n10762 , n2424 );
buf ( n10763 , n2281 );
buf ( n10764 , n2280 );
not ( n10765 , n3260 );
and ( n10766 , n8154 , n5250 );
and ( n10767 , n4112 , n10238 );
or ( n10768 , n10766 , n10767 );
and ( n10769 , n10768 , n5286 );
and ( n10770 , n8165 , n5250 );
and ( n10771 , n4112 , n10238 );
or ( n10772 , n10770 , n10771 );
and ( n10773 , n10772 , n6219 );
and ( n10774 , n8176 , n5250 );
and ( n10775 , n4112 , n10238 );
or ( n10776 , n10774 , n10775 );
and ( n10777 , n10776 , n6711 );
and ( n10778 , n5608 , n5250 );
and ( n10779 , n4112 , n10238 );
or ( n10780 , n10778 , n10779 );
and ( n10781 , n10780 , n6718 );
and ( n10782 , n8188 , n5250 );
and ( n10783 , n4112 , n10238 );
or ( n10784 , n10782 , n10783 );
and ( n10785 , n10784 , n6725 );
and ( n10786 , n4112 , n9116 );
or ( n10787 , n10769 , n10773 , n10777 , n10781 , n10785 , n10786 );
and ( n10788 , n10765 , n10787 );
and ( n10789 , n4112 , n3260 );
or ( n10790 , n10788 , n10789 );
and ( n10791 , n10790 , n2422 );
and ( n10792 , n4112 , n2428 );
or ( n10793 , n10791 , n10792 );
buf ( n10794 , n10793 );
buf ( n10795 , n2424 );
buf ( n10796 , n2281 );
buf ( n10797 , n2280 );
not ( n10798 , n3260 );
and ( n10799 , n8228 , n5250 );
and ( n10800 , n4102 , n10238 );
or ( n10801 , n10799 , n10800 );
and ( n10802 , n10801 , n5286 );
and ( n10803 , n8239 , n5250 );
and ( n10804 , n4102 , n10238 );
or ( n10805 , n10803 , n10804 );
and ( n10806 , n10805 , n6219 );
and ( n10807 , n8250 , n5250 );
and ( n10808 , n4102 , n10238 );
or ( n10809 , n10807 , n10808 );
and ( n10810 , n10809 , n6711 );
and ( n10811 , n5598 , n5250 );
and ( n10812 , n4102 , n10238 );
or ( n10813 , n10811 , n10812 );
and ( n10814 , n10813 , n6718 );
and ( n10815 , n8262 , n5250 );
and ( n10816 , n4102 , n10238 );
or ( n10817 , n10815 , n10816 );
and ( n10818 , n10817 , n6725 );
and ( n10819 , n4102 , n9116 );
or ( n10820 , n10802 , n10806 , n10810 , n10814 , n10818 , n10819 );
and ( n10821 , n10798 , n10820 );
and ( n10822 , n4102 , n3260 );
or ( n10823 , n10821 , n10822 );
and ( n10824 , n10823 , n2422 );
and ( n10825 , n4102 , n2428 );
or ( n10826 , n10824 , n10825 );
buf ( n10827 , n10826 );
buf ( n10828 , n2424 );
buf ( n10829 , n2281 );
buf ( n10830 , n2280 );
not ( n10831 , n3260 );
and ( n10832 , n8302 , n5250 );
and ( n10833 , n4092 , n10238 );
or ( n10834 , n10832 , n10833 );
and ( n10835 , n10834 , n5286 );
and ( n10836 , n8313 , n5250 );
and ( n10837 , n4092 , n10238 );
or ( n10838 , n10836 , n10837 );
and ( n10839 , n10838 , n6219 );
and ( n10840 , n8324 , n5250 );
and ( n10841 , n4092 , n10238 );
or ( n10842 , n10840 , n10841 );
and ( n10843 , n10842 , n6711 );
and ( n10844 , n5588 , n5250 );
and ( n10845 , n4092 , n10238 );
or ( n10846 , n10844 , n10845 );
and ( n10847 , n10846 , n6718 );
and ( n10848 , n8336 , n5250 );
and ( n10849 , n4092 , n10238 );
or ( n10850 , n10848 , n10849 );
and ( n10851 , n10850 , n6725 );
and ( n10852 , n4092 , n9116 );
or ( n10853 , n10835 , n10839 , n10843 , n10847 , n10851 , n10852 );
and ( n10854 , n10831 , n10853 );
and ( n10855 , n4092 , n3260 );
or ( n10856 , n10854 , n10855 );
and ( n10857 , n10856 , n2422 );
and ( n10858 , n4092 , n2428 );
or ( n10859 , n10857 , n10858 );
buf ( n10860 , n10859 );
buf ( n10861 , n2424 );
buf ( n10862 , n2281 );
buf ( n10863 , n2280 );
not ( n10864 , n3260 );
and ( n10865 , n8376 , n5250 );
and ( n10866 , n4082 , n10238 );
or ( n10867 , n10865 , n10866 );
and ( n10868 , n10867 , n5286 );
and ( n10869 , n8387 , n5250 );
and ( n10870 , n4082 , n10238 );
or ( n10871 , n10869 , n10870 );
and ( n10872 , n10871 , n6219 );
and ( n10873 , n8398 , n5250 );
and ( n10874 , n4082 , n10238 );
or ( n10875 , n10873 , n10874 );
and ( n10876 , n10875 , n6711 );
and ( n10877 , n5578 , n5250 );
and ( n10878 , n4082 , n10238 );
or ( n10879 , n10877 , n10878 );
and ( n10880 , n10879 , n6718 );
and ( n10881 , n8410 , n5250 );
and ( n10882 , n4082 , n10238 );
or ( n10883 , n10881 , n10882 );
and ( n10884 , n10883 , n6725 );
and ( n10885 , n4082 , n9116 );
or ( n10886 , n10868 , n10872 , n10876 , n10880 , n10884 , n10885 );
and ( n10887 , n10864 , n10886 );
and ( n10888 , n4082 , n3260 );
or ( n10889 , n10887 , n10888 );
and ( n10890 , n10889 , n2422 );
and ( n10891 , n4082 , n2428 );
or ( n10892 , n10890 , n10891 );
buf ( n10893 , n10892 );
buf ( n10894 , n2424 );
buf ( n10895 , n2281 );
buf ( n10896 , n2280 );
not ( n10897 , n3260 );
and ( n10898 , n8450 , n5250 );
and ( n10899 , n4072 , n10238 );
or ( n10900 , n10898 , n10899 );
and ( n10901 , n10900 , n5286 );
and ( n10902 , n8461 , n5250 );
and ( n10903 , n4072 , n10238 );
or ( n10904 , n10902 , n10903 );
and ( n10905 , n10904 , n6219 );
and ( n10906 , n8472 , n5250 );
and ( n10907 , n4072 , n10238 );
or ( n10908 , n10906 , n10907 );
and ( n10909 , n10908 , n6711 );
and ( n10910 , n5530 , n5250 );
and ( n10911 , n4072 , n10238 );
or ( n10912 , n10910 , n10911 );
and ( n10913 , n10912 , n6718 );
and ( n10914 , n8484 , n5250 );
and ( n10915 , n4072 , n10238 );
or ( n10916 , n10914 , n10915 );
and ( n10917 , n10916 , n6725 );
and ( n10918 , n4072 , n9116 );
or ( n10919 , n10901 , n10905 , n10909 , n10913 , n10917 , n10918 );
and ( n10920 , n10897 , n10919 );
and ( n10921 , n4072 , n3260 );
or ( n10922 , n10920 , n10921 );
and ( n10923 , n10922 , n2422 );
and ( n10924 , n4072 , n2428 );
or ( n10925 , n10923 , n10924 );
buf ( n10926 , n10925 );
buf ( n10927 , n2424 );
buf ( n10928 , n2281 );
buf ( n10929 , n2280 );
not ( n10930 , n3260 );
and ( n10931 , n8524 , n5250 );
and ( n10932 , n4062 , n10238 );
or ( n10933 , n10931 , n10932 );
and ( n10934 , n10933 , n5286 );
and ( n10935 , n8535 , n5250 );
and ( n10936 , n4062 , n10238 );
or ( n10937 , n10935 , n10936 );
and ( n10938 , n10937 , n6219 );
and ( n10939 , n8546 , n5250 );
and ( n10940 , n4062 , n10238 );
or ( n10941 , n10939 , n10940 );
and ( n10942 , n10941 , n6711 );
and ( n10943 , n5527 , n5250 );
and ( n10944 , n4062 , n10238 );
or ( n10945 , n10943 , n10944 );
and ( n10946 , n10945 , n6718 );
and ( n10947 , n8558 , n5250 );
and ( n10948 , n4062 , n10238 );
or ( n10949 , n10947 , n10948 );
and ( n10950 , n10949 , n6725 );
and ( n10951 , n4062 , n9116 );
or ( n10952 , n10934 , n10938 , n10942 , n10946 , n10950 , n10951 );
and ( n10953 , n10930 , n10952 );
and ( n10954 , n4062 , n3260 );
or ( n10955 , n10953 , n10954 );
and ( n10956 , n10955 , n2422 );
and ( n10957 , n4062 , n2428 );
or ( n10958 , n10956 , n10957 );
buf ( n10959 , n10958 );
buf ( n10960 , n2424 );
buf ( n10961 , n2281 );
buf ( n10962 , n2280 );
not ( n10963 , n3260 );
and ( n10964 , n8598 , n5250 );
and ( n10965 , n4052 , n10238 );
or ( n10966 , n10964 , n10965 );
and ( n10967 , n10966 , n5286 );
and ( n10968 , n8609 , n5250 );
and ( n10969 , n4052 , n10238 );
or ( n10970 , n10968 , n10969 );
and ( n10971 , n10970 , n6219 );
and ( n10972 , n8620 , n5250 );
and ( n10973 , n4052 , n10238 );
or ( n10974 , n10972 , n10973 );
and ( n10975 , n10974 , n6711 );
and ( n10976 , n5524 , n5250 );
and ( n10977 , n4052 , n10238 );
or ( n10978 , n10976 , n10977 );
and ( n10979 , n10978 , n6718 );
and ( n10980 , n8632 , n5250 );
and ( n10981 , n4052 , n10238 );
or ( n10982 , n10980 , n10981 );
and ( n10983 , n10982 , n6725 );
and ( n10984 , n4052 , n9116 );
or ( n10985 , n10967 , n10971 , n10975 , n10979 , n10983 , n10984 );
and ( n10986 , n10963 , n10985 );
and ( n10987 , n4052 , n3260 );
or ( n10988 , n10986 , n10987 );
and ( n10989 , n10988 , n2422 );
and ( n10990 , n4052 , n2428 );
or ( n10991 , n10989 , n10990 );
buf ( n10992 , n10991 );
buf ( n10993 , n2424 );
buf ( n10994 , n2281 );
buf ( n10995 , n2280 );
not ( n10996 , n3260 );
and ( n10997 , n8672 , n5250 );
and ( n10998 , n4042 , n10238 );
or ( n10999 , n10997 , n10998 );
and ( n11000 , n10999 , n5286 );
and ( n11001 , n8683 , n5250 );
and ( n11002 , n4042 , n10238 );
or ( n11003 , n11001 , n11002 );
and ( n11004 , n11003 , n6219 );
and ( n11005 , n8694 , n5250 );
and ( n11006 , n4042 , n10238 );
or ( n11007 , n11005 , n11006 );
and ( n11008 , n11007 , n6711 );
and ( n11009 , n5521 , n5250 );
and ( n11010 , n4042 , n10238 );
or ( n11011 , n11009 , n11010 );
and ( n11012 , n11011 , n6718 );
and ( n11013 , n8706 , n5250 );
and ( n11014 , n4042 , n10238 );
or ( n11015 , n11013 , n11014 );
and ( n11016 , n11015 , n6725 );
and ( n11017 , n4042 , n9116 );
or ( n11018 , n11000 , n11004 , n11008 , n11012 , n11016 , n11017 );
and ( n11019 , n10996 , n11018 );
and ( n11020 , n4042 , n3260 );
or ( n11021 , n11019 , n11020 );
and ( n11022 , n11021 , n2422 );
and ( n11023 , n4042 , n2428 );
or ( n11024 , n11022 , n11023 );
buf ( n11025 , n11024 );
buf ( n11026 , n2424 );
buf ( n11027 , n2281 );
buf ( n11028 , n2280 );
not ( n11029 , n3260 );
and ( n11030 , n8746 , n5250 );
and ( n11031 , n4032 , n10238 );
or ( n11032 , n11030 , n11031 );
and ( n11033 , n11032 , n5286 );
and ( n11034 , n8757 , n5250 );
and ( n11035 , n4032 , n10238 );
or ( n11036 , n11034 , n11035 );
and ( n11037 , n11036 , n6219 );
and ( n11038 , n8768 , n5250 );
and ( n11039 , n4032 , n10238 );
or ( n11040 , n11038 , n11039 );
and ( n11041 , n11040 , n6711 );
and ( n11042 , n5518 , n5250 );
and ( n11043 , n4032 , n10238 );
or ( n11044 , n11042 , n11043 );
and ( n11045 , n11044 , n6718 );
and ( n11046 , n8780 , n5250 );
and ( n11047 , n4032 , n10238 );
or ( n11048 , n11046 , n11047 );
and ( n11049 , n11048 , n6725 );
and ( n11050 , n4032 , n9116 );
or ( n11051 , n11033 , n11037 , n11041 , n11045 , n11049 , n11050 );
and ( n11052 , n11029 , n11051 );
and ( n11053 , n4032 , n3260 );
or ( n11054 , n11052 , n11053 );
and ( n11055 , n11054 , n2422 );
and ( n11056 , n4032 , n2428 );
or ( n11057 , n11055 , n11056 );
buf ( n11058 , n11057 );
buf ( n11059 , n2424 );
buf ( n11060 , n2281 );
buf ( n11061 , n2280 );
not ( n11062 , n3260 );
and ( n11063 , n8820 , n5250 );
and ( n11064 , n4022 , n10238 );
or ( n11065 , n11063 , n11064 );
and ( n11066 , n11065 , n5286 );
and ( n11067 , n8831 , n5250 );
and ( n11068 , n4022 , n10238 );
or ( n11069 , n11067 , n11068 );
and ( n11070 , n11069 , n6219 );
and ( n11071 , n8842 , n5250 );
and ( n11072 , n4022 , n10238 );
or ( n11073 , n11071 , n11072 );
and ( n11074 , n11073 , n6711 );
and ( n11075 , n5515 , n5250 );
and ( n11076 , n4022 , n10238 );
or ( n11077 , n11075 , n11076 );
and ( n11078 , n11077 , n6718 );
and ( n11079 , n8854 , n5250 );
and ( n11080 , n4022 , n10238 );
or ( n11081 , n11079 , n11080 );
and ( n11082 , n11081 , n6725 );
and ( n11083 , n4022 , n9116 );
or ( n11084 , n11066 , n11070 , n11074 , n11078 , n11082 , n11083 );
and ( n11085 , n11062 , n11084 );
and ( n11086 , n4022 , n3260 );
or ( n11087 , n11085 , n11086 );
and ( n11088 , n11087 , n2422 );
and ( n11089 , n4022 , n2428 );
or ( n11090 , n11088 , n11089 );
buf ( n11091 , n11090 );
buf ( n11092 , n2424 );
buf ( n11093 , n2281 );
buf ( n11094 , n2280 );
not ( n11095 , n3260 );
and ( n11096 , n8894 , n5250 );
and ( n11097 , n4012 , n10238 );
or ( n11098 , n11096 , n11097 );
and ( n11099 , n11098 , n5286 );
and ( n11100 , n8905 , n5250 );
and ( n11101 , n4012 , n10238 );
or ( n11102 , n11100 , n11101 );
and ( n11103 , n11102 , n6219 );
and ( n11104 , n8916 , n5250 );
and ( n11105 , n4012 , n10238 );
or ( n11106 , n11104 , n11105 );
and ( n11107 , n11106 , n6711 );
and ( n11108 , n5512 , n5250 );
and ( n11109 , n4012 , n10238 );
or ( n11110 , n11108 , n11109 );
and ( n11111 , n11110 , n6718 );
and ( n11112 , n8928 , n5250 );
and ( n11113 , n4012 , n10238 );
or ( n11114 , n11112 , n11113 );
and ( n11115 , n11114 , n6725 );
and ( n11116 , n4012 , n9116 );
or ( n11117 , n11099 , n11103 , n11107 , n11111 , n11115 , n11116 );
and ( n11118 , n11095 , n11117 );
and ( n11119 , n4012 , n3260 );
or ( n11120 , n11118 , n11119 );
and ( n11121 , n11120 , n2422 );
and ( n11122 , n4012 , n2428 );
or ( n11123 , n11121 , n11122 );
buf ( n11124 , n11123 );
buf ( n11125 , n2424 );
buf ( n11126 , n2281 );
buf ( n11127 , n2280 );
not ( n11128 , n3260 );
and ( n11129 , n8968 , n5250 );
and ( n11130 , n4002 , n10238 );
or ( n11131 , n11129 , n11130 );
and ( n11132 , n11131 , n5286 );
and ( n11133 , n8979 , n5250 );
and ( n11134 , n4002 , n10238 );
or ( n11135 , n11133 , n11134 );
and ( n11136 , n11135 , n6219 );
and ( n11137 , n8990 , n5250 );
and ( n11138 , n4002 , n10238 );
or ( n11139 , n11137 , n11138 );
and ( n11140 , n11139 , n6711 );
and ( n11141 , n5509 , n5250 );
and ( n11142 , n4002 , n10238 );
or ( n11143 , n11141 , n11142 );
and ( n11144 , n11143 , n6718 );
and ( n11145 , n9002 , n5250 );
and ( n11146 , n4002 , n10238 );
or ( n11147 , n11145 , n11146 );
and ( n11148 , n11147 , n6725 );
and ( n11149 , n4002 , n9116 );
or ( n11150 , n11132 , n11136 , n11140 , n11144 , n11148 , n11149 );
and ( n11151 , n11128 , n11150 );
and ( n11152 , n4002 , n3260 );
or ( n11153 , n11151 , n11152 );
and ( n11154 , n11153 , n2422 );
and ( n11155 , n4002 , n2428 );
or ( n11156 , n11154 , n11155 );
buf ( n11157 , n11156 );
buf ( n11158 , n2424 );
buf ( n11159 , n2281 );
buf ( n11160 , n2280 );
not ( n11161 , n3260 );
and ( n11162 , n9042 , n5250 );
and ( n11163 , n3992 , n10238 );
or ( n11164 , n11162 , n11163 );
and ( n11165 , n11164 , n5286 );
and ( n11166 , n9053 , n5250 );
and ( n11167 , n3992 , n10238 );
or ( n11168 , n11166 , n11167 );
and ( n11169 , n11168 , n6219 );
and ( n11170 , n9064 , n5250 );
and ( n11171 , n3992 , n10238 );
or ( n11172 , n11170 , n11171 );
and ( n11173 , n11172 , n6711 );
and ( n11174 , n5506 , n5250 );
and ( n11175 , n3992 , n10238 );
or ( n11176 , n11174 , n11175 );
and ( n11177 , n11176 , n6718 );
and ( n11178 , n9076 , n5250 );
and ( n11179 , n3992 , n10238 );
or ( n11180 , n11178 , n11179 );
and ( n11181 , n11180 , n6725 );
and ( n11182 , n3992 , n9116 );
or ( n11183 , n11165 , n11169 , n11173 , n11177 , n11181 , n11182 );
and ( n11184 , n11161 , n11183 );
and ( n11185 , n3992 , n3260 );
or ( n11186 , n11184 , n11185 );
and ( n11187 , n11186 , n2422 );
and ( n11188 , n3992 , n2428 );
or ( n11189 , n11187 , n11188 );
buf ( n11190 , n11189 );
buf ( n11191 , n2424 );
buf ( n11192 , n2281 );
buf ( n11193 , n2280 );
not ( n11194 , n3260 );
and ( n11195 , n10079 , n5250 );
and ( n11196 , n3982 , n10238 );
or ( n11197 , n11195 , n11196 );
and ( n11198 , n11197 , n5286 );
and ( n11199 , n10090 , n5250 );
and ( n11200 , n3982 , n10238 );
or ( n11201 , n11199 , n11200 );
and ( n11202 , n11201 , n6219 );
and ( n11203 , n10101 , n5250 );
and ( n11204 , n3982 , n10238 );
or ( n11205 , n11203 , n11204 );
and ( n11206 , n11205 , n6711 );
and ( n11207 , n5503 , n5250 );
and ( n11208 , n3982 , n10238 );
or ( n11209 , n11207 , n11208 );
and ( n11210 , n11209 , n6718 );
and ( n11211 , n10112 , n5250 );
and ( n11212 , n3982 , n10238 );
or ( n11213 , n11211 , n11212 );
and ( n11214 , n11213 , n6725 );
and ( n11215 , n3982 , n9116 );
or ( n11216 , n11198 , n11202 , n11206 , n11210 , n11214 , n11215 );
and ( n11217 , n11194 , n11216 );
and ( n11218 , n3982 , n3260 );
or ( n11219 , n11217 , n11218 );
and ( n11220 , n11219 , n2422 );
and ( n11221 , n3982 , n2428 );
or ( n11222 , n11220 , n11221 );
buf ( n11223 , n11222 );
buf ( n11224 , n2424 );
buf ( n11225 , n2281 );
buf ( n11226 , n2280 );
not ( n11227 , n3260 );
and ( n11228 , n10148 , n5250 );
and ( n11229 , n3817 , n10238 );
or ( n11230 , n11228 , n11229 );
and ( n11231 , n11230 , n5286 );
and ( n11232 , n10157 , n5250 );
and ( n11233 , n3817 , n10238 );
or ( n11234 , n11232 , n11233 );
and ( n11235 , n11234 , n6219 );
and ( n11236 , n10166 , n5250 );
and ( n11237 , n3817 , n10238 );
or ( n11238 , n11236 , n11237 );
and ( n11239 , n11238 , n6711 );
and ( n11240 , n5500 , n5250 );
and ( n11241 , n3817 , n10238 );
or ( n11242 , n11240 , n11241 );
and ( n11243 , n11242 , n6718 );
and ( n11244 , n10177 , n5250 );
and ( n11245 , n3817 , n10238 );
or ( n11246 , n11244 , n11245 );
and ( n11247 , n11246 , n6725 );
and ( n11248 , n3817 , n9116 );
or ( n11249 , n11231 , n11235 , n11239 , n11243 , n11247 , n11248 );
and ( n11250 , n11227 , n11249 );
and ( n11251 , n3817 , n3260 );
or ( n11252 , n11250 , n11251 );
and ( n11253 , n11252 , n2422 );
and ( n11254 , n3817 , n2428 );
or ( n11255 , n11253 , n11254 );
buf ( n11256 , n11255 );
buf ( n11257 , n2424 );
buf ( n11258 , n2281 );
buf ( n11259 , n2280 );
not ( n11260 , n3260 );
and ( n11261 , n10202 , n5250 );
and ( n11262 , n3767 , n10238 );
or ( n11263 , n11261 , n11262 );
and ( n11264 , n11263 , n5286 );
and ( n11265 , n3767 , n10238 );
and ( n11266 , n11265 , n6219 );
and ( n11267 , n3767 , n10238 );
and ( n11268 , n11267 , n6711 );
and ( n11269 , n5497 , n5250 );
and ( n11270 , n3767 , n10238 );
or ( n11271 , n11269 , n11270 );
and ( n11272 , n11271 , n6718 );
and ( n11273 , n10217 , n5250 );
and ( n11274 , n3767 , n10238 );
or ( n11275 , n11273 , n11274 );
and ( n11276 , n11275 , n6725 );
and ( n11277 , n3767 , n9116 );
or ( n11278 , n11264 , n11266 , n11268 , n11272 , n11276 , n11277 );
and ( n11279 , n11260 , n11278 );
and ( n11280 , n3767 , n3260 );
or ( n11281 , n11279 , n11280 );
and ( n11282 , n11281 , n2422 );
and ( n11283 , n3767 , n2428 );
or ( n11284 , n11282 , n11283 );
buf ( n11285 , n11284 );
buf ( n11286 , n2424 );
buf ( n11287 , n2281 );
buf ( n11288 , n2280 );
not ( n11289 , n3066 );
not ( n11290 , n3259 );
and ( n11291 , n10134 , n5290 );
or ( n11292 , n5153 , n5155 );
or ( n11293 , n11292 , n5288 );
and ( n11294 , n3290 , n11293 );
or ( n11295 , n11291 , n11294 );
and ( n11296 , n11295 , n5286 );
or ( n11297 , n6720 , n6725 );
or ( n11298 , n11297 , n6716 );
or ( n11299 , n11298 , n6717 );
or ( n11300 , n11299 , n6705 );
or ( n11301 , n11300 , n6706 );
or ( n11302 , n11301 , n6213 );
or ( n11303 , n11302 , n6214 );
or ( n11304 , n11303 , n6708 );
or ( n11305 , n11304 , n6216 );
or ( n11306 , n11305 , n6710 );
or ( n11307 , n11306 , n6218 );
or ( n11308 , n11307 , n3631 );
and ( n11309 , n3290 , n11308 );
or ( n11310 , n11296 , n11309 );
and ( n11311 , n11290 , n11310 );
and ( n11312 , n3290 , n3259 );
or ( n11313 , n11311 , n11312 );
and ( n11314 , n11289 , n11313 );
not ( n11315 , n3770 );
and ( n11316 , n11315 , n3819 );
not ( n11317 , n11316 );
and ( n11318 , n11317 , n3770 );
xnor ( n11319 , n3770 , n3819 );
and ( n11320 , n11319 , n11316 );
or ( n11321 , n11318 , n11320 );
xor ( n11322 , n11321 , n5497 );
not ( n11323 , n11322 );
not ( n11324 , n11316 );
and ( n11325 , n11324 , n3819 );
not ( n11326 , n3819 );
and ( n11327 , n11326 , n11316 );
or ( n11328 , n11325 , n11327 );
not ( n11329 , n11328 );
and ( n11330 , n11329 , n5500 );
not ( n11331 , n3984 );
and ( n11332 , n11331 , n5503 );
not ( n11333 , n3994 );
and ( n11334 , n11333 , n5506 );
not ( n11335 , n4004 );
and ( n11336 , n11335 , n5509 );
not ( n11337 , n4014 );
and ( n11338 , n11337 , n5512 );
not ( n11339 , n4024 );
and ( n11340 , n11339 , n5515 );
not ( n11341 , n4034 );
and ( n11342 , n11341 , n5518 );
not ( n11343 , n4044 );
and ( n11344 , n11343 , n5521 );
not ( n11345 , n4054 );
and ( n11346 , n11345 , n5524 );
not ( n11347 , n4064 );
and ( n11348 , n11347 , n5527 );
not ( n11349 , n4074 );
and ( n11350 , n11349 , n5530 );
not ( n11351 , n4084 );
and ( n11352 , n11351 , n5578 );
not ( n11353 , n4094 );
and ( n11354 , n11353 , n5588 );
not ( n11355 , n4104 );
and ( n11356 , n11355 , n5598 );
not ( n11357 , n4114 );
and ( n11358 , n11357 , n5608 );
not ( n11359 , n4124 );
and ( n11360 , n11359 , n5618 );
not ( n11361 , n4134 );
and ( n11362 , n11361 , n5628 );
not ( n11363 , n4144 );
and ( n11364 , n11363 , n5638 );
not ( n11365 , n4154 );
and ( n11366 , n11365 , n5648 );
not ( n11367 , n4164 );
and ( n11368 , n11367 , n5658 );
not ( n11369 , n4174 );
and ( n11370 , n11369 , n5668 );
not ( n11371 , n4184 );
and ( n11372 , n11371 , n5678 );
not ( n11373 , n4194 );
and ( n11374 , n11373 , n5688 );
not ( n11375 , n4204 );
and ( n11376 , n11375 , n5698 );
not ( n11377 , n4214 );
and ( n11378 , n11377 , n5708 );
not ( n11379 , n4224 );
and ( n11380 , n11379 , n5718 );
not ( n11381 , n4234 );
and ( n11382 , n11381 , n5728 );
not ( n11383 , n4244 );
and ( n11384 , n11383 , n5738 );
not ( n11385 , n4258 );
and ( n11386 , n11385 , n5748 );
not ( n11387 , n3785 );
and ( n11388 , n11387 , n5758 );
not ( n11389 , n3795 );
and ( n11390 , n11389 , n5493 );
xnor ( n11391 , n3785 , n5758 );
and ( n11392 , n11390 , n11391 );
or ( n11393 , n11388 , n11392 );
xnor ( n11394 , n4258 , n5748 );
and ( n11395 , n11393 , n11394 );
or ( n11396 , n11386 , n11395 );
xnor ( n11397 , n4244 , n5738 );
and ( n11398 , n11396 , n11397 );
or ( n11399 , n11384 , n11398 );
xnor ( n11400 , n4234 , n5728 );
and ( n11401 , n11399 , n11400 );
or ( n11402 , n11382 , n11401 );
xnor ( n11403 , n4224 , n5718 );
and ( n11404 , n11402 , n11403 );
or ( n11405 , n11380 , n11404 );
xnor ( n11406 , n4214 , n5708 );
and ( n11407 , n11405 , n11406 );
or ( n11408 , n11378 , n11407 );
xnor ( n11409 , n4204 , n5698 );
and ( n11410 , n11408 , n11409 );
or ( n11411 , n11376 , n11410 );
xnor ( n11412 , n4194 , n5688 );
and ( n11413 , n11411 , n11412 );
or ( n11414 , n11374 , n11413 );
xnor ( n11415 , n4184 , n5678 );
and ( n11416 , n11414 , n11415 );
or ( n11417 , n11372 , n11416 );
xnor ( n11418 , n4174 , n5668 );
and ( n11419 , n11417 , n11418 );
or ( n11420 , n11370 , n11419 );
xnor ( n11421 , n4164 , n5658 );
and ( n11422 , n11420 , n11421 );
or ( n11423 , n11368 , n11422 );
xnor ( n11424 , n4154 , n5648 );
and ( n11425 , n11423 , n11424 );
or ( n11426 , n11366 , n11425 );
xnor ( n11427 , n4144 , n5638 );
and ( n11428 , n11426 , n11427 );
or ( n11429 , n11364 , n11428 );
xnor ( n11430 , n4134 , n5628 );
and ( n11431 , n11429 , n11430 );
or ( n11432 , n11362 , n11431 );
xnor ( n11433 , n4124 , n5618 );
and ( n11434 , n11432 , n11433 );
or ( n11435 , n11360 , n11434 );
xnor ( n11436 , n4114 , n5608 );
and ( n11437 , n11435 , n11436 );
or ( n11438 , n11358 , n11437 );
xnor ( n11439 , n4104 , n5598 );
and ( n11440 , n11438 , n11439 );
or ( n11441 , n11356 , n11440 );
xnor ( n11442 , n4094 , n5588 );
and ( n11443 , n11441 , n11442 );
or ( n11444 , n11354 , n11443 );
xnor ( n11445 , n4084 , n5578 );
and ( n11446 , n11444 , n11445 );
or ( n11447 , n11352 , n11446 );
xnor ( n11448 , n4074 , n5530 );
and ( n11449 , n11447 , n11448 );
or ( n11450 , n11350 , n11449 );
xnor ( n11451 , n4064 , n5527 );
and ( n11452 , n11450 , n11451 );
or ( n11453 , n11348 , n11452 );
xnor ( n11454 , n4054 , n5524 );
and ( n11455 , n11453 , n11454 );
or ( n11456 , n11346 , n11455 );
xnor ( n11457 , n4044 , n5521 );
and ( n11458 , n11456 , n11457 );
or ( n11459 , n11344 , n11458 );
xnor ( n11460 , n4034 , n5518 );
and ( n11461 , n11459 , n11460 );
or ( n11462 , n11342 , n11461 );
xnor ( n11463 , n4024 , n5515 );
and ( n11464 , n11462 , n11463 );
or ( n11465 , n11340 , n11464 );
xnor ( n11466 , n4014 , n5512 );
and ( n11467 , n11465 , n11466 );
or ( n11468 , n11338 , n11467 );
xnor ( n11469 , n4004 , n5509 );
and ( n11470 , n11468 , n11469 );
or ( n11471 , n11336 , n11470 );
xnor ( n11472 , n3994 , n5506 );
and ( n11473 , n11471 , n11472 );
or ( n11474 , n11334 , n11473 );
xnor ( n11475 , n3984 , n5503 );
and ( n11476 , n11474 , n11475 );
or ( n11477 , n11332 , n11476 );
xnor ( n11478 , n11328 , n5500 );
and ( n11479 , n11477 , n11478 );
or ( n11480 , n11330 , n11479 );
and ( n11481 , n11323 , n11480 );
not ( n11482 , n5497 );
and ( n11483 , n11482 , n11321 );
and ( n11484 , n11483 , n11322 );
or ( n11485 , n11481 , n11484 );
not ( n11486 , n11485 );
or ( n11487 , n11486 , n3290 );
and ( n11488 , n11487 , n3630 );
or ( n11489 , n11485 , n3290 );
and ( n11490 , n11489 , n3628 );
xor ( n11491 , n3770 , n5497 );
not ( n11492 , n11491 );
not ( n11493 , n5500 );
and ( n11494 , n11493 , n3819 );
not ( n11495 , n5503 );
and ( n11496 , n11495 , n3984 );
not ( n11497 , n5506 );
and ( n11498 , n11497 , n3994 );
not ( n11499 , n5509 );
and ( n11500 , n11499 , n4004 );
not ( n11501 , n5512 );
and ( n11502 , n11501 , n4014 );
not ( n11503 , n5515 );
and ( n11504 , n11503 , n4024 );
not ( n11505 , n5518 );
and ( n11506 , n11505 , n4034 );
not ( n11507 , n5521 );
and ( n11508 , n11507 , n4044 );
not ( n11509 , n5524 );
and ( n11510 , n11509 , n4054 );
not ( n11511 , n5527 );
and ( n11512 , n11511 , n4064 );
not ( n11513 , n5530 );
and ( n11514 , n11513 , n4074 );
not ( n11515 , n5578 );
and ( n11516 , n11515 , n4084 );
not ( n11517 , n5588 );
and ( n11518 , n11517 , n4094 );
not ( n11519 , n5598 );
and ( n11520 , n11519 , n4104 );
not ( n11521 , n5608 );
and ( n11522 , n11521 , n4114 );
not ( n11523 , n5618 );
and ( n11524 , n11523 , n4124 );
not ( n11525 , n5628 );
and ( n11526 , n11525 , n4134 );
not ( n11527 , n5638 );
and ( n11528 , n11527 , n4144 );
not ( n11529 , n5648 );
and ( n11530 , n11529 , n4154 );
not ( n11531 , n5658 );
and ( n11532 , n11531 , n4164 );
not ( n11533 , n5668 );
and ( n11534 , n11533 , n4174 );
not ( n11535 , n5678 );
and ( n11536 , n11535 , n4184 );
not ( n11537 , n5688 );
and ( n11538 , n11537 , n4194 );
not ( n11539 , n5698 );
and ( n11540 , n11539 , n4204 );
not ( n11541 , n5708 );
and ( n11542 , n11541 , n4214 );
not ( n11543 , n5718 );
and ( n11544 , n11543 , n4224 );
not ( n11545 , n5728 );
and ( n11546 , n11545 , n4234 );
not ( n11547 , n5738 );
and ( n11548 , n11547 , n4244 );
not ( n11549 , n5748 );
and ( n11550 , n11549 , n4258 );
not ( n11551 , n5758 );
and ( n11552 , n11551 , n3785 );
not ( n11553 , n5493 );
and ( n11554 , n11553 , n3795 );
xnor ( n11555 , n3785 , n5758 );
and ( n11556 , n11554 , n11555 );
or ( n11557 , n11552 , n11556 );
xnor ( n11558 , n4258 , n5748 );
and ( n11559 , n11557 , n11558 );
or ( n11560 , n11550 , n11559 );
xnor ( n11561 , n4244 , n5738 );
and ( n11562 , n11560 , n11561 );
or ( n11563 , n11548 , n11562 );
xnor ( n11564 , n4234 , n5728 );
and ( n11565 , n11563 , n11564 );
or ( n11566 , n11546 , n11565 );
xnor ( n11567 , n4224 , n5718 );
and ( n11568 , n11566 , n11567 );
or ( n11569 , n11544 , n11568 );
xnor ( n11570 , n4214 , n5708 );
and ( n11571 , n11569 , n11570 );
or ( n11572 , n11542 , n11571 );
xnor ( n11573 , n4204 , n5698 );
and ( n11574 , n11572 , n11573 );
or ( n11575 , n11540 , n11574 );
xnor ( n11576 , n4194 , n5688 );
and ( n11577 , n11575 , n11576 );
or ( n11578 , n11538 , n11577 );
xnor ( n11579 , n4184 , n5678 );
and ( n11580 , n11578 , n11579 );
or ( n11581 , n11536 , n11580 );
xnor ( n11582 , n4174 , n5668 );
and ( n11583 , n11581 , n11582 );
or ( n11584 , n11534 , n11583 );
xnor ( n11585 , n4164 , n5658 );
and ( n11586 , n11584 , n11585 );
or ( n11587 , n11532 , n11586 );
xnor ( n11588 , n4154 , n5648 );
and ( n11589 , n11587 , n11588 );
or ( n11590 , n11530 , n11589 );
xnor ( n11591 , n4144 , n5638 );
and ( n11592 , n11590 , n11591 );
or ( n11593 , n11528 , n11592 );
xnor ( n11594 , n4134 , n5628 );
and ( n11595 , n11593 , n11594 );
or ( n11596 , n11526 , n11595 );
xnor ( n11597 , n4124 , n5618 );
and ( n11598 , n11596 , n11597 );
or ( n11599 , n11524 , n11598 );
xnor ( n11600 , n4114 , n5608 );
and ( n11601 , n11599 , n11600 );
or ( n11602 , n11522 , n11601 );
xnor ( n11603 , n4104 , n5598 );
and ( n11604 , n11602 , n11603 );
or ( n11605 , n11520 , n11604 );
xnor ( n11606 , n4094 , n5588 );
and ( n11607 , n11605 , n11606 );
or ( n11608 , n11518 , n11607 );
xnor ( n11609 , n4084 , n5578 );
and ( n11610 , n11608 , n11609 );
or ( n11611 , n11516 , n11610 );
xnor ( n11612 , n4074 , n5530 );
and ( n11613 , n11611 , n11612 );
or ( n11614 , n11514 , n11613 );
xnor ( n11615 , n4064 , n5527 );
and ( n11616 , n11614 , n11615 );
or ( n11617 , n11512 , n11616 );
xnor ( n11618 , n4054 , n5524 );
and ( n11619 , n11617 , n11618 );
or ( n11620 , n11510 , n11619 );
xnor ( n11621 , n4044 , n5521 );
and ( n11622 , n11620 , n11621 );
or ( n11623 , n11508 , n11622 );
xnor ( n11624 , n4034 , n5518 );
and ( n11625 , n11623 , n11624 );
or ( n11626 , n11506 , n11625 );
xnor ( n11627 , n4024 , n5515 );
and ( n11628 , n11626 , n11627 );
or ( n11629 , n11504 , n11628 );
xnor ( n11630 , n4014 , n5512 );
and ( n11631 , n11629 , n11630 );
or ( n11632 , n11502 , n11631 );
xnor ( n11633 , n4004 , n5509 );
and ( n11634 , n11632 , n11633 );
or ( n11635 , n11500 , n11634 );
xnor ( n11636 , n3994 , n5506 );
and ( n11637 , n11635 , n11636 );
or ( n11638 , n11498 , n11637 );
xnor ( n11639 , n3984 , n5503 );
and ( n11640 , n11638 , n11639 );
or ( n11641 , n11496 , n11640 );
xnor ( n11642 , n3819 , n5500 );
and ( n11643 , n11641 , n11642 );
or ( n11644 , n11494 , n11643 );
and ( n11645 , n11492 , n11644 );
not ( n11646 , n3770 );
and ( n11647 , n11646 , n5497 );
and ( n11648 , n11647 , n11491 );
or ( n11649 , n11645 , n11648 );
or ( n11650 , n11649 , n3290 );
and ( n11651 , n11650 , n3626 );
not ( n11652 , n11649 );
or ( n11653 , n11652 , n3290 );
and ( n11654 , n11653 , n5286 );
xor ( n11655 , n3770 , n5497 );
xor ( n11656 , n3819 , n5500 );
or ( n11657 , n11655 , n11656 );
xor ( n11658 , n3984 , n5503 );
or ( n11659 , n11657 , n11658 );
xor ( n11660 , n3994 , n5506 );
or ( n11661 , n11659 , n11660 );
xor ( n11662 , n4004 , n5509 );
or ( n11663 , n11661 , n11662 );
xor ( n11664 , n4014 , n5512 );
or ( n11665 , n11663 , n11664 );
xor ( n11666 , n4024 , n5515 );
or ( n11667 , n11665 , n11666 );
xor ( n11668 , n4034 , n5518 );
or ( n11669 , n11667 , n11668 );
xor ( n11670 , n4044 , n5521 );
or ( n11671 , n11669 , n11670 );
xor ( n11672 , n4054 , n5524 );
or ( n11673 , n11671 , n11672 );
xor ( n11674 , n4064 , n5527 );
or ( n11675 , n11673 , n11674 );
xor ( n11676 , n4074 , n5530 );
or ( n11677 , n11675 , n11676 );
xor ( n11678 , n4084 , n5578 );
or ( n11679 , n11677 , n11678 );
xor ( n11680 , n4094 , n5588 );
or ( n11681 , n11679 , n11680 );
xor ( n11682 , n4104 , n5598 );
or ( n11683 , n11681 , n11682 );
xor ( n11684 , n4114 , n5608 );
or ( n11685 , n11683 , n11684 );
xor ( n11686 , n4124 , n5618 );
or ( n11687 , n11685 , n11686 );
xor ( n11688 , n4134 , n5628 );
or ( n11689 , n11687 , n11688 );
xor ( n11690 , n4144 , n5638 );
or ( n11691 , n11689 , n11690 );
xor ( n11692 , n4154 , n5648 );
or ( n11693 , n11691 , n11692 );
xor ( n11694 , n4164 , n5658 );
or ( n11695 , n11693 , n11694 );
xor ( n11696 , n4174 , n5668 );
or ( n11697 , n11695 , n11696 );
xor ( n11698 , n4184 , n5678 );
or ( n11699 , n11697 , n11698 );
xor ( n11700 , n4194 , n5688 );
or ( n11701 , n11699 , n11700 );
xor ( n11702 , n4204 , n5698 );
or ( n11703 , n11701 , n11702 );
xor ( n11704 , n4214 , n5708 );
or ( n11705 , n11703 , n11704 );
xor ( n11706 , n4224 , n5718 );
or ( n11707 , n11705 , n11706 );
xor ( n11708 , n4234 , n5728 );
or ( n11709 , n11707 , n11708 );
xor ( n11710 , n4244 , n5738 );
or ( n11711 , n11709 , n11710 );
xor ( n11712 , n4258 , n5748 );
or ( n11713 , n11711 , n11712 );
xor ( n11714 , n3785 , n5758 );
or ( n11715 , n11713 , n11714 );
xor ( n11716 , n3795 , n5493 );
or ( n11717 , n11715 , n11716 );
not ( n11718 , n11717 );
not ( n11719 , n11718 );
or ( n11720 , n11719 , n3290 );
and ( n11721 , n11720 , n6218 );
or ( n11722 , n11718 , n3290 );
and ( n11723 , n11722 , n6710 );
xor ( n11724 , n3770 , n5497 );
not ( n11725 , n11724 );
not ( n11726 , n3819 );
and ( n11727 , n11726 , n5500 );
not ( n11728 , n3984 );
and ( n11729 , n11728 , n5503 );
not ( n11730 , n3994 );
and ( n11731 , n11730 , n5506 );
not ( n11732 , n4004 );
and ( n11733 , n11732 , n5509 );
not ( n11734 , n4014 );
and ( n11735 , n11734 , n5512 );
not ( n11736 , n4024 );
and ( n11737 , n11736 , n5515 );
not ( n11738 , n4034 );
and ( n11739 , n11738 , n5518 );
not ( n11740 , n4044 );
and ( n11741 , n11740 , n5521 );
not ( n11742 , n4054 );
and ( n11743 , n11742 , n5524 );
not ( n11744 , n4064 );
and ( n11745 , n11744 , n5527 );
not ( n11746 , n4074 );
and ( n11747 , n11746 , n5530 );
not ( n11748 , n4084 );
and ( n11749 , n11748 , n5578 );
not ( n11750 , n4094 );
and ( n11751 , n11750 , n5588 );
not ( n11752 , n4104 );
and ( n11753 , n11752 , n5598 );
not ( n11754 , n4114 );
and ( n11755 , n11754 , n5608 );
not ( n11756 , n4124 );
and ( n11757 , n11756 , n5618 );
not ( n11758 , n4134 );
and ( n11759 , n11758 , n5628 );
not ( n11760 , n4144 );
and ( n11761 , n11760 , n5638 );
not ( n11762 , n4154 );
and ( n11763 , n11762 , n5648 );
not ( n11764 , n4164 );
and ( n11765 , n11764 , n5658 );
not ( n11766 , n4174 );
and ( n11767 , n11766 , n5668 );
not ( n11768 , n4184 );
and ( n11769 , n11768 , n5678 );
not ( n11770 , n4194 );
and ( n11771 , n11770 , n5688 );
not ( n11772 , n4204 );
and ( n11773 , n11772 , n5698 );
not ( n11774 , n4214 );
and ( n11775 , n11774 , n5708 );
not ( n11776 , n4224 );
and ( n11777 , n11776 , n5718 );
not ( n11778 , n4234 );
and ( n11779 , n11778 , n5728 );
not ( n11780 , n4244 );
and ( n11781 , n11780 , n5738 );
not ( n11782 , n4258 );
and ( n11783 , n11782 , n5748 );
not ( n11784 , n3785 );
and ( n11785 , n11784 , n5758 );
not ( n11786 , n3795 );
and ( n11787 , n11786 , n5493 );
xnor ( n11788 , n3785 , n5758 );
and ( n11789 , n11787 , n11788 );
or ( n11790 , n11785 , n11789 );
xnor ( n11791 , n4258 , n5748 );
and ( n11792 , n11790 , n11791 );
or ( n11793 , n11783 , n11792 );
xnor ( n11794 , n4244 , n5738 );
and ( n11795 , n11793 , n11794 );
or ( n11796 , n11781 , n11795 );
xnor ( n11797 , n4234 , n5728 );
and ( n11798 , n11796 , n11797 );
or ( n11799 , n11779 , n11798 );
xnor ( n11800 , n4224 , n5718 );
and ( n11801 , n11799 , n11800 );
or ( n11802 , n11777 , n11801 );
xnor ( n11803 , n4214 , n5708 );
and ( n11804 , n11802 , n11803 );
or ( n11805 , n11775 , n11804 );
xnor ( n11806 , n4204 , n5698 );
and ( n11807 , n11805 , n11806 );
or ( n11808 , n11773 , n11807 );
xnor ( n11809 , n4194 , n5688 );
and ( n11810 , n11808 , n11809 );
or ( n11811 , n11771 , n11810 );
xnor ( n11812 , n4184 , n5678 );
and ( n11813 , n11811 , n11812 );
or ( n11814 , n11769 , n11813 );
xnor ( n11815 , n4174 , n5668 );
and ( n11816 , n11814 , n11815 );
or ( n11817 , n11767 , n11816 );
xnor ( n11818 , n4164 , n5658 );
and ( n11819 , n11817 , n11818 );
or ( n11820 , n11765 , n11819 );
xnor ( n11821 , n4154 , n5648 );
and ( n11822 , n11820 , n11821 );
or ( n11823 , n11763 , n11822 );
xnor ( n11824 , n4144 , n5638 );
and ( n11825 , n11823 , n11824 );
or ( n11826 , n11761 , n11825 );
xnor ( n11827 , n4134 , n5628 );
and ( n11828 , n11826 , n11827 );
or ( n11829 , n11759 , n11828 );
xnor ( n11830 , n4124 , n5618 );
and ( n11831 , n11829 , n11830 );
or ( n11832 , n11757 , n11831 );
xnor ( n11833 , n4114 , n5608 );
and ( n11834 , n11832 , n11833 );
or ( n11835 , n11755 , n11834 );
xnor ( n11836 , n4104 , n5598 );
and ( n11837 , n11835 , n11836 );
or ( n11838 , n11753 , n11837 );
xnor ( n11839 , n4094 , n5588 );
and ( n11840 , n11838 , n11839 );
or ( n11841 , n11751 , n11840 );
xnor ( n11842 , n4084 , n5578 );
and ( n11843 , n11841 , n11842 );
or ( n11844 , n11749 , n11843 );
xnor ( n11845 , n4074 , n5530 );
and ( n11846 , n11844 , n11845 );
or ( n11847 , n11747 , n11846 );
xnor ( n11848 , n4064 , n5527 );
and ( n11849 , n11847 , n11848 );
or ( n11850 , n11745 , n11849 );
xnor ( n11851 , n4054 , n5524 );
and ( n11852 , n11850 , n11851 );
or ( n11853 , n11743 , n11852 );
xnor ( n11854 , n4044 , n5521 );
and ( n11855 , n11853 , n11854 );
or ( n11856 , n11741 , n11855 );
xnor ( n11857 , n4034 , n5518 );
and ( n11858 , n11856 , n11857 );
or ( n11859 , n11739 , n11858 );
xnor ( n11860 , n4024 , n5515 );
and ( n11861 , n11859 , n11860 );
or ( n11862 , n11737 , n11861 );
xnor ( n11863 , n4014 , n5512 );
and ( n11864 , n11862 , n11863 );
or ( n11865 , n11735 , n11864 );
xnor ( n11866 , n4004 , n5509 );
and ( n11867 , n11865 , n11866 );
or ( n11868 , n11733 , n11867 );
xnor ( n11869 , n3994 , n5506 );
and ( n11870 , n11868 , n11869 );
or ( n11871 , n11731 , n11870 );
xnor ( n11872 , n3984 , n5503 );
and ( n11873 , n11871 , n11872 );
or ( n11874 , n11729 , n11873 );
xnor ( n11875 , n3819 , n5500 );
and ( n11876 , n11874 , n11875 );
or ( n11877 , n11727 , n11876 );
and ( n11878 , n11725 , n11877 );
not ( n11879 , n5497 );
and ( n11880 , n11879 , n3770 );
and ( n11881 , n11880 , n11724 );
or ( n11882 , n11878 , n11881 );
not ( n11883 , n11882 );
or ( n11884 , n11883 , n3290 );
and ( n11885 , n11884 , n6216 );
or ( n11886 , n11882 , n3290 );
and ( n11887 , n11886 , n6708 );
and ( n11888 , n11486 , n6214 );
and ( n11889 , n11485 , n6213 );
and ( n11890 , n11649 , n6706 );
and ( n11891 , n11652 , n6705 );
and ( n11892 , n11719 , n6717 );
and ( n11893 , n11718 , n6716 );
and ( n11894 , n11883 , n6720 );
and ( n11895 , n11882 , n6725 );
or ( n11896 , n11488 , n11490 , n11651 , n11654 , n11721 , n11723 , n11885 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 );
and ( n11897 , n11896 , n3066 );
or ( n11898 , n11314 , n11897 );
and ( n11899 , n11898 , n2422 );
and ( n11900 , n3290 , n2428 );
or ( n11901 , n11899 , n11900 );
buf ( n11902 , n11901 );
buf ( n11903 , n2424 );
buf ( n11904 , n2281 );
buf ( n11905 , n2280 );
not ( n11906 , n3260 );
and ( n11907 , n3789 , n3631 );
and ( n11908 , n5157 , n5281 );
or ( n11909 , n5251 , n5189 );
buf ( n11910 , n11909 );
and ( n11911 , n3789 , n11910 );
or ( n11912 , n11908 , n11911 );
and ( n11913 , n11912 , n5286 );
and ( n11914 , n6208 , n5281 );
and ( n11915 , n3789 , n11910 );
or ( n11916 , n11914 , n11915 );
and ( n11917 , n11916 , n6219 );
and ( n11918 , n6701 , n5281 );
and ( n11919 , n3789 , n11910 );
or ( n11920 , n11918 , n11919 );
and ( n11921 , n11920 , n6711 );
and ( n11922 , n5493 , n5281 );
and ( n11923 , n3789 , n11910 );
or ( n11924 , n11922 , n11923 );
and ( n11925 , n11924 , n6718 );
and ( n11926 , n3363 , n6720 );
and ( n11927 , n5493 , n5281 );
and ( n11928 , n3789 , n11910 );
or ( n11929 , n11927 , n11928 );
and ( n11930 , n11929 , n6725 );
or ( n11931 , n11907 , n11913 , n11917 , n11921 , n11925 , n11926 , n11930 );
and ( n11932 , n11906 , n11931 );
and ( n11933 , n3789 , n3260 );
or ( n11934 , n11932 , n11933 );
and ( n11935 , n11934 , n2422 );
and ( n11936 , n3789 , n2428 );
or ( n11937 , n11935 , n11936 );
buf ( n11938 , n11937 );
buf ( n11939 , n2424 );
buf ( n11940 , n2281 );
buf ( n11941 , n2280 );
not ( n11942 , n3260 );
and ( n11943 , n3779 , n3631 );
and ( n11944 , n7044 , n5281 );
and ( n11945 , n3779 , n11910 );
or ( n11946 , n11944 , n11945 );
and ( n11947 , n11946 , n5286 );
and ( n11948 , n7055 , n5281 );
and ( n11949 , n3779 , n11910 );
or ( n11950 , n11948 , n11949 );
and ( n11951 , n11950 , n6219 );
and ( n11952 , n7066 , n5281 );
and ( n11953 , n3779 , n11910 );
or ( n11954 , n11952 , n11953 );
and ( n11955 , n11954 , n6711 );
and ( n11956 , n5758 , n5281 );
and ( n11957 , n3779 , n11910 );
or ( n11958 , n11956 , n11957 );
and ( n11959 , n11958 , n6718 );
and ( n11960 , n3776 , n6720 );
and ( n11961 , n7078 , n5281 );
and ( n11962 , n3779 , n11910 );
or ( n11963 , n11961 , n11962 );
and ( n11964 , n11963 , n6725 );
or ( n11965 , n11943 , n11947 , n11951 , n11955 , n11959 , n11960 , n11964 );
and ( n11966 , n11942 , n11965 );
and ( n11967 , n3779 , n3260 );
or ( n11968 , n11966 , n11967 );
and ( n11969 , n11968 , n2422 );
and ( n11970 , n3779 , n2428 );
or ( n11971 , n11969 , n11970 );
buf ( n11972 , n11971 );
buf ( n11973 , n2424 );
buf ( n11974 , n2281 );
buf ( n11975 , n2280 );
not ( n11976 , n3260 );
and ( n11977 , n4252 , n3631 );
and ( n11978 , n7118 , n5281 );
and ( n11979 , n4252 , n11910 );
or ( n11980 , n11978 , n11979 );
and ( n11981 , n11980 , n5286 );
and ( n11982 , n7129 , n5281 );
and ( n11983 , n4252 , n11910 );
or ( n11984 , n11982 , n11983 );
and ( n11985 , n11984 , n6219 );
and ( n11986 , n7140 , n5281 );
and ( n11987 , n4252 , n11910 );
or ( n11988 , n11986 , n11987 );
and ( n11989 , n11988 , n6711 );
and ( n11990 , n5748 , n5281 );
and ( n11991 , n4252 , n11910 );
or ( n11992 , n11990 , n11991 );
and ( n11993 , n11992 , n6718 );
and ( n11994 , n4250 , n6720 );
and ( n11995 , n7152 , n5281 );
and ( n11996 , n4252 , n11910 );
or ( n11997 , n11995 , n11996 );
and ( n11998 , n11997 , n6725 );
or ( n11999 , n11977 , n11981 , n11985 , n11989 , n11993 , n11994 , n11998 );
and ( n12000 , n11976 , n11999 );
and ( n12001 , n4252 , n3260 );
or ( n12002 , n12000 , n12001 );
and ( n12003 , n12002 , n2422 );
and ( n12004 , n4252 , n2428 );
or ( n12005 , n12003 , n12004 );
buf ( n12006 , n12005 );
buf ( n12007 , n2424 );
buf ( n12008 , n2281 );
buf ( n12009 , n2280 );
not ( n12010 , n3260 );
and ( n12011 , n4238 , n3631 );
and ( n12012 , n7192 , n5281 );
and ( n12013 , n4238 , n11910 );
or ( n12014 , n12012 , n12013 );
and ( n12015 , n12014 , n5286 );
and ( n12016 , n7203 , n5281 );
and ( n12017 , n4238 , n11910 );
or ( n12018 , n12016 , n12017 );
and ( n12019 , n12018 , n6219 );
and ( n12020 , n7214 , n5281 );
and ( n12021 , n4238 , n11910 );
or ( n12022 , n12020 , n12021 );
and ( n12023 , n12022 , n6711 );
and ( n12024 , n5738 , n5281 );
and ( n12025 , n4238 , n11910 );
or ( n12026 , n12024 , n12025 );
and ( n12027 , n12026 , n6718 );
and ( n12028 , n4236 , n6720 );
and ( n12029 , n7226 , n5281 );
and ( n12030 , n4238 , n11910 );
or ( n12031 , n12029 , n12030 );
and ( n12032 , n12031 , n6725 );
or ( n12033 , n12011 , n12015 , n12019 , n12023 , n12027 , n12028 , n12032 );
and ( n12034 , n12010 , n12033 );
and ( n12035 , n4238 , n3260 );
or ( n12036 , n12034 , n12035 );
and ( n12037 , n12036 , n2422 );
and ( n12038 , n4238 , n2428 );
or ( n12039 , n12037 , n12038 );
buf ( n12040 , n12039 );
buf ( n12041 , n2424 );
buf ( n12042 , n2281 );
buf ( n12043 , n2280 );
not ( n12044 , n3260 );
and ( n12045 , n4228 , n3631 );
and ( n12046 , n7266 , n5281 );
and ( n12047 , n4228 , n11910 );
or ( n12048 , n12046 , n12047 );
and ( n12049 , n12048 , n5286 );
and ( n12050 , n7277 , n5281 );
and ( n12051 , n4228 , n11910 );
or ( n12052 , n12050 , n12051 );
and ( n12053 , n12052 , n6219 );
and ( n12054 , n7288 , n5281 );
and ( n12055 , n4228 , n11910 );
or ( n12056 , n12054 , n12055 );
and ( n12057 , n12056 , n6711 );
and ( n12058 , n5728 , n5281 );
and ( n12059 , n4228 , n11910 );
or ( n12060 , n12058 , n12059 );
and ( n12061 , n12060 , n6718 );
and ( n12062 , n4226 , n6720 );
and ( n12063 , n7300 , n5281 );
and ( n12064 , n4228 , n11910 );
or ( n12065 , n12063 , n12064 );
and ( n12066 , n12065 , n6725 );
or ( n12067 , n12045 , n12049 , n12053 , n12057 , n12061 , n12062 , n12066 );
and ( n12068 , n12044 , n12067 );
and ( n12069 , n4228 , n3260 );
or ( n12070 , n12068 , n12069 );
and ( n12071 , n12070 , n2422 );
and ( n12072 , n4228 , n2428 );
or ( n12073 , n12071 , n12072 );
buf ( n12074 , n12073 );
buf ( n12075 , n2424 );
buf ( n12076 , n2281 );
buf ( n12077 , n2280 );
not ( n12078 , n3260 );
and ( n12079 , n4218 , n3631 );
and ( n12080 , n7340 , n5281 );
and ( n12081 , n4218 , n11910 );
or ( n12082 , n12080 , n12081 );
and ( n12083 , n12082 , n5286 );
and ( n12084 , n7351 , n5281 );
and ( n12085 , n4218 , n11910 );
or ( n12086 , n12084 , n12085 );
and ( n12087 , n12086 , n6219 );
and ( n12088 , n7362 , n5281 );
and ( n12089 , n4218 , n11910 );
or ( n12090 , n12088 , n12089 );
and ( n12091 , n12090 , n6711 );
and ( n12092 , n5718 , n5281 );
and ( n12093 , n4218 , n11910 );
or ( n12094 , n12092 , n12093 );
and ( n12095 , n12094 , n6718 );
and ( n12096 , n4216 , n6720 );
and ( n12097 , n7374 , n5281 );
and ( n12098 , n4218 , n11910 );
or ( n12099 , n12097 , n12098 );
and ( n12100 , n12099 , n6725 );
or ( n12101 , n12079 , n12083 , n12087 , n12091 , n12095 , n12096 , n12100 );
and ( n12102 , n12078 , n12101 );
and ( n12103 , n4218 , n3260 );
or ( n12104 , n12102 , n12103 );
and ( n12105 , n12104 , n2422 );
and ( n12106 , n4218 , n2428 );
or ( n12107 , n12105 , n12106 );
buf ( n12108 , n12107 );
buf ( n12109 , n2424 );
buf ( n12110 , n2281 );
buf ( n12111 , n2280 );
not ( n12112 , n3260 );
and ( n12113 , n4208 , n3631 );
and ( n12114 , n7414 , n5281 );
and ( n12115 , n4208 , n11910 );
or ( n12116 , n12114 , n12115 );
and ( n12117 , n12116 , n5286 );
and ( n12118 , n7425 , n5281 );
and ( n12119 , n4208 , n11910 );
or ( n12120 , n12118 , n12119 );
and ( n12121 , n12120 , n6219 );
and ( n12122 , n7436 , n5281 );
and ( n12123 , n4208 , n11910 );
or ( n12124 , n12122 , n12123 );
and ( n12125 , n12124 , n6711 );
and ( n12126 , n5708 , n5281 );
and ( n12127 , n4208 , n11910 );
or ( n12128 , n12126 , n12127 );
and ( n12129 , n12128 , n6718 );
and ( n12130 , n4206 , n6720 );
and ( n12131 , n7448 , n5281 );
and ( n12132 , n4208 , n11910 );
or ( n12133 , n12131 , n12132 );
and ( n12134 , n12133 , n6725 );
or ( n12135 , n12113 , n12117 , n12121 , n12125 , n12129 , n12130 , n12134 );
and ( n12136 , n12112 , n12135 );
and ( n12137 , n4208 , n3260 );
or ( n12138 , n12136 , n12137 );
and ( n12139 , n12138 , n2422 );
and ( n12140 , n4208 , n2428 );
or ( n12141 , n12139 , n12140 );
buf ( n12142 , n12141 );
buf ( n12143 , n2424 );
buf ( n12144 , n2281 );
buf ( n12145 , n2280 );
not ( n12146 , n3260 );
and ( n12147 , n4198 , n3631 );
and ( n12148 , n7488 , n5281 );
and ( n12149 , n4198 , n11910 );
or ( n12150 , n12148 , n12149 );
and ( n12151 , n12150 , n5286 );
and ( n12152 , n7499 , n5281 );
and ( n12153 , n4198 , n11910 );
or ( n12154 , n12152 , n12153 );
and ( n12155 , n12154 , n6219 );
and ( n12156 , n7510 , n5281 );
and ( n12157 , n4198 , n11910 );
or ( n12158 , n12156 , n12157 );
and ( n12159 , n12158 , n6711 );
and ( n12160 , n5698 , n5281 );
and ( n12161 , n4198 , n11910 );
or ( n12162 , n12160 , n12161 );
and ( n12163 , n12162 , n6718 );
and ( n12164 , n4196 , n6720 );
and ( n12165 , n7522 , n5281 );
and ( n12166 , n4198 , n11910 );
or ( n12167 , n12165 , n12166 );
and ( n12168 , n12167 , n6725 );
or ( n12169 , n12147 , n12151 , n12155 , n12159 , n12163 , n12164 , n12168 );
and ( n12170 , n12146 , n12169 );
and ( n12171 , n4198 , n3260 );
or ( n12172 , n12170 , n12171 );
and ( n12173 , n12172 , n2422 );
and ( n12174 , n4198 , n2428 );
or ( n12175 , n12173 , n12174 );
buf ( n12176 , n12175 );
buf ( n12177 , n2424 );
buf ( n12178 , n2281 );
buf ( n12179 , n2280 );
not ( n12180 , n3260 );
and ( n12181 , n4188 , n3631 );
and ( n12182 , n7562 , n5281 );
and ( n12183 , n4188 , n11910 );
or ( n12184 , n12182 , n12183 );
and ( n12185 , n12184 , n5286 );
and ( n12186 , n7573 , n5281 );
and ( n12187 , n4188 , n11910 );
or ( n12188 , n12186 , n12187 );
and ( n12189 , n12188 , n6219 );
and ( n12190 , n7584 , n5281 );
and ( n12191 , n4188 , n11910 );
or ( n12192 , n12190 , n12191 );
and ( n12193 , n12192 , n6711 );
and ( n12194 , n5688 , n5281 );
and ( n12195 , n4188 , n11910 );
or ( n12196 , n12194 , n12195 );
and ( n12197 , n12196 , n6718 );
and ( n12198 , n4186 , n6720 );
and ( n12199 , n7596 , n5281 );
and ( n12200 , n4188 , n11910 );
or ( n12201 , n12199 , n12200 );
and ( n12202 , n12201 , n6725 );
or ( n12203 , n12181 , n12185 , n12189 , n12193 , n12197 , n12198 , n12202 );
and ( n12204 , n12180 , n12203 );
and ( n12205 , n4188 , n3260 );
or ( n12206 , n12204 , n12205 );
and ( n12207 , n12206 , n2422 );
and ( n12208 , n4188 , n2428 );
or ( n12209 , n12207 , n12208 );
buf ( n12210 , n12209 );
buf ( n12211 , n2424 );
buf ( n12212 , n2281 );
buf ( n12213 , n2280 );
not ( n12214 , n3260 );
and ( n12215 , n4178 , n3631 );
and ( n12216 , n7636 , n5281 );
and ( n12217 , n4178 , n11910 );
or ( n12218 , n12216 , n12217 );
and ( n12219 , n12218 , n5286 );
and ( n12220 , n7647 , n5281 );
and ( n12221 , n4178 , n11910 );
or ( n12222 , n12220 , n12221 );
and ( n12223 , n12222 , n6219 );
and ( n12224 , n7658 , n5281 );
and ( n12225 , n4178 , n11910 );
or ( n12226 , n12224 , n12225 );
and ( n12227 , n12226 , n6711 );
and ( n12228 , n5678 , n5281 );
and ( n12229 , n4178 , n11910 );
or ( n12230 , n12228 , n12229 );
and ( n12231 , n12230 , n6718 );
and ( n12232 , n4176 , n6720 );
and ( n12233 , n7670 , n5281 );
and ( n12234 , n4178 , n11910 );
or ( n12235 , n12233 , n12234 );
and ( n12236 , n12235 , n6725 );
or ( n12237 , n12215 , n12219 , n12223 , n12227 , n12231 , n12232 , n12236 );
and ( n12238 , n12214 , n12237 );
and ( n12239 , n4178 , n3260 );
or ( n12240 , n12238 , n12239 );
and ( n12241 , n12240 , n2422 );
and ( n12242 , n4178 , n2428 );
or ( n12243 , n12241 , n12242 );
buf ( n12244 , n12243 );
buf ( n12245 , n2424 );
buf ( n12246 , n2281 );
buf ( n12247 , n2280 );
not ( n12248 , n3260 );
and ( n12249 , n4168 , n3631 );
and ( n12250 , n7710 , n5281 );
and ( n12251 , n4168 , n11910 );
or ( n12252 , n12250 , n12251 );
and ( n12253 , n12252 , n5286 );
and ( n12254 , n7721 , n5281 );
and ( n12255 , n4168 , n11910 );
or ( n12256 , n12254 , n12255 );
and ( n12257 , n12256 , n6219 );
and ( n12258 , n7732 , n5281 );
and ( n12259 , n4168 , n11910 );
or ( n12260 , n12258 , n12259 );
and ( n12261 , n12260 , n6711 );
and ( n12262 , n5668 , n5281 );
and ( n12263 , n4168 , n11910 );
or ( n12264 , n12262 , n12263 );
and ( n12265 , n12264 , n6718 );
and ( n12266 , n4166 , n6720 );
and ( n12267 , n7744 , n5281 );
and ( n12268 , n4168 , n11910 );
or ( n12269 , n12267 , n12268 );
and ( n12270 , n12269 , n6725 );
or ( n12271 , n12249 , n12253 , n12257 , n12261 , n12265 , n12266 , n12270 );
and ( n12272 , n12248 , n12271 );
and ( n12273 , n4168 , n3260 );
or ( n12274 , n12272 , n12273 );
and ( n12275 , n12274 , n2422 );
and ( n12276 , n4168 , n2428 );
or ( n12277 , n12275 , n12276 );
buf ( n12278 , n12277 );
buf ( n12279 , n2424 );
buf ( n12280 , n2281 );
buf ( n12281 , n2280 );
not ( n12282 , n3260 );
and ( n12283 , n4158 , n3631 );
and ( n12284 , n7784 , n5281 );
and ( n12285 , n4158 , n11910 );
or ( n12286 , n12284 , n12285 );
and ( n12287 , n12286 , n5286 );
and ( n12288 , n7795 , n5281 );
and ( n12289 , n4158 , n11910 );
or ( n12290 , n12288 , n12289 );
and ( n12291 , n12290 , n6219 );
and ( n12292 , n7806 , n5281 );
and ( n12293 , n4158 , n11910 );
or ( n12294 , n12292 , n12293 );
and ( n12295 , n12294 , n6711 );
and ( n12296 , n5658 , n5281 );
and ( n12297 , n4158 , n11910 );
or ( n12298 , n12296 , n12297 );
and ( n12299 , n12298 , n6718 );
and ( n12300 , n4156 , n6720 );
and ( n12301 , n7818 , n5281 );
and ( n12302 , n4158 , n11910 );
or ( n12303 , n12301 , n12302 );
and ( n12304 , n12303 , n6725 );
or ( n12305 , n12283 , n12287 , n12291 , n12295 , n12299 , n12300 , n12304 );
and ( n12306 , n12282 , n12305 );
and ( n12307 , n4158 , n3260 );
or ( n12308 , n12306 , n12307 );
and ( n12309 , n12308 , n2422 );
and ( n12310 , n4158 , n2428 );
or ( n12311 , n12309 , n12310 );
buf ( n12312 , n12311 );
buf ( n12313 , n2424 );
buf ( n12314 , n2281 );
buf ( n12315 , n2280 );
not ( n12316 , n3260 );
and ( n12317 , n4148 , n3631 );
and ( n12318 , n7858 , n5281 );
and ( n12319 , n4148 , n11910 );
or ( n12320 , n12318 , n12319 );
and ( n12321 , n12320 , n5286 );
and ( n12322 , n7869 , n5281 );
and ( n12323 , n4148 , n11910 );
or ( n12324 , n12322 , n12323 );
and ( n12325 , n12324 , n6219 );
and ( n12326 , n7880 , n5281 );
and ( n12327 , n4148 , n11910 );
or ( n12328 , n12326 , n12327 );
and ( n12329 , n12328 , n6711 );
and ( n12330 , n5648 , n5281 );
and ( n12331 , n4148 , n11910 );
or ( n12332 , n12330 , n12331 );
and ( n12333 , n12332 , n6718 );
and ( n12334 , n4146 , n6720 );
and ( n12335 , n7892 , n5281 );
and ( n12336 , n4148 , n11910 );
or ( n12337 , n12335 , n12336 );
and ( n12338 , n12337 , n6725 );
or ( n12339 , n12317 , n12321 , n12325 , n12329 , n12333 , n12334 , n12338 );
and ( n12340 , n12316 , n12339 );
and ( n12341 , n4148 , n3260 );
or ( n12342 , n12340 , n12341 );
and ( n12343 , n12342 , n2422 );
and ( n12344 , n4148 , n2428 );
or ( n12345 , n12343 , n12344 );
buf ( n12346 , n12345 );
buf ( n12347 , n2424 );
buf ( n12348 , n2281 );
buf ( n12349 , n2280 );
not ( n12350 , n3260 );
and ( n12351 , n4138 , n3631 );
and ( n12352 , n7932 , n5281 );
and ( n12353 , n4138 , n11910 );
or ( n12354 , n12352 , n12353 );
and ( n12355 , n12354 , n5286 );
and ( n12356 , n7943 , n5281 );
and ( n12357 , n4138 , n11910 );
or ( n12358 , n12356 , n12357 );
and ( n12359 , n12358 , n6219 );
and ( n12360 , n7954 , n5281 );
and ( n12361 , n4138 , n11910 );
or ( n12362 , n12360 , n12361 );
and ( n12363 , n12362 , n6711 );
and ( n12364 , n5638 , n5281 );
and ( n12365 , n4138 , n11910 );
or ( n12366 , n12364 , n12365 );
and ( n12367 , n12366 , n6718 );
and ( n12368 , n4136 , n6720 );
and ( n12369 , n7966 , n5281 );
and ( n12370 , n4138 , n11910 );
or ( n12371 , n12369 , n12370 );
and ( n12372 , n12371 , n6725 );
or ( n12373 , n12351 , n12355 , n12359 , n12363 , n12367 , n12368 , n12372 );
and ( n12374 , n12350 , n12373 );
and ( n12375 , n4138 , n3260 );
or ( n12376 , n12374 , n12375 );
and ( n12377 , n12376 , n2422 );
and ( n12378 , n4138 , n2428 );
or ( n12379 , n12377 , n12378 );
buf ( n12380 , n12379 );
buf ( n12381 , n2424 );
buf ( n12382 , n2281 );
buf ( n12383 , n2280 );
not ( n12384 , n3260 );
and ( n12385 , n4128 , n3631 );
and ( n12386 , n8006 , n5281 );
and ( n12387 , n4128 , n11910 );
or ( n12388 , n12386 , n12387 );
and ( n12389 , n12388 , n5286 );
and ( n12390 , n8017 , n5281 );
and ( n12391 , n4128 , n11910 );
or ( n12392 , n12390 , n12391 );
and ( n12393 , n12392 , n6219 );
and ( n12394 , n8028 , n5281 );
and ( n12395 , n4128 , n11910 );
or ( n12396 , n12394 , n12395 );
and ( n12397 , n12396 , n6711 );
and ( n12398 , n5628 , n5281 );
and ( n12399 , n4128 , n11910 );
or ( n12400 , n12398 , n12399 );
and ( n12401 , n12400 , n6718 );
and ( n12402 , n4126 , n6720 );
and ( n12403 , n8040 , n5281 );
and ( n12404 , n4128 , n11910 );
or ( n12405 , n12403 , n12404 );
and ( n12406 , n12405 , n6725 );
or ( n12407 , n12385 , n12389 , n12393 , n12397 , n12401 , n12402 , n12406 );
and ( n12408 , n12384 , n12407 );
and ( n12409 , n4128 , n3260 );
or ( n12410 , n12408 , n12409 );
and ( n12411 , n12410 , n2422 );
and ( n12412 , n4128 , n2428 );
or ( n12413 , n12411 , n12412 );
buf ( n12414 , n12413 );
buf ( n12415 , n2424 );
buf ( n12416 , n2281 );
buf ( n12417 , n2280 );
not ( n12418 , n3260 );
and ( n12419 , n4118 , n3631 );
and ( n12420 , n8080 , n5281 );
and ( n12421 , n4118 , n11910 );
or ( n12422 , n12420 , n12421 );
and ( n12423 , n12422 , n5286 );
and ( n12424 , n8091 , n5281 );
and ( n12425 , n4118 , n11910 );
or ( n12426 , n12424 , n12425 );
and ( n12427 , n12426 , n6219 );
and ( n12428 , n8102 , n5281 );
and ( n12429 , n4118 , n11910 );
or ( n12430 , n12428 , n12429 );
and ( n12431 , n12430 , n6711 );
and ( n12432 , n5618 , n5281 );
and ( n12433 , n4118 , n11910 );
or ( n12434 , n12432 , n12433 );
and ( n12435 , n12434 , n6718 );
and ( n12436 , n4116 , n6720 );
and ( n12437 , n8114 , n5281 );
and ( n12438 , n4118 , n11910 );
or ( n12439 , n12437 , n12438 );
and ( n12440 , n12439 , n6725 );
or ( n12441 , n12419 , n12423 , n12427 , n12431 , n12435 , n12436 , n12440 );
and ( n12442 , n12418 , n12441 );
and ( n12443 , n4118 , n3260 );
or ( n12444 , n12442 , n12443 );
and ( n12445 , n12444 , n2422 );
and ( n12446 , n4118 , n2428 );
or ( n12447 , n12445 , n12446 );
buf ( n12448 , n12447 );
buf ( n12449 , n2424 );
buf ( n12450 , n2281 );
buf ( n12451 , n2280 );
not ( n12452 , n3260 );
and ( n12453 , n4108 , n3631 );
and ( n12454 , n8154 , n5281 );
and ( n12455 , n4108 , n11910 );
or ( n12456 , n12454 , n12455 );
and ( n12457 , n12456 , n5286 );
and ( n12458 , n8165 , n5281 );
and ( n12459 , n4108 , n11910 );
or ( n12460 , n12458 , n12459 );
and ( n12461 , n12460 , n6219 );
and ( n12462 , n8176 , n5281 );
and ( n12463 , n4108 , n11910 );
or ( n12464 , n12462 , n12463 );
and ( n12465 , n12464 , n6711 );
and ( n12466 , n5608 , n5281 );
and ( n12467 , n4108 , n11910 );
or ( n12468 , n12466 , n12467 );
and ( n12469 , n12468 , n6718 );
and ( n12470 , n4106 , n6720 );
and ( n12471 , n8188 , n5281 );
and ( n12472 , n4108 , n11910 );
or ( n12473 , n12471 , n12472 );
and ( n12474 , n12473 , n6725 );
or ( n12475 , n12453 , n12457 , n12461 , n12465 , n12469 , n12470 , n12474 );
and ( n12476 , n12452 , n12475 );
and ( n12477 , n4108 , n3260 );
or ( n12478 , n12476 , n12477 );
and ( n12479 , n12478 , n2422 );
and ( n12480 , n4108 , n2428 );
or ( n12481 , n12479 , n12480 );
buf ( n12482 , n12481 );
buf ( n12483 , n2424 );
buf ( n12484 , n2281 );
buf ( n12485 , n2280 );
not ( n12486 , n3260 );
and ( n12487 , n4098 , n3631 );
and ( n12488 , n8228 , n5281 );
and ( n12489 , n4098 , n11910 );
or ( n12490 , n12488 , n12489 );
and ( n12491 , n12490 , n5286 );
and ( n12492 , n8239 , n5281 );
and ( n12493 , n4098 , n11910 );
or ( n12494 , n12492 , n12493 );
and ( n12495 , n12494 , n6219 );
and ( n12496 , n8250 , n5281 );
and ( n12497 , n4098 , n11910 );
or ( n12498 , n12496 , n12497 );
and ( n12499 , n12498 , n6711 );
and ( n12500 , n5598 , n5281 );
and ( n12501 , n4098 , n11910 );
or ( n12502 , n12500 , n12501 );
and ( n12503 , n12502 , n6718 );
and ( n12504 , n4096 , n6720 );
and ( n12505 , n8262 , n5281 );
and ( n12506 , n4098 , n11910 );
or ( n12507 , n12505 , n12506 );
and ( n12508 , n12507 , n6725 );
or ( n12509 , n12487 , n12491 , n12495 , n12499 , n12503 , n12504 , n12508 );
and ( n12510 , n12486 , n12509 );
and ( n12511 , n4098 , n3260 );
or ( n12512 , n12510 , n12511 );
and ( n12513 , n12512 , n2422 );
and ( n12514 , n4098 , n2428 );
or ( n12515 , n12513 , n12514 );
buf ( n12516 , n12515 );
buf ( n12517 , n2424 );
buf ( n12518 , n2281 );
buf ( n12519 , n2280 );
not ( n12520 , n3260 );
and ( n12521 , n4088 , n3631 );
and ( n12522 , n8302 , n5281 );
and ( n12523 , n4088 , n11910 );
or ( n12524 , n12522 , n12523 );
and ( n12525 , n12524 , n5286 );
and ( n12526 , n8313 , n5281 );
and ( n12527 , n4088 , n11910 );
or ( n12528 , n12526 , n12527 );
and ( n12529 , n12528 , n6219 );
and ( n12530 , n8324 , n5281 );
and ( n12531 , n4088 , n11910 );
or ( n12532 , n12530 , n12531 );
and ( n12533 , n12532 , n6711 );
and ( n12534 , n5588 , n5281 );
and ( n12535 , n4088 , n11910 );
or ( n12536 , n12534 , n12535 );
and ( n12537 , n12536 , n6718 );
and ( n12538 , n4086 , n6720 );
and ( n12539 , n8336 , n5281 );
and ( n12540 , n4088 , n11910 );
or ( n12541 , n12539 , n12540 );
and ( n12542 , n12541 , n6725 );
or ( n12543 , n12521 , n12525 , n12529 , n12533 , n12537 , n12538 , n12542 );
and ( n12544 , n12520 , n12543 );
and ( n12545 , n4088 , n3260 );
or ( n12546 , n12544 , n12545 );
and ( n12547 , n12546 , n2422 );
and ( n12548 , n4088 , n2428 );
or ( n12549 , n12547 , n12548 );
buf ( n12550 , n12549 );
buf ( n12551 , n2424 );
buf ( n12552 , n2281 );
buf ( n12553 , n2280 );
not ( n12554 , n3260 );
and ( n12555 , n4078 , n3631 );
and ( n12556 , n8376 , n5281 );
and ( n12557 , n4078 , n11910 );
or ( n12558 , n12556 , n12557 );
and ( n12559 , n12558 , n5286 );
and ( n12560 , n8387 , n5281 );
and ( n12561 , n4078 , n11910 );
or ( n12562 , n12560 , n12561 );
and ( n12563 , n12562 , n6219 );
and ( n12564 , n8398 , n5281 );
and ( n12565 , n4078 , n11910 );
or ( n12566 , n12564 , n12565 );
and ( n12567 , n12566 , n6711 );
and ( n12568 , n5578 , n5281 );
and ( n12569 , n4078 , n11910 );
or ( n12570 , n12568 , n12569 );
and ( n12571 , n12570 , n6718 );
and ( n12572 , n4076 , n6720 );
and ( n12573 , n8410 , n5281 );
and ( n12574 , n4078 , n11910 );
or ( n12575 , n12573 , n12574 );
and ( n12576 , n12575 , n6725 );
or ( n12577 , n12555 , n12559 , n12563 , n12567 , n12571 , n12572 , n12576 );
and ( n12578 , n12554 , n12577 );
and ( n12579 , n4078 , n3260 );
or ( n12580 , n12578 , n12579 );
and ( n12581 , n12580 , n2422 );
and ( n12582 , n4078 , n2428 );
or ( n12583 , n12581 , n12582 );
buf ( n12584 , n12583 );
buf ( n12585 , n2424 );
buf ( n12586 , n2281 );
buf ( n12587 , n2280 );
not ( n12588 , n3260 );
and ( n12589 , n4068 , n3631 );
and ( n12590 , n8450 , n5281 );
and ( n12591 , n4068 , n11910 );
or ( n12592 , n12590 , n12591 );
and ( n12593 , n12592 , n5286 );
and ( n12594 , n8461 , n5281 );
and ( n12595 , n4068 , n11910 );
or ( n12596 , n12594 , n12595 );
and ( n12597 , n12596 , n6219 );
and ( n12598 , n8472 , n5281 );
and ( n12599 , n4068 , n11910 );
or ( n12600 , n12598 , n12599 );
and ( n12601 , n12600 , n6711 );
and ( n12602 , n5530 , n5281 );
and ( n12603 , n4068 , n11910 );
or ( n12604 , n12602 , n12603 );
and ( n12605 , n12604 , n6718 );
and ( n12606 , n4066 , n6720 );
and ( n12607 , n8484 , n5281 );
and ( n12608 , n4068 , n11910 );
or ( n12609 , n12607 , n12608 );
and ( n12610 , n12609 , n6725 );
or ( n12611 , n12589 , n12593 , n12597 , n12601 , n12605 , n12606 , n12610 );
and ( n12612 , n12588 , n12611 );
and ( n12613 , n4068 , n3260 );
or ( n12614 , n12612 , n12613 );
and ( n12615 , n12614 , n2422 );
and ( n12616 , n4068 , n2428 );
or ( n12617 , n12615 , n12616 );
buf ( n12618 , n12617 );
buf ( n12619 , n2424 );
buf ( n12620 , n2281 );
buf ( n12621 , n2280 );
not ( n12622 , n3260 );
and ( n12623 , n4058 , n3631 );
and ( n12624 , n8524 , n5281 );
and ( n12625 , n4058 , n11910 );
or ( n12626 , n12624 , n12625 );
and ( n12627 , n12626 , n5286 );
and ( n12628 , n8535 , n5281 );
and ( n12629 , n4058 , n11910 );
or ( n12630 , n12628 , n12629 );
and ( n12631 , n12630 , n6219 );
and ( n12632 , n8546 , n5281 );
and ( n12633 , n4058 , n11910 );
or ( n12634 , n12632 , n12633 );
and ( n12635 , n12634 , n6711 );
and ( n12636 , n5527 , n5281 );
and ( n12637 , n4058 , n11910 );
or ( n12638 , n12636 , n12637 );
and ( n12639 , n12638 , n6718 );
and ( n12640 , n4056 , n6720 );
and ( n12641 , n8558 , n5281 );
and ( n12642 , n4058 , n11910 );
or ( n12643 , n12641 , n12642 );
and ( n12644 , n12643 , n6725 );
or ( n12645 , n12623 , n12627 , n12631 , n12635 , n12639 , n12640 , n12644 );
and ( n12646 , n12622 , n12645 );
and ( n12647 , n4058 , n3260 );
or ( n12648 , n12646 , n12647 );
and ( n12649 , n12648 , n2422 );
and ( n12650 , n4058 , n2428 );
or ( n12651 , n12649 , n12650 );
buf ( n12652 , n12651 );
buf ( n12653 , n2424 );
buf ( n12654 , n2281 );
buf ( n12655 , n2280 );
not ( n12656 , n3260 );
and ( n12657 , n4048 , n3631 );
and ( n12658 , n8598 , n5281 );
and ( n12659 , n4048 , n11910 );
or ( n12660 , n12658 , n12659 );
and ( n12661 , n12660 , n5286 );
and ( n12662 , n8609 , n5281 );
and ( n12663 , n4048 , n11910 );
or ( n12664 , n12662 , n12663 );
and ( n12665 , n12664 , n6219 );
and ( n12666 , n8620 , n5281 );
and ( n12667 , n4048 , n11910 );
or ( n12668 , n12666 , n12667 );
and ( n12669 , n12668 , n6711 );
and ( n12670 , n5524 , n5281 );
and ( n12671 , n4048 , n11910 );
or ( n12672 , n12670 , n12671 );
and ( n12673 , n12672 , n6718 );
and ( n12674 , n4046 , n6720 );
and ( n12675 , n8632 , n5281 );
and ( n12676 , n4048 , n11910 );
or ( n12677 , n12675 , n12676 );
and ( n12678 , n12677 , n6725 );
or ( n12679 , n12657 , n12661 , n12665 , n12669 , n12673 , n12674 , n12678 );
and ( n12680 , n12656 , n12679 );
and ( n12681 , n4048 , n3260 );
or ( n12682 , n12680 , n12681 );
and ( n12683 , n12682 , n2422 );
and ( n12684 , n4048 , n2428 );
or ( n12685 , n12683 , n12684 );
buf ( n12686 , n12685 );
buf ( n12687 , n2424 );
buf ( n12688 , n2281 );
buf ( n12689 , n2280 );
not ( n12690 , n3260 );
and ( n12691 , n4038 , n3631 );
and ( n12692 , n8672 , n5281 );
and ( n12693 , n4038 , n11910 );
or ( n12694 , n12692 , n12693 );
and ( n12695 , n12694 , n5286 );
and ( n12696 , n8683 , n5281 );
and ( n12697 , n4038 , n11910 );
or ( n12698 , n12696 , n12697 );
and ( n12699 , n12698 , n6219 );
and ( n12700 , n8694 , n5281 );
and ( n12701 , n4038 , n11910 );
or ( n12702 , n12700 , n12701 );
and ( n12703 , n12702 , n6711 );
and ( n12704 , n5521 , n5281 );
and ( n12705 , n4038 , n11910 );
or ( n12706 , n12704 , n12705 );
and ( n12707 , n12706 , n6718 );
and ( n12708 , n4036 , n6720 );
and ( n12709 , n8706 , n5281 );
and ( n12710 , n4038 , n11910 );
or ( n12711 , n12709 , n12710 );
and ( n12712 , n12711 , n6725 );
or ( n12713 , n12691 , n12695 , n12699 , n12703 , n12707 , n12708 , n12712 );
and ( n12714 , n12690 , n12713 );
and ( n12715 , n4038 , n3260 );
or ( n12716 , n12714 , n12715 );
and ( n12717 , n12716 , n2422 );
and ( n12718 , n4038 , n2428 );
or ( n12719 , n12717 , n12718 );
buf ( n12720 , n12719 );
buf ( n12721 , n2424 );
buf ( n12722 , n2281 );
buf ( n12723 , n2280 );
not ( n12724 , n3260 );
and ( n12725 , n4028 , n3631 );
and ( n12726 , n8746 , n5281 );
and ( n12727 , n4028 , n11910 );
or ( n12728 , n12726 , n12727 );
and ( n12729 , n12728 , n5286 );
and ( n12730 , n8757 , n5281 );
and ( n12731 , n4028 , n11910 );
or ( n12732 , n12730 , n12731 );
and ( n12733 , n12732 , n6219 );
and ( n12734 , n8768 , n5281 );
and ( n12735 , n4028 , n11910 );
or ( n12736 , n12734 , n12735 );
and ( n12737 , n12736 , n6711 );
and ( n12738 , n5518 , n5281 );
and ( n12739 , n4028 , n11910 );
or ( n12740 , n12738 , n12739 );
and ( n12741 , n12740 , n6718 );
and ( n12742 , n4026 , n6720 );
and ( n12743 , n8780 , n5281 );
and ( n12744 , n4028 , n11910 );
or ( n12745 , n12743 , n12744 );
and ( n12746 , n12745 , n6725 );
or ( n12747 , n12725 , n12729 , n12733 , n12737 , n12741 , n12742 , n12746 );
and ( n12748 , n12724 , n12747 );
and ( n12749 , n4028 , n3260 );
or ( n12750 , n12748 , n12749 );
and ( n12751 , n12750 , n2422 );
and ( n12752 , n4028 , n2428 );
or ( n12753 , n12751 , n12752 );
buf ( n12754 , n12753 );
buf ( n12755 , n2424 );
buf ( n12756 , n2281 );
buf ( n12757 , n2280 );
not ( n12758 , n3260 );
and ( n12759 , n4018 , n3631 );
and ( n12760 , n8820 , n5281 );
and ( n12761 , n4018 , n11910 );
or ( n12762 , n12760 , n12761 );
and ( n12763 , n12762 , n5286 );
and ( n12764 , n8831 , n5281 );
and ( n12765 , n4018 , n11910 );
or ( n12766 , n12764 , n12765 );
and ( n12767 , n12766 , n6219 );
and ( n12768 , n8842 , n5281 );
and ( n12769 , n4018 , n11910 );
or ( n12770 , n12768 , n12769 );
and ( n12771 , n12770 , n6711 );
and ( n12772 , n5515 , n5281 );
and ( n12773 , n4018 , n11910 );
or ( n12774 , n12772 , n12773 );
and ( n12775 , n12774 , n6718 );
and ( n12776 , n4016 , n6720 );
and ( n12777 , n8854 , n5281 );
and ( n12778 , n4018 , n11910 );
or ( n12779 , n12777 , n12778 );
and ( n12780 , n12779 , n6725 );
or ( n12781 , n12759 , n12763 , n12767 , n12771 , n12775 , n12776 , n12780 );
and ( n12782 , n12758 , n12781 );
and ( n12783 , n4018 , n3260 );
or ( n12784 , n12782 , n12783 );
and ( n12785 , n12784 , n2422 );
and ( n12786 , n4018 , n2428 );
or ( n12787 , n12785 , n12786 );
buf ( n12788 , n12787 );
buf ( n12789 , n2424 );
buf ( n12790 , n2281 );
buf ( n12791 , n2280 );
not ( n12792 , n3260 );
and ( n12793 , n4008 , n3631 );
and ( n12794 , n8894 , n5281 );
and ( n12795 , n4008 , n11910 );
or ( n12796 , n12794 , n12795 );
and ( n12797 , n12796 , n5286 );
and ( n12798 , n8905 , n5281 );
and ( n12799 , n4008 , n11910 );
or ( n12800 , n12798 , n12799 );
and ( n12801 , n12800 , n6219 );
and ( n12802 , n8916 , n5281 );
and ( n12803 , n4008 , n11910 );
or ( n12804 , n12802 , n12803 );
and ( n12805 , n12804 , n6711 );
and ( n12806 , n5512 , n5281 );
and ( n12807 , n4008 , n11910 );
or ( n12808 , n12806 , n12807 );
and ( n12809 , n12808 , n6718 );
and ( n12810 , n4006 , n6720 );
and ( n12811 , n8928 , n5281 );
and ( n12812 , n4008 , n11910 );
or ( n12813 , n12811 , n12812 );
and ( n12814 , n12813 , n6725 );
or ( n12815 , n12793 , n12797 , n12801 , n12805 , n12809 , n12810 , n12814 );
and ( n12816 , n12792 , n12815 );
and ( n12817 , n4008 , n3260 );
or ( n12818 , n12816 , n12817 );
and ( n12819 , n12818 , n2422 );
and ( n12820 , n4008 , n2428 );
or ( n12821 , n12819 , n12820 );
buf ( n12822 , n12821 );
buf ( n12823 , n2424 );
buf ( n12824 , n2281 );
buf ( n12825 , n2280 );
not ( n12826 , n3260 );
and ( n12827 , n3998 , n3631 );
and ( n12828 , n8968 , n5281 );
and ( n12829 , n3998 , n11910 );
or ( n12830 , n12828 , n12829 );
and ( n12831 , n12830 , n5286 );
and ( n12832 , n8979 , n5281 );
and ( n12833 , n3998 , n11910 );
or ( n12834 , n12832 , n12833 );
and ( n12835 , n12834 , n6219 );
and ( n12836 , n8990 , n5281 );
and ( n12837 , n3998 , n11910 );
or ( n12838 , n12836 , n12837 );
and ( n12839 , n12838 , n6711 );
and ( n12840 , n5509 , n5281 );
and ( n12841 , n3998 , n11910 );
or ( n12842 , n12840 , n12841 );
and ( n12843 , n12842 , n6718 );
and ( n12844 , n3996 , n6720 );
and ( n12845 , n9002 , n5281 );
and ( n12846 , n3998 , n11910 );
or ( n12847 , n12845 , n12846 );
and ( n12848 , n12847 , n6725 );
or ( n12849 , n12827 , n12831 , n12835 , n12839 , n12843 , n12844 , n12848 );
and ( n12850 , n12826 , n12849 );
and ( n12851 , n3998 , n3260 );
or ( n12852 , n12850 , n12851 );
and ( n12853 , n12852 , n2422 );
and ( n12854 , n3998 , n2428 );
or ( n12855 , n12853 , n12854 );
buf ( n12856 , n12855 );
buf ( n12857 , n2424 );
buf ( n12858 , n2281 );
buf ( n12859 , n2280 );
not ( n12860 , n3260 );
and ( n12861 , n3988 , n3631 );
and ( n12862 , n9042 , n5281 );
and ( n12863 , n3988 , n11910 );
or ( n12864 , n12862 , n12863 );
and ( n12865 , n12864 , n5286 );
and ( n12866 , n9053 , n5281 );
and ( n12867 , n3988 , n11910 );
or ( n12868 , n12866 , n12867 );
and ( n12869 , n12868 , n6219 );
and ( n12870 , n9064 , n5281 );
and ( n12871 , n3988 , n11910 );
or ( n12872 , n12870 , n12871 );
and ( n12873 , n12872 , n6711 );
and ( n12874 , n5506 , n5281 );
and ( n12875 , n3988 , n11910 );
or ( n12876 , n12874 , n12875 );
and ( n12877 , n12876 , n6718 );
and ( n12878 , n3986 , n6720 );
and ( n12879 , n9076 , n5281 );
and ( n12880 , n3988 , n11910 );
or ( n12881 , n12879 , n12880 );
and ( n12882 , n12881 , n6725 );
or ( n12883 , n12861 , n12865 , n12869 , n12873 , n12877 , n12878 , n12882 );
and ( n12884 , n12860 , n12883 );
and ( n12885 , n3988 , n3260 );
or ( n12886 , n12884 , n12885 );
and ( n12887 , n12886 , n2422 );
and ( n12888 , n3988 , n2428 );
or ( n12889 , n12887 , n12888 );
buf ( n12890 , n12889 );
buf ( n12891 , n2424 );
buf ( n12892 , n2281 );
buf ( n12893 , n2280 );
not ( n12894 , n3260 );
and ( n12895 , n3978 , n3631 );
and ( n12896 , n10079 , n5281 );
and ( n12897 , n3978 , n11910 );
or ( n12898 , n12896 , n12897 );
and ( n12899 , n12898 , n5286 );
and ( n12900 , n10090 , n5281 );
and ( n12901 , n3978 , n11910 );
or ( n12902 , n12900 , n12901 );
and ( n12903 , n12902 , n6219 );
and ( n12904 , n10101 , n5281 );
and ( n12905 , n3978 , n11910 );
or ( n12906 , n12904 , n12905 );
and ( n12907 , n12906 , n6711 );
and ( n12908 , n5503 , n5281 );
and ( n12909 , n3978 , n11910 );
or ( n12910 , n12908 , n12909 );
and ( n12911 , n12910 , n6718 );
and ( n12912 , n3976 , n6720 );
and ( n12913 , n10112 , n5281 );
and ( n12914 , n3978 , n11910 );
or ( n12915 , n12913 , n12914 );
and ( n12916 , n12915 , n6725 );
or ( n12917 , n12895 , n12899 , n12903 , n12907 , n12911 , n12912 , n12916 );
and ( n12918 , n12894 , n12917 );
and ( n12919 , n3978 , n3260 );
or ( n12920 , n12918 , n12919 );
and ( n12921 , n12920 , n2422 );
and ( n12922 , n3978 , n2428 );
or ( n12923 , n12921 , n12922 );
buf ( n12924 , n12923 );
buf ( n12925 , n2424 );
buf ( n12926 , n2281 );
buf ( n12927 , n2280 );
not ( n12928 , n3260 );
and ( n12929 , n3813 , n3631 );
and ( n12930 , n10148 , n5281 );
and ( n12931 , n3813 , n11910 );
or ( n12932 , n12930 , n12931 );
and ( n12933 , n12932 , n5286 );
and ( n12934 , n10157 , n5281 );
and ( n12935 , n3813 , n11910 );
or ( n12936 , n12934 , n12935 );
and ( n12937 , n12936 , n6219 );
and ( n12938 , n10166 , n5281 );
and ( n12939 , n3813 , n11910 );
or ( n12940 , n12938 , n12939 );
and ( n12941 , n12940 , n6711 );
and ( n12942 , n5500 , n5281 );
and ( n12943 , n3813 , n11910 );
or ( n12944 , n12942 , n12943 );
and ( n12945 , n12944 , n6718 );
and ( n12946 , n10177 , n5281 );
and ( n12947 , n3813 , n11910 );
or ( n12948 , n12946 , n12947 );
and ( n12949 , n12948 , n6725 );
or ( n12950 , n12929 , n12933 , n12937 , n12941 , n12945 , n2424 , n12949 );
and ( n12951 , n12928 , n12950 );
and ( n12952 , n3813 , n3260 );
or ( n12953 , n12951 , n12952 );
and ( n12954 , n12953 , n2422 );
and ( n12955 , n3813 , n2428 );
or ( n12956 , n12954 , n12955 );
buf ( n12957 , n12956 );
buf ( n12958 , n2424 );
buf ( n12959 , n2281 );
buf ( n12960 , n2280 );
not ( n12961 , n3260 );
and ( n12962 , n3635 , n3631 );
and ( n12963 , n10202 , n5281 );
and ( n12964 , n3635 , n11910 );
or ( n12965 , n12963 , n12964 );
and ( n12966 , n12965 , n5286 );
and ( n12967 , n3635 , n11910 );
and ( n12968 , n12967 , n6219 );
and ( n12969 , n3635 , n11910 );
and ( n12970 , n12969 , n6711 );
and ( n12971 , n5497 , n5281 );
and ( n12972 , n3635 , n11910 );
or ( n12973 , n12971 , n12972 );
and ( n12974 , n12973 , n6718 );
and ( n12975 , n10217 , n5281 );
and ( n12976 , n3635 , n11910 );
or ( n12977 , n12975 , n12976 );
and ( n12978 , n12977 , n6725 );
or ( n12979 , n12962 , n12966 , n12968 , n12970 , n12974 , n2424 , n12978 );
and ( n12980 , n12961 , n12979 );
and ( n12981 , n3635 , n3260 );
or ( n12982 , n12980 , n12981 );
and ( n12983 , n12982 , n2422 );
and ( n12984 , n3635 , n2428 );
or ( n12985 , n12983 , n12984 );
buf ( n12986 , n12985 );
buf ( n12987 , n2424 );
buf ( n12988 , n2281 );
buf ( n12989 , n2280 );
not ( n12990 , n3066 );
not ( n12991 , n3259 );
or ( n12992 , n5286 , n3631 );
and ( n12993 , n2352 , n12992 );
xor ( n12994 , n5491 , n3789 );
not ( n12995 , n12994 );
not ( n12996 , n12995 );
and ( n12997 , n5576 , n4078 );
and ( n12998 , n5586 , n4088 );
and ( n12999 , n5596 , n4098 );
and ( n13000 , n5606 , n4108 );
and ( n13001 , n5616 , n4118 );
and ( n13002 , n5626 , n4128 );
and ( n13003 , n5636 , n4138 );
and ( n13004 , n5646 , n4148 );
and ( n13005 , n5656 , n4158 );
and ( n13006 , n5666 , n4168 );
and ( n13007 , n5676 , n4178 );
and ( n13008 , n5686 , n4188 );
and ( n13009 , n5696 , n4198 );
and ( n13010 , n5706 , n4208 );
and ( n13011 , n5716 , n4218 );
and ( n13012 , n5726 , n4228 );
and ( n13013 , n5736 , n4238 );
and ( n13014 , n5746 , n4252 );
and ( n13015 , n5756 , n3779 );
and ( n13016 , n5491 , n3789 );
and ( n13017 , n3779 , n13016 );
and ( n13018 , n5756 , n13016 );
or ( n13019 , n13015 , n13017 , n13018 );
and ( n13020 , n4252 , n13019 );
and ( n13021 , n5746 , n13019 );
or ( n13022 , n13014 , n13020 , n13021 );
and ( n13023 , n4238 , n13022 );
and ( n13024 , n5736 , n13022 );
or ( n13025 , n13013 , n13023 , n13024 );
and ( n13026 , n4228 , n13025 );
and ( n13027 , n5726 , n13025 );
or ( n13028 , n13012 , n13026 , n13027 );
and ( n13029 , n4218 , n13028 );
and ( n13030 , n5716 , n13028 );
or ( n13031 , n13011 , n13029 , n13030 );
and ( n13032 , n4208 , n13031 );
and ( n13033 , n5706 , n13031 );
or ( n13034 , n13010 , n13032 , n13033 );
and ( n13035 , n4198 , n13034 );
and ( n13036 , n5696 , n13034 );
or ( n13037 , n13009 , n13035 , n13036 );
and ( n13038 , n4188 , n13037 );
and ( n13039 , n5686 , n13037 );
or ( n13040 , n13008 , n13038 , n13039 );
and ( n13041 , n4178 , n13040 );
and ( n13042 , n5676 , n13040 );
or ( n13043 , n13007 , n13041 , n13042 );
and ( n13044 , n4168 , n13043 );
and ( n13045 , n5666 , n13043 );
or ( n13046 , n13006 , n13044 , n13045 );
and ( n13047 , n4158 , n13046 );
and ( n13048 , n5656 , n13046 );
or ( n13049 , n13005 , n13047 , n13048 );
and ( n13050 , n4148 , n13049 );
and ( n13051 , n5646 , n13049 );
or ( n13052 , n13004 , n13050 , n13051 );
and ( n13053 , n4138 , n13052 );
and ( n13054 , n5636 , n13052 );
or ( n13055 , n13003 , n13053 , n13054 );
and ( n13056 , n4128 , n13055 );
and ( n13057 , n5626 , n13055 );
or ( n13058 , n13002 , n13056 , n13057 );
and ( n13059 , n4118 , n13058 );
and ( n13060 , n5616 , n13058 );
or ( n13061 , n13001 , n13059 , n13060 );
and ( n13062 , n4108 , n13061 );
and ( n13063 , n5606 , n13061 );
or ( n13064 , n13000 , n13062 , n13063 );
and ( n13065 , n4098 , n13064 );
and ( n13066 , n5596 , n13064 );
or ( n13067 , n12999 , n13065 , n13066 );
and ( n13068 , n4088 , n13067 );
and ( n13069 , n5586 , n13067 );
or ( n13070 , n12998 , n13068 , n13069 );
and ( n13071 , n4078 , n13070 );
and ( n13072 , n5576 , n13070 );
or ( n13073 , n12997 , n13071 , n13072 );
and ( n13074 , n4068 , n13073 );
and ( n13075 , n4058 , n13074 );
and ( n13076 , n4048 , n13075 );
and ( n13077 , n4038 , n13076 );
and ( n13078 , n4028 , n13077 );
and ( n13079 , n4018 , n13078 );
and ( n13080 , n4008 , n13079 );
and ( n13081 , n3998 , n13080 );
and ( n13082 , n3988 , n13081 );
and ( n13083 , n3978 , n13082 );
and ( n13084 , n3813 , n13083 );
xor ( n13085 , n3635 , n13084 );
not ( n13086 , n13085 );
xor ( n13087 , n5756 , n3779 );
xor ( n13088 , n13087 , n13016 );
and ( n13089 , n13086 , n13088 );
not ( n13090 , n13088 );
not ( n13091 , n12994 );
xor ( n13092 , n13090 , n13091 );
and ( n13093 , n13092 , n13085 );
or ( n13094 , n13089 , n13093 );
not ( n13095 , n13094 );
not ( n13096 , n13095 );
or ( n13097 , n12996 , n13096 );
not ( n13098 , n13085 );
xor ( n13099 , n5746 , n4252 );
xor ( n13100 , n13099 , n13019 );
and ( n13101 , n13098 , n13100 );
not ( n13102 , n13100 );
and ( n13103 , n13090 , n13091 );
xor ( n13104 , n13102 , n13103 );
and ( n13105 , n13104 , n13085 );
or ( n13106 , n13101 , n13105 );
not ( n13107 , n13106 );
not ( n13108 , n13107 );
or ( n13109 , n13097 , n13108 );
not ( n13110 , n13085 );
xor ( n13111 , n5736 , n4238 );
xor ( n13112 , n13111 , n13022 );
and ( n13113 , n13110 , n13112 );
not ( n13114 , n13112 );
and ( n13115 , n13102 , n13103 );
xor ( n13116 , n13114 , n13115 );
and ( n13117 , n13116 , n13085 );
or ( n13118 , n13113 , n13117 );
not ( n13119 , n13118 );
not ( n13120 , n13119 );
or ( n13121 , n13109 , n13120 );
not ( n13122 , n13085 );
xor ( n13123 , n5726 , n4228 );
xor ( n13124 , n13123 , n13025 );
and ( n13125 , n13122 , n13124 );
not ( n13126 , n13124 );
and ( n13127 , n13114 , n13115 );
xor ( n13128 , n13126 , n13127 );
and ( n13129 , n13128 , n13085 );
or ( n13130 , n13125 , n13129 );
not ( n13131 , n13130 );
not ( n13132 , n13131 );
or ( n13133 , n13121 , n13132 );
not ( n13134 , n13085 );
xor ( n13135 , n5716 , n4218 );
xor ( n13136 , n13135 , n13028 );
and ( n13137 , n13134 , n13136 );
not ( n13138 , n13136 );
and ( n13139 , n13126 , n13127 );
xor ( n13140 , n13138 , n13139 );
and ( n13141 , n13140 , n13085 );
or ( n13142 , n13137 , n13141 );
not ( n13143 , n13142 );
not ( n13144 , n13143 );
or ( n13145 , n13133 , n13144 );
not ( n13146 , n13085 );
xor ( n13147 , n5706 , n4208 );
xor ( n13148 , n13147 , n13031 );
and ( n13149 , n13146 , n13148 );
not ( n13150 , n13148 );
and ( n13151 , n13138 , n13139 );
xor ( n13152 , n13150 , n13151 );
and ( n13153 , n13152 , n13085 );
or ( n13154 , n13149 , n13153 );
not ( n13155 , n13154 );
not ( n13156 , n13155 );
or ( n13157 , n13145 , n13156 );
not ( n13158 , n13085 );
xor ( n13159 , n5696 , n4198 );
xor ( n13160 , n13159 , n13034 );
and ( n13161 , n13158 , n13160 );
not ( n13162 , n13160 );
and ( n13163 , n13150 , n13151 );
xor ( n13164 , n13162 , n13163 );
and ( n13165 , n13164 , n13085 );
or ( n13166 , n13161 , n13165 );
not ( n13167 , n13166 );
not ( n13168 , n13167 );
or ( n13169 , n13157 , n13168 );
not ( n13170 , n13085 );
xor ( n13171 , n5686 , n4188 );
xor ( n13172 , n13171 , n13037 );
and ( n13173 , n13170 , n13172 );
not ( n13174 , n13172 );
and ( n13175 , n13162 , n13163 );
xor ( n13176 , n13174 , n13175 );
and ( n13177 , n13176 , n13085 );
or ( n13178 , n13173 , n13177 );
not ( n13179 , n13178 );
not ( n13180 , n13179 );
or ( n13181 , n13169 , n13180 );
not ( n13182 , n13085 );
xor ( n13183 , n5676 , n4178 );
xor ( n13184 , n13183 , n13040 );
and ( n13185 , n13182 , n13184 );
not ( n13186 , n13184 );
and ( n13187 , n13174 , n13175 );
xor ( n13188 , n13186 , n13187 );
and ( n13189 , n13188 , n13085 );
or ( n13190 , n13185 , n13189 );
not ( n13191 , n13190 );
not ( n13192 , n13191 );
or ( n13193 , n13181 , n13192 );
not ( n13194 , n13085 );
xor ( n13195 , n5666 , n4168 );
xor ( n13196 , n13195 , n13043 );
and ( n13197 , n13194 , n13196 );
not ( n13198 , n13196 );
and ( n13199 , n13186 , n13187 );
xor ( n13200 , n13198 , n13199 );
and ( n13201 , n13200 , n13085 );
or ( n13202 , n13197 , n13201 );
not ( n13203 , n13202 );
not ( n13204 , n13203 );
or ( n13205 , n13193 , n13204 );
not ( n13206 , n13085 );
xor ( n13207 , n5656 , n4158 );
xor ( n13208 , n13207 , n13046 );
and ( n13209 , n13206 , n13208 );
not ( n13210 , n13208 );
and ( n13211 , n13198 , n13199 );
xor ( n13212 , n13210 , n13211 );
and ( n13213 , n13212 , n13085 );
or ( n13214 , n13209 , n13213 );
not ( n13215 , n13214 );
not ( n13216 , n13215 );
or ( n13217 , n13205 , n13216 );
not ( n13218 , n13085 );
xor ( n13219 , n5646 , n4148 );
xor ( n13220 , n13219 , n13049 );
and ( n13221 , n13218 , n13220 );
not ( n13222 , n13220 );
and ( n13223 , n13210 , n13211 );
xor ( n13224 , n13222 , n13223 );
and ( n13225 , n13224 , n13085 );
or ( n13226 , n13221 , n13225 );
not ( n13227 , n13226 );
not ( n13228 , n13227 );
or ( n13229 , n13217 , n13228 );
not ( n13230 , n13085 );
xor ( n13231 , n5636 , n4138 );
xor ( n13232 , n13231 , n13052 );
and ( n13233 , n13230 , n13232 );
not ( n13234 , n13232 );
and ( n13235 , n13222 , n13223 );
xor ( n13236 , n13234 , n13235 );
and ( n13237 , n13236 , n13085 );
or ( n13238 , n13233 , n13237 );
not ( n13239 , n13238 );
not ( n13240 , n13239 );
or ( n13241 , n13229 , n13240 );
not ( n13242 , n13085 );
xor ( n13243 , n5626 , n4128 );
xor ( n13244 , n13243 , n13055 );
and ( n13245 , n13242 , n13244 );
not ( n13246 , n13244 );
and ( n13247 , n13234 , n13235 );
xor ( n13248 , n13246 , n13247 );
and ( n13249 , n13248 , n13085 );
or ( n13250 , n13245 , n13249 );
not ( n13251 , n13250 );
not ( n13252 , n13251 );
or ( n13253 , n13241 , n13252 );
not ( n13254 , n13085 );
xor ( n13255 , n5616 , n4118 );
xor ( n13256 , n13255 , n13058 );
and ( n13257 , n13254 , n13256 );
not ( n13258 , n13256 );
and ( n13259 , n13246 , n13247 );
xor ( n13260 , n13258 , n13259 );
and ( n13261 , n13260 , n13085 );
or ( n13262 , n13257 , n13261 );
not ( n13263 , n13262 );
not ( n13264 , n13263 );
or ( n13265 , n13253 , n13264 );
not ( n13266 , n13085 );
xor ( n13267 , n5606 , n4108 );
xor ( n13268 , n13267 , n13061 );
and ( n13269 , n13266 , n13268 );
not ( n13270 , n13268 );
and ( n13271 , n13258 , n13259 );
xor ( n13272 , n13270 , n13271 );
and ( n13273 , n13272 , n13085 );
or ( n13274 , n13269 , n13273 );
not ( n13275 , n13274 );
not ( n13276 , n13275 );
or ( n13277 , n13265 , n13276 );
not ( n13278 , n13085 );
xor ( n13279 , n5596 , n4098 );
xor ( n13280 , n13279 , n13064 );
and ( n13281 , n13278 , n13280 );
not ( n13282 , n13280 );
and ( n13283 , n13270 , n13271 );
xor ( n13284 , n13282 , n13283 );
and ( n13285 , n13284 , n13085 );
or ( n13286 , n13281 , n13285 );
not ( n13287 , n13286 );
not ( n13288 , n13287 );
or ( n13289 , n13277 , n13288 );
not ( n13290 , n13085 );
xor ( n13291 , n5586 , n4088 );
xor ( n13292 , n13291 , n13067 );
and ( n13293 , n13290 , n13292 );
not ( n13294 , n13292 );
and ( n13295 , n13282 , n13283 );
xor ( n13296 , n13294 , n13295 );
and ( n13297 , n13296 , n13085 );
or ( n13298 , n13293 , n13297 );
not ( n13299 , n13298 );
not ( n13300 , n13299 );
or ( n13301 , n13289 , n13300 );
not ( n13302 , n13085 );
xor ( n13303 , n5576 , n4078 );
xor ( n13304 , n13303 , n13070 );
and ( n13305 , n13302 , n13304 );
not ( n13306 , n13304 );
and ( n13307 , n13294 , n13295 );
xor ( n13308 , n13306 , n13307 );
and ( n13309 , n13308 , n13085 );
or ( n13310 , n13305 , n13309 );
not ( n13311 , n13310 );
not ( n13312 , n13311 );
or ( n13313 , n13301 , n13312 );
and ( n13314 , n13313 , n13085 );
not ( n13315 , n13314 );
and ( n13316 , n13315 , n12996 );
xor ( n13317 , n12996 , n13085 );
xor ( n13318 , n13317 , n13085 );
and ( n13319 , n13318 , n13314 );
or ( n13320 , n13316 , n13319 );
and ( n13321 , n13320 , n5290 );
xor ( n13322 , n5491 , n3791 );
not ( n13323 , n13322 );
not ( n13324 , n13323 );
and ( n13325 , n5576 , n4080 );
and ( n13326 , n5586 , n4090 );
and ( n13327 , n5596 , n4100 );
and ( n13328 , n5606 , n4110 );
and ( n13329 , n5616 , n4120 );
and ( n13330 , n5626 , n4130 );
and ( n13331 , n5636 , n4140 );
and ( n13332 , n5646 , n4150 );
and ( n13333 , n5656 , n4160 );
and ( n13334 , n5666 , n4170 );
and ( n13335 , n5676 , n4180 );
and ( n13336 , n5686 , n4190 );
and ( n13337 , n5696 , n4200 );
and ( n13338 , n5706 , n4210 );
and ( n13339 , n5716 , n4220 );
and ( n13340 , n5726 , n4230 );
and ( n13341 , n5736 , n4240 );
and ( n13342 , n5746 , n4254 );
and ( n13343 , n5756 , n3781 );
and ( n13344 , n5491 , n3791 );
and ( n13345 , n3781 , n13344 );
and ( n13346 , n5756 , n13344 );
or ( n13347 , n13343 , n13345 , n13346 );
and ( n13348 , n4254 , n13347 );
and ( n13349 , n5746 , n13347 );
or ( n13350 , n13342 , n13348 , n13349 );
and ( n13351 , n4240 , n13350 );
and ( n13352 , n5736 , n13350 );
or ( n13353 , n13341 , n13351 , n13352 );
and ( n13354 , n4230 , n13353 );
and ( n13355 , n5726 , n13353 );
or ( n13356 , n13340 , n13354 , n13355 );
and ( n13357 , n4220 , n13356 );
and ( n13358 , n5716 , n13356 );
or ( n13359 , n13339 , n13357 , n13358 );
and ( n13360 , n4210 , n13359 );
and ( n13361 , n5706 , n13359 );
or ( n13362 , n13338 , n13360 , n13361 );
and ( n13363 , n4200 , n13362 );
and ( n13364 , n5696 , n13362 );
or ( n13365 , n13337 , n13363 , n13364 );
and ( n13366 , n4190 , n13365 );
and ( n13367 , n5686 , n13365 );
or ( n13368 , n13336 , n13366 , n13367 );
and ( n13369 , n4180 , n13368 );
and ( n13370 , n5676 , n13368 );
or ( n13371 , n13335 , n13369 , n13370 );
and ( n13372 , n4170 , n13371 );
and ( n13373 , n5666 , n13371 );
or ( n13374 , n13334 , n13372 , n13373 );
and ( n13375 , n4160 , n13374 );
and ( n13376 , n5656 , n13374 );
or ( n13377 , n13333 , n13375 , n13376 );
and ( n13378 , n4150 , n13377 );
and ( n13379 , n5646 , n13377 );
or ( n13380 , n13332 , n13378 , n13379 );
and ( n13381 , n4140 , n13380 );
and ( n13382 , n5636 , n13380 );
or ( n13383 , n13331 , n13381 , n13382 );
and ( n13384 , n4130 , n13383 );
and ( n13385 , n5626 , n13383 );
or ( n13386 , n13330 , n13384 , n13385 );
and ( n13387 , n4120 , n13386 );
and ( n13388 , n5616 , n13386 );
or ( n13389 , n13329 , n13387 , n13388 );
and ( n13390 , n4110 , n13389 );
and ( n13391 , n5606 , n13389 );
or ( n13392 , n13328 , n13390 , n13391 );
and ( n13393 , n4100 , n13392 );
and ( n13394 , n5596 , n13392 );
or ( n13395 , n13327 , n13393 , n13394 );
and ( n13396 , n4090 , n13395 );
and ( n13397 , n5586 , n13395 );
or ( n13398 , n13326 , n13396 , n13397 );
and ( n13399 , n4080 , n13398 );
and ( n13400 , n5576 , n13398 );
or ( n13401 , n13325 , n13399 , n13400 );
and ( n13402 , n4070 , n13401 );
and ( n13403 , n4060 , n13402 );
and ( n13404 , n4050 , n13403 );
and ( n13405 , n4040 , n13404 );
and ( n13406 , n4030 , n13405 );
and ( n13407 , n4020 , n13406 );
and ( n13408 , n4010 , n13407 );
and ( n13409 , n4000 , n13408 );
and ( n13410 , n3990 , n13409 );
and ( n13411 , n3980 , n13410 );
and ( n13412 , n3815 , n13411 );
xor ( n13413 , n3764 , n13412 );
not ( n13414 , n13413 );
xor ( n13415 , n5756 , n3781 );
xor ( n13416 , n13415 , n13344 );
and ( n13417 , n13414 , n13416 );
not ( n13418 , n13416 );
not ( n13419 , n13322 );
xor ( n13420 , n13418 , n13419 );
and ( n13421 , n13420 , n13413 );
or ( n13422 , n13417 , n13421 );
not ( n13423 , n13422 );
not ( n13424 , n13423 );
or ( n13425 , n13324 , n13424 );
not ( n13426 , n13413 );
xor ( n13427 , n5746 , n4254 );
xor ( n13428 , n13427 , n13347 );
and ( n13429 , n13426 , n13428 );
not ( n13430 , n13428 );
and ( n13431 , n13418 , n13419 );
xor ( n13432 , n13430 , n13431 );
and ( n13433 , n13432 , n13413 );
or ( n13434 , n13429 , n13433 );
not ( n13435 , n13434 );
not ( n13436 , n13435 );
or ( n13437 , n13425 , n13436 );
not ( n13438 , n13413 );
xor ( n13439 , n5736 , n4240 );
xor ( n13440 , n13439 , n13350 );
and ( n13441 , n13438 , n13440 );
not ( n13442 , n13440 );
and ( n13443 , n13430 , n13431 );
xor ( n13444 , n13442 , n13443 );
and ( n13445 , n13444 , n13413 );
or ( n13446 , n13441 , n13445 );
not ( n13447 , n13446 );
not ( n13448 , n13447 );
or ( n13449 , n13437 , n13448 );
not ( n13450 , n13413 );
xor ( n13451 , n5726 , n4230 );
xor ( n13452 , n13451 , n13353 );
and ( n13453 , n13450 , n13452 );
not ( n13454 , n13452 );
and ( n13455 , n13442 , n13443 );
xor ( n13456 , n13454 , n13455 );
and ( n13457 , n13456 , n13413 );
or ( n13458 , n13453 , n13457 );
not ( n13459 , n13458 );
not ( n13460 , n13459 );
or ( n13461 , n13449 , n13460 );
not ( n13462 , n13413 );
xor ( n13463 , n5716 , n4220 );
xor ( n13464 , n13463 , n13356 );
and ( n13465 , n13462 , n13464 );
not ( n13466 , n13464 );
and ( n13467 , n13454 , n13455 );
xor ( n13468 , n13466 , n13467 );
and ( n13469 , n13468 , n13413 );
or ( n13470 , n13465 , n13469 );
not ( n13471 , n13470 );
not ( n13472 , n13471 );
or ( n13473 , n13461 , n13472 );
not ( n13474 , n13413 );
xor ( n13475 , n5706 , n4210 );
xor ( n13476 , n13475 , n13359 );
and ( n13477 , n13474 , n13476 );
not ( n13478 , n13476 );
and ( n13479 , n13466 , n13467 );
xor ( n13480 , n13478 , n13479 );
and ( n13481 , n13480 , n13413 );
or ( n13482 , n13477 , n13481 );
not ( n13483 , n13482 );
not ( n13484 , n13483 );
or ( n13485 , n13473 , n13484 );
not ( n13486 , n13413 );
xor ( n13487 , n5696 , n4200 );
xor ( n13488 , n13487 , n13362 );
and ( n13489 , n13486 , n13488 );
not ( n13490 , n13488 );
and ( n13491 , n13478 , n13479 );
xor ( n13492 , n13490 , n13491 );
and ( n13493 , n13492 , n13413 );
or ( n13494 , n13489 , n13493 );
not ( n13495 , n13494 );
not ( n13496 , n13495 );
or ( n13497 , n13485 , n13496 );
not ( n13498 , n13413 );
xor ( n13499 , n5686 , n4190 );
xor ( n13500 , n13499 , n13365 );
and ( n13501 , n13498 , n13500 );
not ( n13502 , n13500 );
and ( n13503 , n13490 , n13491 );
xor ( n13504 , n13502 , n13503 );
and ( n13505 , n13504 , n13413 );
or ( n13506 , n13501 , n13505 );
not ( n13507 , n13506 );
not ( n13508 , n13507 );
or ( n13509 , n13497 , n13508 );
not ( n13510 , n13413 );
xor ( n13511 , n5676 , n4180 );
xor ( n13512 , n13511 , n13368 );
and ( n13513 , n13510 , n13512 );
not ( n13514 , n13512 );
and ( n13515 , n13502 , n13503 );
xor ( n13516 , n13514 , n13515 );
and ( n13517 , n13516 , n13413 );
or ( n13518 , n13513 , n13517 );
not ( n13519 , n13518 );
not ( n13520 , n13519 );
or ( n13521 , n13509 , n13520 );
not ( n13522 , n13413 );
xor ( n13523 , n5666 , n4170 );
xor ( n13524 , n13523 , n13371 );
and ( n13525 , n13522 , n13524 );
not ( n13526 , n13524 );
and ( n13527 , n13514 , n13515 );
xor ( n13528 , n13526 , n13527 );
and ( n13529 , n13528 , n13413 );
or ( n13530 , n13525 , n13529 );
not ( n13531 , n13530 );
not ( n13532 , n13531 );
or ( n13533 , n13521 , n13532 );
not ( n13534 , n13413 );
xor ( n13535 , n5656 , n4160 );
xor ( n13536 , n13535 , n13374 );
and ( n13537 , n13534 , n13536 );
not ( n13538 , n13536 );
and ( n13539 , n13526 , n13527 );
xor ( n13540 , n13538 , n13539 );
and ( n13541 , n13540 , n13413 );
or ( n13542 , n13537 , n13541 );
not ( n13543 , n13542 );
not ( n13544 , n13543 );
or ( n13545 , n13533 , n13544 );
not ( n13546 , n13413 );
xor ( n13547 , n5646 , n4150 );
xor ( n13548 , n13547 , n13377 );
and ( n13549 , n13546 , n13548 );
not ( n13550 , n13548 );
and ( n13551 , n13538 , n13539 );
xor ( n13552 , n13550 , n13551 );
and ( n13553 , n13552 , n13413 );
or ( n13554 , n13549 , n13553 );
not ( n13555 , n13554 );
not ( n13556 , n13555 );
or ( n13557 , n13545 , n13556 );
not ( n13558 , n13413 );
xor ( n13559 , n5636 , n4140 );
xor ( n13560 , n13559 , n13380 );
and ( n13561 , n13558 , n13560 );
not ( n13562 , n13560 );
and ( n13563 , n13550 , n13551 );
xor ( n13564 , n13562 , n13563 );
and ( n13565 , n13564 , n13413 );
or ( n13566 , n13561 , n13565 );
not ( n13567 , n13566 );
not ( n13568 , n13567 );
or ( n13569 , n13557 , n13568 );
not ( n13570 , n13413 );
xor ( n13571 , n5626 , n4130 );
xor ( n13572 , n13571 , n13383 );
and ( n13573 , n13570 , n13572 );
not ( n13574 , n13572 );
and ( n13575 , n13562 , n13563 );
xor ( n13576 , n13574 , n13575 );
and ( n13577 , n13576 , n13413 );
or ( n13578 , n13573 , n13577 );
not ( n13579 , n13578 );
not ( n13580 , n13579 );
or ( n13581 , n13569 , n13580 );
not ( n13582 , n13413 );
xor ( n13583 , n5616 , n4120 );
xor ( n13584 , n13583 , n13386 );
and ( n13585 , n13582 , n13584 );
not ( n13586 , n13584 );
and ( n13587 , n13574 , n13575 );
xor ( n13588 , n13586 , n13587 );
and ( n13589 , n13588 , n13413 );
or ( n13590 , n13585 , n13589 );
not ( n13591 , n13590 );
not ( n13592 , n13591 );
or ( n13593 , n13581 , n13592 );
not ( n13594 , n13413 );
xor ( n13595 , n5606 , n4110 );
xor ( n13596 , n13595 , n13389 );
and ( n13597 , n13594 , n13596 );
not ( n13598 , n13596 );
and ( n13599 , n13586 , n13587 );
xor ( n13600 , n13598 , n13599 );
and ( n13601 , n13600 , n13413 );
or ( n13602 , n13597 , n13601 );
not ( n13603 , n13602 );
not ( n13604 , n13603 );
or ( n13605 , n13593 , n13604 );
not ( n13606 , n13413 );
xor ( n13607 , n5596 , n4100 );
xor ( n13608 , n13607 , n13392 );
and ( n13609 , n13606 , n13608 );
not ( n13610 , n13608 );
and ( n13611 , n13598 , n13599 );
xor ( n13612 , n13610 , n13611 );
and ( n13613 , n13612 , n13413 );
or ( n13614 , n13609 , n13613 );
not ( n13615 , n13614 );
not ( n13616 , n13615 );
or ( n13617 , n13605 , n13616 );
not ( n13618 , n13413 );
xor ( n13619 , n5586 , n4090 );
xor ( n13620 , n13619 , n13395 );
and ( n13621 , n13618 , n13620 );
not ( n13622 , n13620 );
and ( n13623 , n13610 , n13611 );
xor ( n13624 , n13622 , n13623 );
and ( n13625 , n13624 , n13413 );
or ( n13626 , n13621 , n13625 );
not ( n13627 , n13626 );
not ( n13628 , n13627 );
or ( n13629 , n13617 , n13628 );
not ( n13630 , n13413 );
xor ( n13631 , n5576 , n4080 );
xor ( n13632 , n13631 , n13398 );
and ( n13633 , n13630 , n13632 );
not ( n13634 , n13632 );
and ( n13635 , n13622 , n13623 );
xor ( n13636 , n13634 , n13635 );
and ( n13637 , n13636 , n13413 );
or ( n13638 , n13633 , n13637 );
not ( n13639 , n13638 );
not ( n13640 , n13639 );
or ( n13641 , n13629 , n13640 );
and ( n13642 , n13641 , n13413 );
not ( n13643 , n13642 );
and ( n13644 , n13643 , n13324 );
xor ( n13645 , n13324 , n13413 );
xor ( n13646 , n13645 , n13413 );
and ( n13647 , n13646 , n13642 );
or ( n13648 , n13644 , n13647 );
and ( n13649 , n13648 , n5288 );
and ( n13650 , n5491 , n5153 );
and ( n13651 , n2352 , n5155 );
or ( n13652 , n13321 , n13649 , n13650 , n13651 );
or ( n13653 , n6725 , n6720 );
or ( n13654 , n13653 , n6716 );
or ( n13655 , n13654 , n6717 );
or ( n13656 , n13655 , n6705 );
or ( n13657 , n13656 , n6706 );
or ( n13658 , n13657 , n6213 );
or ( n13659 , n13658 , n6214 );
or ( n13660 , n13659 , n6708 );
or ( n13661 , n13660 , n6216 );
or ( n13662 , n13661 , n6710 );
or ( n13663 , n13662 , n6218 );
and ( n13664 , n13652 , n13663 );
or ( n13665 , n12993 , n13664 );
and ( n13666 , n12991 , n13665 );
and ( n13667 , n2424 , n3259 );
or ( n13668 , n13666 , n13667 );
and ( n13669 , n12990 , n13668 );
and ( n13670 , n13652 , n3066 );
or ( n13671 , n13669 , n13670 );
and ( n13672 , n13671 , n2422 );
not ( n13673 , n3356 );
not ( n13674 , n13673 );
buf ( n13675 , n13674 );
and ( n13676 , n13675 , n2428 );
or ( n13677 , n13672 , n13676 );
buf ( n13678 , n13677 );
buf ( n13679 , n2424 );
buf ( n13680 , n2281 );
buf ( n13681 , n2280 );
not ( n13682 , n3066 );
not ( n13683 , n3259 );
and ( n13684 , n2350 , n12992 );
not ( n13685 , n13314 );
and ( n13686 , n13685 , n13096 );
xor ( n13687 , n13096 , n13085 );
and ( n13688 , n13317 , n13085 );
xor ( n13689 , n13687 , n13688 );
and ( n13690 , n13689 , n13314 );
or ( n13691 , n13686 , n13690 );
and ( n13692 , n13691 , n5290 );
not ( n13693 , n13642 );
and ( n13694 , n13693 , n13424 );
xor ( n13695 , n13424 , n13413 );
and ( n13696 , n13645 , n13413 );
xor ( n13697 , n13695 , n13696 );
and ( n13698 , n13697 , n13642 );
or ( n13699 , n13694 , n13698 );
and ( n13700 , n13699 , n5288 );
and ( n13701 , n5756 , n5153 );
and ( n13702 , n2350 , n5155 );
or ( n13703 , n13692 , n13700 , n13701 , n13702 );
and ( n13704 , n13703 , n13663 );
or ( n13705 , n13684 , n13704 );
and ( n13706 , n13683 , n13705 );
and ( n13707 , n2424 , n3259 );
or ( n13708 , n13706 , n13707 );
and ( n13709 , n13682 , n13708 );
and ( n13710 , n13703 , n3066 );
or ( n13711 , n13709 , n13710 );
and ( n13712 , n13711 , n2422 );
buf ( n13713 , n3772 );
not ( n13714 , n13713 );
not ( n13715 , n13714 );
buf ( n13716 , n13715 );
and ( n13717 , n13716 , n2428 );
or ( n13718 , n13712 , n13717 );
buf ( n13719 , n13718 );
buf ( n13720 , n2424 );
buf ( n13721 , n2281 );
buf ( n13722 , n2280 );
not ( n13723 , n3066 );
not ( n13724 , n3259 );
and ( n13725 , n2348 , n12992 );
not ( n13726 , n13314 );
and ( n13727 , n13726 , n13108 );
xor ( n13728 , n13108 , n13085 );
and ( n13729 , n13687 , n13688 );
xor ( n13730 , n13728 , n13729 );
and ( n13731 , n13730 , n13314 );
or ( n13732 , n13727 , n13731 );
and ( n13733 , n13732 , n5290 );
not ( n13734 , n13642 );
and ( n13735 , n13734 , n13436 );
xor ( n13736 , n13436 , n13413 );
and ( n13737 , n13695 , n13696 );
xor ( n13738 , n13736 , n13737 );
and ( n13739 , n13738 , n13642 );
or ( n13740 , n13735 , n13739 );
and ( n13741 , n13740 , n5288 );
and ( n13742 , n5746 , n5153 );
and ( n13743 , n2348 , n5155 );
or ( n13744 , n13733 , n13741 , n13742 , n13743 );
and ( n13745 , n13744 , n13663 );
or ( n13746 , n13725 , n13745 );
and ( n13747 , n13724 , n13746 );
not ( n13748 , n3789 );
not ( n13749 , n13748 );
not ( n13750 , n3635 );
and ( n13751 , n13750 , n3779 );
not ( n13752 , n3779 );
not ( n13753 , n3789 );
xor ( n13754 , n13752 , n13753 );
and ( n13755 , n13754 , n3635 );
or ( n13756 , n13751 , n13755 );
not ( n13757 , n13756 );
not ( n13758 , n13757 );
or ( n13759 , n13749 , n13758 );
not ( n13760 , n3635 );
and ( n13761 , n13760 , n4252 );
not ( n13762 , n4252 );
and ( n13763 , n13752 , n13753 );
xor ( n13764 , n13762 , n13763 );
and ( n13765 , n13764 , n3635 );
or ( n13766 , n13761 , n13765 );
not ( n13767 , n13766 );
not ( n13768 , n13767 );
or ( n13769 , n13759 , n13768 );
not ( n13770 , n3635 );
and ( n13771 , n13770 , n4238 );
not ( n13772 , n4238 );
and ( n13773 , n13762 , n13763 );
xor ( n13774 , n13772 , n13773 );
and ( n13775 , n13774 , n3635 );
or ( n13776 , n13771 , n13775 );
not ( n13777 , n13776 );
not ( n13778 , n13777 );
or ( n13779 , n13769 , n13778 );
not ( n13780 , n3635 );
and ( n13781 , n13780 , n4228 );
not ( n13782 , n4228 );
and ( n13783 , n13772 , n13773 );
xor ( n13784 , n13782 , n13783 );
and ( n13785 , n13784 , n3635 );
or ( n13786 , n13781 , n13785 );
not ( n13787 , n13786 );
not ( n13788 , n13787 );
or ( n13789 , n13779 , n13788 );
not ( n13790 , n3635 );
and ( n13791 , n13790 , n4218 );
not ( n13792 , n4218 );
and ( n13793 , n13782 , n13783 );
xor ( n13794 , n13792 , n13793 );
and ( n13795 , n13794 , n3635 );
or ( n13796 , n13791 , n13795 );
not ( n13797 , n13796 );
not ( n13798 , n13797 );
or ( n13799 , n13789 , n13798 );
not ( n13800 , n3635 );
and ( n13801 , n13800 , n4208 );
not ( n13802 , n4208 );
and ( n13803 , n13792 , n13793 );
xor ( n13804 , n13802 , n13803 );
and ( n13805 , n13804 , n3635 );
or ( n13806 , n13801 , n13805 );
not ( n13807 , n13806 );
not ( n13808 , n13807 );
or ( n13809 , n13799 , n13808 );
not ( n13810 , n3635 );
and ( n13811 , n13810 , n4198 );
not ( n13812 , n4198 );
and ( n13813 , n13802 , n13803 );
xor ( n13814 , n13812 , n13813 );
and ( n13815 , n13814 , n3635 );
or ( n13816 , n13811 , n13815 );
not ( n13817 , n13816 );
not ( n13818 , n13817 );
or ( n13819 , n13809 , n13818 );
not ( n13820 , n3635 );
and ( n13821 , n13820 , n4188 );
not ( n13822 , n4188 );
and ( n13823 , n13812 , n13813 );
xor ( n13824 , n13822 , n13823 );
and ( n13825 , n13824 , n3635 );
or ( n13826 , n13821 , n13825 );
not ( n13827 , n13826 );
not ( n13828 , n13827 );
or ( n13829 , n13819 , n13828 );
not ( n13830 , n3635 );
and ( n13831 , n13830 , n4178 );
not ( n13832 , n4178 );
and ( n13833 , n13822 , n13823 );
xor ( n13834 , n13832 , n13833 );
and ( n13835 , n13834 , n3635 );
or ( n13836 , n13831 , n13835 );
not ( n13837 , n13836 );
not ( n13838 , n13837 );
or ( n13839 , n13829 , n13838 );
not ( n13840 , n3635 );
and ( n13841 , n13840 , n4168 );
not ( n13842 , n4168 );
and ( n13843 , n13832 , n13833 );
xor ( n13844 , n13842 , n13843 );
and ( n13845 , n13844 , n3635 );
or ( n13846 , n13841 , n13845 );
not ( n13847 , n13846 );
not ( n13848 , n13847 );
or ( n13849 , n13839 , n13848 );
not ( n13850 , n3635 );
and ( n13851 , n13850 , n4158 );
not ( n13852 , n4158 );
and ( n13853 , n13842 , n13843 );
xor ( n13854 , n13852 , n13853 );
and ( n13855 , n13854 , n3635 );
or ( n13856 , n13851 , n13855 );
not ( n13857 , n13856 );
not ( n13858 , n13857 );
or ( n13859 , n13849 , n13858 );
not ( n13860 , n3635 );
and ( n13861 , n13860 , n4148 );
not ( n13862 , n4148 );
and ( n13863 , n13852 , n13853 );
xor ( n13864 , n13862 , n13863 );
and ( n13865 , n13864 , n3635 );
or ( n13866 , n13861 , n13865 );
not ( n13867 , n13866 );
not ( n13868 , n13867 );
or ( n13869 , n13859 , n13868 );
not ( n13870 , n3635 );
and ( n13871 , n13870 , n4138 );
not ( n13872 , n4138 );
and ( n13873 , n13862 , n13863 );
xor ( n13874 , n13872 , n13873 );
and ( n13875 , n13874 , n3635 );
or ( n13876 , n13871 , n13875 );
not ( n13877 , n13876 );
not ( n13878 , n13877 );
or ( n13879 , n13869 , n13878 );
not ( n13880 , n3635 );
and ( n13881 , n13880 , n4128 );
not ( n13882 , n4128 );
and ( n13883 , n13872 , n13873 );
xor ( n13884 , n13882 , n13883 );
and ( n13885 , n13884 , n3635 );
or ( n13886 , n13881 , n13885 );
not ( n13887 , n13886 );
not ( n13888 , n13887 );
or ( n13889 , n13879 , n13888 );
not ( n13890 , n3635 );
and ( n13891 , n13890 , n4118 );
not ( n13892 , n4118 );
and ( n13893 , n13882 , n13883 );
xor ( n13894 , n13892 , n13893 );
and ( n13895 , n13894 , n3635 );
or ( n13896 , n13891 , n13895 );
not ( n13897 , n13896 );
not ( n13898 , n13897 );
or ( n13899 , n13889 , n13898 );
not ( n13900 , n3635 );
and ( n13901 , n13900 , n4108 );
not ( n13902 , n4108 );
and ( n13903 , n13892 , n13893 );
xor ( n13904 , n13902 , n13903 );
and ( n13905 , n13904 , n3635 );
or ( n13906 , n13901 , n13905 );
not ( n13907 , n13906 );
not ( n13908 , n13907 );
or ( n13909 , n13899 , n13908 );
not ( n13910 , n3635 );
and ( n13911 , n13910 , n4098 );
not ( n13912 , n4098 );
and ( n13913 , n13902 , n13903 );
xor ( n13914 , n13912 , n13913 );
and ( n13915 , n13914 , n3635 );
or ( n13916 , n13911 , n13915 );
not ( n13917 , n13916 );
not ( n13918 , n13917 );
or ( n13919 , n13909 , n13918 );
not ( n13920 , n3635 );
and ( n13921 , n13920 , n4088 );
not ( n13922 , n4088 );
and ( n13923 , n13912 , n13913 );
xor ( n13924 , n13922 , n13923 );
and ( n13925 , n13924 , n3635 );
or ( n13926 , n13921 , n13925 );
not ( n13927 , n13926 );
not ( n13928 , n13927 );
or ( n13929 , n13919 , n13928 );
not ( n13930 , n3635 );
and ( n13931 , n13930 , n4078 );
not ( n13932 , n4078 );
and ( n13933 , n13922 , n13923 );
xor ( n13934 , n13932 , n13933 );
and ( n13935 , n13934 , n3635 );
or ( n13936 , n13931 , n13935 );
not ( n13937 , n13936 );
not ( n13938 , n13937 );
or ( n13939 , n13929 , n13938 );
and ( n13940 , n13939 , n3635 );
not ( n13941 , n13940 );
and ( n13942 , n13941 , n13749 );
xor ( n13943 , n13749 , n3635 );
xor ( n13944 , n13943 , n3635 );
and ( n13945 , n13944 , n13940 );
or ( n13946 , n13942 , n13945 );
not ( n13947 , n5491 );
not ( n13948 , n13947 );
xor ( n13949 , n13946 , n13948 );
and ( n13950 , n13949 , n5290 );
not ( n13951 , n3791 );
not ( n13952 , n13951 );
not ( n13953 , n3764 );
and ( n13954 , n13953 , n3781 );
not ( n13955 , n3781 );
not ( n13956 , n3791 );
xor ( n13957 , n13955 , n13956 );
and ( n13958 , n13957 , n3764 );
or ( n13959 , n13954 , n13958 );
not ( n13960 , n13959 );
not ( n13961 , n13960 );
or ( n13962 , n13952 , n13961 );
not ( n13963 , n3764 );
and ( n13964 , n13963 , n4254 );
not ( n13965 , n4254 );
and ( n13966 , n13955 , n13956 );
xor ( n13967 , n13965 , n13966 );
and ( n13968 , n13967 , n3764 );
or ( n13969 , n13964 , n13968 );
not ( n13970 , n13969 );
not ( n13971 , n13970 );
or ( n13972 , n13962 , n13971 );
not ( n13973 , n3764 );
and ( n13974 , n13973 , n4240 );
not ( n13975 , n4240 );
and ( n13976 , n13965 , n13966 );
xor ( n13977 , n13975 , n13976 );
and ( n13978 , n13977 , n3764 );
or ( n13979 , n13974 , n13978 );
not ( n13980 , n13979 );
not ( n13981 , n13980 );
or ( n13982 , n13972 , n13981 );
not ( n13983 , n3764 );
and ( n13984 , n13983 , n4230 );
not ( n13985 , n4230 );
and ( n13986 , n13975 , n13976 );
xor ( n13987 , n13985 , n13986 );
and ( n13988 , n13987 , n3764 );
or ( n13989 , n13984 , n13988 );
not ( n13990 , n13989 );
not ( n13991 , n13990 );
or ( n13992 , n13982 , n13991 );
not ( n13993 , n3764 );
and ( n13994 , n13993 , n4220 );
not ( n13995 , n4220 );
and ( n13996 , n13985 , n13986 );
xor ( n13997 , n13995 , n13996 );
and ( n13998 , n13997 , n3764 );
or ( n13999 , n13994 , n13998 );
not ( n14000 , n13999 );
not ( n14001 , n14000 );
or ( n14002 , n13992 , n14001 );
not ( n14003 , n3764 );
and ( n14004 , n14003 , n4210 );
not ( n14005 , n4210 );
and ( n14006 , n13995 , n13996 );
xor ( n14007 , n14005 , n14006 );
and ( n14008 , n14007 , n3764 );
or ( n14009 , n14004 , n14008 );
not ( n14010 , n14009 );
not ( n14011 , n14010 );
or ( n14012 , n14002 , n14011 );
not ( n14013 , n3764 );
and ( n14014 , n14013 , n4200 );
not ( n14015 , n4200 );
and ( n14016 , n14005 , n14006 );
xor ( n14017 , n14015 , n14016 );
and ( n14018 , n14017 , n3764 );
or ( n14019 , n14014 , n14018 );
not ( n14020 , n14019 );
not ( n14021 , n14020 );
or ( n14022 , n14012 , n14021 );
not ( n14023 , n3764 );
and ( n14024 , n14023 , n4190 );
not ( n14025 , n4190 );
and ( n14026 , n14015 , n14016 );
xor ( n14027 , n14025 , n14026 );
and ( n14028 , n14027 , n3764 );
or ( n14029 , n14024 , n14028 );
not ( n14030 , n14029 );
not ( n14031 , n14030 );
or ( n14032 , n14022 , n14031 );
not ( n14033 , n3764 );
and ( n14034 , n14033 , n4180 );
not ( n14035 , n4180 );
and ( n14036 , n14025 , n14026 );
xor ( n14037 , n14035 , n14036 );
and ( n14038 , n14037 , n3764 );
or ( n14039 , n14034 , n14038 );
not ( n14040 , n14039 );
not ( n14041 , n14040 );
or ( n14042 , n14032 , n14041 );
not ( n14043 , n3764 );
and ( n14044 , n14043 , n4170 );
not ( n14045 , n4170 );
and ( n14046 , n14035 , n14036 );
xor ( n14047 , n14045 , n14046 );
and ( n14048 , n14047 , n3764 );
or ( n14049 , n14044 , n14048 );
not ( n14050 , n14049 );
not ( n14051 , n14050 );
or ( n14052 , n14042 , n14051 );
not ( n14053 , n3764 );
and ( n14054 , n14053 , n4160 );
not ( n14055 , n4160 );
and ( n14056 , n14045 , n14046 );
xor ( n14057 , n14055 , n14056 );
and ( n14058 , n14057 , n3764 );
or ( n14059 , n14054 , n14058 );
not ( n14060 , n14059 );
not ( n14061 , n14060 );
or ( n14062 , n14052 , n14061 );
not ( n14063 , n3764 );
and ( n14064 , n14063 , n4150 );
not ( n14065 , n4150 );
and ( n14066 , n14055 , n14056 );
xor ( n14067 , n14065 , n14066 );
and ( n14068 , n14067 , n3764 );
or ( n14069 , n14064 , n14068 );
not ( n14070 , n14069 );
not ( n14071 , n14070 );
or ( n14072 , n14062 , n14071 );
not ( n14073 , n3764 );
and ( n14074 , n14073 , n4140 );
not ( n14075 , n4140 );
and ( n14076 , n14065 , n14066 );
xor ( n14077 , n14075 , n14076 );
and ( n14078 , n14077 , n3764 );
or ( n14079 , n14074 , n14078 );
not ( n14080 , n14079 );
not ( n14081 , n14080 );
or ( n14082 , n14072 , n14081 );
not ( n14083 , n3764 );
and ( n14084 , n14083 , n4130 );
not ( n14085 , n4130 );
and ( n14086 , n14075 , n14076 );
xor ( n14087 , n14085 , n14086 );
and ( n14088 , n14087 , n3764 );
or ( n14089 , n14084 , n14088 );
not ( n14090 , n14089 );
not ( n14091 , n14090 );
or ( n14092 , n14082 , n14091 );
not ( n14093 , n3764 );
and ( n14094 , n14093 , n4120 );
not ( n14095 , n4120 );
and ( n14096 , n14085 , n14086 );
xor ( n14097 , n14095 , n14096 );
and ( n14098 , n14097 , n3764 );
or ( n14099 , n14094 , n14098 );
not ( n14100 , n14099 );
not ( n14101 , n14100 );
or ( n14102 , n14092 , n14101 );
not ( n14103 , n3764 );
and ( n14104 , n14103 , n4110 );
not ( n14105 , n4110 );
and ( n14106 , n14095 , n14096 );
xor ( n14107 , n14105 , n14106 );
and ( n14108 , n14107 , n3764 );
or ( n14109 , n14104 , n14108 );
not ( n14110 , n14109 );
not ( n14111 , n14110 );
or ( n14112 , n14102 , n14111 );
not ( n14113 , n3764 );
and ( n14114 , n14113 , n4100 );
not ( n14115 , n4100 );
and ( n14116 , n14105 , n14106 );
xor ( n14117 , n14115 , n14116 );
and ( n14118 , n14117 , n3764 );
or ( n14119 , n14114 , n14118 );
not ( n14120 , n14119 );
not ( n14121 , n14120 );
or ( n14122 , n14112 , n14121 );
not ( n14123 , n3764 );
and ( n14124 , n14123 , n4090 );
not ( n14125 , n4090 );
and ( n14126 , n14115 , n14116 );
xor ( n14127 , n14125 , n14126 );
and ( n14128 , n14127 , n3764 );
or ( n14129 , n14124 , n14128 );
not ( n14130 , n14129 );
not ( n14131 , n14130 );
or ( n14132 , n14122 , n14131 );
not ( n14133 , n3764 );
and ( n14134 , n14133 , n4080 );
not ( n14135 , n4080 );
and ( n14136 , n14125 , n14126 );
xor ( n14137 , n14135 , n14136 );
and ( n14138 , n14137 , n3764 );
or ( n14139 , n14134 , n14138 );
not ( n14140 , n14139 );
not ( n14141 , n14140 );
or ( n14142 , n14132 , n14141 );
and ( n14143 , n14142 , n3764 );
not ( n14144 , n14143 );
and ( n14145 , n14144 , n13952 );
xor ( n14146 , n13952 , n3764 );
xor ( n14147 , n14146 , n3764 );
and ( n14148 , n14147 , n14143 );
or ( n14149 , n14145 , n14148 );
xor ( n14150 , n14149 , n13948 );
and ( n14151 , n14150 , n5288 );
or ( n14152 , n5155 , n5153 );
and ( n14153 , n5491 , n14152 );
or ( n14154 , n13950 , n14151 , n14153 );
not ( n14155 , n14154 );
not ( n14156 , n14155 );
buf ( n14157 , n14156 );
and ( n14158 , n14157 , n3259 );
or ( n14159 , n13747 , n14158 );
and ( n14160 , n13723 , n14159 );
and ( n14161 , n13744 , n3066 );
or ( n14162 , n14160 , n14161 );
and ( n14163 , n14162 , n2422 );
buf ( n14164 , n4246 );
not ( n14165 , n14164 );
not ( n14166 , n14165 );
buf ( n14167 , n14166 );
and ( n14168 , n14167 , n2428 );
or ( n14169 , n14163 , n14168 );
buf ( n14170 , n14169 );
buf ( n14171 , n2424 );
buf ( n14172 , n2281 );
buf ( n14173 , n2280 );
not ( n14174 , n3066 );
not ( n14175 , n3259 );
and ( n14176 , n2346 , n12992 );
not ( n14177 , n13314 );
and ( n14178 , n14177 , n13120 );
xor ( n14179 , n13120 , n13085 );
and ( n14180 , n13728 , n13729 );
xor ( n14181 , n14179 , n14180 );
and ( n14182 , n14181 , n13314 );
or ( n14183 , n14178 , n14182 );
and ( n14184 , n14183 , n5290 );
not ( n14185 , n13642 );
and ( n14186 , n14185 , n13448 );
xor ( n14187 , n13448 , n13413 );
and ( n14188 , n13736 , n13737 );
xor ( n14189 , n14187 , n14188 );
and ( n14190 , n14189 , n13642 );
or ( n14191 , n14186 , n14190 );
and ( n14192 , n14191 , n5288 );
and ( n14193 , n5736 , n5153 );
and ( n14194 , n2346 , n5155 );
or ( n14195 , n14184 , n14192 , n14193 , n14194 );
and ( n14196 , n14195 , n13663 );
or ( n14197 , n14176 , n14196 );
and ( n14198 , n14175 , n14197 );
and ( n14199 , n2424 , n3259 );
or ( n14200 , n14198 , n14199 );
and ( n14201 , n14174 , n14200 );
and ( n14202 , n14195 , n3066 );
or ( n14203 , n14201 , n14202 );
and ( n14204 , n14203 , n2422 );
buf ( n14205 , n3946 );
not ( n14206 , n14205 );
not ( n14207 , n14206 );
buf ( n14208 , n14207 );
and ( n14209 , n14208 , n2428 );
or ( n14210 , n14204 , n14209 );
buf ( n14211 , n14210 );
buf ( n14212 , n2424 );
buf ( n14213 , n2281 );
buf ( n14214 , n2280 );
not ( n14215 , n3066 );
not ( n14216 , n3259 );
and ( n14217 , n2344 , n12992 );
not ( n14218 , n13314 );
and ( n14219 , n14218 , n13132 );
xor ( n14220 , n13132 , n13085 );
and ( n14221 , n14179 , n14180 );
xor ( n14222 , n14220 , n14221 );
and ( n14223 , n14222 , n13314 );
or ( n14224 , n14219 , n14223 );
and ( n14225 , n14224 , n5290 );
not ( n14226 , n13642 );
and ( n14227 , n14226 , n13460 );
xor ( n14228 , n13460 , n13413 );
and ( n14229 , n14187 , n14188 );
xor ( n14230 , n14228 , n14229 );
and ( n14231 , n14230 , n13642 );
or ( n14232 , n14227 , n14231 );
and ( n14233 , n14232 , n5288 );
and ( n14234 , n5726 , n5153 );
and ( n14235 , n2344 , n5155 );
or ( n14236 , n14225 , n14233 , n14234 , n14235 );
and ( n14237 , n14236 , n13663 );
or ( n14238 , n14217 , n14237 );
and ( n14239 , n14216 , n14238 );
buf ( n14240 , n14157 );
and ( n14241 , n14240 , n3259 );
or ( n14242 , n14239 , n14241 );
and ( n14243 , n14215 , n14242 );
and ( n14244 , n14236 , n3066 );
or ( n14245 , n14243 , n14244 );
and ( n14246 , n14245 , n2422 );
buf ( n14247 , n3941 );
not ( n14248 , n14247 );
not ( n14249 , n14248 );
buf ( n14250 , n14249 );
and ( n14251 , n14250 , n2428 );
or ( n14252 , n14246 , n14251 );
buf ( n14253 , n14252 );
buf ( n14254 , n2424 );
buf ( n14255 , n2281 );
buf ( n14256 , n2280 );
not ( n14257 , n3066 );
not ( n14258 , n3259 );
and ( n14259 , n2342 , n12992 );
not ( n14260 , n13314 );
and ( n14261 , n14260 , n13144 );
xor ( n14262 , n13144 , n13085 );
and ( n14263 , n14220 , n14221 );
xor ( n14264 , n14262 , n14263 );
and ( n14265 , n14264 , n13314 );
or ( n14266 , n14261 , n14265 );
and ( n14267 , n14266 , n5290 );
not ( n14268 , n13642 );
and ( n14269 , n14268 , n13472 );
xor ( n14270 , n13472 , n13413 );
and ( n14271 , n14228 , n14229 );
xor ( n14272 , n14270 , n14271 );
and ( n14273 , n14272 , n13642 );
or ( n14274 , n14269 , n14273 );
and ( n14275 , n14274 , n5288 );
and ( n14276 , n5716 , n5153 );
and ( n14277 , n2342 , n5155 );
or ( n14278 , n14267 , n14275 , n14276 , n14277 );
and ( n14279 , n14278 , n13663 );
or ( n14280 , n14259 , n14279 );
and ( n14281 , n14258 , n14280 );
and ( n14282 , n2424 , n3259 );
or ( n14283 , n14281 , n14282 );
and ( n14284 , n14257 , n14283 );
and ( n14285 , n14278 , n3066 );
or ( n14286 , n14284 , n14285 );
and ( n14287 , n14286 , n2422 );
buf ( n14288 , n3936 );
not ( n14289 , n14288 );
not ( n14290 , n14289 );
buf ( n14291 , n14290 );
and ( n14292 , n14291 , n2428 );
or ( n14293 , n14287 , n14292 );
buf ( n14294 , n14293 );
buf ( n14295 , n2424 );
buf ( n14296 , n2281 );
buf ( n14297 , n2280 );
not ( n14298 , n3066 );
not ( n14299 , n3259 );
and ( n14300 , n2340 , n12992 );
not ( n14301 , n13314 );
and ( n14302 , n14301 , n13156 );
xor ( n14303 , n13156 , n13085 );
and ( n14304 , n14262 , n14263 );
xor ( n14305 , n14303 , n14304 );
and ( n14306 , n14305 , n13314 );
or ( n14307 , n14302 , n14306 );
and ( n14308 , n14307 , n5290 );
not ( n14309 , n13642 );
and ( n14310 , n14309 , n13484 );
xor ( n14311 , n13484 , n13413 );
and ( n14312 , n14270 , n14271 );
xor ( n14313 , n14311 , n14312 );
and ( n14314 , n14313 , n13642 );
or ( n14315 , n14310 , n14314 );
and ( n14316 , n14315 , n5288 );
and ( n14317 , n5706 , n5153 );
and ( n14318 , n2340 , n5155 );
or ( n14319 , n14308 , n14316 , n14317 , n14318 );
and ( n14320 , n14319 , n13663 );
or ( n14321 , n14300 , n14320 );
and ( n14322 , n14299 , n14321 );
and ( n14323 , n2424 , n3259 );
or ( n14324 , n14322 , n14323 );
and ( n14325 , n14298 , n14324 );
and ( n14326 , n14319 , n3066 );
or ( n14327 , n14325 , n14326 );
and ( n14328 , n14327 , n2422 );
buf ( n14329 , n3931 );
not ( n14330 , n14329 );
not ( n14331 , n14330 );
buf ( n14332 , n14331 );
and ( n14333 , n14332 , n2428 );
or ( n14334 , n14328 , n14333 );
buf ( n14335 , n14334 );
buf ( n14336 , n2424 );
buf ( n14337 , n2281 );
buf ( n14338 , n2280 );
not ( n14339 , n3066 );
not ( n14340 , n3259 );
and ( n14341 , n2338 , n12992 );
not ( n14342 , n13314 );
and ( n14343 , n14342 , n13168 );
xor ( n14344 , n13168 , n13085 );
and ( n14345 , n14303 , n14304 );
xor ( n14346 , n14344 , n14345 );
and ( n14347 , n14346 , n13314 );
or ( n14348 , n14343 , n14347 );
and ( n14349 , n14348 , n5290 );
not ( n14350 , n13642 );
and ( n14351 , n14350 , n13496 );
xor ( n14352 , n13496 , n13413 );
and ( n14353 , n14311 , n14312 );
xor ( n14354 , n14352 , n14353 );
and ( n14355 , n14354 , n13642 );
or ( n14356 , n14351 , n14355 );
and ( n14357 , n14356 , n5288 );
and ( n14358 , n5696 , n5153 );
and ( n14359 , n2338 , n5155 );
or ( n14360 , n14349 , n14357 , n14358 , n14359 );
and ( n14361 , n14360 , n13663 );
or ( n14362 , n14341 , n14361 );
and ( n14363 , n14340 , n14362 );
and ( n14364 , n2424 , n3259 );
or ( n14365 , n14363 , n14364 );
and ( n14366 , n14339 , n14365 );
and ( n14367 , n14360 , n3066 );
or ( n14368 , n14366 , n14367 );
and ( n14369 , n14368 , n2422 );
buf ( n14370 , n3926 );
not ( n14371 , n14370 );
not ( n14372 , n14371 );
buf ( n14373 , n14372 );
and ( n14374 , n14373 , n2428 );
or ( n14375 , n14369 , n14374 );
buf ( n14376 , n14375 );
buf ( n14377 , n2424 );
buf ( n14378 , n2281 );
buf ( n14379 , n2280 );
not ( n14380 , n3066 );
not ( n14381 , n3259 );
and ( n14382 , n2336 , n12992 );
not ( n14383 , n13314 );
and ( n14384 , n14383 , n13180 );
xor ( n14385 , n13180 , n13085 );
and ( n14386 , n14344 , n14345 );
xor ( n14387 , n14385 , n14386 );
and ( n14388 , n14387 , n13314 );
or ( n14389 , n14384 , n14388 );
and ( n14390 , n14389 , n5290 );
not ( n14391 , n13642 );
and ( n14392 , n14391 , n13508 );
xor ( n14393 , n13508 , n13413 );
and ( n14394 , n14352 , n14353 );
xor ( n14395 , n14393 , n14394 );
and ( n14396 , n14395 , n13642 );
or ( n14397 , n14392 , n14396 );
and ( n14398 , n14397 , n5288 );
and ( n14399 , n5686 , n5153 );
and ( n14400 , n2336 , n5155 );
or ( n14401 , n14390 , n14398 , n14399 , n14400 );
and ( n14402 , n14401 , n13663 );
or ( n14403 , n14382 , n14402 );
and ( n14404 , n14381 , n14403 );
and ( n14405 , n2424 , n3259 );
or ( n14406 , n14404 , n14405 );
and ( n14407 , n14380 , n14406 );
and ( n14408 , n14401 , n3066 );
or ( n14409 , n14407 , n14408 );
and ( n14410 , n14409 , n2422 );
buf ( n14411 , n3921 );
not ( n14412 , n14411 );
not ( n14413 , n14412 );
buf ( n14414 , n14413 );
and ( n14415 , n14414 , n2428 );
or ( n14416 , n14410 , n14415 );
buf ( n14417 , n14416 );
buf ( n14418 , n2424 );
buf ( n14419 , n2281 );
buf ( n14420 , n2280 );
not ( n14421 , n3066 );
not ( n14422 , n3259 );
and ( n14423 , n2334 , n12992 );
not ( n14424 , n13314 );
and ( n14425 , n14424 , n13192 );
xor ( n14426 , n13192 , n13085 );
and ( n14427 , n14385 , n14386 );
xor ( n14428 , n14426 , n14427 );
and ( n14429 , n14428 , n13314 );
or ( n14430 , n14425 , n14429 );
and ( n14431 , n14430 , n5290 );
not ( n14432 , n13642 );
and ( n14433 , n14432 , n13520 );
xor ( n14434 , n13520 , n13413 );
and ( n14435 , n14393 , n14394 );
xor ( n14436 , n14434 , n14435 );
and ( n14437 , n14436 , n13642 );
or ( n14438 , n14433 , n14437 );
and ( n14439 , n14438 , n5288 );
and ( n14440 , n5676 , n5153 );
and ( n14441 , n2334 , n5155 );
or ( n14442 , n14431 , n14439 , n14440 , n14441 );
and ( n14443 , n14442 , n13663 );
or ( n14444 , n14423 , n14443 );
and ( n14445 , n14422 , n14444 );
and ( n14446 , n2424 , n3259 );
or ( n14447 , n14445 , n14446 );
and ( n14448 , n14421 , n14447 );
and ( n14449 , n14442 , n3066 );
or ( n14450 , n14448 , n14449 );
and ( n14451 , n14450 , n2422 );
buf ( n14452 , n3916 );
not ( n14453 , n14452 );
not ( n14454 , n14453 );
buf ( n14455 , n14454 );
and ( n14456 , n14455 , n2428 );
or ( n14457 , n14451 , n14456 );
buf ( n14458 , n14457 );
buf ( n14459 , n2424 );
buf ( n14460 , n2281 );
buf ( n14461 , n2280 );
not ( n14462 , n3066 );
not ( n14463 , n3259 );
and ( n14464 , n2332 , n12992 );
not ( n14465 , n13314 );
and ( n14466 , n14465 , n13204 );
xor ( n14467 , n13204 , n13085 );
and ( n14468 , n14426 , n14427 );
xor ( n14469 , n14467 , n14468 );
and ( n14470 , n14469 , n13314 );
or ( n14471 , n14466 , n14470 );
and ( n14472 , n14471 , n5290 );
not ( n14473 , n13642 );
and ( n14474 , n14473 , n13532 );
xor ( n14475 , n13532 , n13413 );
and ( n14476 , n14434 , n14435 );
xor ( n14477 , n14475 , n14476 );
and ( n14478 , n14477 , n13642 );
or ( n14479 , n14474 , n14478 );
and ( n14480 , n14479 , n5288 );
and ( n14481 , n5666 , n5153 );
and ( n14482 , n2332 , n5155 );
or ( n14483 , n14472 , n14480 , n14481 , n14482 );
and ( n14484 , n14483 , n13663 );
or ( n14485 , n14464 , n14484 );
and ( n14486 , n14463 , n14485 );
and ( n14487 , n2424 , n3259 );
or ( n14488 , n14486 , n14487 );
and ( n14489 , n14462 , n14488 );
and ( n14490 , n14483 , n3066 );
or ( n14491 , n14489 , n14490 );
and ( n14492 , n14491 , n2422 );
buf ( n14493 , n3911 );
not ( n14494 , n14493 );
not ( n14495 , n14494 );
buf ( n14496 , n14495 );
and ( n14497 , n14496 , n2428 );
or ( n14498 , n14492 , n14497 );
buf ( n14499 , n14498 );
buf ( n14500 , n2424 );
buf ( n14501 , n2281 );
buf ( n14502 , n2280 );
not ( n14503 , n3066 );
not ( n14504 , n3259 );
and ( n14505 , n2330 , n12992 );
not ( n14506 , n13314 );
and ( n14507 , n14506 , n13216 );
xor ( n14508 , n13216 , n13085 );
and ( n14509 , n14467 , n14468 );
xor ( n14510 , n14508 , n14509 );
and ( n14511 , n14510 , n13314 );
or ( n14512 , n14507 , n14511 );
and ( n14513 , n14512 , n5290 );
not ( n14514 , n13642 );
and ( n14515 , n14514 , n13544 );
xor ( n14516 , n13544 , n13413 );
and ( n14517 , n14475 , n14476 );
xor ( n14518 , n14516 , n14517 );
and ( n14519 , n14518 , n13642 );
or ( n14520 , n14515 , n14519 );
and ( n14521 , n14520 , n5288 );
and ( n14522 , n5656 , n5153 );
and ( n14523 , n2330 , n5155 );
or ( n14524 , n14513 , n14521 , n14522 , n14523 );
and ( n14525 , n14524 , n13663 );
or ( n14526 , n14505 , n14525 );
and ( n14527 , n14504 , n14526 );
and ( n14528 , n2424 , n3259 );
or ( n14529 , n14527 , n14528 );
and ( n14530 , n14503 , n14529 );
and ( n14531 , n14524 , n3066 );
or ( n14532 , n14530 , n14531 );
and ( n14533 , n14532 , n2422 );
buf ( n14534 , n3906 );
not ( n14535 , n14534 );
not ( n14536 , n14535 );
buf ( n14537 , n14536 );
and ( n14538 , n14537 , n2428 );
or ( n14539 , n14533 , n14538 );
buf ( n14540 , n14539 );
buf ( n14541 , n2424 );
buf ( n14542 , n2281 );
buf ( n14543 , n2280 );
not ( n14544 , n3066 );
not ( n14545 , n3259 );
and ( n14546 , n2328 , n12992 );
not ( n14547 , n13314 );
and ( n14548 , n14547 , n13228 );
xor ( n14549 , n13228 , n13085 );
and ( n14550 , n14508 , n14509 );
xor ( n14551 , n14549 , n14550 );
and ( n14552 , n14551 , n13314 );
or ( n14553 , n14548 , n14552 );
and ( n14554 , n14553 , n5290 );
not ( n14555 , n13642 );
and ( n14556 , n14555 , n13556 );
xor ( n14557 , n13556 , n13413 );
and ( n14558 , n14516 , n14517 );
xor ( n14559 , n14557 , n14558 );
and ( n14560 , n14559 , n13642 );
or ( n14561 , n14556 , n14560 );
and ( n14562 , n14561 , n5288 );
and ( n14563 , n5646 , n5153 );
and ( n14564 , n2328 , n5155 );
or ( n14565 , n14554 , n14562 , n14563 , n14564 );
and ( n14566 , n14565 , n13663 );
or ( n14567 , n14546 , n14566 );
and ( n14568 , n14545 , n14567 );
and ( n14569 , n2424 , n3259 );
or ( n14570 , n14568 , n14569 );
and ( n14571 , n14544 , n14570 );
and ( n14572 , n14565 , n3066 );
or ( n14573 , n14571 , n14572 );
and ( n14574 , n14573 , n2422 );
buf ( n14575 , n3901 );
not ( n14576 , n14575 );
not ( n14577 , n14576 );
buf ( n14578 , n14577 );
and ( n14579 , n14578 , n2428 );
or ( n14580 , n14574 , n14579 );
buf ( n14581 , n14580 );
buf ( n14582 , n2424 );
buf ( n14583 , n2281 );
buf ( n14584 , n2280 );
not ( n14585 , n3066 );
not ( n14586 , n3259 );
and ( n14587 , n2326 , n12992 );
not ( n14588 , n13314 );
and ( n14589 , n14588 , n13240 );
xor ( n14590 , n13240 , n13085 );
and ( n14591 , n14549 , n14550 );
xor ( n14592 , n14590 , n14591 );
and ( n14593 , n14592 , n13314 );
or ( n14594 , n14589 , n14593 );
and ( n14595 , n14594 , n5290 );
not ( n14596 , n13642 );
and ( n14597 , n14596 , n13568 );
xor ( n14598 , n13568 , n13413 );
and ( n14599 , n14557 , n14558 );
xor ( n14600 , n14598 , n14599 );
and ( n14601 , n14600 , n13642 );
or ( n14602 , n14597 , n14601 );
and ( n14603 , n14602 , n5288 );
and ( n14604 , n5636 , n5153 );
and ( n14605 , n2326 , n5155 );
or ( n14606 , n14595 , n14603 , n14604 , n14605 );
and ( n14607 , n14606 , n13663 );
or ( n14608 , n14587 , n14607 );
and ( n14609 , n14586 , n14608 );
and ( n14610 , n2424 , n3259 );
or ( n14611 , n14609 , n14610 );
and ( n14612 , n14585 , n14611 );
and ( n14613 , n14606 , n3066 );
or ( n14614 , n14612 , n14613 );
and ( n14615 , n14614 , n2422 );
buf ( n14616 , n3896 );
not ( n14617 , n14616 );
not ( n14618 , n14617 );
buf ( n14619 , n14618 );
and ( n14620 , n14619 , n2428 );
or ( n14621 , n14615 , n14620 );
buf ( n14622 , n14621 );
buf ( n14623 , n2424 );
buf ( n14624 , n2281 );
buf ( n14625 , n2280 );
not ( n14626 , n3066 );
not ( n14627 , n3259 );
and ( n14628 , n2324 , n12992 );
not ( n14629 , n13314 );
and ( n14630 , n14629 , n13252 );
xor ( n14631 , n13252 , n13085 );
and ( n14632 , n14590 , n14591 );
xor ( n14633 , n14631 , n14632 );
and ( n14634 , n14633 , n13314 );
or ( n14635 , n14630 , n14634 );
and ( n14636 , n14635 , n5290 );
not ( n14637 , n13642 );
and ( n14638 , n14637 , n13580 );
xor ( n14639 , n13580 , n13413 );
and ( n14640 , n14598 , n14599 );
xor ( n14641 , n14639 , n14640 );
and ( n14642 , n14641 , n13642 );
or ( n14643 , n14638 , n14642 );
and ( n14644 , n14643 , n5288 );
and ( n14645 , n5626 , n5153 );
and ( n14646 , n2324 , n5155 );
or ( n14647 , n14636 , n14644 , n14645 , n14646 );
and ( n14648 , n14647 , n13663 );
or ( n14649 , n14628 , n14648 );
and ( n14650 , n14627 , n14649 );
and ( n14651 , n2424 , n3259 );
or ( n14652 , n14650 , n14651 );
and ( n14653 , n14626 , n14652 );
and ( n14654 , n14647 , n3066 );
or ( n14655 , n14653 , n14654 );
and ( n14656 , n14655 , n2422 );
buf ( n14657 , n3891 );
not ( n14658 , n14657 );
not ( n14659 , n14658 );
buf ( n14660 , n14659 );
and ( n14661 , n14660 , n2428 );
or ( n14662 , n14656 , n14661 );
buf ( n14663 , n14662 );
buf ( n14664 , n2424 );
buf ( n14665 , n2281 );
buf ( n14666 , n2280 );
not ( n14667 , n3066 );
not ( n14668 , n3259 );
and ( n14669 , n2322 , n12992 );
not ( n14670 , n13314 );
and ( n14671 , n14670 , n13264 );
xor ( n14672 , n13264 , n13085 );
and ( n14673 , n14631 , n14632 );
xor ( n14674 , n14672 , n14673 );
and ( n14675 , n14674 , n13314 );
or ( n14676 , n14671 , n14675 );
and ( n14677 , n14676 , n5290 );
not ( n14678 , n13642 );
and ( n14679 , n14678 , n13592 );
xor ( n14680 , n13592 , n13413 );
and ( n14681 , n14639 , n14640 );
xor ( n14682 , n14680 , n14681 );
and ( n14683 , n14682 , n13642 );
or ( n14684 , n14679 , n14683 );
and ( n14685 , n14684 , n5288 );
and ( n14686 , n5616 , n5153 );
and ( n14687 , n2322 , n5155 );
or ( n14688 , n14677 , n14685 , n14686 , n14687 );
and ( n14689 , n14688 , n13663 );
or ( n14690 , n14669 , n14689 );
and ( n14691 , n14668 , n14690 );
and ( n14692 , n2424 , n3259 );
or ( n14693 , n14691 , n14692 );
and ( n14694 , n14667 , n14693 );
and ( n14695 , n14688 , n3066 );
or ( n14696 , n14694 , n14695 );
and ( n14697 , n14696 , n2422 );
buf ( n14698 , n3886 );
not ( n14699 , n14698 );
not ( n14700 , n14699 );
buf ( n14701 , n14700 );
and ( n14702 , n14701 , n2428 );
or ( n14703 , n14697 , n14702 );
buf ( n14704 , n14703 );
buf ( n14705 , n2424 );
buf ( n14706 , n2281 );
buf ( n14707 , n2280 );
not ( n14708 , n3066 );
not ( n14709 , n3259 );
and ( n14710 , n2320 , n12992 );
not ( n14711 , n13314 );
and ( n14712 , n14711 , n13276 );
xor ( n14713 , n13276 , n13085 );
and ( n14714 , n14672 , n14673 );
xor ( n14715 , n14713 , n14714 );
and ( n14716 , n14715 , n13314 );
or ( n14717 , n14712 , n14716 );
and ( n14718 , n14717 , n5290 );
not ( n14719 , n13642 );
and ( n14720 , n14719 , n13604 );
xor ( n14721 , n13604 , n13413 );
and ( n14722 , n14680 , n14681 );
xor ( n14723 , n14721 , n14722 );
and ( n14724 , n14723 , n13642 );
or ( n14725 , n14720 , n14724 );
and ( n14726 , n14725 , n5288 );
and ( n14727 , n5606 , n5153 );
and ( n14728 , n2320 , n5155 );
or ( n14729 , n14718 , n14726 , n14727 , n14728 );
and ( n14730 , n14729 , n13663 );
or ( n14731 , n14710 , n14730 );
and ( n14732 , n14709 , n14731 );
and ( n14733 , n2424 , n3259 );
or ( n14734 , n14732 , n14733 );
and ( n14735 , n14708 , n14734 );
and ( n14736 , n14729 , n3066 );
or ( n14737 , n14735 , n14736 );
and ( n14738 , n14737 , n2422 );
buf ( n14739 , n3881 );
not ( n14740 , n14739 );
not ( n14741 , n14740 );
buf ( n14742 , n14741 );
and ( n14743 , n14742 , n2428 );
or ( n14744 , n14738 , n14743 );
buf ( n14745 , n14744 );
buf ( n14746 , n2424 );
buf ( n14747 , n2281 );
buf ( n14748 , n2280 );
not ( n14749 , n3066 );
not ( n14750 , n3259 );
and ( n14751 , n2318 , n12992 );
not ( n14752 , n13314 );
and ( n14753 , n14752 , n13288 );
xor ( n14754 , n13288 , n13085 );
and ( n14755 , n14713 , n14714 );
xor ( n14756 , n14754 , n14755 );
and ( n14757 , n14756 , n13314 );
or ( n14758 , n14753 , n14757 );
and ( n14759 , n14758 , n5290 );
not ( n14760 , n13642 );
and ( n14761 , n14760 , n13616 );
xor ( n14762 , n13616 , n13413 );
and ( n14763 , n14721 , n14722 );
xor ( n14764 , n14762 , n14763 );
and ( n14765 , n14764 , n13642 );
or ( n14766 , n14761 , n14765 );
and ( n14767 , n14766 , n5288 );
and ( n14768 , n5596 , n5153 );
and ( n14769 , n2318 , n5155 );
or ( n14770 , n14759 , n14767 , n14768 , n14769 );
and ( n14771 , n14770 , n13663 );
or ( n14772 , n14751 , n14771 );
and ( n14773 , n14750 , n14772 );
and ( n14774 , n2424 , n3259 );
or ( n14775 , n14773 , n14774 );
and ( n14776 , n14749 , n14775 );
and ( n14777 , n14770 , n3066 );
or ( n14778 , n14776 , n14777 );
and ( n14779 , n14778 , n2422 );
buf ( n14780 , n3876 );
not ( n14781 , n14780 );
not ( n14782 , n14781 );
buf ( n14783 , n14782 );
and ( n14784 , n14783 , n2428 );
or ( n14785 , n14779 , n14784 );
buf ( n14786 , n14785 );
buf ( n14787 , n2424 );
buf ( n14788 , n2281 );
buf ( n14789 , n2280 );
not ( n14790 , n3066 );
not ( n14791 , n3259 );
and ( n14792 , n2316 , n12992 );
not ( n14793 , n13314 );
and ( n14794 , n14793 , n13300 );
xor ( n14795 , n13300 , n13085 );
and ( n14796 , n14754 , n14755 );
xor ( n14797 , n14795 , n14796 );
and ( n14798 , n14797 , n13314 );
or ( n14799 , n14794 , n14798 );
and ( n14800 , n14799 , n5290 );
not ( n14801 , n13642 );
and ( n14802 , n14801 , n13628 );
xor ( n14803 , n13628 , n13413 );
and ( n14804 , n14762 , n14763 );
xor ( n14805 , n14803 , n14804 );
and ( n14806 , n14805 , n13642 );
or ( n14807 , n14802 , n14806 );
and ( n14808 , n14807 , n5288 );
and ( n14809 , n5586 , n5153 );
and ( n14810 , n2316 , n5155 );
or ( n14811 , n14800 , n14808 , n14809 , n14810 );
and ( n14812 , n14811 , n13663 );
or ( n14813 , n14792 , n14812 );
and ( n14814 , n14791 , n14813 );
and ( n14815 , n2424 , n3259 );
or ( n14816 , n14814 , n14815 );
and ( n14817 , n14790 , n14816 );
and ( n14818 , n14811 , n3066 );
or ( n14819 , n14817 , n14818 );
and ( n14820 , n14819 , n2422 );
buf ( n14821 , n3871 );
not ( n14822 , n14821 );
not ( n14823 , n14822 );
buf ( n14824 , n14823 );
and ( n14825 , n14824 , n2428 );
or ( n14826 , n14820 , n14825 );
buf ( n14827 , n14826 );
buf ( n14828 , n2424 );
buf ( n14829 , n2281 );
buf ( n14830 , n2280 );
not ( n14831 , n3066 );
not ( n14832 , n3259 );
and ( n14833 , n2314 , n12992 );
not ( n14834 , n13314 );
and ( n14835 , n14834 , n13312 );
xor ( n14836 , n13312 , n13085 );
and ( n14837 , n14795 , n14796 );
xor ( n14838 , n14836 , n14837 );
and ( n14839 , n14838 , n13314 );
or ( n14840 , n14835 , n14839 );
and ( n14841 , n14840 , n5290 );
not ( n14842 , n13642 );
and ( n14843 , n14842 , n13640 );
xor ( n14844 , n13640 , n13413 );
and ( n14845 , n14803 , n14804 );
xor ( n14846 , n14844 , n14845 );
and ( n14847 , n14846 , n13642 );
or ( n14848 , n14843 , n14847 );
and ( n14849 , n14848 , n5288 );
and ( n14850 , n5576 , n5153 );
and ( n14851 , n2314 , n5155 );
or ( n14852 , n14841 , n14849 , n14850 , n14851 );
and ( n14853 , n14852 , n13663 );
or ( n14854 , n14833 , n14853 );
and ( n14855 , n14832 , n14854 );
and ( n14856 , n2424 , n3259 );
or ( n14857 , n14855 , n14856 );
and ( n14858 , n14831 , n14857 );
and ( n14859 , n14852 , n3066 );
or ( n14860 , n14858 , n14859 );
and ( n14861 , n14860 , n2422 );
buf ( n14862 , n3866 );
not ( n14863 , n14862 );
not ( n14864 , n14863 );
buf ( n14865 , n14864 );
and ( n14866 , n14865 , n2428 );
or ( n14867 , n14861 , n14866 );
buf ( n14868 , n14867 );
buf ( n14869 , n2424 );
buf ( n14870 , n2281 );
buf ( n14871 , n2280 );
not ( n14872 , n3259 );
or ( n14873 , n3066 , n14872 );
not ( n14874 , n14873 );
and ( n14875 , n14874 , n3795 );
and ( n14876 , n2416 , n14873 );
or ( n14877 , n14875 , n14876 );
and ( n14878 , n14877 , n2422 );
and ( n14879 , n2416 , n2428 );
or ( n14880 , n14878 , n14879 );
buf ( n14881 , n14880 );
buf ( n14882 , n2424 );
buf ( n14883 , n2281 );
buf ( n14884 , n2280 );
not ( n14885 , n14873 );
and ( n14886 , n14885 , n3785 );
and ( n14887 , n2414 , n14873 );
or ( n14888 , n14886 , n14887 );
and ( n14889 , n14888 , n2422 );
and ( n14890 , n2414 , n2428 );
or ( n14891 , n14889 , n14890 );
buf ( n14892 , n14891 );
buf ( n14893 , n2424 );
buf ( n14894 , n2281 );
buf ( n14895 , n2280 );
not ( n14896 , n14873 );
and ( n14897 , n14896 , n4258 );
and ( n14898 , n2412 , n14873 );
or ( n14899 , n14897 , n14898 );
and ( n14900 , n14899 , n2422 );
and ( n14901 , n2412 , n2428 );
or ( n14902 , n14900 , n14901 );
buf ( n14903 , n14902 );
buf ( n14904 , n2424 );
buf ( n14905 , n2281 );
buf ( n14906 , n2280 );
not ( n14907 , n14873 );
and ( n14908 , n14907 , n4244 );
and ( n14909 , n2410 , n14873 );
or ( n14910 , n14908 , n14909 );
and ( n14911 , n14910 , n2422 );
and ( n14912 , n2410 , n2428 );
or ( n14913 , n14911 , n14912 );
buf ( n14914 , n14913 );
buf ( n14915 , n2424 );
buf ( n14916 , n2281 );
buf ( n14917 , n2280 );
not ( n14918 , n14873 );
and ( n14919 , n14918 , n4234 );
and ( n14920 , n2408 , n14873 );
or ( n14921 , n14919 , n14920 );
and ( n14922 , n14921 , n2422 );
and ( n14923 , n2408 , n2428 );
or ( n14924 , n14922 , n14923 );
buf ( n14925 , n14924 );
buf ( n14926 , n2424 );
buf ( n14927 , n2281 );
buf ( n14928 , n2280 );
not ( n14929 , n14873 );
and ( n14930 , n14929 , n4224 );
and ( n14931 , n2406 , n14873 );
or ( n14932 , n14930 , n14931 );
and ( n14933 , n14932 , n2422 );
and ( n14934 , n2406 , n2428 );
or ( n14935 , n14933 , n14934 );
buf ( n14936 , n14935 );
buf ( n14937 , n2424 );
buf ( n14938 , n2281 );
buf ( n14939 , n2280 );
not ( n14940 , n14873 );
and ( n14941 , n14940 , n4214 );
and ( n14942 , n2404 , n14873 );
or ( n14943 , n14941 , n14942 );
and ( n14944 , n14943 , n2422 );
and ( n14945 , n2404 , n2428 );
or ( n14946 , n14944 , n14945 );
buf ( n14947 , n14946 );
buf ( n14948 , n2424 );
buf ( n14949 , n2281 );
buf ( n14950 , n2280 );
not ( n14951 , n14873 );
and ( n14952 , n14951 , n4204 );
and ( n14953 , n2402 , n14873 );
or ( n14954 , n14952 , n14953 );
and ( n14955 , n14954 , n2422 );
and ( n14956 , n2402 , n2428 );
or ( n14957 , n14955 , n14956 );
buf ( n14958 , n14957 );
buf ( n14959 , n2424 );
buf ( n14960 , n2281 );
buf ( n14961 , n2280 );
not ( n14962 , n14873 );
and ( n14963 , n14962 , n4194 );
and ( n14964 , n2400 , n14873 );
or ( n14965 , n14963 , n14964 );
and ( n14966 , n14965 , n2422 );
and ( n14967 , n2400 , n2428 );
or ( n14968 , n14966 , n14967 );
buf ( n14969 , n14968 );
buf ( n14970 , n2424 );
buf ( n14971 , n2281 );
buf ( n14972 , n2280 );
not ( n14973 , n14873 );
and ( n14974 , n14973 , n4184 );
and ( n14975 , n2398 , n14873 );
or ( n14976 , n14974 , n14975 );
and ( n14977 , n14976 , n2422 );
and ( n14978 , n2398 , n2428 );
or ( n14979 , n14977 , n14978 );
buf ( n14980 , n14979 );
buf ( n14981 , n2424 );
buf ( n14982 , n2281 );
buf ( n14983 , n2280 );
not ( n14984 , n14873 );
and ( n14985 , n14984 , n4174 );
and ( n14986 , n2396 , n14873 );
or ( n14987 , n14985 , n14986 );
and ( n14988 , n14987 , n2422 );
and ( n14989 , n2396 , n2428 );
or ( n14990 , n14988 , n14989 );
buf ( n14991 , n14990 );
buf ( n14992 , n2424 );
buf ( n14993 , n2281 );
buf ( n14994 , n2280 );
not ( n14995 , n14873 );
and ( n14996 , n14995 , n4164 );
and ( n14997 , n2394 , n14873 );
or ( n14998 , n14996 , n14997 );
and ( n14999 , n14998 , n2422 );
and ( n15000 , n2394 , n2428 );
or ( n15001 , n14999 , n15000 );
buf ( n15002 , n15001 );
buf ( n15003 , n2424 );
buf ( n15004 , n2281 );
buf ( n15005 , n2280 );
not ( n15006 , n14873 );
and ( n15007 , n15006 , n4154 );
and ( n15008 , n2392 , n14873 );
or ( n15009 , n15007 , n15008 );
and ( n15010 , n15009 , n2422 );
and ( n15011 , n2392 , n2428 );
or ( n15012 , n15010 , n15011 );
buf ( n15013 , n15012 );
buf ( n15014 , n2424 );
buf ( n15015 , n2281 );
buf ( n15016 , n2280 );
not ( n15017 , n14873 );
and ( n15018 , n15017 , n4144 );
and ( n15019 , n2390 , n14873 );
or ( n15020 , n15018 , n15019 );
and ( n15021 , n15020 , n2422 );
and ( n15022 , n2390 , n2428 );
or ( n15023 , n15021 , n15022 );
buf ( n15024 , n15023 );
buf ( n15025 , n2424 );
buf ( n15026 , n2281 );
buf ( n15027 , n2280 );
not ( n15028 , n14873 );
and ( n15029 , n15028 , n4134 );
and ( n15030 , n2388 , n14873 );
or ( n15031 , n15029 , n15030 );
and ( n15032 , n15031 , n2422 );
and ( n15033 , n2388 , n2428 );
or ( n15034 , n15032 , n15033 );
buf ( n15035 , n15034 );
buf ( n15036 , n2424 );
buf ( n15037 , n2281 );
buf ( n15038 , n2280 );
not ( n15039 , n14873 );
and ( n15040 , n15039 , n4124 );
and ( n15041 , n2386 , n14873 );
or ( n15042 , n15040 , n15041 );
and ( n15043 , n15042 , n2422 );
and ( n15044 , n2386 , n2428 );
or ( n15045 , n15043 , n15044 );
buf ( n15046 , n15045 );
buf ( n15047 , n2424 );
buf ( n15048 , n2281 );
buf ( n15049 , n2280 );
not ( n15050 , n14873 );
and ( n15051 , n15050 , n4114 );
and ( n15052 , n2384 , n14873 );
or ( n15053 , n15051 , n15052 );
and ( n15054 , n15053 , n2422 );
and ( n15055 , n2384 , n2428 );
or ( n15056 , n15054 , n15055 );
buf ( n15057 , n15056 );
buf ( n15058 , n2424 );
buf ( n15059 , n2281 );
buf ( n15060 , n2280 );
not ( n15061 , n14873 );
and ( n15062 , n15061 , n4104 );
and ( n15063 , n2382 , n14873 );
or ( n15064 , n15062 , n15063 );
and ( n15065 , n15064 , n2422 );
and ( n15066 , n2382 , n2428 );
or ( n15067 , n15065 , n15066 );
buf ( n15068 , n15067 );
buf ( n15069 , n2424 );
buf ( n15070 , n2281 );
buf ( n15071 , n2280 );
not ( n15072 , n14873 );
and ( n15073 , n15072 , n4094 );
and ( n15074 , n2380 , n14873 );
or ( n15075 , n15073 , n15074 );
and ( n15076 , n15075 , n2422 );
and ( n15077 , n2380 , n2428 );
or ( n15078 , n15076 , n15077 );
buf ( n15079 , n15078 );
buf ( n15080 , n2424 );
buf ( n15081 , n2281 );
buf ( n15082 , n2280 );
not ( n15083 , n14873 );
and ( n15084 , n15083 , n4084 );
and ( n15085 , n2378 , n14873 );
or ( n15086 , n15084 , n15085 );
and ( n15087 , n15086 , n2422 );
and ( n15088 , n2378 , n2428 );
or ( n15089 , n15087 , n15088 );
buf ( n15090 , n15089 );
buf ( n15091 , n2424 );
buf ( n15092 , n2281 );
buf ( n15093 , n2280 );
not ( n15094 , n14873 );
and ( n15095 , n15094 , n4074 );
and ( n15096 , n2376 , n14873 );
or ( n15097 , n15095 , n15096 );
and ( n15098 , n15097 , n2422 );
and ( n15099 , n2376 , n2428 );
or ( n15100 , n15098 , n15099 );
buf ( n15101 , n15100 );
buf ( n15102 , n2424 );
buf ( n15103 , n2281 );
buf ( n15104 , n2280 );
not ( n15105 , n14873 );
and ( n15106 , n15105 , n4064 );
and ( n15107 , n2374 , n14873 );
or ( n15108 , n15106 , n15107 );
and ( n15109 , n15108 , n2422 );
and ( n15110 , n2374 , n2428 );
or ( n15111 , n15109 , n15110 );
buf ( n15112 , n15111 );
buf ( n15113 , n2424 );
buf ( n15114 , n2281 );
buf ( n15115 , n2280 );
not ( n15116 , n14873 );
and ( n15117 , n15116 , n4054 );
and ( n15118 , n2372 , n14873 );
or ( n15119 , n15117 , n15118 );
and ( n15120 , n15119 , n2422 );
and ( n15121 , n2372 , n2428 );
or ( n15122 , n15120 , n15121 );
buf ( n15123 , n15122 );
buf ( n15124 , n2424 );
buf ( n15125 , n2281 );
buf ( n15126 , n2280 );
not ( n15127 , n14873 );
and ( n15128 , n15127 , n4044 );
and ( n15129 , n2370 , n14873 );
or ( n15130 , n15128 , n15129 );
and ( n15131 , n15130 , n2422 );
and ( n15132 , n2370 , n2428 );
or ( n15133 , n15131 , n15132 );
buf ( n15134 , n15133 );
buf ( n15135 , n2424 );
buf ( n15136 , n2281 );
buf ( n15137 , n2280 );
not ( n15138 , n14873 );
and ( n15139 , n15138 , n4034 );
and ( n15140 , n2368 , n14873 );
or ( n15141 , n15139 , n15140 );
and ( n15142 , n15141 , n2422 );
and ( n15143 , n2368 , n2428 );
or ( n15144 , n15142 , n15143 );
buf ( n15145 , n15144 );
buf ( n15146 , n2424 );
buf ( n15147 , n2281 );
buf ( n15148 , n2280 );
not ( n15149 , n14873 );
and ( n15150 , n15149 , n4024 );
and ( n15151 , n2366 , n14873 );
or ( n15152 , n15150 , n15151 );
and ( n15153 , n15152 , n2422 );
and ( n15154 , n2366 , n2428 );
or ( n15155 , n15153 , n15154 );
buf ( n15156 , n15155 );
buf ( n15157 , n2424 );
buf ( n15158 , n2281 );
buf ( n15159 , n2280 );
not ( n15160 , n14873 );
and ( n15161 , n15160 , n4014 );
and ( n15162 , n2364 , n14873 );
or ( n15163 , n15161 , n15162 );
and ( n15164 , n15163 , n2422 );
and ( n15165 , n2364 , n2428 );
or ( n15166 , n15164 , n15165 );
buf ( n15167 , n15166 );
buf ( n15168 , n2424 );
buf ( n15169 , n2281 );
buf ( n15170 , n2280 );
not ( n15171 , n14873 );
and ( n15172 , n15171 , n4004 );
and ( n15173 , n2362 , n14873 );
or ( n15174 , n15172 , n15173 );
and ( n15175 , n15174 , n2422 );
and ( n15176 , n2362 , n2428 );
or ( n15177 , n15175 , n15176 );
buf ( n15178 , n15177 );
buf ( n15179 , n2424 );
buf ( n15180 , n2281 );
buf ( n15181 , n2280 );
not ( n15182 , n14873 );
and ( n15183 , n15182 , n3994 );
and ( n15184 , n2360 , n14873 );
or ( n15185 , n15183 , n15184 );
and ( n15186 , n15185 , n2422 );
and ( n15187 , n2360 , n2428 );
or ( n15188 , n15186 , n15187 );
buf ( n15189 , n15188 );
buf ( n15190 , n2424 );
buf ( n15191 , n2281 );
buf ( n15192 , n2280 );
not ( n15193 , n14873 );
and ( n15194 , n15193 , n3984 );
and ( n15195 , n2358 , n14873 );
or ( n15196 , n15194 , n15195 );
and ( n15197 , n15196 , n2422 );
and ( n15198 , n2358 , n2428 );
or ( n15199 , n15197 , n15198 );
buf ( n15200 , n15199 );
buf ( n15201 , n2424 );
buf ( n15202 , n2281 );
buf ( n15203 , n2280 );
not ( n15204 , n14873 );
and ( n15205 , n15204 , n3819 );
and ( n15206 , n2356 , n14873 );
or ( n15207 , n15205 , n15206 );
and ( n15208 , n15207 , n2422 );
and ( n15209 , n2356 , n2428 );
or ( n15210 , n15208 , n15209 );
buf ( n15211 , n15210 );
buf ( n15212 , n2424 );
buf ( n15213 , n2281 );
buf ( n15214 , n2280 );
not ( n15215 , n14873 );
and ( n15216 , n15215 , n3770 );
and ( n15217 , n2354 , n14873 );
or ( n15218 , n15216 , n15217 );
and ( n15219 , n15218 , n2422 );
and ( n15220 , n2354 , n2428 );
or ( n15221 , n15219 , n15220 );
buf ( n15222 , n15221 );
buf ( n15223 , n2424 );
buf ( n15224 , n2281 );
buf ( n15225 , n2280 );
not ( n15226 , n3066 );
and ( n15227 , n5291 , n13663 );
not ( n15228 , n3259 );
and ( n15229 , n15227 , n15228 );
and ( n15230 , n15226 , n15229 );
and ( n15231 , n5291 , n3066 );
or ( n15232 , n15230 , n15231 );
and ( n15233 , n15232 , n2422 );
or ( n15234 , n15233 , n2428 );
buf ( n15235 , n15234 );
buf ( n15236 , n2424 );
buf ( n15237 , n2281 );
buf ( n15238 , n2280 );
not ( n15239 , n14873 );
and ( n15240 , n3259 , n15239 );
and ( n15241 , n15240 , n2422 );
buf ( n15242 , n15241 );
endmodule

