//
// Conformal-LEC Version 15.10-d003 ( 23-Apr-2015) ( 64 bit executable)
//
module top ( 
    n0 , 
    n1 , 
    n2 , 
    n3 , 
    n4 , 
    n5 , 
    n6 , 
    n7 , 
    n8 , 
    n9 , 
    n10 , 
    n11 , 
    n12 , 
    n13 , 
    n14 , 
    n15 , 
    n16 , 
    n17 , 
    n18 , 
    n19 , 
    n20 , 
    n21 , 
    n22 , 
    n23 , 
    n24 , 
    n25 , 
    n26 , 
    n27 , 
    n28 , 
    n29 , 
    n30 , 
    n31 , 
    n32 , 
    n33 , 
    n34 , 
    n35 , 
    n36 , 
    n37 , 
    n38 , 
    n39 , 
    n40 , 
    n41 , 
    n42 , 
    n43 , 
    n44 , 
    n45 , 
    n46 , 
    n47 , 
    n48 , 
    n49 , 
    n50 , 
    n51 , 
    n52 , 
    n53 , 
    n54 , 
    n55 , 
    n56 , 
    n57 , 
    n58 , 
    n59 , 
    n60 , 
    n61 , 
    n62 , 
    n63 , 
    n64 , 
    n65 , 
    n66 , 
    n67 , 
    n68 , 
    n69 , 
    n70 , 
    n71 , 
    n72 , 
    n73 , 
    n74 , 
    n75 , 
    n76 , 
    n77 , 
    n78 , 
    n79 , 
    n80 , 
    n81 , 
    n82 , 
    n83 , 
    n84 , 
    n85 , 
    n86 , 
    n87 , 
    n88 , 
    n89 , 
    n90 , 
    n91 , 
    n92 , 
    n93 , 
    n94 , 
    n95 , 
    n96 , 
    n97 , 
    n98 , 
    n99 , 
    n100 , 
    n101 , 
    n102 , 
    n103 , 
    n104 , 
    n105 , 
    n106 , 
    n107 , 
    n108 , 
    n109 , 
    n110 , 
    n111 , 
    n112 , 
    n113 , 
    n114 , 
    n115 , 
    n116 , 
    n117 , 
    n118 , 
    n119 , 
    n120 , 
    n121 , 
    n122 , 
    n123 , 
    n124 , 
    n125 , 
    n126 , 
    n127 , 
    n128 , 
    n129 , 
    n130 , 
    n131 , 
    n132 , 
    n133 , 
    n134 , 
    n135 , 
    n136 , 
    n137 , 
    n138 , 
    n139 , 
    n140 , 
    n141 , 
    n142 , 
    n143 , 
    n144 , 
    n145 , 
    n146 , 
    n147 , 
    n148 , 
    n149 , 
    n150 , 
    n151 , 
    n152 , 
    n153 , 
    n154 , 
    n155 , 
    n156 , 
    n157 , 
    n158 , 
    n159 , 
    n160 , 
    n161 , 
    n162 , 
    n163 , 
    n164 , 
    n165 , 
    n166 , 
    n167 , 
    n168 , 
    n169 , 
    n170 , 
    n171 , 
    n172 , 
    n173 , 
    n174 , 
    n175 , 
    n176 , 
    n177 , 
    n178 , 
    n179 , 
    n180 , 
    n181 , 
    n182 , 
    n183 , 
    n184 , 
    n185 , 
    n186 , 
    n187 , 
    n188 , 
    n189 , 
    n190 , 
    n191 , 
    n192 , 
    n193 , 
    n194 , 
    n195 , 
    n196 , 
    n197 , 
    n198 , 
    n199 , 
    n200 , 
    n201 , 
    n202 , 
    n203 , 
    n204 , 
    n205 , 
    n206 , 
    n207 , 
    n208 , 
    n209 , 
    n210 , 
    n211 , 
    n212 , 
    n213 , 
    n214 , 
    n215 , 
    n216 , 
    n217 , 
    n218 , 
    n219 , 
    n220 , 
    n221 , 
    n222 , 
    n223 , 
    n224 , 
    n225 , 
    n226 , 
    n227 , 
    n228 , 
    n229 , 
    n230 , 
    n231 , 
    n232 , 
    n233 , 
    n234 , 
    n235 , 
    n236 , 
    n237 , 
    n238 , 
    n239 , 
    n240 , 
    n241 , 
    n242 , 
    n243 , 
    n244 , 
    n245 , 
    n246 , 
    n247 , 
    n248 , 
    n249 , 
    n250 , 
    n251 , 
    n252 , 
    n253 , 
    n254 , 
    n255 , 
    n256 , 
    n257 , 
    n258 , 
    n259 , 
    n260 , 
    n261 , 
    n262 , 
    n263 , 
    n264 , 
    n265 , 
    n266 , 
    n267 , 
    n268 , 
    n269 , 
    n270 , 
    n271 , 
    n272 , 
    n273 , 
    n274 , 
    n275 , 
    n276 , 
    n277 , 
    n278 , 
    n279 , 
    n280 , 
    n281 , 
    n282 , 
    n283 , 
    n284 , 
    n285 , 
    n286 , 
    n287 , 
    n288 , 
    n289 , 
    n290 , 
    n291 , 
    n292 , 
    n293 , 
    n294 , 
    n295 , 
    n296 , 
    n297 , 
    n298 , 
    n299 , 
    n300 , 
    n301 , 
    n302 , 
    n303 , 
    n304 , 
    n305 , 
    n306 , 
    n307 , 
    n308 , 
    n309 , 
    n310 , 
    n311 , 
    n312 , 
    n313 , 
    n314 , 
    n315 , 
    n316 , 
    n317 , 
    n318 , 
    n319 , 
    n320 , 
    n321 , 
    n322 , 
    n323 , 
    n324 , 
    n325 , 
    n326 , 
    n327 , 
    n328 , 
    n329 , 
    n330 , 
    n331 , 
    n332 , 
    n333 , 
    n334 , 
    n335 , 
    n336 , 
    n337 , 
    n338 , 
    n339 , 
    n340 , 
    n341 , 
    n342 , 
    n343 , 
    n344 , 
    n345 , 
    n346 , 
    n347 , 
    n348 , 
    n349 , 
    n350 , 
    n351 , 
    n352 , 
    n353 , 
    n354 , 
    n355 , 
    n356 , 
    n357 , 
    n358 , 
    n359 , 
    n360 , 
    n361 , 
    n362 , 
    n363 , 
    n364 , 
    n365 , 
    n366 , 
    n367 , 
    n368 , 
    n369 , 
    n370 , 
    n371 , 
    n372 , 
    n373 , 
    n374 , 
    n375 , 
    n376 , 
    n377 , 
    n378 , 
    n379 , 
    n380 , 
    n381 , 
    n382 , 
    n383 , 
    n384 , 
    n385 , 
    n386 , 
    n387 , 
    n388 , 
    n389 , 
    n390 , 
    n391 , 
    n392 , 
    n393 , 
    n394 , 
    n395 , 
    n396 , 
    n397 , 
    n398 , 
    n399 , 
    n400 , 
    n401 , 
    n402 , 
    n403 , 
    n404 , 
    n405 , 
    n406 , 
    n407 , 
    n408 , 
    n409 , 
    n410 , 
    n411 , 
    n412 , 
    n413 , 
    n414 , 
    n415 , 
    n416 , 
    n417 , 
    n418 , 
    n419 , 
    n420 , 
    n421 , 
    n422 , 
    n423 , 
    n424 , 
    n425 , 
    n426 , 
    n427 , 
    n428 , 
    n429 , 
    n430 , 
    n431 , 
    n432 , 
    n433 , 
    n434 , 
    n435 , 
    n436 , 
    n437 , 
    n438 , 
    n439 , 
    n440 , 
    n441 , 
    n442 , 
    n443 , 
    n444 , 
    n445 , 
    n446 , 
    n447 , 
    n448 , 
    n449 , 
    n450 , 
    n451 , 
    n452 , 
    n453 , 
    n454 , 
    n455 , 
    n456 , 
    n457 , 
    n458 , 
    n459 , 
    n460 , 
    n461 , 
    n462 , 
    n463 , 
    n464 , 
    n465 , 
    n466 , 
    n467 , 
    n468 , 
    n469 , 
    n470 , 
    n471 , 
    n472 , 
    n473 , 
    n474 , 
    n475 , 
    n476 , 
    n477 , 
    n478 , 
    n479 , 
    n480 , 
    n481 , 
    n482 , 
    n483 , 
    n484 , 
    n485 , 
    n486 , 
    n487 , 
    n488 , 
    n489 , 
    n490 , 
    n491 , 
    n492 , 
    n493 , 
    n494 , 
    n495 , 
    n496 , 
    n497 , 
    n498 , 
    n499 , 
    n500 , 
    n501 , 
    n502 , 
    n503 , 
    n504 , 
    n505 , 
    n506 , 
    n507 , 
    n508 , 
    n509 , 
    n510 , 
    n511 , 
    n512 , 
    n513 , 
    n514 , 
    n515 , 
    n516 , 
    n517 , 
    n518 , 
    n519 , 
    n520 , 
    n521 , 
    n522 , 
    n523 , 
    n524 , 
    n525 , 
    n526 , 
    n527 , 
    n528 , 
    n529 , 
    n530 , 
    n531 , 
    n532 , 
    n533 , 
    n534 , 
    n535 , 
    n536 , 
    n537 , 
    n538 , 
    n539 , 
    n540 , 
    n541 , 
    n542 , 
    n543 , 
    n544 , 
    n545 , 
    n546 , 
    n547 , 
    n548 , 
    n549 , 
    n550 , 
    n551 , 
    n552 , 
    n553 , 
    n554 , 
    n555 , 
    n556 , 
    n557 , 
    n558 , 
    n559 , 
    n560 , 
    n561 , 
    n562 , 
    n563 , 
    n564 , 
    n565 , 
    n566 , 
    n567 , 
    n568 , 
    n569 , 
    n570 , 
    n571 , 
    n572 , 
    n573 , 
    n574 , 
    n575 , 
    n576 , 
    n577 , 
    n578 , 
    n579 , 
    n580 , 
    n581 , 
    n582 , 
    n583 , 
    n584 , 
    n585 , 
    n586 , 
    n587 , 
    n588 , 
    n589 , 
    n590 , 
    n591 , 
    n592 , 
    n593 , 
    n594 , 
    n595 , 
    n596 , 
    n597 , 
    n598 , 
    n599 , 
    n600 , 
    n601 , 
    n602 , 
    n603 , 
    n604 , 
    n605 , 
    n606 , 
    n607 , 
    n608 , 
    n609 , 
    n610 , 
    n611 , 
    n612 , 
    n613 , 
    n614 , 
    n615 , 
    n616 , 
    n617 , 
    n618 , 
    n619 , 
    n620 , 
    n621 , 
    n622 , 
    n623 , 
    n624 , 
    n625 , 
    n626 , 
    n627 , 
    n628 , 
    n629 , 
    n630 , 
    n631 , 
    n632 , 
    n633 , 
    n634 , 
    n635 , 
    n636 , 
    n637 , 
    n638 , 
    n639 , 
    n640 , 
    n641 , 
    n642 , 
    n643 , 
    n644 , 
    n645 , 
    n646 , 
    n647 , 
    n648 , 
    n649 , 
    n650 , 
    n651 , 
    n652 , 
    n653 , 
    n654 , 
    n655 , 
    n656 , 
    n657 , 
    n658 , 
    n659 , 
    n660 , 
    n661 , 
    n662 , 
    n663 , 
    n664 , 
    n665 , 
    n666 , 
    n667 , 
    n668 , 
    n669 , 
    n670 , 
    n671 , 
    n672 , 
    n673 , 
    n674 , 
    n675 , 
    n676 , 
    n677 , 
    n678 , 
    n679 , 
    n680 , 
    n681 , 
    n682 , 
    n683 , 
    n684 , 
    n685 , 
    n686 , 
    n687 , 
    n688 , 
    n689 , 
    n690 , 
    n691 , 
    n692 , 
    n693 , 
    n694 , 
    n695 , 
    n696 , 
    n697 , 
    n698 , 
    n699 , 
    n700 , 
    n701 , 
    n702 , 
    n703 , 
    n704 , 
    n705 , 
    n706 , 
    n707 , 
    n708 , 
    n709 , 
    n710 , 
    n711 , 
    n712 , 
    n713 , 
    n714 , 
    n715 , 
    n716 , 
    n717 , 
    n718 , 
    n719 , 
    n720 , 
    n721 , 
    n722 , 
    n723 , 
    n724 , 
    n725 , 
    n726 , 
    n727 , 
    n728 , 
    n729 , 
    n730 , 
    n731 , 
    n732 , 
    n733 , 
    n734 , 
    n735 , 
    n736 , 
    n737 , 
    n738 , 
    n739 , 
    n740 , 
    n741 , 
    n742 , 
    n743 , 
    n744 , 
    n745 , 
    n746 , 
    n747 , 
    n748 , 
    n749 , 
    n750 , 
    n751 , 
    n752 , 
    n753 , 
    n754 , 
    n755 , 
    n756 , 
    n757 , 
    n758 , 
    n759 , 
    n760 , 
    n761 , 
    n762 , 
    n763 , 
    n764 , 
    n765 , 
    n766 , 
    n767 , 
    n768 , 
    n769 , 
    n770 , 
    n771 , 
    n772 , 
    n773 , 
    n774 , 
    n775 , 
    n776 , 
    n777 , 
    n778 , 
    n779 , 
    n780 , 
    n781 , 
    n782 , 
    n783 , 
    n784 , 
    n785 , 
    n786 , 
    n787 , 
    n788 , 
    n789 , 
    n790 , 
    n791 , 
    n792 , 
    n793 , 
    n794 , 
    n795 , 
    n796 , 
    n797 , 
    n798 , 
    n799 , 
    n800 , 
    n801 , 
    n802 , 
    n803 , 
    n804 , 
    n805 , 
    n806 , 
    n807 , 
    n808 , 
    n809 , 
    n810 , 
    n811 , 
    n812 , 
    n813 , 
    n814 , 
    n815 , 
    n816 , 
    n817 , 
    n818 , 
    n819 , 
    n820 , 
    n821 , 
    n822 , 
    n823 , 
    n824 , 
    n825 , 
    n826 , 
    n827 , 
    n828 , 
    n829 , 
    n830 , 
    n831 , 
    n832 , 
    n833 , 
    n834 , 
    n835 , 
    n836 , 
    n837 , 
    n838 , 
    n839 , 
    n840 , 
    n841 , 
    n842 , 
    n843 , 
    n844 , 
    n845 , 
    n846 , 
    n847 , 
    n848 , 
    n849 , 
    n850 , 
    n851 , 
    n852 , 
    n853 , 
    n854 , 
    n855 , 
    n856 , 
    n857 , 
    n858 , 
    n859 , 
    n860 , 
    n861 , 
    n862 , 
    n863 , 
    n864 , 
    n865 , 
    n866 , 
    n867 , 
    n868 , 
    n869 , 
    n870 , 
    n871 , 
    n872 , 
    n873 , 
    n874 , 
    n875 , 
    n876 , 
    n877 , 
    n878 , 
    n879 , 
    n880 , 
    n881 , 
    n882 , 
    n883 , 
    n884 , 
    n885 , 
    n886 , 
    n887 , 
    n888 , 
    n889 , 
    n890 , 
    n891 , 
    n892 , 
    n893 , 
    n894 , 
    n895 , 
    n896 , 
    n897 , 
    n898 , 
    n899 , 
    n900 , 
    n901 , 
    n902 , 
    n903 , 
    n904 , 
    n905 , 
    n906 , 
    n907 , 
    n908 , 
    n909 , 
    n910 , 
    n911 , 
    n912 , 
    n913 , 
    n914 , 
    n915 , 
    n916 , 
    n917 , 
    n918 , 
    n919 , 
    n920 , 
    n921 , 
    n922 , 
    n923 , 
    n924 , 
    n925 , 
    n926 , 
    n927 , 
    n928 , 
    n929 , 
    n930 , 
    n931 , 
    n932 , 
    n933 , 
    n934 , 
    n935 , 
    n936 , 
    n937 , 
    n938 , 
    n939 , 
    n940 , 
    n941 , 
    n942 , 
    n943 , 
    n944 , 
    n945 , 
    n946 , 
    n947 , 
    n948 , 
    n949 , 
    n950 , 
    n951 , 
    n952 , 
    n953 , 
    n954 , 
    n955 , 
    n956 , 
    n957 , 
    n958 , 
    n959 , 
    n960 , 
    n961 , 
    n962 , 
    n963 , 
    n964 , 
    n965 , 
    n966 , 
    n967 , 
    n968 , 
    n969 , 
    n970 , 
    n971 , 
    n972 , 
    n973 , 
    n974 , 
    n975 , 
    n976 , 
    n977 , 
    n978 , 
    n979 , 
    n980 , 
    n981 , 
    n982 , 
    n983 , 
    n984 , 
    n985 , 
    n986 , 
    n987 , 
    n988 , 
    n989 , 
    n990 , 
    n991 , 
    n992 , 
    n993 , 
    n994 , 
    n995 , 
    n996 , 
    n997 , 
    n998 , 
    n999 , 
    n1000 , 
    n1001 , 
    n1002 , 
    n1003 , 
    n1004 , 
    n1005 , 
    n1006 , 
    n1007 , 
    n1008 , 
    n1009 , 
    n1010 , 
    n1011 , 
    n1012 , 
    n1013 , 
    n1014 , 
    n1015 , 
    n1016 , 
    n1017 , 
    n1018 , 
    n1019 , 
    n1020 , 
    n1021 , 
    n1022 , 
    n1023 , 
    n1024 , 
    n1025 , 
    n1026 , 
    n1027 , 
    n1028 , 
    n1029 , 
    n1030 , 
    n1031 , 
    n1032 , 
    n1033 , 
    n1034 , 
    n1035 , 
    n1036 , 
    n1037 , 
    n1038 , 
    n1039 , 
    n1040 , 
    n1041 , 
    n1042 , 
    n1043 , 
    n1044 , 
    n1045 , 
    n1046 , 
    n1047 , 
    n1048 , 
    n1049 , 
    n1050 , 
    n1051 , 
    n1052 , 
    n1053 , 
    n1054 , 
    n1055 , 
    n1056 , 
    n1057 , 
    n1058 , 
    n1059 , 
    n1060 , 
    n1061 , 
    n1062 , 
    n1063 , 
    n1064 , 
    n1065 , 
    n1066 , 
    n1067 , 
    n1068 , 
    n1069 , 
    n1070 , 
    n1071 , 
    n1072 , 
    n1073 , 
    n1074 , 
    n1075 , 
    n1076 , 
    n1077 , 
    n1078 , 
    n1079 , 
    n1080 , 
    n1081 , 
    n1082 , 
    n1083 , 
    n1084 , 
    n1085 , 
    n1086 , 
    n1087 , 
    n1088 , 
    n1089 , 
    n1090 , 
    n1091 , 
    n1092 , 
    n1093 , 
    n1094 , 
    n1095 , 
    n1096 , 
    n1097 , 
    n1098 , 
    n1099 , 
    n1100 , 
    n1101 , 
    n1102 , 
    n1103 , 
    n1104 , 
    n1105 , 
    n1106 , 
    n1107 , 
    n1108 , 
    n1109 , 
    n1110 , 
    n1111 , 
    n1112 , 
    n1113 , 
    n1114 , 
    n1115 , 
    n1116 , 
    n1117 , 
    n1118 , 
    n1119 , 
    n1120 , 
    n1121 , 
    n1122 , 
    n1123 , 
    n1124 , 
    n1125 , 
    n1126 , 
    n1127 , 
    n1128 , 
    n1129 , 
    n1130 , 
    n1131 , 
    n1132 , 
    n1133 , 
    n1134 , 
    n1135 , 
    n1136 , 
    n1137 , 
    n1138 , 
    n1139 , 
    n1140 , 
    n1141 , 
    n1142 , 
    n1143 , 
    n1144 , 
    n1145 , 
    n1146 , 
    n1147 , 
    n1148 , 
    n1149 , 
    n1150 , 
    n1151 , 
    n1152 , 
    n1153 , 
    n1154 , 
    n1155 , 
    n1156 , 
    n1157 , 
    n1158 , 
    n1159 , 
    n1160 , 
    n1161 , 
    n1162 , 
    n1163 , 
    n1164 , 
    n1165 , 
    n1166 , 
    n1167 , 
    n1168 , 
    n1169 , 
    n1170 , 
    n1171 , 
    n1172 , 
    n1173 , 
    n1174 , 
    n1175 , 
    n1176 , 
    n1177 , 
    n1178 , 
    n1179 , 
    n1180 , 
    n1181 , 
    n1182 , 
    n1183 , 
    n1184 , 
    n1185 , 
    n1186 , 
    n1187 , 
    n1188 , 
    n1189 , 
    n1190 , 
    n1191 , 
    n1192 , 
    n1193 , 
    n1194 , 
    n1195 , 
    n1196 , 
    n1197 , 
    n1198 , 
    n1199 , 
    n1200 , 
    n1201 , 
    n1202 , 
    n1203 , 
    n1204 , 
    n1205 , 
    n1206 , 
    n1207 , 
    n1208 , 
    n1209 , 
    n1210 , 
    n1211 , 
    n1212 , 
    n1213 , 
    n1214 , 
    n1215 , 
    n1216 , 
    n1217 , 
    n1218 , 
    n1219 , 
    n1220 , 
    n1221 , 
    n1222 , 
    n1223 , 
    n1224 , 
    n1225 , 
    n1226 , 
    n1227 , 
    n1228 , 
    n1229 , 
    n1230 , 
    n1231 , 
    n1232 , 
    n1233 , 
    n1234 , 
    n1235 , 
    n1236 , 
    n1237 , 
    n1238 , 
    n1239 , 
    n1240 , 
    n1241 , 
    n1242 , 
    n1243 , 
    n1244 , 
    n1245 , 
    n1246 , 
    n1247 , 
    n1248 , 
    n1249 , 
    n1250 , 
    n1251 , 
    n1252 , 
    n1253 , 
    n1254 , 
    n1255 , 
    n1256 , 
    n1257 , 
    n1258 , 
    n1259 , 
    n1260 , 
    n1261 , 
    n1262 , 
    n1263 , 
    n1264 , 
    n1265 , 
    n1266 , 
    n1267 , 
    n1268 , 
    n1269 , 
    n1270 , 
    n1271 , 
    n1272 , 
    n1273 , 
    n1274 , 
    n1275 , 
    n1276 , 
    n1277 , 
    n1278 , 
    n1279 , 
    n1280 , 
    n1281 , 
    n1282 , 
    n1283 , 
    n1284 , 
    n1285 , 
    n1286 , 
    n1287 , 
    n1288 , 
    n1289 , 
    n1290 , 
    n1291 , 
    n1292 , 
    n1293 , 
    n1294 , 
    n1295 , 
    n1296 , 
    n1297 , 
    n1298 , 
    n1299 , 
    n1300 , 
    n1301 , 
    n1302 , 
    n1303 , 
    n1304 , 
    n1305 , 
    n1306 , 
    n1307 , 
    n1308 , 
    n1309 , 
    n1310 , 
    n1311 , 
    n1312 , 
    n1313 , 
    n1314 , 
    n1315 , 
    n1316 , 
    n1317 , 
    n1318 , 
    n1319 , 
    n1320 , 
    n1321 , 
    n1322 , 
    n1323 , 
    n1324 , 
    n1325 , 
    n1326 , 
    n1327 , 
    n1328 , 
    n1329 , 
    n1330 , 
    n1331 , 
    n1332 , 
    n1333 , 
    n1334 , 
    n1335 , 
    n1336 , 
    n1337 , 
    n1338 , 
    n1339 , 
    n1340 , 
    n1341 , 
    n1342 , 
    n1343 , 
    n1344 , 
    n1345 , 
    n1346 , 
    n1347 , 
    n1348 , 
    n1349 , 
    n1350 , 
    n1351 , 
    n1352 , 
    n1353 , 
    n1354 , 
    n1355 , 
    n1356 , 
    n1357 , 
    n1358 , 
    n1359 , 
    n1360 , 
    n1361 , 
    n1362 , 
    n1363 , 
    n1364 , 
    n1365 , 
    n1366 , 
    n1367 , 
    n1368 , 
    n1369 , 
    n1370 , 
    n1371 , 
    n1372 , 
    n1373 , 
    n1374 , 
    n1375 , 
    n1376 , 
    n1377 , 
    n1378 , 
    n1379 , 
    n1380 , 
    n1381 , 
    n1382 , 
    n1383 , 
    n1384 , 
    n1385 , 
    n1386 , 
    n1387 , 
    n1388 , 
    n1389 , 
    n1390 , 
    n1391 , 
    n1392 , 
    n1393 , 
    n1394 , 
    n1395 , 
    n1396 , 
    n1397 , 
    n1398 , 
    n1399 , 
    n1400 , 
    n1401 , 
    n1402 , 
    n1403 , 
    n1404 , 
    n1405 , 
    n1406 , 
    n1407 , 
    n1408 , 
    n1409 , 
    n1410 , 
    n1411 , 
    n1412 , 
    n1413 , 
    n1414 , 
    n1415 , 
    n1416 , 
    n1417 , 
    n1418 , 
    n1419 , 
    n1420 , 
    n1421 , 
    n1422 , 
    n1423 , 
    n1424 , 
    n1425 , 
    n1426 , 
    n1427 , 
    n1428 , 
    n1429 , 
    n1430 , 
    n1431 , 
    n1432 , 
    n1433 , 
    n1434 , 
    n1435 , 
    n1436 , 
    n1437 , 
    n1438 , 
    n1439 , 
    n1440 , 
    n1441 , 
    n1442 , 
    n1443 , 
    n1444 , 
    n1445 , 
    n1446 , 
    n1447 , 
    n1448 , 
    n1449 , 
    n1450 , 
    n1451 , 
    n1452 , 
    n1453 , 
    n1454 , 
    n1455 , 
    n1456 , 
    n1457 , 
    n1458 , 
    n1459 , 
    n1460 , 
    n1461 , 
    n1462 , 
    n1463 , 
    n1464 , 
    n1465 , 
    n1466 , 
    n1467 , 
    n1468 , 
    n1469 , 
    n1470 , 
    n1471 , 
    n1472 , 
    n1473 , 
    n1474 , 
    n1475 , 
    n1476 , 
    n1477 , 
    n1478 , 
    n1479 , 
    n1480 , 
    n1481 , 
    n1482 , 
    n1483 , 
    n1484 , 
    n1485 , 
    n1486 , 
    n1487 , 
    n1488 , 
    n1489 , 
    n1490 , 
    n1491 , 
    n1492 , 
    n1493 , 
    n1494 , 
    n1495 , 
    n1496 , 
    n1497 , 
    n1498 , 
    n1499 , 
    n1500 , 
    n1501 , 
    n1502 , 
    n1503 , 
    n1504 , 
    n1505 , 
    n1506 , 
    n1507 , 
    n1508 , 
    n1509 , 
    n1510 , 
    n1511 , 
    n1512 , 
    n1513 , 
    n1514 , 
    n1515 , 
    n1516 , 
    n1517 , 
    n1518 , 
    n1519 , 
    n1520 , 
    n1521 , 
    n1522 , 
    n1523 , 
    n1524 , 
    n1525 , 
    n1526 , 
    n1527 , 
    n1528 , 
    n1529 , 
    n1530 , 
    n1531 , 
    n1532 , 
    n1533 , 
    n1534 , 
    n1535 , 
    n1536 , 
    n1537 , 
    n1538 , 
    n1539 , 
    n1540 , 
    n1541 , 
    n1542 , 
    n1543 , 
    n1544 , 
    n1545 , 
    n1546 , 
    n1547 , 
    n1548 , 
    n1549 , 
    n1550 , 
    n1551 , 
    n1552 , 
    n1553 , 
    n1554 , 
    n1555 , 
    n1556 , 
    n1557 , 
    n1558 , 
    n1559 , 
    n1560 , 
    n1561 , 
    n1562 , 
    n1563 , 
    n1564 , 
    n1565 , 
    n1566 , 
    n1567 , 
    n1568 , 
    n1569 , 
    n1570 , 
    n1571 , 
    n1572 , 
    n1573 , 
    n1574 , 
    n1575 , 
    n1576 , 
    n1577 , 
    n1578 , 
    n1579 , 
    n1580 , 
    n1581 , 
    n1582 , 
    n1583 , 
    n1584 , 
    n1585 , 
    n1586 , 
    n1587 , 
    n1588 , 
    n1589 , 
    n1590 , 
    n1591 , 
    n1592 , 
    n1593 , 
    n1594 , 
    n1595 , 
    n1596 , 
    n1597 , 
    n1598 , 
    n1599 , 
    n1600 , 
    n1601 , 
    n1602 , 
    n1603 , 
    n1604 , 
    n1605 , 
    n1606 , 
    n1607 , 
    n1608 , 
    n1609 , 
    n1610 , 
    n1611 , 
    n1612 , 
    n1613 , 
    n1614 , 
    n1615 , 
    n1616 , 
    n1617 , 
    n1618 , 
    n1619 , 
    n1620 , 
    n1621 , 
    n1622 , 
    n1623 , 
    n1624 , 
    n1625 , 
    n1626 , 
    n1627 , 
    n1628 , 
    n1629 , 
    n1630 , 
    n1631 , 
    n1632 , 
    n1633 , 
    n1634 , 
    n1635 , 
    n1636 , 
    n1637 , 
    n1638 , 
    n1639 , 
    n1640 , 
    n1641 , 
    n1642 , 
    n1643 , 
    n1644 , 
    n1645 , 
    n1646 , 
    n1647 , 
    n1648 , 
    n1649 , 
    n1650 , 
    n1651 , 
    n1652 , 
    n1653 , 
    n1654 , 
    n1655 , 
    n1656 , 
    n1657 , 
    n1658 , 
    n1659 , 
    n1660 , 
    n1661 , 
    n1662 , 
    n1663 , 
    n1664 , 
    n1665 , 
    n1666 , 
    n1667 , 
    n1668 , 
    n1669 , 
    n1670 , 
    n1671 , 
    n1672 , 
    n1673 , 
    n1674 , 
    n1675 , 
    n1676 , 
    n1677 , 
    n1678 , 
    n1679 , 
    n1680 , 
    n1681 , 
    n1682 , 
    n1683 , 
    n1684 , 
    n1685 , 
    n1686 , 
    n1687 , 
    n1688 , 
    n1689 , 
    n1690 , 
    n1691 , 
    n1692 , 
    n1693 , 
    n1694 , 
    n1695 , 
    n1696 , 
    n1697 , 
    n1698 , 
    n1699 , 
    n1700 , 
    n1701 , 
    n1702 , 
    n1703 , 
    n1704 , 
    n1705 , 
    n1706 , 
    n1707 , 
    n1708 , 
    n1709 , 
    n1710 , 
    n1711 , 
    n1712 , 
    n1713 , 
    n1714 , 
    n1715 , 
    n1716 , 
    n1717 , 
    n1718 , 
    n1719 , 
    n1720 , 
    n1721 , 
    n1722 , 
    n1723 , 
    n1724 , 
    n1725 , 
    n1726 , 
    n1727 , 
    n1728 , 
    n1729 , 
    n1730 , 
    n1731 , 
    n1732 , 
    n1733 , 
    n1734 , 
    n1735 , 
    n1736 , 
    n1737 , 
    n1738 , 
    n1739 , 
    n1740 , 
    n1741 , 
    n1742 , 
    n1743 , 
    n1744 , 
    n1745 , 
    n1746 , 
    n1747 , 
    n1748 , 
    n1749 , 
    n1750 , 
    n1751 , 
    n1752 , 
    n1753 , 
    n1754 , 
    n1755 , 
    n1756 , 
    n1757 , 
    n1758 , 
    n1759 , 
    n1760 , 
    n1761 , 
    n1762 , 
    n1763 , 
    n1764 , 
    n1765 , 
    n1766 , 
    n1767 , 
    n1768 , 
    n1769 , 
    n1770 , 
    n1771 , 
    n1772 , 
    n1773 , 
    n1774 , 
    n1775 , 
    n1776 , 
    n1777 , 
    n1778 , 
    n1779 , 
    n1780 , 
    n1781 , 
    n1782 , 
    n1783 , 
    n1784 , 
    n1785 , 
    n1786 , 
    n1787 , 
    n1788 , 
    n1789 , 
    n1790 , 
    n1791 , 
    n1792 , 
    n1793 , 
    n1794 , 
    n1795 , 
    n1796 , 
    n1797 , 
    n1798 , 
    n1799 , 
    n1800 , 
    n1801 , 
    n1802 , 
    n1803 , 
    n1804 , 
    n1805 , 
    n1806 , 
    n1807 , 
    n1808 , 
    n1809 , 
    n1810 , 
    n1811 , 
    n1812 , 
    n1813 , 
    n1814 , 
    n1815 , 
    n1816 , 
    n1817 , 
    n1818 , 
    n1819 , 
    n1820 , 
    n1821 , 
    n1822 , 
    n1823 , 
    n1824 , 
    n1825 , 
    n1826 , 
    n1827 , 
    n1828 , 
    n1829 , 
    n1830 , 
    n1831 , 
    n1832 , 
    n1833 , 
    n1834 , 
    n1835 , 
    n1836 , 
    n1837 , 
    n1838 , 
    n1839 , 
    n1840 , 
    n1841 , 
    n1842 , 
    n1843 , 
    n1844 , 
    n1845 , 
    n1846 , 
    n1847 , 
    n1848 , 
    n1849 , 
    n1850 , 
    n1851 , 
    n1852 , 
    n1853 , 
    n1854 , 
    n1855 , 
    n1856 , 
    n1857 , 
    n1858 , 
    n1859 , 
    n1860 , 
    n1861 , 
    n1862 , 
    n1863 , 
    n1864 , 
    n1865 , 
    n1866 , 
    n1867 , 
    n1868 , 
    n1869 , 
    n1870 , 
    n1871 , 
    n1872 , 
    n1873 , 
    n1874 , 
    n1875 , 
    n1876 , 
    n1877 , 
    n1878 , 
    n1879 , 
    n1880 , 
    n1881 , 
    n1882 , 
    n1883 , 
    n1884 , 
    n1885 , 
    n1886 , 
    n1887 , 
    n1888 , 
    n1889 , 
    n1890 , 
    n1891 , 
    n1892 , 
    n1893 , 
    n1894 , 
    n1895 , 
    n1896 , 
    n1897 , 
    n1898 , 
    n1899 , 
    n1900 , 
    n1901 , 
    n1902 , 
    n1903 , 
    n1904 , 
    n1905 , 
    n1906 , 
    n1907 , 
    n1908 , 
    n1909 , 
    n1910 , 
    n1911 , 
    n1912 , 
    n1913 , 
    n1914 , 
    n1915 , 
    n1916 , 
    n1917 , 
    n1918 , 
    n1919 , 
    n1920 , 
    n1921 , 
    n1922 , 
    n1923 , 
    n1924 , 
    n1925 , 
    n1926 , 
    n1927 , 
    n1928 , 
    n1929 , 
    n1930 , 
    n1931 , 
    n1932 , 
    n1933 , 
    n1934 , 
    n1935 , 
    n1936 , 
    n1937 , 
    n1938 , 
    n1939 , 
    n1940 , 
    n1941 , 
    n1942 , 
    n1943 , 
    n1944 , 
    n1945 , 
    n1946 , 
    n1947 , 
    n1948 , 
    n1949 , 
    n1950 , 
    n1951 , 
    n1952 , 
    n1953 , 
    n1954 , 
    n1955 , 
    n1956 , 
    n1957 , 
    n1958 , 
    n1959 , 
    n1960 , 
    n1961 , 
    n1962 , 
    n1963 , 
    n1964 , 
    n1965 , 
    n1966 , 
    n1967 , 
    n1968 , 
    n1969 , 
    n1970 , 
    n1971 , 
    n1972 , 
    n1973 , 
    n1974 , 
    n1975 , 
    n1976 , 
    n1977 , 
    n1978 , 
    n1979 , 
    n1980 , 
    n1981 , 
    n1982 , 
    n1983 , 
    n1984 , 
    n1985 , 
    n1986 , 
    n1987 , 
    n1988 , 
    n1989 , 
    n1990 , 
    n1991 , 
    n1992 , 
    n1993 , 
    n1994 , 
    n1995 , 
    n1996 , 
    n1997 , 
    n1998 , 
    n1999 , 
    n2000 , 
    n2001 , 
    n2002 , 
    n2003 , 
    n2004 , 
    n2005 , 
    n2006 , 
    n2007 , 
    n2008 , 
    n2009 , 
    n2010 , 
    n2011 , 
    n2012 , 
    n2013 , 
    n2014 , 
    n2015 , 
    n2016 , 
    n2017 , 
    n2018 , 
    n2019 , 
    n2020 , 
    n2021 , 
    n2022 , 
    n2023 , 
    n2024 , 
    n2025 , 
    n2026 , 
    n2027 , 
    n2028 , 
    n2029 , 
    n2030 , 
    n2031 , 
    n2032 , 
    n2033 , 
    n2034 , 
    n2035 , 
    n2036 , 
    n2037 , 
    n2038 , 
    n2039 , 
    n2040 , 
    n2041 , 
    n2042 , 
    n2043 , 
    n2044 , 
    n2045 , 
    n2046 , 
    n2047 , 
    n2048 , 
    n2049 , 
    n2050 , 
    n2051 , 
    n2052 , 
    n2053 , 
    n2054 , 
    n2055 , 
    n2056 , 
    n2057 , 
    n2058 , 
    n2059 , 
    n2060 , 
    n2061 , 
    n2062 , 
    n2063 , 
    n2064 , 
    n2065 , 
    n2066 , 
    n2067 , 
    n2068 , 
    n2069 , 
    n2070 , 
    n2071 , 
    n2072 , 
    n2073 , 
    n2074 , 
    n2075 , 
    n2076 , 
    n2077 , 
    n2078 , 
    n2079 , 
    n2080 , 
    n2081 , 
    n2082 , 
    n2083 , 
    n2084 , 
    n2085 , 
    n2086 , 
    n2087 , 
    n2088 , 
    n2089 , 
    n2090 , 
    n2091 , 
    n2092 , 
    n2093 , 
    n2094 , 
    n2095 , 
    n2096 , 
    n2097 , 
    n2098 , 
    n2099 , 
    n2100 , 
    n2101 , 
    n2102 , 
    n2103 , 
    n2104 , 
    n2105 , 
    n2106 , 
    n2107 , 
    n2108 , 
    n2109 , 
    n2110 , 
    n2111 , 
    n2112 , 
    n2113 , 
    n2114 , 
    n2115 , 
    n2116 , 
    n2117 , 
    n2118 , 
    n2119 , 
    n2120 , 
    n2121 , 
    n2122 , 
    n2123 , 
    n2124 , 
    n2125 , 
    n2126 , 
    n2127 , 
    n2128 , 
    n2129 , 
    n2130 , 
    n2131 , 
    n2132 , 
    n2133 , 
    n2134 , 
    n2135 , 
    n2136 , 
    n2137 , 
    n2138 , 
    n2139 , 
    n2140 , 
    n2141 , 
    n2142 , 
    n2143 , 
    n2144 , 
    n2145 , 
    n2146 , 
    n2147 , 
    n2148 , 
    n2149 , 
    n2150 , 
    n2151 , 
    n2152 , 
    n2153 , 
    n2154 , 
    n2155 , 
    n2156 , 
    n2157 , 
    n2158 , 
    n2159 , 
    n2160 , 
    n2161 , 
    n2162 , 
    n2163 , 
    n2164 , 
    n2165 , 
    n2166 , 
    n2167 , 
    n2168 , 
    n2169 , 
    n2170 , 
    n2171 , 
    n2172 , 
    n2173 , 
    n2174 , 
    n2175 , 
    n2176 , 
    n2177 , 
    n2178 , 
    n2179 , 
    n2180 , 
    n2181 , 
    n2182 , 
    n2183 , 
    n2184 , 
    n2185 , 
    n2186 , 
    n2187 , 
    n2188 , 
    n2189 , 
    n2190 , 
    n2191 , 
    n2192 , 
    n2193 , 
    n2194 , 
    n2195 , 
    n2196 , 
    n2197 , 
    n2198 , 
    n2199 , 
    n2200 , 
    n2201 , 
    n2202 , 
    n2203 , 
    n2204 , 
    n2205 , 
    n2206 , 
    n2207 , 
    n2208 , 
    n2209 , 
    n2210 , 
    n2211 , 
    n2212 , 
    n2213 , 
    n2214 , 
    n2215 , 
    n2216 , 
    n2217 , 
    n2218 , 
    n2219 , 
    n2220 , 
    n2221 , 
    n2222 , 
    n2223 , 
    n2224 , 
    n2225 , 
    n2226 , 
    n2227 , 
    n2228 , 
    n2229 , 
    n2230 , 
    n2231 , 
    n2232 , 
    n2233 , 
    n2234 , 
    n2235 , 
    n2236 , 
    n2237 , 
    n2238 , 
    n2239 , 
    n2240 , 
    n2241 , 
    n2242 , 
    n2243 , 
    n2244 , 
    n2245 , 
    n2246 , 
    n2247 , 
    n2248 , 
    n2249 , 
    n2250 , 
    n2251 , 
    n2252 , 
    n2253 , 
    n2254 , 
    n2255 , 
    n2256 , 
    n2257 , 
    n2258 , 
    n2259 , 
    n2260 , 
    n2261 , 
    n2262 , 
    n2263 , 
    n2264 , 
    n2265 , 
    n2266 , 
    n2267 , 
    n2268 , 
    n2269 , 
    n2270 , 
    n2271 , 
    n2272 , 
    n2273 , 
    n2274 , 
    n2275 , 
    n2276 , 
    n2277 , 
    n2278 , 
    n2279 , 
    n2280 , 
    n2281 , 
    n2282 , 
    n2283 , 
    n2284 , 
    n2285 , 
    n2286 , 
    n2287 , 
    n2288 , 
    n2289 , 
    n2290 , 
    n2291 , 
    n2292 , 
    n2293 , 
    n2294 , 
    n2295 , 
    n2296 , 
    n2297 , 
    n2298 , 
    n2299 , 
    n2300 , 
    n2301 , 
    n2302 , 
    n2303 , 
    n2304 , 
    n2305 , 
    n2306 , 
    n2307 , 
    n2308 , 
    n2309 , 
    n2310 , 
    n2311 , 
    n2312 , 
    n2313 , 
    n2314 , 
    n2315 , 
    n2316 , 
    n2317 , 
    n2318 , 
    n2319 , 
    n2320 , 
    n2321 , 
    n2322 , 
    n2323 , 
    n2324 , 
    n2325 , 
    n2326 , 
    n2327 , 
    n2328 , 
    n2329 , 
    n2330 , 
    n2331 , 
    n2332 , 
    n2333 , 
    n2334 , 
    n2335 , 
    n2336 , 
    n2337 , 
    n2338 , 
    n2339 , 
    n2340 , 
    n2341 , 
    n2342 , 
    n2343 , 
    n2344 , 
    n2345 , 
    n2346 , 
    n2347 , 
    n2348 , 
    n2349 , 
    n2350 , 
    n2351 , 
    n2352 , 
    n2353 , 
    n2354 , 
    n2355 , 
    n2356 , 
    n2357 , 
    n2358 , 
    n2359 , 
    n2360 , 
    n2361 , 
    n2362 , 
    n2363 , 
    n2364 , 
    n2365 , 
    n2366 , 
    n2367 , 
    n2368 , 
    n2369 , 
    n2370 , 
    n2371 , 
    n2372 , 
    n2373 , 
    n2374 , 
    n2375 , 
    n2376 , 
    n2377 , 
    n2378 , 
    n2379 , 
    n2380 , 
    n2381 , 
    n2382 , 
    n2383 , 
    n2384 , 
    n2385 , 
    n2386 , 
    n2387 , 
    n2388 , 
    n2389 , 
    n2390 , 
    n2391 , 
    n2392 , 
    n2393 , 
    n2394 , 
    n2395 , 
    n2396 , 
    n2397 , 
    n2398 , 
    n2399 , 
    n2400 , 
    n2401 , 
    n2402 , 
    n2403 , 
    n2404 , 
    n2405 , 
    n2406 , 
    n2407 , 
    n2408 , 
    n2409 , 
    n2410 , 
    n2411 , 
    n2412 , 
    n2413 , 
    n2414 , 
    n2415 , 
    n2416 , 
    n2417 , 
    n2418 , 
    n2419 , 
    n2420 , 
    n2421 , 
    n2422 , 
    n2423 , 
    n2424 , 
    n2425 , 
    n2426 , 
    n2427 , 
    n2428 , 
    n2429 , 
    n2430 , 
    n2431 , 
    n2432 , 
    n2433 , 
    n2434 , 
    n2435 , 
    n2436 , 
    n2437 , 
    n2438 , 
    n2439 , 
    n2440 , 
    n2441 , 
    n2442 , 
    n2443 , 
    n2444 , 
    n2445 , 
    n2446 , 
    n2447 , 
    n2448 , 
    n2449 , 
    n2450 , 
    n2451 , 
    n2452 , 
    n2453 , 
    n2454 , 
    n2455 , 
    n2456 , 
    n2457 , 
    n2458 , 
    n2459 , 
    n2460 , 
    n2461 , 
    n2462 , 
    n2463 , 
    n2464 , 
    n2465 , 
    n2466 , 
    n2467 , 
    n2468 , 
    n2469 , 
    n2470 , 
    n2471 , 
    n2472 , 
    n2473 , 
    n2474 , 
    n2475 , 
    n2476 , 
    n2477 , 
    n2478 , 
    n2479 , 
    n2480 , 
    n2481 , 
    n2482 , 
    n2483 , 
    n2484 , 
    n2485 , 
    n2486 , 
    n2487 , 
    n2488 , 
    n2489 , 
    n2490 , 
    n2491 , 
    n2492 , 
    n2493 , 
    n2494 , 
    n2495 , 
    n2496 , 
    n2497 , 
    n2498 , 
    n2499 , 
    n2500 , 
    n2501 , 
    n2502 , 
    n2503 , 
    n2504 , 
    n2505 , 
    n2506 , 
    n2507 , 
    n2508 , 
    n2509 , 
    n2510 , 
    n2511 , 
    n2512 , 
    n2513 , 
    n2514 , 
    n2515 , 
    n2516 , 
    n2517 , 
    n2518 , 
    n2519 , 
    n2520 , 
    n2521 , 
    n2522 , 
    n2523 , 
    n2524 , 
    n2525 , 
    n2526 , 
    n2527 , 
    n2528 , 
    n2529 , 
    n2530 , 
    n2531 , 
    n2532 , 
    n2533 , 
    n2534 , 
    n2535 , 
    n2536 , 
    n2537 , 
    n2538 , 
    n2539 , 
    n2540 , 
    n2541 , 
    n2542 , 
    n2543 , 
    n2544 , 
    n2545 , 
    n2546 , 
    n2547 , 
    n2548 , 
    n2549 , 
    n2550 , 
    n2551 , 
    n2552 , 
    n2553 , 
    n2554 , 
    n2555 , 
    n2556 , 
    n2557 , 
    n2558 , 
    n2559 , 
    n2560 , 
    n2561 , 
    n2562 , 
    n2563 , 
    n2564 , 
    n2565 , 
    n2566 , 
    n2567 , 
    n2568 , 
    n2569 , 
    n2570 , 
    n2571 , 
    n2572 , 
    n2573 , 
    n2574 , 
    n2575 , 
    n2576 , 
    n2577 , 
    n2578 , 
    n2579 , 
    n2580 , 
    n2581 , 
    n2582 , 
    n2583 , 
    n2584 , 
    n2585 , 
    n2586 , 
    n2587 , 
    n2588 , 
    n2589 , 
    n2590 , 
    n2591 , 
    n2592 , 
    n2593 , 
    n2594 , 
    n2595 , 
    n2596 , 
    n2597 , 
    n2598 , 
    n2599 , 
    n2600 , 
    n2601 , 
    n2602 , 
    n2603 , 
    n2604 , 
    n2605 , 
    n2606 , 
    n2607 , 
    n2608 , 
    n2609 , 
    n2610 , 
    n2611 , 
    n2612 , 
    n2613 , 
    n2614 , 
    n2615 , 
    n2616 , 
    n2617 , 
    n2618 , 
    n2619 , 
    n2620 , 
    n2621 , 
    n2622 , 
    n2623 , 
    n2624 , 
    n2625 , 
    n2626 , 
    n2627 , 
    n2628 , 
    n2629 , 
    n2630 , 
    n2631 , 
    n2632 , 
    n2633 , 
    n2634 , 
    n2635 , 
    n2636 , 
    n2637 , 
    n2638 , 
    n2639 , 
    n2640 , 
    n2641 , 
    n2642 , 
    n2643 , 
    n2644 , 
    n2645 , 
    n2646 , 
    n2647 , 
    n2648 , 
    n2649 , 
    n2650 , 
    n2651 , 
    n2652 , 
    n2653 , 
    n2654 , 
    n2655 , 
    n2656 , 
    n2657 , 
    n2658 , 
    n2659 , 
    n2660 , 
    n2661 , 
    n2662 , 
    n2663 , 
    n2664 , 
    n2665 , 
    n2666 , 
    n2667 , 
    n2668 , 
    n2669 , 
    n2670 , 
    n2671 , 
    n2672 , 
    n2673 , 
    n2674 , 
    n2675 , 
    n2676 , 
    n2677 , 
    n2678 , 
    n2679 , 
    n2680 , 
    n2681 , 
    n2682 , 
    n2683 , 
    n2684 , 
    n2685 , 
    n2686 , 
    n2687 , 
    n2688 , 
    n2689 , 
    n2690 , 
    n2691 , 
    n2692 , 
    n2693 , 
    n2694 , 
    n2695 , 
    n2696 , 
    n2697 , 
    n2698 , 
    n2699 , 
    n2700 , 
    n2701 , 
    n2702 , 
    n2703 , 
    n2704 , 
    n2705 , 
    n2706 , 
    n2707 , 
    n2708 , 
    n2709 , 
    n2710 , 
    n2711 , 
    n2712 , 
    n2713 , 
    n2714 , 
    n2715 , 
    n2716 , 
    n2717 , 
    n2718 , 
    n2719 , 
    n2720 , 
    n2721 , 
    n2722 , 
    n2723 , 
    n2724 , 
    n2725 , 
    n2726 , 
    n2727 , 
    n2728 , 
    n2729 , 
    n2730 , 
    n2731 , 
    n2732 , 
    n2733 , 
    n2734 , 
    n2735 , 
    n2736 , 
    n2737 , 
    n2738 , 
    n2739 , 
    n2740 , 
    n2741 , 
    n2742 , 
    n2743 , 
    n2744 , 
    n2745 , 
    n2746 , 
    n2747 , 
    n2748 , 
    n2749 , 
    n2750 , 
    n2751 , 
    n2752 , 
    n2753 , 
    n2754 , 
    n2755 , 
    n2756 , 
    n2757 , 
    n2758 , 
    n2759 , 
    n2760 , 
    n2761 , 
    n2762 , 
    n2763 , 
    n2764 , 
    n2765 , 
    n2766 , 
    n2767 , 
    n2768 , 
    n2769 , 
    n2770 , 
    n2771 , 
    n2772 , 
    n2773 , 
    n2774 , 
    n2775 , 
    n2776 , 
    n2777 , 
    n2778 , 
    n2779 , 
    n2780 , 
    n2781 , 
    n2782 , 
    n2783 , 
    n2784 , 
    n2785 , 
    n2786 , 
    n2787 , 
    n2788 , 
    n2789 , 
    n2790 , 
    n2791 , 
    n2792 , 
    n2793 , 
    n2794 , 
    n2795 , 
    n2796 , 
    n2797 , 
    n2798 , 
    n2799 , 
    n2800 , 
    n2801 , 
    n2802 , 
    n2803 , 
    n2804 , 
    n2805 , 
    n2806 , 
    n2807 , 
    n2808 , 
    n2809 , 
    n2810 , 
    n2811 , 
    n2812 , 
    n2813 , 
    n2814 , 
    n2815 , 
    n2816 , 
    n2817 , 
    n2818 , 
    n2819 , 
    n2820 , 
    n2821 , 
    n2822 , 
    n2823 , 
    n2824 , 
    n2825 , 
    n2826 , 
    n2827 , 
    n2828 , 
    n2829 , 
    n2830 , 
    n2831 , 
    n2832 , 
    n2833 , 
    n2834 , 
    n2835 , 
    n2836 , 
    n2837 , 
    n2838 , 
    n2839 , 
    n2840 , 
    n2841 , 
    n2842 , 
    n2843 , 
    n2844 , 
    n2845 , 
    n2846 , 
    n2847 , 
    n2848 , 
    n2849 , 
    n2850 , 
    n2851 , 
    n2852 , 
    n2853 , 
    n2854 , 
    n2855 , 
    n2856 , 
    n2857 , 
    n2858 , 
    n2859 , 
    n2860 , 
    n2861 , 
    n2862 , 
    n2863 , 
    n2864 , 
    n2865 , 
    n2866 , 
    n2867 , 
    n2868 , 
    n2869 , 
    n2870 , 
    n2871 , 
    n2872 , 
    n2873 , 
    n2874 , 
    n2875 , 
    n2876 , 
    n2877 , 
    n2878 , 
    n2879 , 
    n2880 , 
    n2881 , 
    n2882 , 
    n2883 , 
    n2884 , 
    n2885 , 
    n2886 , 
    n2887 , 
    n2888 , 
    n2889 , 
    n2890 , 
    n2891 , 
    n2892 , 
    n2893 , 
    n2894 , 
    n2895 , 
    n2896 , 
    n2897 , 
    n2898 , 
    n2899 , 
    n2900 , 
    n2901 , 
    n2902 , 
    n2903 , 
    n2904 , 
    n2905 , 
    n2906 , 
    n2907 , 
    n2908 , 
    n2909 , 
    n2910 , 
    n2911 , 
    n2912 , 
    n2913 , 
    n2914 , 
    n2915 , 
    n2916 , 
    n2917 , 
    n2918 , 
    n2919 , 
    n2920 , 
    n2921 , 
    n2922 , 
    n2923 , 
    n2924 , 
    n2925 , 
    n2926 , 
    n2927 , 
    n2928 , 
    n2929 , 
    n2930 , 
    n2931 , 
    n2932 , 
    n2933 , 
    n2934 , 
    n2935 , 
    n2936 , 
    n2937 , 
    n2938 , 
    n2939 , 
    n2940 , 
    n2941 , 
    n2942 , 
    n2943 , 
    n2944 , 
    n2945 , 
    n2946 , 
    n2947 , 
    n2948 , 
    n2949 , 
    n2950 , 
    n2951 , 
    n2952 , 
    n2953 , 
    n2954 , 
    n2955 , 
    n2956 , 
    n2957 , 
    n2958 , 
    n2959 , 
    n2960 , 
    n2961 , 
    n2962 , 
    n2963 , 
    n2964 , 
    n2965 , 
    n2966 , 
    n2967 , 
    n2968 , 
    n2969 , 
    n2970 , 
    n2971 , 
    n2972 , 
    n2973 , 
    n2974 , 
    n2975 , 
    n2976 , 
    n2977 , 
    n2978 , 
    n2979 , 
    n2980 , 
    n2981 , 
    n2982 , 
    n2983 , 
    n2984 , 
    n2985 , 
    n2986 , 
    n2987 , 
    n2988 , 
    n2989 , 
    n2990 , 
    n2991 , 
    n2992 , 
    n2993 , 
    n2994 , 
    n2995 , 
    n2996 , 
    n2997 , 
    n2998 , 
    n2999 , 
    n3000 , 
    n3001 , 
    n3002 , 
    n3003 , 
    n3004 , 
    n3005 , 
    n3006 , 
    n3007 , 
    n3008 , 
    n3009 , 
    n3010 , 
    n3011 , 
    n3012 , 
    n3013 , 
    n3014 , 
    n3015 , 
    n3016 , 
    n3017 , 
    n3018 , 
    n3019 , 
    n3020 , 
    n3021 , 
    n3022 , 
    n3023 , 
    n3024 , 
    n3025 , 
    n3026 , 
    n3027 , 
    n3028 , 
    n3029 , 
    n3030 , 
    n3031 , 
    n3032 , 
    n3033 , 
    n3034 , 
    n3035 , 
    n3036 , 
    n3037 , 
    n3038 , 
    n3039 , 
    n3040 , 
    n3041 , 
    n3042 , 
    n3043 , 
    n3044 , 
    n3045 , 
    n3046 , 
    n3047 , 
    n3048 , 
    n3049 , 
    n3050 , 
    n3051 , 
    n3052 , 
    n3053 , 
    n3054 , 
    n3055 , 
    n3056 , 
    n3057 , 
    n3058 , 
    n3059 , 
    n3060 , 
    n3061 , 
    n3062 , 
    n3063 , 
    n3064 , 
    n3065 , 
    n3066 , 
    n3067 , 
    n3068 , 
    n3069 , 
    n3070 , 
    n3071 , 
    n3072 , 
    n3073 , 
    n3074 , 
    n3075 , 
    n3076 , 
    n3077 , 
    n3078 , 
    n3079 , 
    n3080 , 
    n3081 , 
    n3082 , 
    n3083 , 
    n3084 , 
    n3085 , 
    n3086 , 
    n3087 , 
    n3088 , 
    n3089 , 
    n3090 , 
    n3091 , 
    n3092 , 
    n3093 , 
    n3094 , 
    n3095 , 
    n3096 , 
    n3097 , 
    n3098 , 
    n3099 , 
    n3100 , 
    n3101 , 
    n3102 , 
    n3103 , 
    n3104 , 
    n3105 , 
    n3106 , 
    n3107 , 
    n3108 , 
    n3109 , 
    n3110 , 
    n3111 , 
    n3112 , 
    n3113 , 
    n3114 , 
    n3115 , 
    n3116 , 
    n3117 , 
    n3118 , 
    n3119 , 
    n3120 , 
    n3121 , 
    n3122 , 
    n3123 );
input  n0 , 
    n1 , 
    n2 , 
    n3 , 
    n4 , 
    n5 , 
    n6 , 
    n7 , 
    n8 , 
    n9 , 
    n10 , 
    n11 , 
    n12 , 
    n13 , 
    n14 , 
    n15 , 
    n16 , 
    n17 , 
    n18 , 
    n19 , 
    n20 , 
    n21 , 
    n22 , 
    n23 , 
    n24 , 
    n25 , 
    n26 , 
    n27 , 
    n28 , 
    n29 , 
    n30 , 
    n31 , 
    n32 , 
    n33 , 
    n34 , 
    n35 , 
    n36 , 
    n37 , 
    n38 , 
    n39 , 
    n40 , 
    n41 , 
    n42 , 
    n43 , 
    n44 , 
    n45 , 
    n46 , 
    n47 , 
    n48 , 
    n49 , 
    n50 , 
    n51 , 
    n52 , 
    n53 , 
    n54 , 
    n55 , 
    n56 , 
    n57 , 
    n58 , 
    n59 , 
    n60 , 
    n61 , 
    n62 , 
    n63 , 
    n64 , 
    n65 , 
    n66 , 
    n67 , 
    n68 , 
    n69 , 
    n70 , 
    n71 , 
    n72 , 
    n73 , 
    n74 , 
    n75 , 
    n76 , 
    n77 , 
    n78 , 
    n79 , 
    n80 , 
    n81 , 
    n82 , 
    n83 , 
    n84 , 
    n85 , 
    n86 , 
    n87 , 
    n88 , 
    n89 , 
    n90 , 
    n91 , 
    n92 , 
    n93 , 
    n94 , 
    n95 , 
    n96 , 
    n97 , 
    n98 , 
    n99 , 
    n100 , 
    n101 , 
    n102 , 
    n103 , 
    n104 , 
    n105 , 
    n106 , 
    n107 , 
    n108 , 
    n109 , 
    n110 , 
    n111 , 
    n112 , 
    n113 , 
    n114 , 
    n115 , 
    n116 , 
    n117 , 
    n118 , 
    n119 , 
    n120 , 
    n121 , 
    n122 , 
    n123 , 
    n124 , 
    n125 , 
    n126 , 
    n127 , 
    n128 , 
    n129 , 
    n130 , 
    n131 , 
    n132 , 
    n133 , 
    n134 , 
    n135 , 
    n136 , 
    n137 , 
    n138 , 
    n139 , 
    n140 , 
    n141 , 
    n142 , 
    n143 , 
    n144 , 
    n145 , 
    n146 , 
    n147 , 
    n148 , 
    n149 , 
    n150 , 
    n151 , 
    n152 , 
    n153 , 
    n154 , 
    n155 , 
    n156 , 
    n157 , 
    n158 , 
    n159 , 
    n160 , 
    n161 , 
    n162 , 
    n163 , 
    n164 , 
    n165 , 
    n166 , 
    n167 , 
    n168 , 
    n169 , 
    n170 , 
    n171 , 
    n172 , 
    n173 , 
    n174 , 
    n175 , 
    n176 , 
    n177 , 
    n178 , 
    n179 , 
    n180 , 
    n181 , 
    n182 , 
    n183 , 
    n184 , 
    n185 , 
    n186 , 
    n187 , 
    n188 , 
    n189 , 
    n190 , 
    n191 , 
    n192 , 
    n193 , 
    n194 , 
    n195 , 
    n196 , 
    n197 , 
    n198 , 
    n199 , 
    n200 , 
    n201 , 
    n202 , 
    n203 , 
    n204 , 
    n205 , 
    n206 , 
    n207 , 
    n208 , 
    n209 , 
    n210 , 
    n211 , 
    n212 , 
    n213 , 
    n214 , 
    n215 , 
    n216 , 
    n217 , 
    n218 , 
    n219 , 
    n220 , 
    n221 , 
    n222 , 
    n223 , 
    n224 , 
    n225 , 
    n226 , 
    n227 , 
    n228 , 
    n229 , 
    n230 , 
    n231 , 
    n232 , 
    n233 , 
    n234 , 
    n235 , 
    n236 , 
    n237 , 
    n238 , 
    n239 , 
    n240 , 
    n241 , 
    n242 , 
    n243 , 
    n244 , 
    n245 , 
    n246 , 
    n247 , 
    n248 , 
    n249 , 
    n250 , 
    n251 , 
    n252 , 
    n253 , 
    n254 , 
    n255 , 
    n256 , 
    n257 , 
    n258 , 
    n259 , 
    n260 , 
    n261 , 
    n262 , 
    n263 , 
    n264 , 
    n265 , 
    n266 , 
    n267 , 
    n268 , 
    n269 , 
    n270 , 
    n271 , 
    n272 , 
    n273 , 
    n274 , 
    n275 , 
    n276 , 
    n277 , 
    n278 , 
    n279 , 
    n280 , 
    n281 , 
    n282 , 
    n283 , 
    n284 , 
    n285 , 
    n286 , 
    n287 , 
    n288 , 
    n289 , 
    n290 , 
    n291 , 
    n292 , 
    n293 , 
    n294 , 
    n295 , 
    n296 , 
    n297 , 
    n298 , 
    n299 , 
    n300 , 
    n301 , 
    n302 , 
    n303 , 
    n304 , 
    n305 , 
    n306 , 
    n307 , 
    n308 , 
    n309 , 
    n310 , 
    n311 , 
    n312 , 
    n313 , 
    n314 , 
    n315 , 
    n316 , 
    n317 , 
    n318 , 
    n319 , 
    n320 , 
    n321 , 
    n322 , 
    n323 , 
    n324 , 
    n325 , 
    n326 , 
    n327 , 
    n328 , 
    n329 , 
    n330 , 
    n331 , 
    n332 , 
    n333 , 
    n334 , 
    n335 , 
    n336 , 
    n337 , 
    n338 , 
    n339 , 
    n340 , 
    n341 , 
    n342 , 
    n343 , 
    n344 , 
    n345 , 
    n346 , 
    n347 , 
    n348 , 
    n349 , 
    n350 , 
    n351 , 
    n352 , 
    n353 , 
    n354 , 
    n355 , 
    n356 , 
    n357 , 
    n358 , 
    n359 , 
    n360 , 
    n361 , 
    n362 , 
    n363 , 
    n364 , 
    n365 , 
    n366 , 
    n367 , 
    n368 , 
    n369 , 
    n370 , 
    n371 , 
    n372 , 
    n373 , 
    n374 , 
    n375 , 
    n376 , 
    n377 , 
    n378 , 
    n379 , 
    n380 , 
    n381 , 
    n382 , 
    n383 , 
    n384 , 
    n385 , 
    n386 , 
    n387 , 
    n388 , 
    n389 , 
    n390 , 
    n391 , 
    n392 , 
    n393 , 
    n394 , 
    n395 , 
    n396 , 
    n397 , 
    n398 , 
    n399 , 
    n400 , 
    n401 , 
    n402 , 
    n403 , 
    n404 , 
    n405 , 
    n406 , 
    n407 , 
    n408 , 
    n409 , 
    n410 , 
    n411 , 
    n412 , 
    n413 , 
    n414 , 
    n415 , 
    n416 , 
    n417 , 
    n418 , 
    n419 , 
    n420 , 
    n421 , 
    n422 , 
    n423 , 
    n424 , 
    n425 , 
    n426 , 
    n427 , 
    n428 , 
    n429 , 
    n430 , 
    n431 , 
    n432 , 
    n433 , 
    n434 , 
    n435 , 
    n436 , 
    n437 , 
    n438 , 
    n439 , 
    n440 , 
    n441 , 
    n442 , 
    n443 , 
    n444 , 
    n445 , 
    n446 , 
    n447 , 
    n448 , 
    n449 , 
    n450 , 
    n451 , 
    n452 , 
    n453 , 
    n454 , 
    n455 , 
    n456 , 
    n457 , 
    n458 , 
    n459 , 
    n460 , 
    n461 , 
    n462 , 
    n463 , 
    n464 , 
    n465 , 
    n466 , 
    n467 , 
    n468 , 
    n469 , 
    n470 , 
    n471 , 
    n472 , 
    n473 , 
    n474 , 
    n475 , 
    n476 , 
    n477 , 
    n478 , 
    n479 , 
    n480 , 
    n481 , 
    n482 , 
    n483 , 
    n484 , 
    n485 , 
    n486 , 
    n487 , 
    n488 , 
    n489 , 
    n490 , 
    n491 , 
    n492 , 
    n493 , 
    n494 , 
    n495 , 
    n496 , 
    n497 , 
    n498 , 
    n499 , 
    n500 , 
    n501 , 
    n502 , 
    n503 , 
    n504 , 
    n505 , 
    n506 , 
    n507 , 
    n508 , 
    n509 , 
    n510 , 
    n511 , 
    n512 , 
    n513 , 
    n514 , 
    n515 , 
    n516 , 
    n517 , 
    n518 , 
    n519 , 
    n520 , 
    n521 , 
    n522 , 
    n523 , 
    n524 , 
    n525 , 
    n526 , 
    n527 , 
    n528 , 
    n529 , 
    n530 , 
    n531 , 
    n532 , 
    n533 , 
    n534 , 
    n535 , 
    n536 , 
    n537 , 
    n538 , 
    n539 , 
    n540 , 
    n541 , 
    n542 , 
    n543 , 
    n544 , 
    n545 , 
    n546 , 
    n547 , 
    n548 , 
    n549 , 
    n550 , 
    n551 , 
    n552 , 
    n553 , 
    n554 , 
    n555 , 
    n556 , 
    n557 , 
    n558 , 
    n559 , 
    n560 , 
    n561 , 
    n562 , 
    n563 , 
    n564 , 
    n565 , 
    n566 , 
    n567 , 
    n568 , 
    n569 , 
    n570 , 
    n571 , 
    n572 , 
    n573 , 
    n574 , 
    n575 , 
    n576 , 
    n577 , 
    n578 , 
    n579 , 
    n580 , 
    n581 , 
    n582 , 
    n583 , 
    n584 , 
    n585 , 
    n586 , 
    n587 , 
    n588 , 
    n589 , 
    n590 , 
    n591 , 
    n592 , 
    n593 , 
    n594 , 
    n595 , 
    n596 , 
    n597 , 
    n598 , 
    n599 , 
    n600 , 
    n601 , 
    n602 , 
    n603 , 
    n604 , 
    n605 , 
    n606 , 
    n607 , 
    n608 , 
    n609 , 
    n610 , 
    n611 , 
    n612 , 
    n613 , 
    n614 , 
    n615 , 
    n616 , 
    n617 , 
    n618 , 
    n619 , 
    n620 , 
    n621 , 
    n622 , 
    n623 , 
    n624 , 
    n625 , 
    n626 , 
    n627 , 
    n628 , 
    n629 , 
    n630 , 
    n631 , 
    n632 , 
    n633 , 
    n634 , 
    n635 , 
    n636 , 
    n637 , 
    n638 , 
    n639 , 
    n640 , 
    n641 , 
    n642 , 
    n643 , 
    n644 , 
    n645 , 
    n646 , 
    n647 , 
    n648 , 
    n649 ;
output 
    n650 , 
    n651 , 
    n652 , 
    n653 , 
    n654 , 
    n655 , 
    n656 , 
    n657 , 
    n658 , 
    n659 , 
    n660 , 
    n661 , 
    n662 , 
    n663 , 
    n664 , 
    n665 , 
    n666 , 
    n667 , 
    n668 , 
    n669 , 
    n670 , 
    n671 , 
    n672 , 
    n673 , 
    n674 , 
    n675 , 
    n676 , 
    n677 , 
    n678 , 
    n679 , 
    n680 , 
    n681 , 
    n682 , 
    n683 , 
    n684 , 
    n685 , 
    n686 , 
    n687 , 
    n688 , 
    n689 , 
    n690 , 
    n691 , 
    n692 , 
    n693 , 
    n694 , 
    n695 , 
    n696 , 
    n697 , 
    n698 , 
    n699 , 
    n700 , 
    n701 , 
    n702 , 
    n703 , 
    n704 , 
    n705 , 
    n706 , 
    n707 , 
    n708 , 
    n709 , 
    n710 , 
    n711 , 
    n712 , 
    n713 , 
    n714 , 
    n715 , 
    n716 , 
    n717 , 
    n718 , 
    n719 , 
    n720 , 
    n721 , 
    n722 , 
    n723 , 
    n724 , 
    n725 , 
    n726 , 
    n727 , 
    n728 , 
    n729 , 
    n730 , 
    n731 , 
    n732 , 
    n733 , 
    n734 , 
    n735 , 
    n736 , 
    n737 , 
    n738 , 
    n739 , 
    n740 , 
    n741 , 
    n742 , 
    n743 , 
    n744 , 
    n745 , 
    n746 , 
    n747 , 
    n748 , 
    n749 , 
    n750 , 
    n751 , 
    n752 , 
    n753 , 
    n754 , 
    n755 , 
    n756 , 
    n757 , 
    n758 , 
    n759 , 
    n760 , 
    n761 , 
    n762 , 
    n763 , 
    n764 , 
    n765 , 
    n766 , 
    n767 , 
    n768 , 
    n769 , 
    n770 , 
    n771 , 
    n772 , 
    n773 , 
    n774 , 
    n775 , 
    n776 , 
    n777 , 
    n778 , 
    n779 , 
    n780 , 
    n781 , 
    n782 , 
    n783 , 
    n784 , 
    n785 , 
    n786 , 
    n787 , 
    n788 , 
    n789 , 
    n790 , 
    n791 , 
    n792 , 
    n793 , 
    n794 , 
    n795 , 
    n796 , 
    n797 , 
    n798 , 
    n799 , 
    n800 , 
    n801 , 
    n802 , 
    n803 , 
    n804 , 
    n805 , 
    n806 , 
    n807 , 
    n808 , 
    n809 , 
    n810 , 
    n811 , 
    n812 , 
    n813 , 
    n814 , 
    n815 , 
    n816 , 
    n817 , 
    n818 , 
    n819 , 
    n820 , 
    n821 , 
    n822 , 
    n823 , 
    n824 , 
    n825 , 
    n826 , 
    n827 , 
    n828 , 
    n829 , 
    n830 , 
    n831 , 
    n832 , 
    n833 , 
    n834 , 
    n835 , 
    n836 , 
    n837 , 
    n838 , 
    n839 , 
    n840 , 
    n841 , 
    n842 , 
    n843 , 
    n844 , 
    n845 , 
    n846 , 
    n847 , 
    n848 , 
    n849 , 
    n850 , 
    n851 , 
    n852 , 
    n853 , 
    n854 , 
    n855 , 
    n856 , 
    n857 , 
    n858 , 
    n859 , 
    n860 , 
    n861 , 
    n862 , 
    n863 , 
    n864 , 
    n865 , 
    n866 , 
    n867 , 
    n868 , 
    n869 , 
    n870 , 
    n871 , 
    n872 , 
    n873 , 
    n874 , 
    n875 , 
    n876 , 
    n877 , 
    n878 , 
    n879 , 
    n880 , 
    n881 , 
    n882 , 
    n883 , 
    n884 , 
    n885 , 
    n886 , 
    n887 , 
    n888 , 
    n889 , 
    n890 , 
    n891 , 
    n892 , 
    n893 , 
    n894 , 
    n895 , 
    n896 , 
    n897 , 
    n898 , 
    n899 , 
    n900 , 
    n901 , 
    n902 , 
    n903 , 
    n904 , 
    n905 , 
    n906 , 
    n907 , 
    n908 , 
    n909 , 
    n910 , 
    n911 , 
    n912 , 
    n913 , 
    n914 , 
    n915 , 
    n916 , 
    n917 , 
    n918 , 
    n919 , 
    n920 , 
    n921 , 
    n922 , 
    n923 , 
    n924 , 
    n925 , 
    n926 , 
    n927 , 
    n928 , 
    n929 , 
    n930 , 
    n931 , 
    n932 , 
    n933 , 
    n934 , 
    n935 , 
    n936 , 
    n937 , 
    n938 , 
    n939 , 
    n940 , 
    n941 , 
    n942 , 
    n943 , 
    n944 , 
    n945 , 
    n946 , 
    n947 , 
    n948 , 
    n949 , 
    n950 , 
    n951 , 
    n952 , 
    n953 , 
    n954 , 
    n955 , 
    n956 , 
    n957 , 
    n958 , 
    n959 , 
    n960 , 
    n961 , 
    n962 , 
    n963 , 
    n964 , 
    n965 , 
    n966 , 
    n967 , 
    n968 , 
    n969 , 
    n970 , 
    n971 , 
    n972 , 
    n973 , 
    n974 , 
    n975 , 
    n976 , 
    n977 , 
    n978 , 
    n979 , 
    n980 , 
    n981 , 
    n982 , 
    n983 , 
    n984 , 
    n985 , 
    n986 , 
    n987 , 
    n988 , 
    n989 , 
    n990 , 
    n991 , 
    n992 , 
    n993 , 
    n994 , 
    n995 , 
    n996 , 
    n997 , 
    n998 , 
    n999 , 
    n1000 , 
    n1001 , 
    n1002 , 
    n1003 , 
    n1004 , 
    n1005 , 
    n1006 , 
    n1007 , 
    n1008 , 
    n1009 , 
    n1010 , 
    n1011 , 
    n1012 , 
    n1013 , 
    n1014 , 
    n1015 , 
    n1016 , 
    n1017 , 
    n1018 , 
    n1019 , 
    n1020 , 
    n1021 , 
    n1022 , 
    n1023 , 
    n1024 , 
    n1025 , 
    n1026 , 
    n1027 , 
    n1028 , 
    n1029 , 
    n1030 , 
    n1031 , 
    n1032 , 
    n1033 , 
    n1034 , 
    n1035 , 
    n1036 , 
    n1037 , 
    n1038 , 
    n1039 , 
    n1040 , 
    n1041 , 
    n1042 , 
    n1043 , 
    n1044 , 
    n1045 , 
    n1046 , 
    n1047 , 
    n1048 , 
    n1049 , 
    n1050 , 
    n1051 , 
    n1052 , 
    n1053 , 
    n1054 , 
    n1055 , 
    n1056 , 
    n1057 , 
    n1058 , 
    n1059 , 
    n1060 , 
    n1061 , 
    n1062 , 
    n1063 , 
    n1064 , 
    n1065 , 
    n1066 , 
    n1067 , 
    n1068 , 
    n1069 , 
    n1070 , 
    n1071 , 
    n1072 , 
    n1073 , 
    n1074 , 
    n1075 , 
    n1076 , 
    n1077 , 
    n1078 , 
    n1079 , 
    n1080 , 
    n1081 , 
    n1082 , 
    n1083 , 
    n1084 , 
    n1085 , 
    n1086 , 
    n1087 , 
    n1088 , 
    n1089 , 
    n1090 , 
    n1091 , 
    n1092 , 
    n1093 , 
    n1094 , 
    n1095 , 
    n1096 , 
    n1097 , 
    n1098 , 
    n1099 , 
    n1100 , 
    n1101 , 
    n1102 , 
    n1103 , 
    n1104 , 
    n1105 , 
    n1106 , 
    n1107 , 
    n1108 , 
    n1109 , 
    n1110 , 
    n1111 , 
    n1112 , 
    n1113 , 
    n1114 , 
    n1115 , 
    n1116 , 
    n1117 , 
    n1118 , 
    n1119 , 
    n1120 , 
    n1121 , 
    n1122 , 
    n1123 , 
    n1124 , 
    n1125 , 
    n1126 , 
    n1127 , 
    n1128 , 
    n1129 , 
    n1130 , 
    n1131 , 
    n1132 , 
    n1133 , 
    n1134 , 
    n1135 , 
    n1136 , 
    n1137 , 
    n1138 , 
    n1139 , 
    n1140 , 
    n1141 , 
    n1142 , 
    n1143 , 
    n1144 , 
    n1145 , 
    n1146 , 
    n1147 , 
    n1148 , 
    n1149 , 
    n1150 , 
    n1151 , 
    n1152 , 
    n1153 , 
    n1154 , 
    n1155 , 
    n1156 , 
    n1157 , 
    n1158 , 
    n1159 , 
    n1160 , 
    n1161 , 
    n1162 , 
    n1163 , 
    n1164 , 
    n1165 , 
    n1166 , 
    n1167 , 
    n1168 , 
    n1169 , 
    n1170 , 
    n1171 , 
    n1172 , 
    n1173 , 
    n1174 , 
    n1175 , 
    n1176 , 
    n1177 , 
    n1178 , 
    n1179 , 
    n1180 , 
    n1181 , 
    n1182 , 
    n1183 , 
    n1184 , 
    n1185 , 
    n1186 , 
    n1187 , 
    n1188 , 
    n1189 , 
    n1190 , 
    n1191 , 
    n1192 , 
    n1193 , 
    n1194 , 
    n1195 , 
    n1196 , 
    n1197 , 
    n1198 , 
    n1199 , 
    n1200 , 
    n1201 , 
    n1202 , 
    n1203 , 
    n1204 , 
    n1205 , 
    n1206 , 
    n1207 , 
    n1208 , 
    n1209 , 
    n1210 , 
    n1211 , 
    n1212 , 
    n1213 , 
    n1214 , 
    n1215 , 
    n1216 , 
    n1217 , 
    n1218 , 
    n1219 , 
    n1220 , 
    n1221 , 
    n1222 , 
    n1223 , 
    n1224 , 
    n1225 , 
    n1226 , 
    n1227 , 
    n1228 , 
    n1229 , 
    n1230 , 
    n1231 , 
    n1232 , 
    n1233 , 
    n1234 , 
    n1235 , 
    n1236 , 
    n1237 , 
    n1238 , 
    n1239 , 
    n1240 , 
    n1241 , 
    n1242 , 
    n1243 , 
    n1244 , 
    n1245 , 
    n1246 , 
    n1247 , 
    n1248 , 
    n1249 , 
    n1250 , 
    n1251 , 
    n1252 , 
    n1253 , 
    n1254 , 
    n1255 , 
    n1256 , 
    n1257 , 
    n1258 , 
    n1259 , 
    n1260 , 
    n1261 , 
    n1262 , 
    n1263 , 
    n1264 , 
    n1265 , 
    n1266 , 
    n1267 , 
    n1268 , 
    n1269 , 
    n1270 , 
    n1271 , 
    n1272 , 
    n1273 , 
    n1274 , 
    n1275 , 
    n1276 , 
    n1277 , 
    n1278 , 
    n1279 , 
    n1280 , 
    n1281 , 
    n1282 , 
    n1283 , 
    n1284 , 
    n1285 , 
    n1286 , 
    n1287 , 
    n1288 , 
    n1289 , 
    n1290 , 
    n1291 , 
    n1292 , 
    n1293 , 
    n1294 , 
    n1295 , 
    n1296 , 
    n1297 , 
    n1298 , 
    n1299 , 
    n1300 , 
    n1301 , 
    n1302 , 
    n1303 , 
    n1304 , 
    n1305 , 
    n1306 , 
    n1307 , 
    n1308 , 
    n1309 , 
    n1310 , 
    n1311 , 
    n1312 , 
    n1313 , 
    n1314 , 
    n1315 , 
    n1316 , 
    n1317 , 
    n1318 , 
    n1319 , 
    n1320 , 
    n1321 , 
    n1322 , 
    n1323 , 
    n1324 , 
    n1325 , 
    n1326 , 
    n1327 , 
    n1328 , 
    n1329 , 
    n1330 , 
    n1331 , 
    n1332 , 
    n1333 , 
    n1334 , 
    n1335 , 
    n1336 , 
    n1337 , 
    n1338 , 
    n1339 , 
    n1340 , 
    n1341 , 
    n1342 , 
    n1343 , 
    n1344 , 
    n1345 , 
    n1346 , 
    n1347 , 
    n1348 , 
    n1349 , 
    n1350 , 
    n1351 , 
    n1352 , 
    n1353 , 
    n1354 , 
    n1355 , 
    n1356 , 
    n1357 , 
    n1358 , 
    n1359 , 
    n1360 , 
    n1361 , 
    n1362 , 
    n1363 , 
    n1364 , 
    n1365 , 
    n1366 , 
    n1367 , 
    n1368 , 
    n1369 , 
    n1370 , 
    n1371 , 
    n1372 , 
    n1373 , 
    n1374 , 
    n1375 , 
    n1376 , 
    n1377 , 
    n1378 , 
    n1379 , 
    n1380 , 
    n1381 , 
    n1382 , 
    n1383 , 
    n1384 , 
    n1385 , 
    n1386 , 
    n1387 , 
    n1388 , 
    n1389 , 
    n1390 , 
    n1391 , 
    n1392 , 
    n1393 , 
    n1394 , 
    n1395 , 
    n1396 , 
    n1397 , 
    n1398 , 
    n1399 , 
    n1400 , 
    n1401 , 
    n1402 , 
    n1403 , 
    n1404 , 
    n1405 , 
    n1406 , 
    n1407 , 
    n1408 , 
    n1409 , 
    n1410 , 
    n1411 , 
    n1412 , 
    n1413 , 
    n1414 , 
    n1415 , 
    n1416 , 
    n1417 , 
    n1418 , 
    n1419 , 
    n1420 , 
    n1421 , 
    n1422 , 
    n1423 , 
    n1424 , 
    n1425 , 
    n1426 , 
    n1427 , 
    n1428 , 
    n1429 , 
    n1430 , 
    n1431 , 
    n1432 , 
    n1433 , 
    n1434 , 
    n1435 , 
    n1436 , 
    n1437 , 
    n1438 , 
    n1439 , 
    n1440 , 
    n1441 , 
    n1442 , 
    n1443 , 
    n1444 , 
    n1445 , 
    n1446 , 
    n1447 , 
    n1448 , 
    n1449 , 
    n1450 , 
    n1451 , 
    n1452 , 
    n1453 , 
    n1454 , 
    n1455 , 
    n1456 , 
    n1457 , 
    n1458 , 
    n1459 , 
    n1460 , 
    n1461 , 
    n1462 , 
    n1463 , 
    n1464 , 
    n1465 , 
    n1466 , 
    n1467 , 
    n1468 , 
    n1469 , 
    n1470 , 
    n1471 , 
    n1472 , 
    n1473 , 
    n1474 , 
    n1475 , 
    n1476 , 
    n1477 , 
    n1478 , 
    n1479 , 
    n1480 , 
    n1481 , 
    n1482 , 
    n1483 , 
    n1484 , 
    n1485 , 
    n1486 , 
    n1487 , 
    n1488 , 
    n1489 , 
    n1490 , 
    n1491 , 
    n1492 , 
    n1493 , 
    n1494 , 
    n1495 , 
    n1496 , 
    n1497 , 
    n1498 , 
    n1499 , 
    n1500 , 
    n1501 , 
    n1502 , 
    n1503 , 
    n1504 , 
    n1505 , 
    n1506 , 
    n1507 , 
    n1508 , 
    n1509 , 
    n1510 , 
    n1511 , 
    n1512 , 
    n1513 , 
    n1514 , 
    n1515 , 
    n1516 , 
    n1517 , 
    n1518 , 
    n1519 , 
    n1520 , 
    n1521 , 
    n1522 , 
    n1523 , 
    n1524 , 
    n1525 , 
    n1526 , 
    n1527 , 
    n1528 , 
    n1529 , 
    n1530 , 
    n1531 , 
    n1532 , 
    n1533 , 
    n1534 , 
    n1535 , 
    n1536 , 
    n1537 , 
    n1538 , 
    n1539 , 
    n1540 , 
    n1541 , 
    n1542 , 
    n1543 , 
    n1544 , 
    n1545 , 
    n1546 , 
    n1547 , 
    n1548 , 
    n1549 , 
    n1550 , 
    n1551 , 
    n1552 , 
    n1553 , 
    n1554 , 
    n1555 , 
    n1556 , 
    n1557 , 
    n1558 , 
    n1559 , 
    n1560 , 
    n1561 , 
    n1562 , 
    n1563 , 
    n1564 , 
    n1565 , 
    n1566 , 
    n1567 , 
    n1568 , 
    n1569 , 
    n1570 , 
    n1571 , 
    n1572 , 
    n1573 , 
    n1574 , 
    n1575 , 
    n1576 , 
    n1577 , 
    n1578 , 
    n1579 , 
    n1580 , 
    n1581 , 
    n1582 , 
    n1583 , 
    n1584 , 
    n1585 , 
    n1586 , 
    n1587 , 
    n1588 , 
    n1589 , 
    n1590 , 
    n1591 , 
    n1592 , 
    n1593 , 
    n1594 , 
    n1595 , 
    n1596 , 
    n1597 , 
    n1598 , 
    n1599 , 
    n1600 , 
    n1601 , 
    n1602 , 
    n1603 , 
    n1604 , 
    n1605 , 
    n1606 , 
    n1607 , 
    n1608 , 
    n1609 , 
    n1610 , 
    n1611 , 
    n1612 , 
    n1613 , 
    n1614 , 
    n1615 , 
    n1616 , 
    n1617 , 
    n1618 , 
    n1619 , 
    n1620 , 
    n1621 , 
    n1622 , 
    n1623 , 
    n1624 , 
    n1625 , 
    n1626 , 
    n1627 , 
    n1628 , 
    n1629 , 
    n1630 , 
    n1631 , 
    n1632 , 
    n1633 , 
    n1634 , 
    n1635 , 
    n1636 , 
    n1637 , 
    n1638 , 
    n1639 , 
    n1640 , 
    n1641 , 
    n1642 , 
    n1643 , 
    n1644 , 
    n1645 , 
    n1646 , 
    n1647 , 
    n1648 , 
    n1649 , 
    n1650 , 
    n1651 , 
    n1652 , 
    n1653 , 
    n1654 , 
    n1655 , 
    n1656 , 
    n1657 , 
    n1658 , 
    n1659 , 
    n1660 , 
    n1661 , 
    n1662 , 
    n1663 , 
    n1664 , 
    n1665 , 
    n1666 , 
    n1667 , 
    n1668 , 
    n1669 , 
    n1670 , 
    n1671 , 
    n1672 , 
    n1673 , 
    n1674 , 
    n1675 , 
    n1676 , 
    n1677 , 
    n1678 , 
    n1679 , 
    n1680 , 
    n1681 , 
    n1682 , 
    n1683 , 
    n1684 , 
    n1685 , 
    n1686 , 
    n1687 , 
    n1688 , 
    n1689 , 
    n1690 , 
    n1691 , 
    n1692 , 
    n1693 , 
    n1694 , 
    n1695 , 
    n1696 , 
    n1697 , 
    n1698 , 
    n1699 , 
    n1700 , 
    n1701 , 
    n1702 , 
    n1703 , 
    n1704 , 
    n1705 , 
    n1706 , 
    n1707 , 
    n1708 , 
    n1709 , 
    n1710 , 
    n1711 , 
    n1712 , 
    n1713 , 
    n1714 , 
    n1715 , 
    n1716 , 
    n1717 , 
    n1718 , 
    n1719 , 
    n1720 , 
    n1721 , 
    n1722 , 
    n1723 , 
    n1724 , 
    n1725 , 
    n1726 , 
    n1727 , 
    n1728 , 
    n1729 , 
    n1730 , 
    n1731 , 
    n1732 , 
    n1733 , 
    n1734 , 
    n1735 , 
    n1736 , 
    n1737 , 
    n1738 , 
    n1739 , 
    n1740 , 
    n1741 , 
    n1742 , 
    n1743 , 
    n1744 , 
    n1745 , 
    n1746 , 
    n1747 , 
    n1748 , 
    n1749 , 
    n1750 , 
    n1751 , 
    n1752 , 
    n1753 , 
    n1754 , 
    n1755 , 
    n1756 , 
    n1757 , 
    n1758 , 
    n1759 , 
    n1760 , 
    n1761 , 
    n1762 , 
    n1763 , 
    n1764 , 
    n1765 , 
    n1766 , 
    n1767 , 
    n1768 , 
    n1769 , 
    n1770 , 
    n1771 , 
    n1772 , 
    n1773 , 
    n1774 , 
    n1775 , 
    n1776 , 
    n1777 , 
    n1778 , 
    n1779 , 
    n1780 , 
    n1781 , 
    n1782 , 
    n1783 , 
    n1784 , 
    n1785 , 
    n1786 , 
    n1787 , 
    n1788 , 
    n1789 , 
    n1790 , 
    n1791 , 
    n1792 , 
    n1793 , 
    n1794 , 
    n1795 , 
    n1796 , 
    n1797 , 
    n1798 , 
    n1799 , 
    n1800 , 
    n1801 , 
    n1802 , 
    n1803 , 
    n1804 , 
    n1805 , 
    n1806 , 
    n1807 , 
    n1808 , 
    n1809 , 
    n1810 , 
    n1811 , 
    n1812 , 
    n1813 , 
    n1814 , 
    n1815 , 
    n1816 , 
    n1817 , 
    n1818 , 
    n1819 , 
    n1820 , 
    n1821 , 
    n1822 , 
    n1823 , 
    n1824 , 
    n1825 , 
    n1826 , 
    n1827 , 
    n1828 , 
    n1829 , 
    n1830 , 
    n1831 , 
    n1832 , 
    n1833 , 
    n1834 , 
    n1835 , 
    n1836 , 
    n1837 , 
    n1838 , 
    n1839 , 
    n1840 , 
    n1841 , 
    n1842 , 
    n1843 , 
    n1844 , 
    n1845 , 
    n1846 , 
    n1847 , 
    n1848 , 
    n1849 , 
    n1850 , 
    n1851 , 
    n1852 , 
    n1853 , 
    n1854 , 
    n1855 , 
    n1856 , 
    n1857 , 
    n1858 , 
    n1859 , 
    n1860 , 
    n1861 , 
    n1862 , 
    n1863 , 
    n1864 , 
    n1865 , 
    n1866 , 
    n1867 , 
    n1868 , 
    n1869 , 
    n1870 , 
    n1871 , 
    n1872 , 
    n1873 , 
    n1874 , 
    n1875 , 
    n1876 , 
    n1877 , 
    n1878 , 
    n1879 , 
    n1880 , 
    n1881 , 
    n1882 , 
    n1883 , 
    n1884 , 
    n1885 , 
    n1886 , 
    n1887 , 
    n1888 , 
    n1889 , 
    n1890 , 
    n1891 , 
    n1892 , 
    n1893 , 
    n1894 , 
    n1895 , 
    n1896 , 
    n1897 , 
    n1898 , 
    n1899 , 
    n1900 , 
    n1901 , 
    n1902 , 
    n1903 , 
    n1904 , 
    n1905 , 
    n1906 , 
    n1907 , 
    n1908 , 
    n1909 , 
    n1910 , 
    n1911 , 
    n1912 , 
    n1913 , 
    n1914 , 
    n1915 , 
    n1916 , 
    n1917 , 
    n1918 , 
    n1919 , 
    n1920 , 
    n1921 , 
    n1922 , 
    n1923 , 
    n1924 , 
    n1925 , 
    n1926 , 
    n1927 , 
    n1928 , 
    n1929 , 
    n1930 , 
    n1931 , 
    n1932 , 
    n1933 , 
    n1934 , 
    n1935 , 
    n1936 , 
    n1937 , 
    n1938 , 
    n1939 , 
    n1940 , 
    n1941 , 
    n1942 , 
    n1943 , 
    n1944 , 
    n1945 , 
    n1946 , 
    n1947 , 
    n1948 , 
    n1949 , 
    n1950 , 
    n1951 , 
    n1952 , 
    n1953 , 
    n1954 , 
    n1955 , 
    n1956 , 
    n1957 , 
    n1958 , 
    n1959 , 
    n1960 , 
    n1961 , 
    n1962 , 
    n1963 , 
    n1964 , 
    n1965 , 
    n1966 , 
    n1967 , 
    n1968 , 
    n1969 , 
    n1970 , 
    n1971 , 
    n1972 , 
    n1973 , 
    n1974 , 
    n1975 , 
    n1976 , 
    n1977 , 
    n1978 , 
    n1979 , 
    n1980 , 
    n1981 , 
    n1982 , 
    n1983 , 
    n1984 , 
    n1985 , 
    n1986 , 
    n1987 , 
    n1988 , 
    n1989 , 
    n1990 , 
    n1991 , 
    n1992 , 
    n1993 , 
    n1994 , 
    n1995 , 
    n1996 , 
    n1997 , 
    n1998 , 
    n1999 , 
    n2000 , 
    n2001 , 
    n2002 , 
    n2003 , 
    n2004 , 
    n2005 , 
    n2006 , 
    n2007 , 
    n2008 , 
    n2009 , 
    n2010 , 
    n2011 , 
    n2012 , 
    n2013 , 
    n2014 , 
    n2015 , 
    n2016 , 
    n2017 , 
    n2018 , 
    n2019 , 
    n2020 , 
    n2021 , 
    n2022 , 
    n2023 , 
    n2024 , 
    n2025 , 
    n2026 , 
    n2027 , 
    n2028 , 
    n2029 , 
    n2030 , 
    n2031 , 
    n2032 , 
    n2033 , 
    n2034 , 
    n2035 , 
    n2036 , 
    n2037 , 
    n2038 , 
    n2039 , 
    n2040 , 
    n2041 , 
    n2042 , 
    n2043 , 
    n2044 , 
    n2045 , 
    n2046 , 
    n2047 , 
    n2048 , 
    n2049 , 
    n2050 , 
    n2051 , 
    n2052 , 
    n2053 , 
    n2054 , 
    n2055 , 
    n2056 , 
    n2057 , 
    n2058 , 
    n2059 , 
    n2060 , 
    n2061 , 
    n2062 , 
    n2063 , 
    n2064 , 
    n2065 , 
    n2066 , 
    n2067 , 
    n2068 , 
    n2069 , 
    n2070 , 
    n2071 , 
    n2072 , 
    n2073 , 
    n2074 , 
    n2075 , 
    n2076 , 
    n2077 , 
    n2078 , 
    n2079 , 
    n2080 , 
    n2081 , 
    n2082 , 
    n2083 , 
    n2084 , 
    n2085 , 
    n2086 , 
    n2087 , 
    n2088 , 
    n2089 , 
    n2090 , 
    n2091 , 
    n2092 , 
    n2093 , 
    n2094 , 
    n2095 , 
    n2096 , 
    n2097 , 
    n2098 , 
    n2099 , 
    n2100 , 
    n2101 , 
    n2102 , 
    n2103 , 
    n2104 , 
    n2105 , 
    n2106 , 
    n2107 , 
    n2108 , 
    n2109 , 
    n2110 , 
    n2111 , 
    n2112 , 
    n2113 , 
    n2114 , 
    n2115 , 
    n2116 , 
    n2117 , 
    n2118 , 
    n2119 , 
    n2120 , 
    n2121 , 
    n2122 , 
    n2123 , 
    n2124 , 
    n2125 , 
    n2126 , 
    n2127 , 
    n2128 , 
    n2129 , 
    n2130 , 
    n2131 , 
    n2132 , 
    n2133 , 
    n2134 , 
    n2135 , 
    n2136 , 
    n2137 , 
    n2138 , 
    n2139 , 
    n2140 , 
    n2141 , 
    n2142 , 
    n2143 , 
    n2144 , 
    n2145 , 
    n2146 , 
    n2147 , 
    n2148 , 
    n2149 , 
    n2150 , 
    n2151 , 
    n2152 , 
    n2153 , 
    n2154 , 
    n2155 , 
    n2156 , 
    n2157 , 
    n2158 , 
    n2159 , 
    n2160 , 
    n2161 , 
    n2162 , 
    n2163 , 
    n2164 , 
    n2165 , 
    n2166 , 
    n2167 , 
    n2168 , 
    n2169 , 
    n2170 , 
    n2171 , 
    n2172 , 
    n2173 , 
    n2174 , 
    n2175 , 
    n2176 , 
    n2177 , 
    n2178 , 
    n2179 , 
    n2180 , 
    n2181 , 
    n2182 , 
    n2183 , 
    n2184 , 
    n2185 , 
    n2186 , 
    n2187 , 
    n2188 , 
    n2189 , 
    n2190 , 
    n2191 , 
    n2192 , 
    n2193 , 
    n2194 , 
    n2195 , 
    n2196 , 
    n2197 , 
    n2198 , 
    n2199 , 
    n2200 , 
    n2201 , 
    n2202 , 
    n2203 , 
    n2204 , 
    n2205 , 
    n2206 , 
    n2207 , 
    n2208 , 
    n2209 , 
    n2210 , 
    n2211 , 
    n2212 , 
    n2213 , 
    n2214 , 
    n2215 , 
    n2216 , 
    n2217 , 
    n2218 , 
    n2219 , 
    n2220 , 
    n2221 , 
    n2222 , 
    n2223 , 
    n2224 , 
    n2225 , 
    n2226 , 
    n2227 , 
    n2228 , 
    n2229 , 
    n2230 , 
    n2231 , 
    n2232 , 
    n2233 , 
    n2234 , 
    n2235 , 
    n2236 , 
    n2237 , 
    n2238 , 
    n2239 , 
    n2240 , 
    n2241 , 
    n2242 , 
    n2243 , 
    n2244 , 
    n2245 , 
    n2246 , 
    n2247 , 
    n2248 , 
    n2249 , 
    n2250 , 
    n2251 , 
    n2252 , 
    n2253 , 
    n2254 , 
    n2255 , 
    n2256 , 
    n2257 , 
    n2258 , 
    n2259 , 
    n2260 , 
    n2261 , 
    n2262 , 
    n2263 , 
    n2264 , 
    n2265 , 
    n2266 , 
    n2267 , 
    n2268 , 
    n2269 , 
    n2270 , 
    n2271 , 
    n2272 , 
    n2273 , 
    n2274 , 
    n2275 , 
    n2276 , 
    n2277 , 
    n2278 , 
    n2279 , 
    n2280 , 
    n2281 , 
    n2282 , 
    n2283 , 
    n2284 , 
    n2285 , 
    n2286 , 
    n2287 , 
    n2288 , 
    n2289 , 
    n2290 , 
    n2291 , 
    n2292 , 
    n2293 , 
    n2294 , 
    n2295 , 
    n2296 , 
    n2297 , 
    n2298 , 
    n2299 , 
    n2300 , 
    n2301 , 
    n2302 , 
    n2303 , 
    n2304 , 
    n2305 , 
    n2306 , 
    n2307 , 
    n2308 , 
    n2309 , 
    n2310 , 
    n2311 , 
    n2312 , 
    n2313 , 
    n2314 , 
    n2315 , 
    n2316 , 
    n2317 , 
    n2318 , 
    n2319 , 
    n2320 , 
    n2321 , 
    n2322 , 
    n2323 , 
    n2324 , 
    n2325 , 
    n2326 , 
    n2327 , 
    n2328 , 
    n2329 , 
    n2330 , 
    n2331 , 
    n2332 , 
    n2333 , 
    n2334 , 
    n2335 , 
    n2336 , 
    n2337 , 
    n2338 , 
    n2339 , 
    n2340 , 
    n2341 , 
    n2342 , 
    n2343 , 
    n2344 , 
    n2345 , 
    n2346 , 
    n2347 , 
    n2348 , 
    n2349 , 
    n2350 , 
    n2351 , 
    n2352 , 
    n2353 , 
    n2354 , 
    n2355 , 
    n2356 , 
    n2357 , 
    n2358 , 
    n2359 , 
    n2360 , 
    n2361 , 
    n2362 , 
    n2363 , 
    n2364 , 
    n2365 , 
    n2366 , 
    n2367 , 
    n2368 , 
    n2369 , 
    n2370 , 
    n2371 , 
    n2372 , 
    n2373 , 
    n2374 , 
    n2375 , 
    n2376 , 
    n2377 , 
    n2378 , 
    n2379 , 
    n2380 , 
    n2381 , 
    n2382 , 
    n2383 , 
    n2384 , 
    n2385 , 
    n2386 , 
    n2387 , 
    n2388 , 
    n2389 , 
    n2390 , 
    n2391 , 
    n2392 , 
    n2393 , 
    n2394 , 
    n2395 , 
    n2396 , 
    n2397 , 
    n2398 , 
    n2399 , 
    n2400 , 
    n2401 , 
    n2402 , 
    n2403 , 
    n2404 , 
    n2405 , 
    n2406 , 
    n2407 , 
    n2408 , 
    n2409 , 
    n2410 , 
    n2411 , 
    n2412 , 
    n2413 , 
    n2414 , 
    n2415 , 
    n2416 , 
    n2417 , 
    n2418 , 
    n2419 , 
    n2420 , 
    n2421 , 
    n2422 , 
    n2423 , 
    n2424 , 
    n2425 , 
    n2426 , 
    n2427 , 
    n2428 , 
    n2429 , 
    n2430 , 
    n2431 , 
    n2432 , 
    n2433 , 
    n2434 , 
    n2435 , 
    n2436 , 
    n2437 , 
    n2438 , 
    n2439 , 
    n2440 , 
    n2441 , 
    n2442 , 
    n2443 , 
    n2444 , 
    n2445 , 
    n2446 , 
    n2447 , 
    n2448 , 
    n2449 , 
    n2450 , 
    n2451 , 
    n2452 , 
    n2453 , 
    n2454 , 
    n2455 , 
    n2456 , 
    n2457 , 
    n2458 , 
    n2459 , 
    n2460 , 
    n2461 , 
    n2462 , 
    n2463 , 
    n2464 , 
    n2465 , 
    n2466 , 
    n2467 , 
    n2468 , 
    n2469 , 
    n2470 , 
    n2471 , 
    n2472 , 
    n2473 , 
    n2474 , 
    n2475 , 
    n2476 , 
    n2477 , 
    n2478 , 
    n2479 , 
    n2480 , 
    n2481 , 
    n2482 , 
    n2483 , 
    n2484 , 
    n2485 , 
    n2486 , 
    n2487 , 
    n2488 , 
    n2489 , 
    n2490 , 
    n2491 , 
    n2492 , 
    n2493 , 
    n2494 , 
    n2495 , 
    n2496 , 
    n2497 , 
    n2498 , 
    n2499 , 
    n2500 , 
    n2501 , 
    n2502 , 
    n2503 , 
    n2504 , 
    n2505 , 
    n2506 , 
    n2507 , 
    n2508 , 
    n2509 , 
    n2510 , 
    n2511 , 
    n2512 , 
    n2513 , 
    n2514 , 
    n2515 , 
    n2516 , 
    n2517 , 
    n2518 , 
    n2519 , 
    n2520 , 
    n2521 , 
    n2522 , 
    n2523 , 
    n2524 , 
    n2525 , 
    n2526 , 
    n2527 , 
    n2528 , 
    n2529 , 
    n2530 , 
    n2531 , 
    n2532 , 
    n2533 , 
    n2534 , 
    n2535 , 
    n2536 , 
    n2537 , 
    n2538 , 
    n2539 , 
    n2540 , 
    n2541 , 
    n2542 , 
    n2543 , 
    n2544 , 
    n2545 , 
    n2546 , 
    n2547 , 
    n2548 , 
    n2549 , 
    n2550 , 
    n2551 , 
    n2552 , 
    n2553 , 
    n2554 , 
    n2555 , 
    n2556 , 
    n2557 , 
    n2558 , 
    n2559 , 
    n2560 , 
    n2561 , 
    n2562 , 
    n2563 , 
    n2564 , 
    n2565 , 
    n2566 , 
    n2567 , 
    n2568 , 
    n2569 , 
    n2570 , 
    n2571 , 
    n2572 , 
    n2573 , 
    n2574 , 
    n2575 , 
    n2576 , 
    n2577 , 
    n2578 , 
    n2579 , 
    n2580 , 
    n2581 , 
    n2582 , 
    n2583 , 
    n2584 , 
    n2585 , 
    n2586 , 
    n2587 , 
    n2588 , 
    n2589 , 
    n2590 , 
    n2591 , 
    n2592 , 
    n2593 , 
    n2594 , 
    n2595 , 
    n2596 , 
    n2597 , 
    n2598 , 
    n2599 , 
    n2600 , 
    n2601 , 
    n2602 , 
    n2603 , 
    n2604 , 
    n2605 , 
    n2606 , 
    n2607 , 
    n2608 , 
    n2609 , 
    n2610 , 
    n2611 , 
    n2612 , 
    n2613 , 
    n2614 , 
    n2615 , 
    n2616 , 
    n2617 , 
    n2618 , 
    n2619 , 
    n2620 , 
    n2621 , 
    n2622 , 
    n2623 , 
    n2624 , 
    n2625 , 
    n2626 , 
    n2627 , 
    n2628 , 
    n2629 , 
    n2630 , 
    n2631 , 
    n2632 , 
    n2633 , 
    n2634 , 
    n2635 , 
    n2636 , 
    n2637 , 
    n2638 , 
    n2639 , 
    n2640 , 
    n2641 , 
    n2642 , 
    n2643 , 
    n2644 , 
    n2645 , 
    n2646 , 
    n2647 , 
    n2648 , 
    n2649 , 
    n2650 , 
    n2651 , 
    n2652 , 
    n2653 , 
    n2654 , 
    n2655 , 
    n2656 , 
    n2657 , 
    n2658 , 
    n2659 , 
    n2660 , 
    n2661 , 
    n2662 , 
    n2663 , 
    n2664 , 
    n2665 , 
    n2666 , 
    n2667 , 
    n2668 , 
    n2669 , 
    n2670 , 
    n2671 , 
    n2672 , 
    n2673 , 
    n2674 , 
    n2675 , 
    n2676 , 
    n2677 , 
    n2678 , 
    n2679 , 
    n2680 , 
    n2681 , 
    n2682 , 
    n2683 , 
    n2684 , 
    n2685 , 
    n2686 , 
    n2687 , 
    n2688 , 
    n2689 , 
    n2690 , 
    n2691 , 
    n2692 , 
    n2693 , 
    n2694 , 
    n2695 , 
    n2696 , 
    n2697 , 
    n2698 , 
    n2699 , 
    n2700 , 
    n2701 , 
    n2702 , 
    n2703 , 
    n2704 , 
    n2705 , 
    n2706 , 
    n2707 , 
    n2708 , 
    n2709 , 
    n2710 , 
    n2711 , 
    n2712 , 
    n2713 , 
    n2714 , 
    n2715 , 
    n2716 , 
    n2717 , 
    n2718 , 
    n2719 , 
    n2720 , 
    n2721 , 
    n2722 , 
    n2723 , 
    n2724 , 
    n2725 , 
    n2726 , 
    n2727 , 
    n2728 , 
    n2729 , 
    n2730 , 
    n2731 , 
    n2732 , 
    n2733 , 
    n2734 , 
    n2735 , 
    n2736 , 
    n2737 , 
    n2738 , 
    n2739 , 
    n2740 , 
    n2741 , 
    n2742 , 
    n2743 , 
    n2744 , 
    n2745 , 
    n2746 , 
    n2747 , 
    n2748 , 
    n2749 , 
    n2750 , 
    n2751 , 
    n2752 , 
    n2753 , 
    n2754 , 
    n2755 , 
    n2756 , 
    n2757 , 
    n2758 , 
    n2759 , 
    n2760 , 
    n2761 , 
    n2762 , 
    n2763 , 
    n2764 , 
    n2765 , 
    n2766 , 
    n2767 , 
    n2768 , 
    n2769 , 
    n2770 , 
    n2771 , 
    n2772 , 
    n2773 , 
    n2774 , 
    n2775 , 
    n2776 , 
    n2777 , 
    n2778 , 
    n2779 , 
    n2780 , 
    n2781 , 
    n2782 , 
    n2783 , 
    n2784 , 
    n2785 , 
    n2786 , 
    n2787 , 
    n2788 , 
    n2789 , 
    n2790 , 
    n2791 , 
    n2792 , 
    n2793 , 
    n2794 , 
    n2795 , 
    n2796 , 
    n2797 , 
    n2798 , 
    n2799 , 
    n2800 , 
    n2801 , 
    n2802 , 
    n2803 , 
    n2804 , 
    n2805 , 
    n2806 , 
    n2807 , 
    n2808 , 
    n2809 , 
    n2810 , 
    n2811 , 
    n2812 , 
    n2813 , 
    n2814 , 
    n2815 , 
    n2816 , 
    n2817 , 
    n2818 , 
    n2819 , 
    n2820 , 
    n2821 , 
    n2822 , 
    n2823 , 
    n2824 , 
    n2825 , 
    n2826 , 
    n2827 , 
    n2828 , 
    n2829 , 
    n2830 , 
    n2831 , 
    n2832 , 
    n2833 , 
    n2834 , 
    n2835 , 
    n2836 , 
    n2837 , 
    n2838 , 
    n2839 , 
    n2840 , 
    n2841 , 
    n2842 , 
    n2843 , 
    n2844 , 
    n2845 , 
    n2846 , 
    n2847 , 
    n2848 , 
    n2849 , 
    n2850 , 
    n2851 , 
    n2852 , 
    n2853 , 
    n2854 , 
    n2855 , 
    n2856 , 
    n2857 , 
    n2858 , 
    n2859 , 
    n2860 , 
    n2861 , 
    n2862 , 
    n2863 , 
    n2864 , 
    n2865 , 
    n2866 , 
    n2867 , 
    n2868 , 
    n2869 , 
    n2870 , 
    n2871 , 
    n2872 , 
    n2873 , 
    n2874 , 
    n2875 , 
    n2876 , 
    n2877 , 
    n2878 , 
    n2879 , 
    n2880 , 
    n2881 , 
    n2882 , 
    n2883 , 
    n2884 , 
    n2885 , 
    n2886 , 
    n2887 , 
    n2888 , 
    n2889 , 
    n2890 , 
    n2891 , 
    n2892 , 
    n2893 , 
    n2894 , 
    n2895 , 
    n2896 , 
    n2897 , 
    n2898 , 
    n2899 , 
    n2900 , 
    n2901 , 
    n2902 , 
    n2903 , 
    n2904 , 
    n2905 , 
    n2906 , 
    n2907 , 
    n2908 , 
    n2909 , 
    n2910 , 
    n2911 , 
    n2912 , 
    n2913 , 
    n2914 , 
    n2915 , 
    n2916 , 
    n2917 , 
    n2918 , 
    n2919 , 
    n2920 , 
    n2921 , 
    n2922 , 
    n2923 , 
    n2924 , 
    n2925 , 
    n2926 , 
    n2927 , 
    n2928 , 
    n2929 , 
    n2930 , 
    n2931 , 
    n2932 , 
    n2933 , 
    n2934 , 
    n2935 , 
    n2936 , 
    n2937 , 
    n2938 , 
    n2939 , 
    n2940 , 
    n2941 , 
    n2942 , 
    n2943 , 
    n2944 , 
    n2945 , 
    n2946 , 
    n2947 , 
    n2948 , 
    n2949 , 
    n2950 , 
    n2951 , 
    n2952 , 
    n2953 , 
    n2954 , 
    n2955 , 
    n2956 , 
    n2957 , 
    n2958 , 
    n2959 , 
    n2960 , 
    n2961 , 
    n2962 , 
    n2963 , 
    n2964 , 
    n2965 , 
    n2966 , 
    n2967 , 
    n2968 , 
    n2969 , 
    n2970 , 
    n2971 , 
    n2972 , 
    n2973 , 
    n2974 , 
    n2975 , 
    n2976 , 
    n2977 , 
    n2978 , 
    n2979 , 
    n2980 , 
    n2981 , 
    n2982 , 
    n2983 , 
    n2984 , 
    n2985 , 
    n2986 , 
    n2987 , 
    n2988 , 
    n2989 , 
    n2990 , 
    n2991 , 
    n2992 , 
    n2993 , 
    n2994 , 
    n2995 , 
    n2996 , 
    n2997 , 
    n2998 , 
    n2999 , 
    n3000 , 
    n3001 , 
    n3002 , 
    n3003 , 
    n3004 , 
    n3005 , 
    n3006 , 
    n3007 , 
    n3008 , 
    n3009 , 
    n3010 , 
    n3011 , 
    n3012 , 
    n3013 , 
    n3014 , 
    n3015 , 
    n3016 , 
    n3017 , 
    n3018 , 
    n3019 , 
    n3020 , 
    n3021 , 
    n3022 , 
    n3023 , 
    n3024 , 
    n3025 , 
    n3026 , 
    n3027 , 
    n3028 , 
    n3029 , 
    n3030 , 
    n3031 , 
    n3032 , 
    n3033 , 
    n3034 , 
    n3035 , 
    n3036 , 
    n3037 , 
    n3038 , 
    n3039 , 
    n3040 , 
    n3041 , 
    n3042 , 
    n3043 , 
    n3044 , 
    n3045 , 
    n3046 , 
    n3047 , 
    n3048 , 
    n3049 , 
    n3050 , 
    n3051 , 
    n3052 , 
    n3053 , 
    n3054 , 
    n3055 , 
    n3056 , 
    n3057 , 
    n3058 , 
    n3059 , 
    n3060 , 
    n3061 , 
    n3062 , 
    n3063 , 
    n3064 , 
    n3065 , 
    n3066 , 
    n3067 , 
    n3068 , 
    n3069 , 
    n3070 , 
    n3071 , 
    n3072 , 
    n3073 , 
    n3074 , 
    n3075 , 
    n3076 , 
    n3077 , 
    n3078 , 
    n3079 , 
    n3080 , 
    n3081 , 
    n3082 , 
    n3083 , 
    n3084 , 
    n3085 , 
    n3086 , 
    n3087 , 
    n3088 , 
    n3089 , 
    n3090 , 
    n3091 , 
    n3092 , 
    n3093 , 
    n3094 , 
    n3095 , 
    n3096 , 
    n3097 , 
    n3098 , 
    n3099 , 
    n3100 , 
    n3101 , 
    n3102 , 
    n3103 , 
    n3104 , 
    n3105 , 
    n3106 , 
    n3107 , 
    n3108 , 
    n3109 , 
    n3110 , 
    n3111 , 
    n3112 , 
    n3113 , 
    n3114 , 
    n3115 , 
    n3116 , 
    n3117 , 
    n3118 , 
    n3119 , 
    n3120 , 
    n3121 , 
    n3122 , 
    n3123 ;

wire  C0 , C1 , RI21a19c60_2 , 
    RI21a5daf0_1 , 
    RI2107e620_463 , 
    RI21a139f0_68 , 
    RI21084368_418 , 
    RI21079850_497 , 
    RI21a12820_78 , 
    RI210beb08_292 , 
    RI21a12898_77 , 
    RI210beb80_291 , 
    RI21a12910_76 , 
    RI210bf3f0_290 , 
    RI21a12988_75 , 
    RI210bf468_289 , 
    RI21a13090_74 , 
    RI210bf4e0_288 , 
    RI21a13108_73 , 
    RI210bf558_287 , 
    RI21a13180_72 , 
    RI210bfdc8_286 , 
    RI21a131f8_71 , 
    RI210bfe40_285 , 
    RI21a13270_70 , 
    RI210bfeb8_284 , 
    RI21a132e8_69 , 
    RI210bff30_283 , 
    RI21a116c8_87 , 
    RI210bd6e0_301 , 
    RI21a11dd0_86 , 
    RI210bd758_300 , 
    RI21a11e48_85 , 
    RI210bd7d0_299 , 
    RI21a11ec0_84 , 
    RI210be040_298 , 
    RI21a11f38_83 , 
    RI210be0b8_297 , 
    RI21a11fb0_82 , 
    RI210be130_296 , 
    RI21a12028_81 , 
    RI210be1a8_295 , 
    RI21a12730_80 , 
    RI210bea18_294 , 
    RI21a127a8_79 , 
    RI210bea90_293 , 
    RI21077f00_507 , 
    RI21077f78_506 , 
    RI21078a40_505 , 
    RI21078ab8_504 , 
    RI21078b30_503 , 
    RI21078ba8_502 , 
    RI21078c20_501 , 
    RI21078c98_500 , 
    RI21079760_499 , 
    RI210797d8_498 , 
    RI21077078_516 , 
    RI210770f0_515 , 
    RI21077168_514 , 
    RI210771e0_513 , 
    RI21077258_512 , 
    RI21077d20_511 , 
    RI21077d98_510 , 
    RI21077e10_509 , 
    RI21077e88_508 , 
    RI2107a660_489 , 
    RI2107a6d8_488 , 
    RI2107b218_486 , 
    RI2107b290_485 , 
    RI2107b308_484 , 
    RI2107b380_483 , 
    RI2107b3f8_482 , 
    RI2107bec0_481 , 
    RI2107bf38_480 , 
    RI2107bfb0_479 , 
    RI2107c028_478 , 
    RI2107c0a0_477 , 
    RI2107cbe0_475 , 
    RI2107cc58_474 , 
    RI2107ccd0_473 , 
    RI2107cd48_472 , 
    RI2107cdc0_471 , 
    RI2107ce38_470 , 
    RI2107d900_469 , 
    RI2107d978_468 , 
    RI2107d9f0_467 , 
    RI2107da68_466 , 
    RI210798c8_496 , 
    RI21079940_495 , 
    RI210799b8_494 , 
    RI2107a480_493 , 
    RI2107a4f8_492 , 
    RI2107a570_491 , 
    RI2107a5e8_490 , 
    RI2107b1a0_487 , 
    RI2107c118_476 , 
    RI2106bde0_608 , 
    GI20478f00_682 , 
    RI2106c0b0_602 , 
    RI2106c128_601 , 
    RI2106c1a0_600 , 
    RI2106c218_599 , 
    RI2106c290_598 , 
    RI2106a238_641 , 
    RI2106a2b0_640 , 
    RI2106a328_639 , 
    RI2106a3a0_638 , 
    RI2106a490_636 , 
    RI2106a508_635 , 
    RI2106a580_634 , 
    RI2106c308_597 , 
    RI2106a5f8_633 , 
    RI2106a670_632 , 
    RI2106a6e8_631 , 
    RI2106a760_630 , 
    RI2106a7d8_629 , 
    RI2106ae68_628 , 
    RI21069a40_645 , 
    RI2106bed0_606 , 
    RI21069ab8_644 , 
    RI2106bf48_605 , 
    RI2106bfc0_604 , 
    RI2106c038_603 , 
    RI2106a148_643 , 
    RI2106a1c0_642 , 
    RI2106a418_637 , 
    RI2106c380_596 , 
    RI2106cbf0_591 , 
    RI2106dd48_567 , 
    RI21073040_543 , 
    RI2106cd58_588 , 
    RI2106deb0_564 , 
    RI21073c70_539 , 
    RI2106cdd0_587 , 
    RI2106df28_563 , 
    RI21073ce8_538 , 
    RI2106ce48_586 , 
    RI2106dfa0_562 , 
    RI21073d60_537 , 
    RI2106cec0_585 , 
    RI2106e018_561 , 
    RI21073dd8_536 , 
    RI2106cf38_584 , 
    RI2106e090_560 , 
    RI210748a0_535 , 
    RI2106cfb0_583 , 
    RI2106e108_559 , 
    RI21074918_534 , 
    RI2106d028_582 , 
    RI21070a48_558 , 
    RI21074990_533 , 
    RI2106d0a0_581 , 
    RI21070ac0_557 , 
    RI21074a08_532 , 
    RI2106d118_580 , 
    RI21071588_556 , 
    RI21074a80_531 , 
    RI2106b138_622 , 
    RI2106b4f8_614 , 
    RI210755c0_529 , 
    RI2106b1b0_621 , 
    RI2106b570_613 , 
    RI21075638_528 , 
    RI2106b228_620 , 
    RI2106bc00_612 , 
    RI210756b0_527 , 
    RI2106d190_579 , 
    RI21071600_555 , 
    RI21075728_526 , 
    RI2106d208_578 , 
    RI21071678_554 , 
    RI210757a0_525 , 
    RI2106d898_577 , 
    RI2106bc78_611 , 
    RI21075818_524 , 
    RI2106d910_576 , 
    RI2106bcf0_610 , 
    RI210762e0_523 , 
    RI2106d988_575 , 
    RI210716f0_553 , 
    RI21076358_522 , 
    RI2106da00_574 , 
    RI210721b8_552 , 
    RI210763d0_521 , 
    RI2106da78_573 , 
    RI2106bd68_609 , 
    RI21076448_520 , 
    RI2106ca10_595 , 
    RI2106db68_571 , 
    RI210722a8_550 , 
    RI2106ca88_594 , 
    RI2106dbe0_570 , 
    RI21072320_549 , 
    RI2106aee0_627 , 
    RI2106dc58_569 , 
    RI21072398_548 , 
    RI2106af58_626 , 
    RI2106dcd0_568 , 
    RI21072e60_547 , 
    RI2106cb00_593 , 
    RI2106b2a0_619 , 
    RI21072ed8_546 , 
    RI2106afd0_625 , 
    RI2106b318_618 , 
    RI21072f50_545 , 
    RI2106cb78_592 , 
    RI2106b390_617 , 
    RI21072fc8_544 , 
    RI2106b048_624 , 
    RI2106b408_616 , 
    RI21073b80_541 , 
    RI2106b0c0_623 , 
    RI2106b480_615 , 
    RI21074af8_530 , 
    RI2106daf0_572 , 
    RI21072230_551 , 
    RI210764c0_519 , 
    RI2107dae0_465 , 
    RI2106cc68_590 , 
    RI2106ddc0_566 , 
    RI210730b8_542 , 
    RI21a0e608_121 , 
    RI210b87a8_334 , 
    RI21a19a08_3 , 
    RI21a0f058_113 , 
    RI210b9b58_326 , 
    RI21a0f0d0_112 , 
    RI210b9bd0_325 , 
    RI21a0f850_110 , 
    RI210b9c48_324 , 
    RI21a0f8c8_109 , 
    RI210b9cc0_323 , 
    RI21a0f940_108 , 
    RI210ba530_322 , 
    RI21a0f9b8_107 , 
    RI210ba5a8_321 , 
    RI21a0fa30_106 , 
    RI210ba620_320 , 
    RI21a0faa8_105 , 
    RI210ba698_319 , 
    RI21a101b0_104 , 
    RI210baf08_318 , 
    RI21a10228_103 , 
    RI210baf80_317 , 
    RI21a102a0_102 , 
    RI210baff8_316 , 
    RI21a10318_101 , 
    RI210bb070_315 , 
    RI21a10390_100 , 
    RI210bb8e0_314 , 
    RI21a10408_99 , 
    RI210bb958_313 , 
    RI21a10b10_98 , 
    RI210bb9d0_312 , 
    RI21a10b88_97 , 
    RI210bba48_311 , 
    RI21a10c00_96 , 
    RI210bc2b8_310 , 
    RI21a10c78_95 , 
    RI210bc330_309 , 
    RI21a10cf0_94 , 
    RI210bc3a8_308 , 
    RI21a10d68_93 , 
    RI210bc420_307 , 
    RI21a11470_92 , 
    RI210bcc90_306 , 
    RI21a114e8_91 , 
    RI210bcd08_305 , 
    RI21a0e680_120 , 
    RI210b8820_333 , 
    RI21a0e6f8_119 , 
    RI210b8898_332 , 
    RI21a0e770_118 , 
    RI210b8910_331 , 
    RI21a0e7e8_117 , 
    RI210b9180_330 , 
    RI21a0eef0_116 , 
    RI210b91f8_329 , 
    RI21a0ef68_115 , 
    RI210b9270_328 , 
    RI21a0efe0_114 , 
    RI210b92e8_327 , 
    RI21a0f148_111 , 
    RI21084278_420 , 
    RI210cfcc8_237 , 
    RI210842f0_419 , 
    RI21a11560_90 , 
    RI210bcd80_304 , 
    RI21a19990_4 , 
    RI2106cce0_589 , 
    RI2106de38_565 , 
    RI21073bf8_540 , 
    RI21a19918_5 , 
    RI21a198a0_6 , 
    RI21a19828_7 , 
    RI21a197b0_8 , 
    RI21a190a8_9 , 
    RI21a19030_10 , 
    RI21a18fb8_11 , 
    RI21a18f40_12 , 
    RI21a18ec8_13 , 
    RI21a18e50_14 , 
    RI21a18748_15 , 
    RI21a186d0_16 , 
    RI21a18658_17 , 
    RI21a185e0_18 , 
    RI21a18568_19 , 
    RI21a184f0_20 , 
    RI21a17de8_21 , 
    RI21a17d70_22 , 
    RI21a17cf8_23 , 
    RI21a17c80_24 , 
    RI21a17c08_25 , 
    RI21a17b90_26 , 
    RI21a17488_27 , 
    RI21a17410_28 , 
    RI21a17398_29 , 
    RI21a17320_30 , 
    RI21a172a8_31 , 
    RI21a17230_32 , 
    RI21a16b28_33 , 
    RI21a16ab0_34 , 
    RI2106be58_607 , 
    RI21a14440_60 , 
    RI21a144b8_59 , 
    RI21a145a8_57 , 
    RI21a14cb0_56 , 
    RI21a14d28_55 , 
    RI21a14da0_54 , 
    RI21a14e18_53 , 
    RI21a14e90_52 , 
    RI21a14f08_51 , 
    RI21a15610_50 , 
    RI21a15688_49 , 
    RI21a15700_48 , 
    RI21a157f0_46 , 
    RI21a15868_45 , 
    RI21a15f70_44 , 
    RI21a15fe8_43 , 
    RI21a16060_42 , 
    RI21a160d8_41 , 
    RI21a16150_40 , 
    RI21a161c8_39 , 
    RI21a168d0_38 , 
    RI21a16948_37 , 
    RI21a13a68_67 , 
    RI21a13ae0_66 , 
    RI21a13b58_65 , 
    RI21a13bd0_64 , 
    RI21a13c48_63 , 
    RI21a14350_62 , 
    RI21a143c8_61 , 
    RI21a14530_58 , 
    RI21a15778_47 , 
    RI21a169c0_36 , 
    RI210d6910_193 , 
    RI210cdfb8_248 , 
    GI2046a680_186 , 
    RI210d2d88_218 , 
    RI210d10f0_228 , 
    RI210d1078_229 , 
    RI210d1000_230 , 
    RI210d0790_231 , 
    RI210d0718_232 , 
    RI210d06a0_233 , 
    RI210d0628_234 , 
    RI210cfdb8_235 , 
    RI210d4228_208 , 
    RI210d41b0_209 , 
    RI210d4138_210 , 
    RI210d38c8_211 , 
    RI210d3850_212 , 
    RI210d37d8_213 , 
    RI210d3760_214 , 
    RI210d2ef0_215 , 
    RI210d2e78_216 , 
    RI210d2e00_217 , 
    RI210d2518_219 , 
    RI210d24a0_220 , 
    RI210d2428_221 , 
    RI210d23b0_222 , 
    RI210d1b40_223 , 
    RI210d1ac8_224 , 
    RI210d1a50_225 , 
    RI210d19d8_226 , 
    RI210d1168_227 , 
    RI210d8ff8_178 , 
    RI21a0b7a0_150 , 
    RI21a0e590_122 , 
    RI210d55d8_200 , 
    RI210da3a8_170 , 
    RI21a0c178_143 , 
    RI210d73d8_187 , 
    RI21a0a6c0_158 , 
    RI21a0d438_131 , 
    RI210d5ec0_198 , 
    RI210da498_168 , 
    RI21a0c268_141 , 
    RI210d5560_201 , 
    RI210d9b38_171 , 
    RI21a0c100_144 , 
    RI210d54e8_202 , 
    RI210d9ac0_172 , 
    RI210cf2f0_241 , 
    RI210d4c78_203 , 
    RI210d9a48_173 , 
    RI21a0c088_145 , 
    RI210d4c00_204 , 
    RI210d99d0_174 , 
    RI21a0c010_146 , 
    RI210d4b88_205 , 
    RI210d9160_175 , 
    RI21a0b908_147 , 
    RI210d4b10_206 , 
    RI210d90e8_176 , 
    RI21a0b890_148 , 
    RI210d42a0_207 , 
    RI210d9070_177 , 
    RI21a0b818_149 , 
    RI210d8788_179 , 
    RI21a0b728_151 , 
    RI21a0de88_123 , 
    RI210d8710_180 , 
    RI21a0b6b0_152 , 
    RI21a0de10_124 , 
    RI210d8698_181 , 
    RI21a0afa8_153 , 
    RI21a0dd98_125 , 
    RI210d8620_182 , 
    RI21a0af30_154 , 
    RI21a0dd20_126 , 
    RI210d7db0_183 , 
    RI21a0aeb8_155 , 
    RI21a0dca8_127 , 
    RI210d7d38_184 , 
    RI21a0ae40_156 , 
    RI21a0dc30_128 , 
    RI210ce8a0_246 , 
    RI210cf278_242 , 
    RI21a0d528_129 , 
    RI210d7cc0_185 , 
    RI210cea08_243 , 
    RI210cfc50_238 , 
    RI210ce030_247 , 
    RI21a0adc8_157 , 
    RI21a0d4b0_130 , 
    RI210d7c48_186 , 
    RI210ce990_244 , 
    RI210cf3e0_239 , 
    RI210d7360_188 , 
    RI210ce918_245 , 
    RI210cf368_240 , 
    RI210d72e8_189 , 
    RI21a0a648_159 , 
    RI21a0d3c0_132 , 
    RI210d7270_190 , 
    RI21a0a5d0_160 , 
    RI21a0d348_133 , 
    RI210d6a00_191 , 
    RI21a0a558_161 , 
    RI21a0d2d0_134 , 
    RI210d6988_192 , 
    RI21a09e50_162 , 
    RI21a0cbc8_135 , 
    RI21a09dd8_163 , 
    RI21a0cb50_136 , 
    RI210d6898_194 , 
    RI21a09478_164 , 
    RI21a0cad8_137 , 
    RI210d6028_195 , 
    RI210dadf8_165 , 
    RI21a0ca60_138 , 
    RI210d5fb0_196 , 
    RI210dad80_166 , 
    RI21a0c9e8_139 , 
    RI21a16a38_35 , 
    RI210d5650_199 , 
    RI210da420_169 , 
    RI21a0c1f0_142 , 
    RI210d5f38_197 , 
    RI210da510_167 , 
    RI21a0c970_140 , 
    RI21a11650_88 , 
    RI21a115d8_89 , 
    RI210cfd40_236 , 
    RI210c9b48_275 , 
    RI210ca3b8_274 , 
    RI210ca4a8_272 , 
    RI210ca520_271 , 
    RI210cad90_270 , 
    RI210cae08_269 , 
    RI210cae80_268 , 
    RI210caef8_267 , 
    RI210cb768_266 , 
    RI210cb7e0_265 , 
    RI210cb858_264 , 
    RI210cb8d0_263 , 
    RI210cc1b8_261 , 
    RI210cc230_260 , 
    RI210cc2a8_259 , 
    RI210ccb18_258 , 
    RI210ccb90_257 , 
    RI210ccc08_256 , 
    RI210ccc80_255 , 
    RI210cd4f0_254 , 
    RI210cd568_253 , 
    RI210cd5e0_252 , 
    RI210c07a0_282 , 
    RI210c0818_281 , 
    RI210c2078_280 , 
    RI210c9170_279 , 
    RI210c91e8_278 , 
    RI210c9a58_277 , 
    RI210c9ad0_276 , 
    RI210ca430_273 , 
    RI210cc140_262 , 
    RI210cd658_251 , 
    RI2107f4a8_454 , 
    RI210aeb90_395 , 
    GI20471ac0_434 , 
    RI2107f340_457 , 
    RI2107e878_458 , 
    RI21084f20_415 , 
    RI21084458_416 , 
    RI2107e800_459 , 
    RI2107e788_460 , 
    RI2107e710_461 , 
    RI2107e698_462 , 
    RI210843e0_417 , 
    RI210a63a0_396 , 
    RI21086e10_397 , 
    RI21086bb8_398 , 
    RI21086b40_399 , 
    RI21086ac8_400 , 
    RI21086a50_401 , 
    RI210869d8_402 , 
    RI21086960_403 , 
    RI21085e98_404 , 
    RI21085e20_405 , 
    RI21085da8_406 , 
    RI21085d30_407 , 
    RI21085cb8_408 , 
    RI21085c40_409 , 
    RI21085178_410 , 
    RI21085100_411 , 
    RI21085088_412 , 
    RI21085010_413 , 
    RI21084f98_414 , 
    RI210b2538_374 , 
    RI210b43b0_360 , 
    RI210b7f38_335 , 
    RI210afec8_388 , 
    RI210b2628_372 , 
    RI210b4d88_356 , 
    RI21081b18_438 , 
    RI210b6b88_343 , 
    RI210b07b0_386 , 
    RI21081aa0_439 , 
    RI210b5670_354 , 
    RI210afe50_389 , 
    RI21080fd8_440 , 
    RI21083648_424 , 
    RI2107f3b8_456 , 
    RI21080f60_441 , 
    RI210835d0_425 , 
    RI210afdd8_390 , 
    RI21080ee8_442 , 
    RI210b4d10_357 , 
    RI210af568_391 , 
    RI21080e70_443 , 
    RI210b4c98_358 , 
    RI210af4f0_392 , 
    RI21080df8_444 , 
    RI21083558_426 , 
    RI210af478_393 , 
    RI21080d80_445 , 
    RI210834e0_427 , 
    RI210aec08_394 , 
    RI210b25b0_373 , 
    RI210b4428_359 , 
    RI210b1cc8_375 , 
    RI21082a18_428 , 
    RI210b7ec0_336 , 
    RI210802b8_446 , 
    RI210829a0_429 , 
    RI210b7e48_337 , 
    RI21080240_447 , 
    RI21082928_430 , 
    RI210b7dd0_338 , 
    RI210801c8_448 , 
    RI210828b0_431 , 
    RI210b7560_339 , 
    RI21080150_449 , 
    RI21082838_432 , 
    RI210b74e8_340 , 
    RI210800d8_450 , 
    RI210827c0_433 , 
    RI210b7470_341 , 
    RI21080060_451 , 
    RI21081cf8_434 , 
    RI21084200_421 , 
    RI2107f598_452 , 
    RI21081c80_435 , 
    RI21083738_422 , 
    RI210b1c50_376 , 
    RI21081c08_436 , 
    RI210836c0_423 , 
    RI2107f520_453 , 
    RI21081b90_437 , 
    RI210b73f8_342 , 
    RI2107f430_455 , 
    RI210b4338_361 , 
    RI210b6b10_344 , 
    RI210b1bd8_377 , 
    RI210b42c0_362 , 
    RI210b6a98_345 , 
    RI210b1b60_378 , 
    RI210b3a50_363 , 
    RI210b6a20_346 , 
    RI210b12f0_379 , 
    RI210b39d8_364 , 
    RI210b61b0_347 , 
    RI210b1278_380 , 
    RI210b3960_365 , 
    RI210b6138_348 , 
    RI210b1200_381 , 
    RI210b38e8_366 , 
    RI210b60c0_349 , 
    RI210b1188_382 , 
    RI210b3078_367 , 
    RI210b6048_350 , 
    RI210b0918_383 , 
    RI210b3000_368 , 
    RI210b57d8_351 , 
    RI210b08a0_384 , 
    RI210b2f88_369 , 
    RI210b5760_352 , 
    RI210cdec8_250 , 
    RI210aff40_387 , 
    RI210b26a0_371 , 
    RI210b4e00_355 , 
    RI210b0828_385 , 
    RI210b2f10_370 , 
    RI210b56e8_353 , 
    RI210bd668_302 , 
    RI210bcdf8_303 , 
    RI21077000_517 , 
    RI21076538_518 , 
    RI210cdf40_249 , 
    RI2107db58_464 , 
    RI21069950_647 , 
    RI210699c8_646 , 
    R_61e_1dfaf3c8 , 
    R_8f7_1e09b6c8 , 
    R_714_1dfb8888 , 
    R_951_1e17ef68 , 
    R_28c_1d9fb268 , 
    R_9be_1e183888 , 
    R_9ab_1e1827a8 , 
    R_30f_1d9d04a8 , 
    R_959_1e17f468 , 
    R_b13_1e6b0908 , 
    R_519_1dda4b48 , 
    R_92d_1e09d888 , 
    R_c06_1e6bafe8 , 
    R_8c6_1e099d28 , 
    R_845_1e094788 , 
    R_414_1d9da7c8 , 
    R_313_1d9d0728 , 
    R_518_1dda4aa8 , 
    R_9d9_1e184468 , 
    R_4dd_1dda25c8 , 
    R_59f_1dda9f08 , 
    R_517_1dda4a08 , 
    R_509_1dda4148 , 
    R_508_1dda40a8 , 
    R_401_1d9d9be8 , 
    R_5f9_1ddad748 , 
    R_6ef_1dfb7168 , 
    R_a30_1e187ac8 , 
    R_2b0_1d9fc8e8 , 
    R_77c_1dfbc988 , 
    R_8f1_1e09b308 , 
    R_36a_1d9d4288 , 
    R_507_1dda4008 , 
    R_516_1dda4e68 , 
    R_98e_1e181a88 , 
    R_8d5_1e09a188 , 
    R_498_1dd9faa8 , 
    R_68b_1dfb32e8 , 
    R_773_1dfbc3e8 , 
    R_45b_1d9dd428 , 
    R_48d_1dd9f3c8 , 
    R_5ff_1ddadb08 , 
    R_705_1dfb7f28 , 
    R_644_1dfb0688 , 
    R_63a_1dfb0548 , 
    R_ac7_1e18d928 , 
    R_320_1d9d0f48 , 
    R_737_1dfb9e68 , 
    R_506_1dda4468 , 
    R_647_1dfb0868 , 
    R_b86_1e6bb4e8 , 
    R_883_1e096e48 , 
    R_6a8_1dfb4508 , 
    R_aa5_1e18c3e8 , 
    R_440_1d9dc348 , 
    R_2f9_1d9cf6e8 , 
    R_69c_1dfb3d88 , 
    R_65d_1dfb1628 , 
    R_b0c_1e6b04a8 , 
    R_b20_1e6b1128 , 
    R_a2e_1e189788 , 
    R_905_1e09bf88 , 
    R_a57_1e189328 , 
    R_5f8_1ddad6a8 , 
    R_54c_1dda6b28 , 
    R_bd2_1e6b32e8 , 
    R_aca_1e6ae068 , 
    R_58b_1dda9288 , 
    R_2e3_1d9ce928 , 
    R_3e2_1d9d8d88 , 
    R_8f6_1e09bb28 , 
    R_331_1d9d19e8 , 
    R_97d_1e180ae8 , 
    R_5cd_1ddabbc8 , 
    R_45c_1d9dd4c8 , 
    R_999_1e181c68 , 
    R_b99_1e6b5cc8 , 
    R_948_1e17e9c8 , 
    R_97e_1e181308 , 
    R_ab0_1e18cac8 , 
    R_bb8_1e6b7028 , 
    R_489_1dd9f148 , 
    R_4b6_1dda1268 , 
    R_63f_1dfb0368 , 
    R_3e7_1d9d8ba8 , 
    R_2bd_1d9fd108 , 
    R_81b_1e092d48 , 
    R_b54_1e6b31a8 , 
    R_4df_1dda2708 , 
    R_bab_1e6b6808 , 
    R_431_1d9db9e8 , 
    R_2f2_1d9cf788 , 
    R_601_1ddadc48 , 
    R_6e7_1dfb6c68 , 
    R_bdf_1e6b8888 , 
    R_656_1dfb1bc8 , 
    R_4e0_1dda27a8 , 
    R_4de_1dda2b68 , 
    R_a4e_1e189288 , 
    R_8e1_1e09a908 , 
    R_8f0_1e09b268 , 
    R_299_1d9fba88 , 
    R_292_1d9fb628 , 
    R_4e1_1dda2848 , 
    R_a7f_1e18ac28 , 
    R_c04_1e6b9fa8 , 
    R_3ef_1d9d90a8 , 
    R_5de_1dd9f1e8 , 
    R_878_1e096768 , 
    R_720_1dfb9008 , 
    R_ad6_1e6ae7e8 , 
    R_9a2_1e182708 , 
    R_630_1dfafa08 , 
    R_52f_1dda5908 , 
    R_7a9_1e08e608 , 
    R_976_1e180b88 , 
    R_439_1d9dbee8 , 
    R_604_1ddade28 , 
    R_530_1dda59a8 , 
    R_52e_1dda5d68 , 
    R_7ed_1e091088 , 
    R_3f2_1d9d4c88 , 
    R_3d4_1d9d7fc8 , 
    R_84a_1e094fa8 , 
    R_2de_1d9ceb08 , 
    R_690_1dfb3608 , 
    R_4cd_1dda1bc8 , 
    R_531_1dda5a48 , 
    R_b34_1e6b1da8 , 
    R_5f7_1ddad608 , 
    R_806_1e092528 , 
    R_a5b_1e1895a8 , 
    R_718_1dfb8b08 , 
    R_695_1dfb3928 , 
    R_7af_1e08e9c8 , 
    R_62b_1dfaf6e8 , 
    R_904_1e09bee8 , 
    R_501_1dda3c48 , 
    R_585_1dda8ec8 , 
    R_9cd_1e183ce8 , 
    R_78c_1dfbd388 , 
    R_392_1d9d5b88 , 
    R_4b4_1dda0c28 , 
    R_b44_1e6b27a8 , 
    R_969_1e17fe68 , 
    R_40d_1d9da368 , 
    R_627_1dfaf468 , 
    R_67a_1dfadfc8 , 
    R_45d_1d9dd568 , 
    R_7c1_1e08f508 , 
    R_552_1dda73e8 , 
    R_2bf_1d9fd248 , 
    R_5d4_1ddac028 , 
    R_b77_1e6b4788 , 
    R_3fa_1d9db088 , 
    R_6aa_1dfb4b48 , 
    R_82a_1e093ba8 , 
    R_3aa_1d9d6a88 , 
    R_300_1d9cfb48 , 
    R_405_1d9d9e68 , 
    R_953_1e17f0a8 , 
    R_3cf_1d9d7ca8 , 
    R_ac1_1e18d568 , 
    R_61c_1dfaed88 , 
    R_a99_1e18bc68 , 
    R_4ae_1dda0fe8 , 
    R_aec_1e6af0a8 , 
    R_af8_1e6af828 , 
    R_762_1dfbbe48 , 
    R_3a8_1d9d6448 , 
    R_4ca_1dda1ee8 , 
    R_6b7_1dfb4e68 , 
    R_57c_1dda8928 , 
    R_52b_1dda5688 , 
    R_8ef_1e09b1c8 , 
    R_8c5_1e099788 , 
    R_8ab_1e098748 , 
    R_71c_1dfb8d88 , 
    R_388_1d9d5048 , 
    R_b6e_1e6b46e8 , 
    R_9cc_1e183c48 , 
    R_65b_1dfb14e8 , 
    R_bbd_1e6b7348 , 
    R_3b2_1d9d6f88 , 
    R_862_1e095ea8 , 
    R_4a5_1dda02c8 , 
    R_90f_1e09c5c8 , 
    R_702_1dfb8248 , 
    R_29f_1d9fbe48 , 
    R_72b_1dfb96e8 , 
    R_6f4_1dfb7488 , 
    R_5f2_1dda8a68 , 
    R_a64_1e189b48 , 
    R_2e9_1d9cece8 , 
    R_683_1dfb2de8 , 
    R_2fd_1d9cf968 , 
    R_8b2_1e0990a8 , 
    R_5f0_1ddad1a8 , 
    R_bac_1e6b68a8 , 
    R_642_1dfb0a48 , 
    R_5f6_1d9fbda8 , 
    R_568_1dda7ca8 , 
    R_409_1d9da0e8 , 
    R_5a8_1ddaa4a8 , 
    R_5e3_1ddac988 , 
    R_96b_1e17ffa8 , 
    R_bca_1e6b14e8 , 
    R_3b8_1d9d6e48 , 
    R_789_1dfbd1a8 , 
    R_86a_1e0963a8 , 
    R_416_1ddabc68 , 
    R_903_1e09be48 , 
    R_a2d_1e1878e8 , 
    R_9cb_1e183ba8 , 
    R_59b_1dda9c88 , 
    R_a4c_1e188c48 , 
    R_79c_1dfbdd88 , 
    R_888_1e097168 , 
    R_2a7_1d9fc348 , 
    R_7f3_1e091448 , 
    R_73c_1dfba188 , 
    R_bd1_1e6b7fc8 , 
    R_4a6_1dda0868 , 
    R_3dd_1d9d8568 , 
    R_346_1d9d2c08 , 
    R_4c4_1dda1628 , 
    R_b15_1e6b0a48 , 
    R_5ec_1ddacf28 , 
    R_bb4_1e6b6da8 , 
    R_bed_1e6b9148 , 
    R_7bf_1e08f3c8 , 
    R_344_1d9d25c8 , 
    R_c0b_1e6ba408 , 
    R_6a5_1dfb4328 , 
    R_b8c_1e6b54a8 , 
    R_3a1_1d9d5fe8 , 
    R_7ea_1e09d928 , 
    R_46e_1dd9e568 , 
    R_8ee_1e09b628 , 
    R_697_1dfb3a68 , 
    R_77f_1dfbcb68 , 
    R_391_1d9d55e8 , 
    R_746_1dfb6448 , 
    R_b3b_1e6b2208 , 
    R_7f1_1e091308 , 
    R_410_1d9da548 , 
    R_700_1dfb7c08 , 
    R_58f_1dda9508 , 
    R_582_1dda91e8 , 
    R_793_1dfbd7e8 , 
    R_847_1e0948c8 , 
    R_95e_1e17fc88 , 
    R_560_1dda77a8 , 
    R_9ca_1e184008 , 
    R_397_1d9d59a8 , 
    R_46b_1d9dde28 , 
    R_44e_1d9fc028 , 
    R_6cc_1dfb5b88 , 
    R_62e_1dfafdc8 , 
    R_2b1_1d9fc988 , 
    R_6f9_1dfb77a8 , 
    R_af5_1e6af648 , 
    R_b81_1e6b4dc8 , 
    R_427_1d9db3a8 , 
    R_547_1dda6808 , 
    R_c1d_1e6baf48 , 
    R_a2c_1e187848 , 
    R_355_1d9d3068 , 
    R_857_1e0952c8 , 
    R_413_1d9da728 , 
    R_afa_1e6afe68 , 
    R_adc_1e6ae6a8 , 
    R_5fc_1ddad928 , 
    R_c24_1e6bb3a8 , 
    R_421_1d9dafe8 , 
    R_892_1e17e608 , 
    R_70b_1dfb82e8 , 
    R_aad_1e18c8e8 , 
    R_3ca_1d9d8108 , 
    R_7ac_1e08e7e8 , 
    R_8da_1e09a9a8 , 
    R_400_1d9d9b48 , 
    R_bb0_1e6b6b28 , 
    R_893_1e097848 , 
    R_902_1e09c2a8 , 
    R_a93_1e18b8a8 , 
    R_8cd_1e099c88 , 
    R_861_1e095908 , 
    R_3ea_1d9d9288 , 
    R_915_1e09c988 , 
    R_844_1e0946e8 , 
    R_677_1dfb2668 , 
    R_602_1dfae248 , 
    R_39c_1d9d5cc8 , 
    R_be3_1e6b8b08 , 
    R_bea_1e6b9468 , 
    R_993_1e1818a8 , 
    R_bad_1e6b6948 , 
    R_88d_1e097488 , 
    R_5a2_1ddaa5e8 , 
    R_655_1dfb1128 , 
    R_4ad_1dda07c8 , 
    R_493_1dd9f788 , 
    R_894_1e0978e8 , 
    R_668_1dfb1d08 , 
    R_730_1dfb9a08 , 
    R_7dc_1e0905e8 , 
    R_abd_1e18d2e8 , 
    R_662_1dfb1e48 , 
    R_a7c_1e18aa48 , 
    R_5cf_1ddabd08 , 
    R_328_1d9d1448 , 
    R_741_1dfba4a8 , 
    R_9a6_1e182988 , 
    R_36d_1d9d3f68 , 
    R_308_1d9d0048 , 
    R_95b_1e17f5a8 , 
    R_b63_1e6b3b08 , 
    R_2da_1d9ce888 , 
    R_5dc_1ddac528 , 
    R_49f_1dd9ff08 , 
    R_895_1e097988 , 
    R_761_1dfbb8a8 , 
    R_2e4_1d9ce9c8 , 
    R_ab5_1e18cde8 , 
    R_c28_1e6bb628 , 
    R_8d4_1e09a0e8 , 
    R_a8c_1e18b448 , 
    R_597_1dda9a08 , 
    R_5c4_1ddab628 , 
    R_384_1d9d4dc8 , 
    R_31c_1d9d0cc8 , 
    R_987_1e181128 , 
    R_b2e_1e6b1ee8 , 
    R_2f3_1d9cf328 , 
    R_6cf_1dfb5d68 , 
    R_6e4_1dfb6a88 , 
    R_357_1d9d31a8 , 
    R_3c1_1d9d73e8 , 
    R_5e7_1ddacc08 , 
    R_974_1e180548 , 
    R_61a_1dfaf148 , 
    R_3f8_1d9d9648 , 
    R_802_1e0922a8 , 
    R_593_1dda9788 , 
    R_a69_1e189e68 , 
    R_a87_1e18b128 , 
    R_a5d_1e1896e8 , 
    R_a2b_1e1877a8 , 
    R_671_1dfb22a8 , 
    R_4cf_1dda1d08 , 
    R_420_1d9daf48 , 
    R_6bc_1dfb5188 , 
    R_43f_1d9dc2a8 , 
    R_692_1dfb3c48 , 
    R_80b_1e092348 , 
    R_882_1e0972a8 , 
    R_871_1e096308 , 
    R_2c2_1d9fd928 , 
    R_2ce_1d9cfa08 , 
    R_a9c_1e18be48 , 
    R_768_1dfbbd08 , 
    R_56d_1dda7fc8 , 
    R_34c_1d9d2ac8 , 
    R_b8f_1e6b5688 , 
    R_b07_1e6b0188 , 
    R_6b5_1dfb4d28 , 
    R_5ae_1ddaad68 , 
    R_2df_1d9ce6a8 , 
    R_674_1dfb2488 , 
    R_608_1dfae108 , 
    R_ad3_1e6ae108 , 
    R_505_1dda3ec8 , 
    R_8bf_1e0993c8 , 
    R_542_1dda69e8 , 
    R_7f6_1e091b28 , 
    R_504_1dda3e28 , 
    R_8a7_1e0984c8 , 
    R_76a_1dfbc5c8 , 
    R_937_1e09dec8 , 
    R_6fb_1dfb78e8 , 
    R_3b0_1d9d6948 , 
    R_2c0_1d9fd2e8 , 
    R_37c_1d9d48c8 , 
    R_782_1dfbd248 , 
    R_503_1dda3d88 , 
    R_82e_1e093e28 , 
    R_8bb_1e099148 , 
    R_430_1d9db948 , 
    R_5cb_1ddaba88 , 
    R_ae6_1e6af1e8 , 
    R_7a3_1e08e248 , 
    R_b78_1e6b4828 , 
    R_bc9_1e6b7ac8 , 
    R_380_1d9d4b48 , 
    R_33d_1d9d2168 , 
    R_8e0_1e09a868 , 
    R_3c7_1d9d77a8 , 
    R_2b2_1d9fcf28 , 
    R_618_1dfaeb08 , 
    R_823_1e093248 , 
    R_89e_1e098428 , 
    R_502_1dda41e8 , 
    R_b6f_1e6b4288 , 
    R_c00_1e6b9d28 , 
    R_98d_1e1814e8 , 
    R_28b_1d9fb1c8 , 
    R_a55_1e1891e8 , 
    R_3c4_1d9d75c8 , 
    R_40c_1d9da2c8 , 
    R_2d2_1d9ce388 , 
    R_c21_1e6bb1c8 , 
    R_b3d_1e6b2348 , 
    R_877_1e0966c8 , 
    R_855_1e095188 , 
    R_41d_1d9dad68 , 
    R_438_1d9dbe48 , 
    R_2d6_1d9ce608 , 
    R_7da_1e0909a8 , 
    R_6f6_1dfb7ac8 , 
    R_9aa_1e182e88 , 
    R_b47_1e6b2988 , 
    R_a2a_1e6b3ce8 , 
    R_41f_1d9daea8 , 
    R_ae4_1e6aeba8 , 
    R_a79_1e18a868 , 
    R_3a3_1d9d6128 , 
    R_5bd_1ddab1c8 , 
    R_301_1d9cfbe8 , 
    R_298_1d9fb9e8 , 
    R_bb9_1e6b70c8 , 
    R_82d_1e093888 , 
    R_404_1d9d9dc8 , 
    R_a62_1e189f08 , 
    R_93c_1e17e248 , 
    R_62d_1dfaf828 , 
    R_579_1dda8748 , 
    R_452_1ddac3e8 , 
    R_54d_1dda6bc8 , 
    R_4d9_1dda2348 , 
    R_4d4_1dda2028 , 
    R_6c1_1dfb54a8 , 
    R_379_1d9d46e8 , 
    R_34e_1d9d3108 , 
    R_94a_1e097ca8 , 
    R_74b_1dfbaae8 , 
    R_ade_1e6aece8 , 
    R_79f_1e08dfc8 , 
    R_797_1dfbda68 , 
    R_943_1e17e6a8 , 
    R_653_1dfb0fe8 , 
    R_3d8_1d9d8248 , 
    R_b61_1e6b39c8 , 
    R_bc4_1e6b77a8 , 
    R_a02_1e186308 , 
    R_368_1d9d3c48 , 
    R_35e_1d9d3b08 , 
    R_7fe_1e092028 , 
    R_499_1dd9fb48 , 
    R_680_1dfb2c08 , 
    R_2a8_1d9fc3e8 , 
    R_6ec_1dfb6f88 , 
    R_776_1dfbcac8 , 
    R_b5e_1e6b0368 , 
    R_635_1dfafd28 , 
    R_7fa_1e091da8 , 
    R_af7_1e6af788 , 
    R_8c4_1e0996e8 , 
    R_408_1d9da048 , 
    R_ab9_1e18d068 , 
    R_6a2_1dfb61c8 , 
    R_291_1d9fb588 , 
    R_7b8_1e08ef68 , 
    R_8b6_1e08e6a8 , 
    R_48a_1dda0d68 , 
    R_6c7_1dfb5868 , 
    R_c10_1e6ba728 , 
    R_bf1_1e6b93c8 , 
    R_4d6_1dd9e2e8 , 
    R_5b3_1ddaab88 , 
    R_771_1dfbc2a8 , 
    R_af1_1e6af3c8 , 
    R_6e1_1dfb68a8 , 
    R_a9f_1e18c028 , 
    R_b17_1e6b0b88 , 
    R_b30_1e6b1b28 , 
    R_bde_1e6b37e8 , 
    R_998_1e181bc8 , 
    R_a4a_1e189008 , 
    R_48e_1dd9f968 , 
    R_688_1dfb3108 , 
    R_810_1e092668 , 
    R_75c_1dfbb588 , 
    R_3bb_1d9d7028 , 
    R_c2e_1e17f008 , 
    R_5d2_1d9db308 , 
    R_32e_1d9d1d08 , 
    R_580_1dda8ba8 , 
    R_453_1d9dcf28 , 
    R_83a_1e0913a8 , 
    R_41e_1d9dc988 , 
    R_97c_1e180a48 , 
    R_5b8_1ddaaea8 , 
    R_363_1d9d3928 , 
    R_94e_1ddadce8 , 
    R_7c4_1e08f6e8 , 
    R_52c_1dda5728 , 
    R_aa2_1e18c708 , 
    R_625_1dfaf328 , 
    R_4b7_1dda0e08 , 
    R_55d_1dda75c8 , 
    R_b0e_1e6b0ae8 , 
    R_425_1d9db268 , 
    R_30c_1d9d02c8 , 
    R_3db_1d9d8428 , 
    R_a48_1e1889c8 , 
    R_aaf_1e18ca28 , 
    R_5ad_1ddaa7c8 , 
    R_589_1dda9148 , 
    R_338_1d9d1e48 , 
    R_832_1e0940a8 , 
    R_790_1dfbd608 , 
    R_318_1d9d0a48 , 
    R_869_1e095e08 , 
    R_6d3_1dfb5fe8 , 
    R_60c_1dfae388 , 
    R_56a_1dda82e8 , 
    R_887_1e0970c8 , 
    R_815_1e092988 , 
    R_66b_1dfb1ee8 , 
    R_a34_1e187d48 , 
    R_40f_1d9da4a8 , 
    R_ac3_1e18d6a8 , 
    R_324_1d9d11c8 , 
    R_614_1dfae888 , 
    R_752_1dfbb448 , 
    R_4c0_1dda13a8 , 
    R_7d9_1e090408 , 
    R_ad0_1e18dec8 , 
    R_bee_1e6b96e8 , 
    R_736_1dfba2c8 , 
    R_727_1dfb9468 , 
    R_a8a_1e18b808 , 
    R_933_1e09dc48 , 
    R_8b1_1e098b08 , 
    R_606_1dfae4c8 , 
    R_927_1e09d4c8 , 
    R_a7a_1e18ae08 , 
    R_333_1d9d1b28 , 
    R_968_1e17fdc8 , 
    R_574_1dda8428 , 
    R_836_1e094328 , 
    R_757_1dfbb268 , 
    R_2db_1d9ce428 , 
    R_af4_1e6af5a8 , 
    R_454_1d9dcfc8 , 
    R_412_1d9dab88 , 
    R_709_1dfb81a8 , 
    R_8a4_1e0982e8 , 
    R_c1b_1e6bae08 , 
    R_846_1e094d28 , 
    R_3ff_1d9d9aa8 , 
    R_76e_1dfbdec8 , 
    R_33f_1d9d22a8 , 
    R_4af_1dda0908 , 
    R_a67_1e189d28 , 
    R_616_1dfaeec8 , 
    R_b49_1e6b2ac8 , 
    R_2f4_1d9cf3c8 , 
    R_426_1d9db808 , 
    R_2e5_1d9cea68 , 
    R_bb5_1e6b6e48 , 
    R_7b6_1e08f328 , 
    R_751_1dfbaea8 , 
    R_bd0_1e6b7f28 , 
    R_610_1dfae608 , 
    R_918_1e09cb68 , 
    R_35c_1d9d34c8 , 
    R_924_1e09d2e8 , 
    R_912_1e09cca8 , 
    R_77d_1dfbca28 , 
    R_774_1dfbc488 , 
    R_a71_1e18a368 , 
    R_32d_1d9d1768 , 
    R_99d_1e181ee8 , 
    R_87d_1e096a88 , 
    R_472_1dd9e7e8 , 
    R_b2a_1e6b1c68 , 
    R_56f_1dda8108 , 
    R_b87_1e6b5188 , 
    R_921_1e09d108 , 
    R_375_1d9d4468 , 
    R_576_1dda8ce8 , 
    R_b82_1e6b5368 , 
    R_39e_1d9d6308 , 
    R_856_1e095728 , 
    R_6c2_1dfb5a48 , 
    R_2c3_1d9fd4c8 , 
    R_90b_1e09c348 , 
    R_92f_1e09d9c8 , 
    R_38e_1d9d5908 , 
    R_b9e_1e18d388 , 
    R_8cc_1e099be8 , 
    R_860_1e095868 , 
    R_c09_1e6ba2c8 , 
    R_b09_1e6b02c8 , 
    R_521_1dda5048 , 
    R_b4a_1e6b3068 , 
    R_88c_1e0973e8 , 
    R_520_1dda4fa8 , 
    R_8b5_1e098d88 , 
    R_b5d_1e6b3748 , 
    R_843_1e094648 , 
    R_633_1dfafbe8 , 
    R_7c2_1e08faa8 , 
    R_6d8_1dfb6308 , 
    R_38d_1d9d5368 , 
    R_7e7_1e090cc8 , 
    R_bfc_1e6b9aa8 , 
    R_841_1e094508 , 
    R_a96_1e18bf88 , 
    R_7e5_1e090b88 , 
    R_51f_1dda4f08 , 
    R_949_1e17ea68 , 
    R_b5a_1e6b3a68 , 
    R_2e0_1d9ce748 , 
    R_acd_1e18dce8 , 
    R_70f_1dfb8568 , 
    R_c15_1e6baa48 , 
    R_310_1d9d0548 , 
    R_bf5_1e6b9648 , 
    R_314_1d9d07c8 , 
    R_6af_1dfb4968 , 
    R_445_1d9dc668 , 
    R_658_1dfb1308 , 
    R_a6c_1e18a048 , 
    R_2c1_1d9fd388 , 
    R_2b3_1d9fcac8 , 
    R_6de_1dfb6bc8 , 
    R_9b9_1e183068 , 
    R_6ad_1dfb4828 , 
    R_548_1dda68a8 , 
    R_4c9_1dda1948 , 
    R_51e_1dda5368 , 
    R_96a_1e180408 , 
    R_455_1d9dd068 , 
    R_8d3_1e09a048 , 
    R_bb1_1e6b6bc8 , 
    R_7d7_1e0902c8 , 
    R_6a0_1dfb4008 , 
    R_b79_1e6b48c8 , 
    R_565_1dda7ac8 , 
    R_586_1dda9468 , 
    R_4a7_1dda0408 , 
    R_b70_1e6b4328 , 
    R_661_1dfb18a8 , 
    R_2d3_1d9fdec8 , 
    R_ad9_1e6ae4c8 , 
    R_a85_1e18afe8 , 
    R_a77_1e18a728 , 
    R_2d7_1d9ce1a8 , 
    R_7b3_1e08ec48 , 
    R_870_1e096268 , 
    R_43e_1d9dc708 , 
    R_6db_1dfb64e8 , 
    R_807_1e0920c8 , 
    R_a74_1e18a548 , 
    R_bf9_1e6b98c8 , 
    R_321_1d9d0fe8 , 
    R_a53_1e1890a8 , 
    R_4e3_1dda2988 , 
    R_831_1e093b08 , 
    R_66e_1dfb25c8 , 
    R_ac6_1e18dd88 , 
    R_55a_1dda78e8 , 
    R_4c6_1dda1c68 , 
    R_4e4_1dda2a28 , 
    R_4e2_1dda2de8 , 
    R_c22_1e6b55e8 , 
    R_92c_1e09d7e8 , 
    R_7c9_1e08fa08 , 
    R_623_1dfaf1e8 , 
    R_b58_1e6b3428 , 
    R_370_1d9d4148 , 
    R_3be_1d9d7708 , 
    R_4e5_1dda2ac8 , 
    R_a03_1e185ea8 , 
    R_c12_1e6bad68 , 
    R_456_1d9dd608 , 
    R_bf2_1e6b9968 , 
    R_6a7_1dfb4468 , 
    R_c30_1e6bbb28 , 
    R_40b_1d9da228 , 
    R_42f_1d9db8a8 , 
    R_68d_1dfb3428 , 
    R_735_1dfb9d28 , 
    R_78d_1dfbd428 , 
    R_8df_1e09a7c8 , 
    R_41c_1d9dacc8 , 
    R_46f_1dd9e108 , 
    R_2a9_1d9fc488 , 
    R_81e_1e093428 , 
    R_5e0_1ddac7a8 , 
    R_462_1d9ddd88 , 
    R_60a_1dfae748 , 
    R_5a7_1ddaa408 , 
    R_403_1d9d9d28 , 
    R_2c6_1d9fdba8 , 
    R_7e3_1e090a48 , 
    R_7ee_1e09c528 , 
    R_706_1dfb84c8 , 
    R_c17_1e6bab88 , 
    R_c1f_1e6bb088 , 
    R_b93_1e6b5908 , 
    R_854_1e0950e8 , 
    R_b9f_1e6b6088 , 
    R_8e5_1e09ab88 , 
    R_437_1d9dbda8 , 
    R_612_1dfaec48 , 
    R_816_1e0931a8 , 
    R_b19_1e6b0cc8 , 
    R_73b_1dfba0e8 , 
    R_a44_1e188748 , 
    R_93e_1e17e888 , 
    R_67c_1dfb2988 , 
    R_992_1e181d08 , 
    R_494_1dd9f828 , 
    R_3e0_1d9d8748 , 
    R_7a7_1e08e4c8 , 
    R_876_1e096b28 , 
    R_543_1dda6588 , 
    R_8ae_1dfbc0c8 , 
    R_351_1d9d2de8 , 
    R_457_1d9dd1a8 , 
    R_bf6_1e6b3f68 , 
    R_a38_1e187fc8 , 
    R_6f1_1dfb72a8 , 
    R_b3e_1e6b28e8 , 
    R_53e_1dda6768 , 
    R_ac0_1e18d4c8 , 
    R_763_1dfbb9e8 , 
    R_c26_1e6b8ce8 , 
    R_650_1dfb0e08 , 
    R_361_1d9d37e8 , 
    R_aaa_1e187e88 , 
    R_b10_1e6b0728 , 
    R_b2c_1e6b18a8 , 
    R_5a1_1ddaa048 , 
    R_be7_1e6b8d88 , 
    R_b26_1e6b19e8 , 
    R_4a0_1dd9ffa8 , 
    R_95a_1e17fa08 , 
    R_909_1e09c208 , 
    R_463_1d9dd928 , 
    R_407_1d9d9fa8 , 
    R_5c5_1ddab6c8 , 
    R_986_1e181588 , 
    R_515_1dda48c8 , 
    R_5c1_1ddab448 , 
    R_297_1d9fb948 , 
    R_514_1dda4828 , 
    R_b4c_1e6b2ca8 , 
    R_973_1e1804a8 , 
    R_60e_1dfae9c8 , 
    R_7d4_1e0900e8 , 
    R_7c7_1e08f8c8 , 
    R_513_1dda4788 , 
    R_65f_1dfb1768 , 
    R_9b5_1e182de8 , 
    R_2ee_1d9cf508 , 
    R_91b_1e09cd48 , 
    R_af6_1e6afbe8 , 
    R_83d_1e094288 , 
    R_8c3_1e099648 , 
    R_458_1d9dd248 , 
    R_512_1dda4be8 , 
    R_ba6_1e6b69e8 , 
    R_5e5_1ddacac8 , 
    R_57b_1dda8888 , 
    R_aeb_1e6af008 , 
    R_7f4_1e0914e8 , 
    R_a46_1e188d88 , 
    R_b8d_1e6b5548 , 
    R_562_1dda7de8 , 
    R_745_1dfba728 , 
    R_557_1dda7208 , 
    R_464_1d9dd9c8 , 
    R_835_1e093d88 , 
    R_49a_1dda00e8 , 
    R_7d1_1e08ff08 , 
    R_911_1e09c708 , 
    R_6e9_1dfb6da8 , 
    R_723_1dfb91e8 , 
    R_a95_1e18b9e8 , 
    R_58d_1dda93c8 , 
    R_a89_1e18b268 , 
    R_780_1dfbcc08 , 
    R_740_1dfba408 , 
    R_72f_1dfb9968 , 
    R_828_1e093568 , 
    R_89c_1e097de8 , 
    R_a32_1e188108 , 
    R_840_1e094468 , 
    R_b37_1e6b1f88 , 
    R_9db_1e1845a8 , 
    R_b22_1e6b1768 , 
    R_9dc_1e184648 , 
    R_9da_1e184a08 , 
    R_794_1dfbd888 , 
    R_33a_1d9d2488 , 
    R_424_1d9db1c8 , 
    R_2dc_1d9ce4c8 , 
    R_a6f_1e18a228 , 
    R_98c_1e181448 , 
    R_6b6_1dfb52c8 , 
    R_908_1e09c168 , 
    R_9dd_1e1846e8 , 
    R_965_1e17fbe8 , 
    R_28a_1d9fb128 , 
    R_529_1dda5548 , 
    R_40e_1d9da908 , 
    R_bcd_1e6b7d48 , 
    R_476_1dd9ea68 , 
    R_393_1d9d5728 , 
    R_a40_1e1884c8 , 
    R_528_1dda54a8 , 
    R_2fa_1d9d0188 , 
    R_a3c_1e188248 , 
    R_868_1e095d68 , 
    R_2cf_1d9fdc48 , 
    R_2c4_1d9fd568 , 
    R_7cc_1e08fbe8 , 
    R_8fd_1e09ba88 , 
    R_3d5_1d9d8068 , 
    R_b64_1e6b3ba8 , 
    R_527_1dda5408 , 
    R_9d1_1e183f68 , 
    R_46c_1d9ddec8 , 
    R_2f5_1d9cf468 , 
    R_839_1e094008 , 
    R_554_1dda7028 , 
    R_3ab_1d9d6628 , 
    R_459_1d9dd2e8 , 
    R_b4f_1e6b2e88 , 
    R_886_1e097528 , 
    R_3e5_1d9d8a68 , 
    R_52d_1dda57c8 , 
    R_290_1d9fb4e8 , 
    R_b7a_1e18cc08 , 
    R_526_1dda5ae8 , 
    R_79a_1e098e28 , 
    R_ba0_1e6b6128 , 
    R_6d1_1dfb5ea8 , 
    R_713_1dfb87e8 , 
    R_685_1dfb2f28 , 
    R_3fe_1d9d9f08 , 
    R_638_1dfaff08 , 
    R_465_1d9dda68 , 
    R_b91_1e6b57c8 , 
    R_b53_1e6b3108 , 
    R_8ad_1e098888 , 
    R_59e_1dd9e068 , 
    R_9c5_1e1837e8 , 
    R_3a9_1d9d64e8 , 
    R_3b3_1d9d6b28 , 
    R_2b4_1d9fcb68 , 
    R_af3_1e6af508 , 
    R_4f9_1dda3748 , 
    R_a90_1e18b6c8 , 
    R_389_1d9d50e8 , 
    R_a6a_1e18a408 , 
    R_b1b_1e6b0e08 , 
    R_4f8_1dda36a8 , 
    R_b66_1e6b9be8 , 
    R_9d0_1e183ec8 , 
    R_2e1_1d9ce7e8 , 
    R_7d2_1e0904a8 , 
    R_803_1e091e48 , 
    R_91e_1e09d428 , 
    R_4f7_1dda3608 , 
    R_ab4_1e18cd48 , 
    R_6ee_1dfb75c8 , 
    R_c05_1e6ba048 , 
    R_704_1dfb7e88 , 
    R_353_1d9d2f28 , 
    R_ba7_1e6b6588 , 
    R_87c_1e0969e8 , 
    R_3f5_1d9d9468 , 
    R_abc_1e18d248 , 
    R_a83_1e18aea8 , 
    R_b40_1e6b2528 , 
    R_a06_1e186588 , 
    R_907_1e09c0c8 , 
    R_664_1dfb1a88 , 
    R_b71_1e6b43c8 , 
    R_4f6_1ddad2e8 , 
    R_8b9_1e099008 , 
    R_971_1e180368 , 
    R_64e_1dfb11c8 , 
    R_679_1dfb27a8 , 
    R_80c_1e0923e8 , 
    R_347_1d9d27a8 , 
    R_b28_1e6b1628 , 
    R_7cf_1e08fdc8 , 
    R_8fc_1e09b9e8 , 
    R_72d_1dfb9828 , 
    R_9c4_1e183748 , 
    R_997_1e181b28 , 
    R_85f_1e0957c8 , 
    R_2d4_1d9cdfc8 , 
    R_48f_1dd9f508 , 
    R_adb_1e6ae608 , 
    R_3b9_1d9d6ee8 , 
    R_a51_1e188f68 , 
    R_8cb_1e099b48 , 
    R_2d8_1d9ce248 , 
    R_a72_1e18a908 , 
    R_7f7_1e0916c8 , 
    R_4b5_1dda0cc8 , 
    R_88b_1e097348 , 
    R_aa7_1e18c528 , 
    R_699_1dfb3ba8 , 
    R_68a_1dfb3748 , 
    R_9cf_1e183e28 , 
    R_345_1d9d2668 , 
    R_76b_1dfbbee8 , 
    R_7aa_1e099328 , 
    R_5e9_1ddacd48 , 
    R_a04_1e185f48 , 
    R_36b_1d9d3e28 , 
    R_444_1d9dc5c8 , 
    R_842_1e094aa8 , 
    R_58a_1dda96e8 , 
    R_97b_1e1809a8 , 
    R_5bc_1ddab128 , 
    R_ae9_1e6aeec8 , 
    R_74e_1dfbc348 , 
    R_69b_1dfb3ce8 , 
    R_783_1dfbcde8 , 
    R_64d_1dfb0c28 , 
    R_938_1e17dfc8 , 
    R_7bd_1e08f288 , 
    R_7ca_1e08ffa8 , 
    R_482_1ddac668 , 
    R_2c7_1d9fd748 , 
    R_621_1dfaf0a8 , 
    R_9c3_1e1836a8 , 
    R_309_1d9d00e8 , 
    R_5f1_1ddad248 , 
    R_4b8_1dda0ea8 , 
    R_bcf_1e6b7e88 , 
    R_824_1e0932e8 , 
    R_6e6_1dfb70c8 , 
    R_7a4_1e08e2e8 , 
    R_59d_1dda9dc8 , 
    R_769_1dfbbda8 , 
    R_38a_1d9d5688 , 
    R_4cb_1dda1a88 , 
    R_8d9_1e09a408 , 
    R_8d2_1e09a4a8 , 
    R_b24_1e6b13a8 , 
    R_4ba_1d9d9a08 , 
    R_bdd_1e6b8748 , 
    R_398_1d9d5a48 , 
    R_31d_1d9d0d68 , 
    R_47a_1dd9ece8 , 
    R_2ca_1d9ce108 , 
    R_b03_1e6aff08 , 
    R_2a0_1d9fbee8 , 
    R_71f_1dfb8f68 , 
    R_950_1e17eec8 , 
    R_9ce_1e184288 , 
    R_aae_1e6b6c68 , 
    R_b39_1e6b20c8 , 
    R_906_1e090ea8 , 
    R_786_1dfbd4c8 , 
    R_81c_1e092de8 , 
    R_94b_1e17eba8 , 
    R_8fb_1e09b948 , 
    R_3cb_1d9d7a28 , 
    R_86f_1e0961c8 , 
    R_584_1dda8e28 , 
    R_40a_1d9da688 , 
    R_954_1e17f148 , 
    R_944_1e17e748 , 
    R_bc8_1e6b7a28 , 
    R_9a1_1e182168 , 
    R_c02_1e6ba5e8 , 
    R_967_1e17fd28 , 
    R_7ff_1e091bc8 , 
    R_329_1d9d14e8 , 
    R_ba1_1e6b61c8 , 
    R_717_1dfb8a68 , 
    R_aa1_1e18c168 , 
    R_591_1dda9648 , 
    R_99c_1e181e48 , 
    R_a42_1e188b08 , 
    R_ba8_1e6b6628 , 
    R_ae1_1e6ae9c8 , 
    R_9c2_1e183b08 , 
    R_6bb_1dfb50e8 , 
    R_41b_1d9dac28 , 
    R_93d_1e17e2e8 , 
    R_5b2_1ddaafe8 , 
    R_5d6_1d9dd388 , 
    R_402_1d9da188 , 
    R_4b0_1dda09a8 , 
    R_549_1dda6948 , 
    R_53a_1dda64e8 , 
    R_70d_1dfb8428 , 
    R_aa4_1e18c348 , 
    R_798_1dfbdb08 , 
    R_7fb_1e091948 , 
    R_32a_1d9d1a88 , 
    R_a36_1e188388 , 
    R_5ed_1ddacfc8 , 
    R_b9a_1e6b6268 , 
    R_c07_1e6ba188 , 
    R_47e_1dd9ef68 , 
    R_ad2_1e6ae568 , 
    R_39d_1d9d5d68 , 
    R_83f_1e0943c8 , 
    R_7eb_1e090f48 , 
    R_42e_1d9dbd08 , 
    R_b51_1e6b2fc8 , 
    R_6b4_1dfb4c88 , 
    R_694_1dfb3888 , 
    R_68f_1dfb3568 , 
    R_777_1dfbc668 , 
    R_7b0_1e08ea68 , 
    R_7a0_1e08e068 , 
    R_75e_1dfbbbc8 , 
    R_5b7_1ddaae08 , 
    R_63d_1dfb0228 , 
    R_636_1dfb02c8 , 
    R_8de_1e09ac28 , 
    R_2ef_1d9cf0a8 , 
    R_302_1d9d4508 , 
    R_9b8_1e182fc8 , 
    R_4b2_1dda14e8 , 
    R_8e4_1e09aae8 , 
    R_3de_1d9d8b08 , 
    R_ab8_1e18cfc8 , 
    R_71b_1dfb8ce8 , 
    R_c0c_1e6ba4a8 , 
    R_c2b_1e6bb808 , 
    R_5ac_1ddaa728 , 
    R_853_1e095048 , 
    R_2aa_1d9fca28 , 
    R_385_1d9d4e68 , 
    R_436_1d9dc208 , 
    R_a60_1e1898c8 , 
    R_7bb_1e08f148 , 
    R_811_1e092708 , 
    R_4c5_1dda16c8 , 
    R_406_1d9da408 , 
    R_473_1dd9e388 , 
    R_8aa_1e098ba8 , 
    R_b7e_1e6b50e8 , 
    R_7b5_1e08ed88 , 
    R_5fb_1ddad888 , 
    R_34d_1d9d2b68 , 
    R_ae3_1e6aeb08 , 
    R_6f3_1dfb73e8 , 
    R_82b_1e093748 , 
    R_72a_1dfbacc8 , 
    R_bc3_1e6b7708 , 
    R_8fa_1e09bda8 , 
    R_567_1dda7c08 , 
    R_89f_1e097fc8 , 
    R_3ed_1d9d8f68 , 
    R_599_1dda9b48 , 
    R_851_1e094f08 , 
    R_2dd_1d9ce568 , 
    R_4a8_1dda04a8 , 
    R_8a9_1e098608 , 
    R_366_1d9d4008 , 
    R_376_1ddad568 , 
    R_75d_1dfbb628 , 
    R_59a_1ddaa0e8 , 
    R_4c2_1dda19e8 , 
    R_8be_1e08eba8 , 
    R_2c5_1d9fd608 , 
    R_595_1dda98c8 , 
    R_446_1d9dd108 , 
    R_6c5_1dfb5728 , 
    R_5d8_1ddac2a8 , 
    R_682_1dfb3248 , 
    R_64b_1dfb0ae8 , 
    R_791_1dfbd6a8 , 
    R_b7b_1e6b4a08 , 
    R_3b1_1d9d69e8 , 
    R_7e9_1e090e08 , 
    R_beb_1e6b9008 , 
    R_6c0_1dfb5408 , 
    R_8ba_1e0995a8 , 
    R_a8e_1e17f508 , 
    R_3c8_1d9d7848 , 
    R_be4_1e6b8ba8 , 
    R_544_1dda6628 , 
    R_53f_1dda6308 , 
    R_90e_1e09ca28 , 
    R_381_1d9d4be8 , 
    R_a3e_1e188888 , 
    R_6fd_1dfb7a28 , 
    R_a3a_1e188608 , 
    R_8c2_1e099aa8 , 
    R_af0_1e6af328 , 
    R_296_1d9fb8a8 , 
    R_b12_1e6b0d68 , 
    R_ba9_1e6b66c8 , 
    R_b1d_1e6b0f48 , 
    R_2b5_1d9fcc08 , 
    R_6ff_1dfb7b68 , 
    R_a98_1e18bbc8 , 
    R_58e_1dda9968 , 
    R_753_1dfbafe8 , 
    R_3c5_1d9d7668 , 
    R_447_1d9dc7a8 , 
    R_61f_1dfaef68 , 
    R_54e_1dda28e8 , 
    R_6f8_1dfb7708 , 
    R_3a4_1d9d61c8 , 
    R_423_1d9db128 , 
    R_6a4_1dfb4288 , 
    R_b9b_1e6b5e08 , 
    R_a07_1e186128 , 
    R_55f_1dda7708 , 
    R_79d_1dfbde28 , 
    R_66d_1dfb2028 , 
    R_5e2_1ddacde8 , 
    R_48b_1dd9f288 , 
    R_5ee_1dda3a68 , 
    R_6c6_1dfb2d48 , 
    R_3e3_1d9d8928 , 
    R_b83_1e6b4f08 , 
    R_533_1dda5b88 , 
    R_42d_1d9db768 , 
    R_7e0_1e090868 , 
    R_696_1dfb3ec8 , 
    R_3f9_1d9d96e8 , 
    R_b88_1e6b5228 , 
    R_758_1dfbb308 , 
    R_3d2_1d9d8388 , 
    R_534_1dda5c28 , 
    R_532_1d9d1308 , 
    R_867_1e095cc8 , 
    R_2b6_1d9fd1a8 , 
    R_775_1dfbc528 , 
    R_3e8_1d9d8c48 , 
    R_4d0_1dda1da8 , 
    R_30d_1d9d0368 , 
    R_4e7_1dda2c08 , 
    R_70a_1dfb8748 , 
    R_a58_1e1893c8 , 
    R_4e8_1dda2ca8 , 
    R_4e6_1dda3068 , 
    R_535_1dda5cc8 , 
    R_5ea_1dda37e8 , 
    R_929_1e09d608 , 
    R_448_1d9dc848 , 
    R_b0b_1e6b0408 , 
    R_319_1d9d0ae8 , 
    R_985_1e180fe8 , 
    R_32f_1d9d18a8 , 
    R_4e9_1dda2d48 , 
    R_b1f_1e6b1088 , 
    R_495_1dd9f8c8 , 
    R_63b_1dfb00e8 , 
    R_536_1dda6268 , 
    R_3d9_1d9d82e8 , 
    R_a4f_1e188e28 , 
    R_470_1dd9e1a8 , 
    R_2d5_1d9ce068 , 
    R_3f0_1d9d9148 , 
    R_acf_1e18de28 , 
    R_ac2_1e18db08 , 
    R_9b4_1e182d48 , 
    R_a05_1e185fe8 , 
    R_2d9_1d9ce2e8 , 
    R_8ed_1e09b088 , 
    R_3f3_1d9d9328 , 
    R_af2_1e6af968 , 
    R_44d_1d9dcb68 , 
    R_645_1dfb0728 , 
    R_648_1dfb0908 , 
    R_4a1_1dda0048 , 
    R_749_1dfba9a8 , 
    R_2c8_1d9fd7e8 , 
    R_3bc_1d9d70c8 , 
    R_3f6_1ddad7e8 , 
    R_596_1dda9e68 , 
    R_c01_1e6b9dc8 , 
    R_734_1dfb9c88 , 
    R_5a5_1ddaa2c8 , 
    R_6e3_1dfb69e8 , 
    R_914_1e09c8e8 , 
    R_43d_1d9dc168 , 
    R_2cb_1d9fd9c8 , 
    R_3d0_1d9d7d48 , 
    R_b67_1e6b3d88 , 
    R_b01_1e6afdc8 , 
    R_37d_1d9d4968 , 
    R_a80_1e18acc8 , 
    R_9bd_1e1832e8 , 
    R_339_1d9d1ee8 , 
    R_7ad_1e08e888 , 
    R_972_1e180908 , 
    R_a22_1e184788 , 
    R_486_1ddacb68 , 
    R_5d5_1ddac0c8 , 
    R_592_1dda9be8 , 
    R_449_1d9dc8e8 , 
    R_87b_1e096948 , 
    R_8f5_1e09b588 , 
    R_35a_1d9d3888 , 
    R_37a_1ddab9e8 , 
    R_991_1e181768 , 
    R_62a_1dfb1448 , 
    R_808_1e092168 , 
    R_3a6_1d9d6808 , 
    R_b95_1e6b5a48 , 
    R_83e_1e17e108 , 
    R_386_1d9d5408 , 
    R_90d_1e09c488 , 
    R_931_1e09db08 , 
    R_ac9_1e18da68 , 
    R_a31_1e187b68 , 
    R_640_1dfb0408 , 
    R_667_1dfb1c68 , 
    R_6cb_1dfb5ae8 , 
    R_74a_1e17f288 , 
    R_676_1dfb2ac8 , 
    R_372_1d9d4788 , 
    R_56c_1dda7f28 , 
    R_334_1d9d1bc8 , 
    R_31e_1d9fc528 , 
    R_981_1e180d68 , 
    R_8ca_1e099fa8 , 
    R_85e_1e095c28 , 
    R_bbe_1e6af6e8 , 
    R_49b_1dd9fc88 , 
    R_73a_1dfba548 , 
    R_5fe_1dfaf8c8 , 
    R_98b_1e1813a8 , 
    R_88e_1e097a28 , 
    R_28f_1d9fb448 , 
    R_9bc_1e183248 , 
    R_5db_1ddac488 , 
    R_88a_1e08ee28 , 
    R_5a6_1ddaa868 , 
    R_443_1d9dc528 , 
    R_a0a_1e186808 , 
    R_358_1d9d3248 , 
    R_88f_1e0975c8 , 
    R_acc_1e18dc48 , 
    R_aac_1e18c848 , 
    R_2a2_1d9fde28 , 
    R_8a5_1e098388 , 
    R_8ec_1e09afe8 , 
    R_289_1d9fb088 , 
    R_340_1d9d2348 , 
    R_c2d_1e6bb948 , 
    R_964_1e17fb48 , 
    R_85d_1e095688 , 
    R_6fa_1dfb7d48 , 
    R_4d5_1dda20c8 , 
    R_a5a_1e18b308 , 
    R_7de_1e090c28 , 
    R_605_1ddadec8 , 
    R_311_1d9d05e8 , 
    R_8a6_1e098928 , 
    R_a2f_1e187a28 , 
    R_81f_1e092fc8 , 
    R_3b6_1d9d7208 , 
    R_315_1d9d0868 , 
    R_93f_1e17e428 , 
    R_5b1_1ddaaa48 , 
    R_631_1dfafaa8 , 
    R_890_1e097668 , 
    R_670_1dfb2208 , 
    R_b9c_1e6b5ea8 , 
    R_8e9_1e09ae08 , 
    R_932_1e093928 , 
    R_817_1e092ac8 , 
    R_b60_1e6b3928 , 
    R_979_1e180868 , 
    R_8d8_1e09a368 , 
    R_628_1dfaf508 , 
    R_729_1dfb95a8 , 
    R_a92_1e18bd08 , 
    R_b33_1e6b1d08 , 
    R_2ab_1d9fc5c8 , 
    R_5e6_1dd9f6e8 , 
    R_5c0_1ddab3a8 , 
    R_600_1ddadba8 , 
    R_8f4_1e09b4e8 , 
    R_29d_1d9fbd08 , 
    R_c11_1e6ba7c8 , 
    R_4d7_1dda2208 , 
    R_b43_1e6b2708 , 
    R_881_1e096d08 , 
    R_891_1e097708 , 
    R_8b4_1e098ce8 , 
    R_6ac_1dfb4788 , 
    R_2f0_1d9cf148 , 
    R_ad8_1e6ae428 , 
    R_9bb_1e1831a8 , 
    R_bd9_1e6b84c8 , 
    R_39f_1d9d5ea8 , 
    R_a5e_1e189c88 , 
    R_303_1d9cfd28 , 
    R_6ae_1dfb4dc8 , 
    R_477_1dd9e608 , 
    R_6d2_1e0981a8 , 
    R_38f_1d9d54a8 , 
    R_4d2_1dda23e8 , 
    R_82f_1e0939c8 , 
    R_61d_1dfaee28 , 
    R_673_1dfb23e8 , 
    R_578_1dda86a8 , 
    R_a65_1e189be8 , 
    R_9a5_1e1823e8 , 
    R_744_1dfba688 , 
    R_bfe_1e6ba0e8 , 
    R_86e_1e096628 , 
    R_6ce_1e0945a8 , 
    R_9df_1e184828 , 
    R_571_1dda8248 , 
    R_9e0_1e1848c8 , 
    R_9de_1e184c88 , 
    R_41a_1ddabee8 , 
    R_36e_1d9d1588 , 
    R_6b9_1dfb4fa8 , 
    R_b72_1e6b4968 , 
    R_73f_1dfba368 , 
    R_a4d_1e188ce8 , 
    R_9e1_1e184968 , 
    R_2d0_1d9fdce8 , 
    R_72e_1dfb9dc8 , 
    R_c25_1e6bb448 , 
    R_8eb_1e09af48 , 
    R_6eb_1dfb6ee8 , 
    R_764_1dfbba88 , 
    R_9b1_1e182b68 , 
    R_970_1e1802c8 , 
    R_bce_1e6b82e8 , 
    R_325_1d9d1268 , 
    R_65c_1dfb1588 , 
    R_643_1dfb05e8 , 
    R_abf_1e18d428 , 
    R_a9b_1e18bda8 , 
    R_b7c_1e6b4aa8 , 
    R_9ba_1e183608 , 
    R_bef_1e6b9288 , 
    R_b14_1e6b09a8 , 
    R_996_1e181f88 , 
    R_812_1e092ca8 , 
    R_4a2_1dda05e8 , 
    R_6e0_1dfb6808 , 
    R_490_1dd9f5a8 , 
    R_711_1dfb86a8 , 
    R_a86_1e18ba88 , 
    R_342_1d9d2988 , 
    R_c0e_1e6baae8 , 
    R_8e3_1e09aa48 , 
    R_646_1dfb0cc8 , 
    R_74d_1dfbac28 , 
    R_67f_1dfb2b68 , 
    R_34f_1d9d2ca8 , 
    R_8f3_1e09b448 , 
    R_bdc_1e6b86a8 , 
    R_57f_1dda8b08 , 
    R_77a_1dfbcd48 , 
    R_4c1_1dda1448 , 
    R_b8e_1e6b5ae8 , 
    R_c29_1e6bb6c8 , 
    R_875_1e096588 , 
    R_852_1e0954a8 , 
    R_6a6_1dfb48c8 , 
    R_76f_1dfbc168 , 
    R_984_1e180f48 , 
    R_39a_1d9d6088 , 
    R_35f_1d9d36a8 , 
    R_5d0_1ddabda8 , 
    R_b65_1e6b3c48 , 
    R_92b_1e09d748 , 
    R_3eb_1d9d8e28 , 
    R_53b_1dda6088 , 
    R_97a_1e180e08 , 
    R_369_1d9d3ce8 , 
    R_7f5_1e091588 , 
    R_588_1dda90a8 , 
    R_b6a_1e6b4468 , 
    R_435_1d9dbc68 , 
    R_a08_1e1861c8 , 
    R_7ef_1e0911c8 , 
    R_781_1dfbcca8 , 
    R_55c_1dda7528 , 
    R_3bf_1d9d72a8 , 
    R_850_1e094e68 , 
    R_2ea_1d9cf288 , 
    R_687_1dfb3068 , 
    R_795_1dfbd928 , 
    R_382_1d9d5188 , 
    R_63e_1dfb07c8 , 
    R_2b7_1d9fcd48 , 
    R_9b0_1e182ac8 , 
    R_6dd_1dfb6628 , 
    R_4be_1dda1768 , 
    R_bfd_1e6b9b48 , 
    R_b0d_1e6b0548 , 
    R_b9d_1e6b5f48 , 
    R_b3a_1e6b2668 , 
    R_4b9_1dda0f48 , 
    R_4bb_1dda1088 , 
    R_9a0_1e1820c8 , 
    R_83b_1e094148 , 
    R_8ea_1e09b3a8 , 
    R_b21_1e6b11c8 , 
    R_62f_1dfaf968 , 
    R_91d_1e09ce88 , 
    R_483_1dd9ed88 , 
    R_7c0_1e08f468 , 
    R_bd5_1e6b8248 , 
    R_364_1d9d39c8 , 
    R_322_1d9d2e88 , 
    R_326_1d9d1808 , 
    R_99b_1e181da8 , 
    R_961_1e17f968 , 
    R_726_1dfb98c8 , 
    R_a7d_1e18aae8 , 
    R_826_1e09de28 , 
    R_89a_1dfb4648 , 
    R_511_1dda4648 , 
    R_2fb_1d9cf828 , 
    R_b5c_1e6b36a8 , 
    R_8b0_1e098a68 , 
    R_708_1dfb8108 , 
    R_603_1ddadd88 , 
    R_804_1e091ee8 , 
    R_573_1dda8388 , 
    R_a56_1e189a08 , 
    R_510_1dda45a8 , 
    R_833_1e093c48 , 
    R_8c1_1e099508 , 
    R_966_1e180188 , 
    R_46d_1dd9dfc8 , 
    R_bcc_1e6b7ca8 , 
    R_47b_1dd9e888 , 
    R_aea_1e6af468 , 
    R_8d1_1e099f08 , 
    R_57a_1ddaa368 , 
    R_8f2_1e09b8a8 , 
    R_b35_1e6b1e48 , 
    R_b05_1e6b0048 , 
    R_aa9_1e18c668 , 
    R_9b7_1e182f28 , 
    R_3ae_1d9d6d08 , 
    R_50f_1dda4508 , 
    R_a23_1e1872a8 , 
    R_2c9_1d9fd888 , 
    R_5c6_1d9d7e88 , 
    R_8bd_1e099288 , 
    R_4b1_1dda0a48 , 
    R_b45_1e6b2848 , 
    R_422_1d9db588 , 
    R_2cc_1d9fda68 , 
    R_9d5_1e1841e8 , 
    R_37e_1d9d4f08 , 
    R_42c_1d9db6c8 , 
    R_a7e_1e18b088 , 
    R_a8d_1e18b4e8 , 
    R_50e_1dda4968 , 
    R_626_1dfafb48 , 
    R_5cc_1ddabb28 , 
    R_295_1d9fb808 , 
    R_a9e_1e18c488 , 
    R_80d_1e092488 , 
    R_9af_1e182a28 , 
    R_946_1e17ed88 , 
    R_a5c_1e189648 , 
    R_5bb_1ddab088 , 
    R_3e6_1d9d9008 , 
    R_ab3_1e18cca8 , 
    R_a1e_1e187488 , 
    R_66a_1dfb2348 , 
    R_7f8_1e091768 , 
    R_56e_1dda8568 , 
    R_3c2_1d9d7988 , 
    R_837_1e093ec8 , 
    R_866_1e096128 , 
    R_65a_1dfb1948 , 
    R_4aa_1dda0ae8 , 
    R_540_1dda63a8 , 
    R_61b_1dfaece8 , 
    R_78a_1dfbd748 , 
    R_76c_1dfbbf88 , 
    R_4c7_1dda1808 , 
    R_47f_1dd9eb08 , 
    R_34a_1d9d4a08 , 
    R_b57_1e6b3388 , 
    R_545_1dda66c8 , 
    R_c13_1e6ba908 , 
    R_44c_1d9dcac8 , 
    R_a0b_1e1863a8 , 
    R_6d5_1dfb6128 , 
    R_bf3_1e6b9508 , 
    R_3ee_1d9d9508 , 
    R_6d7_1dfb6268 , 
    R_3d6_1d9d9788 , 
    R_b06_1e6b05e8 , 
    R_9d4_1e184148 , 
    R_33b_1d9d2028 , 
    R_739_1dfb9fa8 , 
    R_a0e_1e186a88 , 
    R_7dd_1e090688 , 
    R_54f_1dda6d08 , 
    R_926_1e09dba8 , 
    R_abb_1e18d1a8 , 
    R_70e_1dfb89c8 , 
    R_ba2_1e6b6768 , 
    R_917_1e09cac8 , 
    R_923_1e09d248 , 
    R_784_1dfbce88 , 
    R_920_1e09d068 , 
    R_564_1dda7a28 , 
    R_9a9_1e182668 , 
    R_bfa_1e6b9e68 , 
    R_62c_1dfaf788 , 
    R_8c9_1e099a08 , 
    R_43c_1d9dc0c8 , 
    R_b00_1e6afd28 , 
    R_35d_1d9d3568 , 
    R_c18_1e6bac28 , 
    R_306_1d9d0408 , 
    R_939_1e17e068 , 
    R_474_1dd9e428 , 
    R_4a9_1dda0548 , 
    R_2ac_1d9fc668 , 
    R_609_1dfae1a8 , 
    R_94c_1e17ec48 , 
    R_90a_1e09c7a8 , 
    R_92e_1e0918a8 , 
    R_7be_1e08f828 , 
    R_825_1e093388 , 
    R_559_1dda7348 , 
    R_bf7_1e6b9788 , 
    R_87a_1e096da8 , 
    R_9d3_1e1840a8 , 
    R_394_1d9d57c8 , 
    R_31a_1d9d1088 , 
    R_69f_1dfb3f68 , 
    R_787_1dfbd068 , 
    R_a63_1e189aa8 , 
    R_9ae_1e183388 , 
    R_945_1e17e7e8 , 
    R_537_1dda5e08 , 
    R_725_1dfb9328 , 
    R_b68_1e6b3e28 , 
    R_7a5_1e08e388 , 
    R_4eb_1dda2e88 , 
    R_619_1dfaeba8 , 
    R_800_1e091c68 , 
    R_be8_1e6b8e28 , 
    R_4ec_1dda2f28 , 
    R_4ea_1dda32e8 , 
    R_2f1_1d9cf1e8 , 
    R_5d3_1ddabf88 , 
    R_6da_1dfb6948 , 
    R_5b6_1ddab268 , 
    R_3ac_1d9d66c8 , 
    R_983_1e180ea8 , 
    R_b73_1e6b4508 , 
    R_4ed_1dda2fc8 , 
    R_ada_1e6aea68 , 
    R_7fc_1e0919e8 , 
    R_b3c_1e6b22a8 , 
    R_304_1d9cfdc8 , 
    R_5ab_1ddaa688 , 
    R_85c_1e0955e8 , 
    R_442_1d9dcc08 , 
    R_3ce_1d9d8608 , 
    R_ad5_1e6ae248 , 
    R_ae8_1e6aee28 , 
    R_3b4_1d9d6bc8 , 
    R_8b8_1e098f68 , 
    R_b46_1e6b2de8 , 
    R_8e8_1e09ad68 , 
    R_bbf_1e6b7488 , 
    R_799_1dfbdba8 , 
    R_778_1dfbc708 , 
    R_a4b_1e188ba8 , 
    R_51d_1dda4dc8 , 
    R_657_1dfb1268 , 
    R_9d2_1e17f788 , 
    R_348_1d9d2848 , 
    R_51c_1dda4d28 , 
    R_8d7_1e09a2c8 , 
    R_9b3_1e182ca8 , 
    R_7db_1e090548 , 
    R_715_1dfb8928 , 
    R_68c_1dfb3388 , 
    R_880_1e096c68 , 
    R_29c_1d9fbc68 , 
    R_b7d_1e6b4b48 , 
    R_51b_1dda4c88 , 
    R_bba_1e6b7668 , 
    R_3dc_1d9d84c8 , 
    R_5a0_1dda9fa8 , 
    R_75f_1dfbb768 , 
    R_b7f_1e6b4c88 , 
    R_b16_1e6b0fe8 , 
    R_ba3_1e6b6308 , 
    R_654_1dfb1088 , 
    R_bc7_1e6b7988 , 
    R_2a3_1d9fc0c8 , 
    R_6f0_1dfb7208 , 
    R_7a1_1e08e108 , 
    R_371_1d9d41e8 , 
    R_51a_1dda50e8 , 
    R_ab7_1e18cf28 , 
    R_7e6_1e099828 , 
    R_b6b_1e6b4008 , 
    R_9ad_1e1828e8 , 
    R_935_1e09dd88 , 
    R_b8a_1e6bb768 , 
    R_69d_1dfb3e28 , 
    R_45e_1d9ddb08 , 
    R_a1a_1e187208 , 
    R_a49_1e188a68 , 
    R_a09_1e186268 , 
    R_496_1dd9fe68 , 
    R_336_1d9d2208 , 
    R_5df_1ddac708 , 
    R_5c7_1ddab808 , 
    R_990_1e1816c8 , 
    R_6c9_1dfb59a8 , 
    R_2eb_1d9cee28 , 
    R_2b8_1d9fcde8 , 
    R_ae0_1e6ae928 , 
    R_b2f_1e6b1a88 , 
    R_84d_1e094c88 , 
    R_a12_1e186d08 , 
    R_74f_1dfbad68 , 
    R_a35_1e187de8 , 
    R_28e_1d9fb3a8 , 
    R_81a_1e0936a8 , 
    R_487_1dd9f008 , 
    R_c1c_1e6baea8 , 
    R_7a8_1e08e568 , 
    R_471_1dd9e248 , 
    R_766_1e0986a8 , 
    R_38b_1d9d5228 , 
    R_a7b_1e18a9a8 , 
    R_b52_1e6b8568 , 
    R_9ff_1e185c28 , 
    R_7b9_1e08f008 , 
    R_67b_1dfb28e8 , 
    R_a00_1e185cc8 , 
    R_9fe_1e6bb9e8 , 
    R_980_1e180cc8 , 
    R_874_1e0964e8 , 
    R_49c_1dd9fd28 , 
    R_58c_1dda9328 , 
    R_45f_1d9dd6a8 , 
    R_98a_1e181808 , 
    R_8e2_1e09aea8 , 
    R_6ba_1dfb5548 , 
    R_bd8_1e6b8428 , 
    R_a8b_1e18b3a8 , 
    R_a01_1e185d68 , 
    R_6b3_1dfb4be8 , 
    R_60d_1dfae428 , 
    R_6e8_1dfb6d08 , 
    R_399_1d9d5ae8 , 
    R_a16_1e186f88 , 
    R_bc2_1e6b7b68 , 
    R_32b_1d9d1628 , 
    R_434_1d9dbbc8 , 
    R_a24_1e187348 , 
    R_377_1d9d45a8 , 
    R_3cc_1d9d7ac8 , 
    R_a68_1e189dc8 , 
    R_963_1e17faa8 , 
    R_7c5_1e08f788 , 
    R_615_1dfae928 , 
    R_8a2_1dfb9b48 , 
    R_722_1dfb9648 , 
    R_288_1d9f96e8 , 
    R_556_1dda7668 , 
    R_748_1dfba908 , 
    R_865_1e095b88 , 
    R_607_1dfae068 , 
    R_691_1dfb36a8 , 
    R_978_1e1807c8 , 
    R_84f_1e094dc8 , 
    R_2cd_1d9fdb08 , 
    R_ae2_1e6aef68 , 
    R_a1f_1e187028 , 
    R_721_1dfb90a8 , 
    R_733_1dfb9be8 , 
    R_9e3_1e184aa8 , 
    R_9e4_1e184b48 , 
    R_c23_1e6bb308 , 
    R_9e2_1e184f08 , 
    R_7ae_1dfbb1c8 , 
    R_91a_1e09d1a8 , 
    R_b84_1e6b4fa8 , 
    R_b92_1e181088 , 
    R_ba4_1e6b63a8 , 
    R_754_1dfbb088 , 
    R_5a4_1ddaa228 , 
    R_9a4_1e182348 , 
    R_b08_1e6b0228 , 
    R_9e5_1e184be8 , 
    R_617_1dfaea68 , 
    R_5ce_1ddac168 , 
    R_b89_1e6b52c8 , 
    R_7b2_1e09b128 , 
    R_460_1d9dd748 , 
    R_5e4_1ddaca28 , 
    R_30a_1d9d0688 , 
    R_a0c_1e186448 , 
    R_910_1e09c668 , 
    R_553_1dda6f88 , 
    R_86d_1e096088 , 
    R_a0f_1e186628 , 
    R_719_1dfb8ba8 , 
    R_b48_1e6b2a28 , 
    R_316_1d9d0e08 , 
    R_901_1e09bd08 , 
    R_611_1dfae6a8 , 
    R_ac5_1e18d7e8 , 
    R_6c4_1dfb5688 , 
    R_53c_1dda6128 , 
    R_712_1dfb8c48 , 
    R_2f6_1d9cfc88 , 
    R_829_1e093608 , 
    R_89d_1e097e88 , 
    R_8d0_1e099e68 , 
    R_8ac_1e0987e8 , 
    R_8a0_1e098068 , 
    R_aef_1e6af288 , 
    R_759_1dfbb3a8 , 
    R_a6d_1e18a0e8 , 
    R_6bf_1dfb5368 , 
    R_982_1e182c08 , 
    R_bdb_1e6b8608 , 
    R_684_1dfb2e88 , 
    R_7b7_1e08eec8 , 
    R_478_1dd9e6a8 , 
    R_be1_1e6b89c8 , 
    R_b55_1e6b3248 , 
    R_79b_1dfbdce8 , 
    R_c27_1e6bb588 , 
    R_96f_1e180228 , 
    R_42b_1d9db628 , 
    R_6cd_1dfb5c28 , 
    R_652_1dfb16c8 , 
    R_71d_1dfb8e28 , 
    R_703_1dfb7de8 , 
    R_a54_1e189148 , 
    R_4a3_1dda0188 , 
    R_634_1dfafc88 , 
    R_2ad_1d9fc708 , 
    R_4cc_1dda1b28 , 
    R_2a1_1d9fbf88 , 
    R_93a_1e0977a8 , 
    R_a78_1e18a7c8 , 
    R_c03_1e6b9f08 , 
    R_72c_1dfb9788 , 
    R_809_1e092208 , 
    R_5b0_1ddaa9a8 , 
    R_44b_1d9dca28 , 
    R_952_1ddab768 , 
    R_899_1e097c08 , 
    R_bd4_1e6b81a8 , 
    R_a94_1e18b948 , 
    R_6b1_1dfb4aa8 , 
    R_491_1dd9f648 , 
    R_5ca_1d9dae08 , 
    R_6f5_1dfb7528 , 
    R_9c9_1e183a68 , 
    R_75a_1dfbb948 , 
    R_461_1d9dd7e8 , 
    R_7c3_1e08f648 , 
    R_569_1dda7d48 , 
    R_a75_1e18a5e8 , 
    R_7ec_1e090fe8 , 
    R_c20_1e6bb128 , 
    R_96d_1e1800e8 , 
    R_54a_1dda6ee8 , 
    R_b31_1e6b1bc8 , 
    R_5bf_1ddab308 , 
    R_900_1e09bc68 , 
    R_b74_1e6b45a8 , 
    R_940_1e17e4c8 , 
    R_8dd_1e09a688 , 
    R_a88_1e18b1c8 , 
    R_743_1dfba5e8 , 
    R_2d1_1d9fdd88 , 
    R_4b3_1dda0b88 , 
    R_48c_1dd9f328 , 
    R_419_1d9daae8 , 
    R_2ba_1d9fd428 , 
    R_898_1e097b68 , 
    R_354_1d9d2fc8 , 
    R_3c9_1d9d78e8 , 
    R_afd_1e6afb48 , 
    R_698_1dfb3b08 , 
    R_8c8_1e099968 , 
    R_aff_1e6afc88 , 
    R_59c_1dda9d28 , 
    R_43b_1d9dc028 , 
    R_3e1_1d9d87e8 , 
    R_7d8_1e090368 , 
    R_624_1dfaf288 , 
    R_ace_1e6ae2e8 , 
    R_294_1d9fb768 , 
    R_818_1e092b68 , 
    R_9c8_1e1839c8 , 
    R_5c8_1ddab8a8 , 
    R_c2f_1e6bba88 , 
    R_ba5_1e6b6448 , 
    R_6d0_1dfb5e08 , 
    R_820_1e093068 , 
    R_30e_1d9d0908 , 
    R_99f_1e182028 , 
    R_73e_1dfba7c8 , 
    R_4ef_1dda3108 , 
    R_451_1d9dcde8 , 
    R_678_1dfb2708 , 
    R_663_1dfb19e8 , 
    R_5fa_1e091128 , 
    R_312_1d9d0b88 , 
    R_a45_1e1887e8 , 
    R_b18_1e6b0c28 , 
    R_4f0_1dda31a8 , 
    R_4ee_1dda3568 , 
    R_7ab_1e08e748 , 
    R_305_1d9cfe68 , 
    R_955_1e17f1e8 , 
    R_373_1d9d4328 , 
    R_a39_1e188068 , 
    R_669_1dfb1da8 , 
    R_3a5_1d9d6268 , 
    R_c0d_1e6ba548 , 
    R_4f1_1dda3248 , 
    R_541_1dda6448 , 
    R_69a_1dfb4148 , 
    R_b90_1e6b5728 , 
    R_99a_1e182208 , 
    R_960_1e17f8c8 , 
    R_6a9_1dfb45a8 , 
    R_4bc_1dda1128 , 
    R_897_1e097ac8 , 
    R_701_1dfb7ca8 , 
    R_36c_1d9d3ec8 , 
    R_60b_1dfae2e8 , 
    R_583_1dda8d88 , 
    R_330_1d9d1948 , 
    R_bb6_1e6b73e8 , 
    R_71e_1dfb93c8 , 
    R_590_1dda95a8 , 
    R_29e_1dda2668 , 
    R_b0f_1e6b0688 , 
    R_a1b_1e186da8 , 
    R_550_1dda6da8 , 
    R_ac8_1e18d9c8 , 
    R_a9d_1e18bee8 , 
    R_561_1dda7848 , 
    R_80e_1e092a28 , 
    R_9b6_1e187708 , 
    R_5e8_1ddacca8 , 
    R_613_1dfae7e8 , 
    R_b6c_1e6b40a8 , 
    R_3d3_1d9d7f28 , 
    R_31f_1d9d0ea8 , 
    R_9c7_1e183928 , 
    R_5dd_1ddac5c8 , 
    R_78e_1dfbd9c8 , 
    R_a13_1e1868a8 , 
    R_70c_1dfb8388 , 
    R_885_1e096f88 , 
    R_85b_1e095548 , 
    R_8ff_1e09bbc8 , 
    R_716_1dfb8ec8 , 
    R_2b9_1d9fce88 , 
    R_b69_1e6b3ec8 , 
    R_356_1d9d3608 , 
    R_2e6_1d9cf008 , 
    R_484_1dd9ee28 , 
    R_2ec_1d9ceec8 , 
    R_acb_1e18dba8 , 
    R_813_1e092848 , 
    R_4c3_1dda1588 , 
    R_a47_1e188928 , 
    R_81d_1e092e88 , 
    R_8e7_1e09acc8 , 
    R_5ef_1ddad108 , 
    R_896_1e094828 , 
    R_bec_1e6b90a8 , 
    R_b2b_1e6b1808 , 
    R_4ab_1dda0688 , 
    R_7e4_1e090ae8 , 
    R_a33_1e187ca8 , 
    R_47c_1dd9e928 , 
    R_8d6_1e09a728 , 
    R_87f_1e096bc8 , 
    R_5b5_1ddaacc8 , 
    R_651_1dfb0ea8 , 
    R_3da_1d9d8888 , 
    R_538_1dda5ea8 , 
    R_675_1dfb2528 , 
    R_60f_1dfae568 , 
    R_29b_1d9fbbc8 , 
    R_aa6_1e18c988 , 
    R_3bd_1d9d7168 , 
    R_be5_1e6b8c48 , 
    R_c0a_1e6ba868 , 
    R_5f5_1ddad4c8 , 
    R_b4b_1e6b2c08 , 
    R_7b1_1e08eb08 , 
    R_95d_1e17f6e8 , 
    R_a17_1e186b28 , 
    R_a29_1e187668 , 
    R_71a_1dfb9148 , 
    R_693_1dfb37e8 , 
    R_77b_1dfbc8e8 , 
    R_9c6_1e183d88 , 
    R_3a7_1d9d63a8 , 
    R_bc0_1e6b7528 , 
    R_68e_1dfb39c8 , 
    R_335_1d9d1c68 , 
    R_5eb_1ddace88 , 
    R_ad7_1e6ae388 , 
    R_765_1dfbbb28 , 
    R_387_1d9d4fa8 , 
    R_9a8_1e1825c8 , 
    R_632_1dfb0048 , 
    R_6e5_1dfb6b28 , 
    R_772_1dfbc848 , 
    R_995_1e1819e8 , 
    R_7d6_1e090728 , 
    R_598_1dda9aa8 , 
    R_a70_1e18a2c8 , 
    R_a25_1e1873e8 , 
    R_bbb_1e6b7208 , 
    R_6f2_1dfb7848 , 
    R_a41_1e188568 , 
    R_a66_1e18a188 , 
    R_a3d_1e1882e8 , 
    R_341_1d9d23e8 , 
    R_594_1dda9828 , 
    R_4fe_1dda5868 , 
    R_480_1dd9eba8 , 
    R_6ab_1dfb46e8 , 
    R_84c_1e094be8 , 
    R_660_1dfb1808 , 
    R_a20_1e1870c8 , 
    R_abe_1e6b64e8 , 
    R_566_1dda8068 , 
    R_7c8_1e08f968 , 
    R_5c2_1d9fc2a8 , 
    R_989_1e181268 , 
    R_8a8_1e098568 , 
    R_2a4_1d9fc168 , 
    R_7d5_1e090188 , 
    R_8fe_1e09c028 , 
    R_3b7_1d9d6da8 , 
    R_6b8_1dfb4f08 , 
    R_8b3_1e098c48 , 
    R_94f_1e17ee28 , 
    R_9fb_1e1859a8 , 
    R_a10_1e1866c8 , 
    R_b36_1e6b23e8 , 
    R_aa0_1e18c0c8 , 
    R_c1a_1e6bb268 , 
    R_82c_1e0937e8 , 
    R_4d1_1dda1e48 , 
    R_6fc_1dfb7988 , 
    R_9fa_1e185e08 , 
    R_9fc_1e185a48 , 
    R_a0d_1e1864e8 , 
    R_be2_1e6b8f68 , 
    R_b02_1e6b8068 , 
    R_a28_1e1875c8 , 
    R_4fd_1dda39c8 , 
    R_5fd_1ddad9c8 , 
    R_873_1e096448 , 
    R_9fd_1e185ae8 , 
    R_a6b_1e189fa8 , 
    R_aa3_1e18c2a8 , 
    R_738_1dfb9f08 , 
    R_805_1e091f88 , 
    R_2f7_1d9cf5a8 , 
    R_5ba_1ddab4e8 , 
    R_57d_1dda89c8 , 
    R_475_1dd9e4c8 , 
    R_433_1d9dbb28 , 
    R_aed_1e6af148 , 
    R_4fc_1dda3928 , 
    R_3a0_1d9d5f48 , 
    R_3f7_1d9d95a8 , 
    R_367_1d9d3ba8 , 
    R_947_1e17e928 , 
    R_b1a_1e6b1268 , 
    R_525_1dda52c8 , 
    R_50d_1dda43c8 , 
    R_390_1d9d5548 , 
    R_6fe_1dfb7fc8 , 
    R_6f7_1dfb7668 , 
    R_2ae_1d9fcca8 , 
    R_864_1e095ae8 , 
    R_9e7_1e184d28 , 
    R_524_1dda5228 , 
    R_50c_1dda4328 , 
    R_9e6_1e185188 , 
    R_9e8_1e184dc8 , 
    R_9b2_1e183108 , 
    R_7e2_1dfbaf48 , 
    R_622_1dfaf648 , 
    R_b4e_1e184508 , 
    R_a91_1e18b768 , 
    R_a84_1e18af48 , 
    R_4ce_1dda2168 , 
    R_bb2_1e6b7168 , 
    R_523_1dda5188 , 
    R_50b_1dda4288 , 
    R_9e9_1e184e68 , 
    R_4f3_1dda3388 , 
    R_4fb_1dda3888 , 
    R_4f2_1ddad068 , 
    R_4f4_1dda3428 , 
    R_55e_1dda7b68 , 
    R_84e_1e095228 , 
    R_a76_1e18ab88 , 
    R_5c9_1ddab948 , 
    R_343_1d9d2528 , 
    R_a73_1e18a4a8 , 
    R_7cd_1e08fc88 , 
    R_522_1dda55e8 , 
    R_50a_1dda46e8 , 
    R_4f5_1dda34c8 , 
    R_396_1d9d5e08 , 
    R_7f9_1e091808 , 
    R_681_1dfb2ca8 , 
    R_37b_1d9d4828 , 
    R_639_1dfaffa8 , 
    R_76d_1dfbc028 , 
    R_78b_1dfbd2e8 , 
    R_6a3_1dfb41e8 , 
    R_9ac_1e182848 , 
    R_86c_1e095fe8 , 
    R_c08_1e6ba228 , 
    R_2fc_1d9cf8c8 , 
    R_7f0_1e091268 , 
    R_c31_1e6bbbc8 , 
    R_a52_1e189508 , 
    R_ab2_1e18d108 , 
    R_28d_1d9fb308 , 
    R_bcb_1e6b7c08 , 
    R_4fa_1dda3f68 , 
    R_2bb_1d9fcfc8 , 
    R_b3f_1e6b2488 , 
    R_a27_1e187528 , 
    R_362_1d9d3d88 , 
    R_497_1dd9fa08 , 
    R_64f_1dfb0d68 , 
    R_bd7_1e6b8388 , 
    R_b75_1e6b4648 , 
    R_98f_1e181628 , 
    R_6ed_1dfb7028 , 
    R_7d3_1e090048 , 
    R_b27_1e6b1588 , 
    R_39b_1d9d5c28 , 
    R_8cf_1e099dc8 , 
    R_689_1dfb31a8 , 
    R_7c6_1e08fd28 , 
    R_b2d_1e6b1948 , 
    R_92a_1e092f28 , 
    R_66c_1dfb1f88 , 
    R_956_1e6b00e8 , 
    R_b96_1e18ce88 , 
    R_bae_1e6b6ee8 , 
    R_94d_1e17ece8 , 
    R_785_1dfbcf28 , 
    R_6e2_1dfb6e48 , 
    R_65e_1dfb5cc8 , 
    R_42a_1d9dba88 , 
    R_7e8_1e090d68 , 
    R_b4d_1e6b2d48 , 
    R_bff_1e6b9c88 , 
    R_3c0_1d9d7348 , 
    R_44a_1d9dce88 , 
    R_2fe_1d9cff08 , 
    R_383_1d9d4d28 , 
    R_928_1e09d568 , 
    R_488_1dd9f0a8 , 
    R_5aa_1ddaaae8 , 
    R_3fd_1d9d9968 , 
    R_7d0_1e08fe68 , 
    R_7b4_1e08ece8 , 
    R_4d8_1dda22a8 , 
    R_418_1d9daa48 , 
    R_a43_1e1886a8 , 
    R_327_1d9d13a8 , 
    R_849_1e094a08 , 
    R_b5f_1e6b3888 , 
    R_4d3_1dda1f88 , 
    R_a97_1e18bb28 , 
    R_aba_1e18d608 , 
    R_ab1_1e18cb68 , 
    R_97f_1e180c28 , 
    R_788_1dfbd108 , 
    R_a1c_1e186e48 , 
    R_b11_1e6b07c8 , 
    R_a37_1e187f28 , 
    R_801_1e091d08 , 
    R_581_1dda8c48 , 
    R_49d_1dd9fdc8 , 
    R_56b_1dda7e88 , 
    R_4da_1dda3ce8 , 
    R_7f2_1e09d6a8 , 
    R_53d_1dda61c8 , 
    R_3df_1d9d86a8 , 
    R_429_1d9db4e8 , 
    R_8dc_1e09a5e8 , 
    R_a14_1e186948 , 
    R_9d6_1e186088 , 
    R_add_1e6ae748 , 
    R_b6d_1e6b4148 , 
    R_c1e_1e6b4e68 , 
    R_7fd_1e091a88 , 
    R_859_1e095408 , 
    R_b23_1e6b1308 , 
    R_afc_1e6afaa8 , 
    R_913_1e09c848 , 
    R_450_1d9dcd48 , 
    R_7cb_1e08fb48 , 
    R_b38_1e6b2028 , 
    R_a26_1e187988 , 
    R_74c_1dfbab88 , 
    R_35b_1d9d3428 , 
    R_962_1e17ff08 , 
    R_2e7_1d9ceba8 , 
    R_8c0_1e099468 , 
    R_8c7_1e0998c8 , 
    R_afe_1e6b5d68 , 
    R_977_1e180728 , 
    R_925_1e09d388 , 
    R_919_1e09cc08 , 
    R_728_1dfb9508 , 
    R_43a_1d9dc488 , 
    R_bf0_1e6b9328 , 
    R_9a3_1e1822a8 , 
    R_3af_1d9d68a8 , 
    R_930_1e09da68 , 
    R_90c_1e09c3e8 , 
    R_5a9_1ddaa548 , 
    R_659_1dfb13a8 , 
    R_c0f_1e6ba688 , 
    R_307_1d9cffa8 , 
    R_8bc_1e0991e8 , 
    R_2ed_1d9cef68 , 
    R_770_1dfbc208 , 
    R_34b_1d9d2a28 , 
    R_37f_1d9d4aa8 , 
    R_5f4_1ddad428 , 
    R_779_1dfbc7a8 , 
    R_46a_1dd9f468 , 
    R_be0_1e6b8928 , 
    R_bd3_1e6b8108 , 
    R_466_1d9d9c88 , 
    R_77e_1dfbcfc8 , 
    R_575_1dda84c8 , 
    R_4ff_1dda3b08 , 
    R_a18_1e186bc8 , 
    R_bda_1e6b8a68 , 
    R_31b_1d9d0c28 , 
    R_3c6_1d9d7c08 , 
    R_792_1dfbdc48 , 
    R_54b_1dda6a88 , 
    R_6bd_1dfb5228 , 
    R_b50_1e6b2f28 , 
    R_a61_1e189968 , 
    R_b8b_1e6b5408 , 
    R_b80_1e6b4d28 , 
    R_33c_1d9d20c8 , 
    R_3c3_1d9d7528 , 
    R_666_1dfb20c8 , 
    R_c2a_1e6bbc68 , 
    R_359_1d9d32e8 , 
    R_415_1d9da868 , 
    R_5da_1ddac8e8 , 
    R_577_1dda8608 , 
    R_637_1dfafe68 , 
    R_9f7_1e185728 , 
    R_570_1dda81a8 , 
    R_9f6_1e185b88 , 
    R_9f8_1e1857c8 , 
    R_a6e_1e18a688 , 
    R_73d_1dfba228 , 
    R_293_1d9fb6c8 , 
    R_884_1e096ee8 , 
    R_3a2_1d9d6588 , 
    R_9f9_1e185868 , 
    R_957_1e17f328 , 
    R_ab6_1e6b5fe8 , 
    R_760_1dfbb808 , 
    R_a21_1e187168 , 
    R_bb7_1e6b6f88 , 
    R_9eb_1e184fa8 , 
    R_a3f_1e188428 , 
    R_747_1dfba868 , 
    R_4bf_1dda1308 , 
    R_3d7_1d9d81a8 , 
    R_4a4_1dda0228 , 
    R_441_1d9dc3e8 , 
    R_7ce_1e090228 , 
    R_85a_1e0959a8 , 
    R_66f_1dfb2168 , 
    R_9ea_1e185408 , 
    R_9ec_1e185048 , 
    R_a3b_1e1881a8 , 
    R_ad4_1e6ae1a8 , 
    R_b94_1e6b59a8 , 
    R_467_1d9ddba8 , 
    R_96e_1e180688 , 
    R_323_1d9d1128 , 
    R_6ea_1dfb7348 , 
    R_6ca_1dfb5f48 , 
    R_9ed_1e1850e8 , 
    R_ae7_1e6aed88 , 
    R_830_1e093a68 , 
    R_6d9_1dfb63a8 , 
    R_8e6_1e08f0a8 , 
    R_6a1_1dfb40a8 , 
    R_710_1dfb8608 , 
    R_b41_1e6b25c8 , 
    R_732_1dfba048 , 
    R_6df_1dfb6768 , 
    R_a11_1e186768 , 
    R_a8f_1e18b628 , 
    R_b97_1e6b5b88 , 
    R_bc6_1e6b7de8 , 
    R_4db_1dda2488 , 
    R_9d7_1e184328 , 
    R_b29_1e6b16c8 , 
    R_57e_1dda8f68 , 
    R_29a_1d9fbb28 , 
    R_36f_1d9d40a8 , 
    R_3e4_1d9d89c8 , 
    R_7bc_1e08f1e8 , 
    R_87e_1e097028 , 
    R_b1c_1e6b0ea8 , 
    R_aab_1e18c7a8 , 
    R_96c_1e180048 , 
    R_551_1dda6e48 , 
    R_6d4_1dfb6088 , 
    R_2af_1d9fc848 , 
    R_479_1dd9e748 , 
    R_5a3_1ddaa188 , 
    R_672_1dfb2848 , 
    R_587_1dda9008 , 
    R_767_1dfbbc68 , 
    R_395_1d9d5868 , 
    R_3e9_1d9d8ce8 , 
    R_2f8_1d9cf648 , 
    R_64c_1dfb0b88 , 
    R_5e1_1ddac848 , 
    R_3fc_1d9d98c8 , 
    R_468_1d9ddc48 , 
    R_3ba_1d9d7488 , 
    R_55b_1dda7488 , 
    R_67e_1dfb2fc8 , 
    R_8b7_1e098ec8 , 
    R_879_1e096808 , 
    R_b5b_1e6b3608 , 
    R_a82_1e18b588 , 
    R_ae5_1e6aec48 , 
    R_84b_1e094b48 , 
    R_99e_1e182488 , 
    R_6dc_1dfb6588 , 
    R_3ad_1d9d6768 , 
    R_a59_1e189468 , 
    R_b62_1e6ba368 , 
    R_731_1dfb9aa8 , 
    R_3f1_1d9d91e8 , 
    R_620_1dfaf008 , 
    R_67d_1dfb2a28 , 
    R_adf_1e6ae888 , 
    R_349_1d9d28e8 , 
    R_3d1_1d9d7de8 , 
    R_3f4_1d9d93c8 , 
    R_80a_1e0927a8 , 
    R_350_1d9d2d48 , 
    R_a50_1e188ec8 , 
    R_bc1_1e6b75c8 , 
    R_b85_1e6b5048 , 
    R_5d7_1ddac208 , 
    R_7a2_1ddada68 , 
    R_539_1dda5f48 , 
    R_bbc_1e6b72a8 , 
    R_c14_1e6ba9a8 , 
    R_6c8_1dfb5908 , 
    R_4c8_1dda18a8 , 
    R_360_1d9d3748 , 
    R_2e2_1d9ced88 , 
    R_936_1e17e388 , 
    R_9f3_1e1854a8 , 
    R_b25_1e6b1448 , 
    R_b0a_1e6b0868 , 
    R_b56_1e6b87e8 , 
    R_bf4_1e6b95a8 , 
    R_95f_1e17f828 , 
    R_3b5_1d9d6c68 , 
    R_52a_1dda5fe8 , 
    R_9f2_1e185908 , 
    R_9f4_1e185548 , 
    R_686_1dfb34c8 , 
    R_2bc_1d9fd068 , 
    R_7a6_1e08e928 , 
    R_9ef_1e185228 , 
    R_b1e_1e6b78e8 , 
    R_bfb_1e6b9a08 , 
    R_378_1d9d4648 , 
    R_9ee_1e185688 , 
    R_9f0_1e1852c8 , 
    R_9f5_1e1855e8 , 
    R_4bd_1dda11c8 , 
    R_5af_1ddaa908 , 
    R_822_1e097f28 , 
    R_872_1e0968a8 , 
    R_9f1_1e185368 , 
    R_337_1d9d1da8 , 
    R_707_1dfb8068 , 
    R_755_1dfbb128 , 
    R_8f9_1e09b808 , 
    R_432_1d9dbf88 , 
    R_8af_1e0989c8 , 
    R_bc5_1e6b7848 , 
    R_934_1e09dce8 , 
    R_469_1d9ddce8 , 
    R_572_1dda87e8 , 
    R_863_1e095a48 , 
    R_958_1e17f3c8 , 
    R_742_1dfbaa48 , 
    R_2a5_1d9fc208 , 
    R_a9a_1e18c208 , 
    R_af9_1e6af8c8 , 
    R_9c1_1e183568 , 
    R_83c_1e0941e8 , 
    R_a81_1e18ad68 , 
    R_c19_1e6bacc8 , 
    R_91c_1e09cde8 , 
    R_4ac_1dda0728 , 
    R_bf8_1e6b9828 , 
    R_5be_1dda7168 , 
    R_93b_1e17e1a8 , 
    R_63c_1dfb0188 , 
    R_7e1_1e090908 , 
    R_7ba_1e08f5a8 , 
    R_6b2_1dfb5048 , 
    R_4dc_1dda2528 , 
    R_79e_1e08e428 , 
    R_492_1dd9fbe8 , 
    R_750_1dfbae08 , 
    R_9d8_1e1843c8 , 
    R_365_1d9d3a68 , 
    R_994_1e181948 , 
    R_95c_1e17f648 , 
    R_2ff_1d9cfaa8 , 
    R_89b_1e097d48 , 
    R_827_1e0934c8 , 
    R_332_1d9d1f88 , 
    R_9a7_1e182528 , 
    R_834_1e093ce8 , 
    R_30b_1d9d0228 , 
    R_86b_1e095f48 , 
    R_649_1dfb09a8 , 
    R_a1d_1e186ee8 , 
    R_b59_1e6b34c8 , 
    R_bb3_1e6b6d08 , 
    R_796_1e08e1a8 , 
    R_941_1e17e568 , 
    R_be9_1e6b8ec8 , 
    R_485_1dd9eec8 , 
    R_317_1d9d09a8 , 
    R_8a3_1e098248 , 
    R_49e_1dda0368 , 
    R_9c0_1e1834c8 , 
    R_32c_1d9d16c8 , 
    R_6d6_1dfb66c8 , 
    R_a15_1e1869e8 , 
    R_33e_1d9d2708 , 
    R_38c_1d9d52c8 , 
    R_75b_1dfbb4e8 , 
    R_ac4_1e18d748 , 
    R_5d9_1ddac348 , 
    R_546_1dda6c68 , 
    R_2be_1d9fd6a8 , 
    R_b76_1e6b4be8 , 
    R_975_1e1805e8 , 
    R_5c3_1ddab588 , 
    R_500_1dda3ba8 , 
    R_889_1e097208 , 
    R_988_1e1811c8 , 
    R_c2c_1e6bb8a8 , 
    R_b98_1e6b5c28 , 
    R_47d_1dd9e9c8 , 
    R_417_1d9da9a8 , 
    R_819_1e092c08 , 
    R_8f8_1e09b768 , 
    R_942_1e17eb08 , 
    R_ad1_1e6adfc8 , 
    R_8ce_1e09a228 , 
    R_563_1dda7988 , 
    R_2e8_1d9cec48 , 
    R_838_1e093f68 , 
    R_aee_1e187c08 , 
    R_641_1dfb04a8 , 
    R_c16_1e6b41e8 , 
    R_6c3_1dfb55e8 , 
    R_5f3_1ddad388 , 
    R_558_1dda72a8 , 
    R_821_1e093108 , 
    R_a5f_1e189828 , 
    R_3cd_1d9d7b68 , 
    R_80f_1e0925c8 , 
    R_724_1dfb9288 , 
    R_848_1e094968 , 
    R_9bf_1e183428 , 
    R_a19_1e186c68 , 
    R_baf_1e6b6a88 , 
    R_64a_1dfb0f48 , 
    R_aa8_1e18c5c8 , 
    R_6be_1dfb57c8 , 
    R_481_1dd9ec48 , 
    R_428_1d9db448 , 
    R_be6_1e6b91e8 , 
    R_44f_1d9dcca8 , 
    R_5b4_1ddaac28 , 
    R_629_1dfaf5a8 , 
    R_78f_1dfbd568 , 
    R_91f_1e09cfc8 , 
    R_858_1e095368 , 
    R_afb_1e6afa08 , 
    R_3fb_1d9d9828 , 
    R_922_1e091628 , 
    R_916_1e09cf28 , 
    R_8a1_1e098108 , 
    R_8db_1e09a548 , 
    R_b32_1e6b2168 , 
    R_411_1d9da5e8 , 
    R_6b0_1dfb4a08 , 
    R_5d1_1ddabe48 , 
    R_7df_1e0907c8 , 
    R_b04_1e6affa8 , 
    R_45a_1d9dd888 , 
    R_814_1e0928e8 , 
    R_665_1dfb1b28 , 
    R_69e_1dfb43c8 , 
    R_b42_1e6b2b68 , 
    R_555_1dda70c8 , 
    R_374_1d9d43c8 , 
    R_352_1d9d3388 , 
    R_2a6_1d9fc7a8 , 
    R_756_1dfbb6c8 , 
    R_bd6_1e6b3568 , 
    R_baa_1e18d888 , 
    R_5b9_1ddaaf48 , 
    R_3ec_1d9d8ec8;
wire n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , 
     n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , 
     n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , 
     n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , 
     n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , 
     n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , 
     n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , 
     n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , 
     n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , 
     n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , 
     n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , 
     n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , 
     n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , 
     n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , 
     n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , 
     n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , 
     n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , 
     n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , 
     n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , 
     n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , 
     n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , 
     n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , 
     n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , 
     n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , 
     n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , 
     n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , 
     n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , 
     n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , 
     n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , 
     n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , 
     n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , 
     n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , 
     n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , 
     n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , 
     n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , 
     n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , 
     n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , 
     n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , 
     n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , 
     n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , 
     n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , 
     n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , 
     n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , 
     n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , 
     n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , 
     n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , 
     n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , 
     n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , 
     n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , 
     n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , 
     n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , 
     n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , 
     n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , 
     n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , 
     n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , 
     n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , 
     n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , 
     n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , 
     n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , 
     n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , 
     n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , 
     n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , 
     n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , 
     n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , 
     n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , 
     n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , 
     n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , 
     n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , 
     n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , 
     n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , 
     n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , 
     n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , 
     n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , 
     n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , 
     n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , 
     n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , 
     n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , 
     n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , 
     n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , 
     n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , 
     n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , 
     n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , 
     n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , 
     n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , 
     n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , 
     n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , 
     n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , 
     n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , 
     n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , 
     n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , 
     n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , 
     n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , 
     n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , 
     n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , 
     n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , 
     n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , 
     n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , 
     n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , 
     n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , 
     n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , 
     n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , 
     n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , 
     n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , 
     n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , 
     n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , 
     n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , 
     n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , 
     n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , 
     n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , 
     n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , 
     n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , 
     n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , 
     n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , 
     n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , 
     n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , 
     n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , 
     n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , 
     n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , 
     n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , 
     n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , 
     n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , 
     n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , 
     n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , 
     n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , 
     n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , 
     n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , 
     n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , 
     n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , 
     n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , 
     n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , 
     n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , 
     n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , 
     n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , 
     n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , 
     n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , 
     n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , 
     n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , 
     n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , 
     n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , 
     n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , 
     n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , 
     n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , 
     n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , 
     n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , 
     n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , 
     n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , 
     n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , 
     n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , 
     n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , 
     n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , 
     n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , 
     n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , 
     n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , 
     n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , 
     n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , 
     n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , 
     n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , 
     n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , 
     n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , 
     n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , 
     n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , 
     n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , 
     n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , 
     n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , 
     n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , 
     n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , 
     n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , 
     n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , 
     n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , 
     n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , 
     n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , 
     n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , 
     n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , 
     n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , 
     n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , 
     n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , 
     n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , 
     n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , 
     n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , 
     n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , 
     n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , 
     n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , 
     n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , 
     n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , 
     n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , 
     n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , 
     n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , 
     n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , 
     n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , 
     n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , 
     n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , 
     n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , 
     n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , 
     n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , 
     n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , 
     n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , 
     n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , 
     n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , 
     n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , 
     n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , 
     n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , 
     n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , 
     n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , 
     n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , 
     n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , 
     n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , 
     n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , 
     n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , 
     n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , 
     n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , 
     n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , 
     n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , 
     n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , 
     n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , 
     n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , 
     n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , 
     n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , 
     n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , 
     n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , 
     n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , 
     n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , 
     n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , 
     n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , 
     n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , 
     n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , 
     n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , 
     n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , 
     n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , 
     n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , 
     n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , 
     n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , 
     n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , 
     n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , 
     n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , 
     n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , 
     n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , 
     n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , 
     n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , 
     n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , 
     n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , 
     n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , 
     n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , 
     n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , 
     n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , 
     n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , 
     n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , 
     n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , 
     n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , 
     n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , 
     n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , 
     n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , 
     n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , 
     n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , 
     n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , 
     n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , 
     n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , 
     n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , 
     n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , 
     n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , 
     n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , 
     n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , 
     n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , 
     n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , 
     n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , 
     n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , 
     n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , 
     n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , 
     n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , 
     n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , 
     n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , 
     n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , 
     n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , 
     n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , 
     n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , 
     n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , 
     n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , 
     n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , 
     n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , 
     n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , 
     n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , 
     n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , 
     n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , 
     n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , 
     n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , 
     n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , 
     n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , 
     n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , 
     n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , 
     n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , 
     n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , 
     n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , 
     n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , 
     n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , 
     n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , 
     n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , 
     n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , 
     n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , 
     n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , 
     n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , 
     n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , 
     n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , 
     n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , 
     n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , 
     n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , 
     n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , 
     n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , 
     n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , 
     n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , 
     n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , 
     n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , 
     n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , 
     n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , 
     n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , 
     n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , 
     n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , 
     n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , 
     n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , 
     n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , 
     n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , 
     n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , 
     n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , 
     n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , 
     n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , 
     n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , 
     n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , 
     n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , 
     n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , 
     n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , 
     n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , 
     n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , 
     n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , 
     n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , 
     n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , 
     n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , 
     n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , 
     n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , 
     n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , 
     n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , 
     n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , 
     n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , 
     n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , 
     n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , 
     n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , 
     n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , 
     n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , 
     n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , 
     n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , 
     n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , 
     n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , 
     n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , 
     n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , 
     n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , 
     n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , 
     n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , 
     n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , 
     n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , 
     n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , 
     n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , 
     n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , 
     n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , 
     n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , 
     n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , 
     n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , 
     n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , 
     n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , 
     n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , 
     n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , 
     n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , 
     n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , 
     n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , 
     n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , 
     n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , 
     n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , 
     n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , 
     n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , 
     n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , 
     n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , 
     n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , 
     n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , 
     n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , 
     n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , 
     n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , 
     n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , 
     n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , 
     n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , 
     n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , 
     n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , 
     n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , 
     n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , 
     n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , 
     n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , 
     n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , 
     n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , 
     n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , 
     n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , 
     n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , 
     n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , 
     n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , 
     n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , 
     n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , 
     n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , 
     n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , 
     n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , 
     n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , 
     n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , 
     n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , 
     n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , 
     n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , 
     n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , 
     n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , 
     n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , 
     n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , 
     n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , 
     n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , 
     n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , 
     n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , 
     n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , 
     n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , 
     n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , 
     n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , 
     n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , 
     n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , 
     n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , 
     n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , 
     n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , 
     n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , 
     n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , 
     n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , 
     n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , 
     n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , 
     n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , 
     n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , 
     n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , 
     n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , 
     n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , 
     n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , 
     n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , 
     n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , 
     n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , 
     n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , 
     n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , 
     n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , 
     n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , 
     n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , 
     n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , 
     n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , 
     n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , 
     n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , 
     n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , 
     n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , 
     n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , 
     n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , 
     n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , 
     n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , 
     n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , 
     n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , 
     n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , 
     n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , 
     n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , 
     n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , 
     n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , 
     n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , 
     n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , 
     n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , 
     n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , 
     n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , 
     n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , 
     n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , 
     n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , 
     n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , 
     n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , 
     n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , 
     n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , 
     n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , 
     n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , 
     n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , 
     n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , 
     n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , 
     n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , 
     n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , 
     n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , 
     n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , 
     n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , 
     n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , 
     n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , 
     n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , 
     n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , 
     n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , 
     n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , 
     n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , 
     n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , 
     n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , 
     n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , 
     n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , 
     n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , 
     n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , 
     n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , 
     n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , 
     n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , 
     n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , 
     n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , 
     n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , 
     n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , 
     n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , 
     n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , 
     n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , 
     n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , 
     n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , 
     n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , 
     n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , 
     n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , 
     n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , 
     n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , 
     n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , 
     n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , 
     n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , 
     n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , 
     n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , 
     n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , 
     n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , 
     n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , 
     n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , 
     n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , 
     n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , 
     n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , 
     n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , 
     n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , 
     n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , 
     n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , 
     n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , 
     n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , 
     n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , 
     n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , 
     n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , 
     n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , 
     n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , 
     n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , 
     n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , 
     n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , 
     n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , 
     n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , 
     n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , 
     n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , 
     n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , 
     n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , 
     n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , 
     n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , 
     n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , 
     n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , 
     n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , 
     n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , 
     n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , 
     n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , 
     n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , 
     n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , 
     n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , 
     n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , 
     n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , 
     n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , 
     n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , 
     n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , 
     n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , 
     n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , 
     n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , 
     n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , 
     n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , 
     n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , 
     n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , 
     n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , 
     n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , 
     n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , 
     n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , 
     n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , 
     n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , 
     n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , 
     n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , 
     n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , 
     n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , 
     n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , 
     n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , 
     n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , 
     n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , 
     n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , 
     n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , 
     n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , 
     n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , 
     n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , 
     n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , 
     n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , 
     n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , 
     n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , 
     n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , 
     n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , 
     n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , 
     n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , 
     n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , 
     n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , 
     n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , 
     n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , 
     n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , 
     n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , 
     n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , 
     n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , 
     n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , 
     n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , 
     n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , 
     n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , 
     n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , 
     n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , 
     n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , 
     n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , 
     n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , 
     n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , 
     n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , 
     n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , 
     n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , 
     n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , 
     n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , 
     n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , 
     n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , 
     n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , 
     n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , 
     n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , 
     n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , 
     n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , 
     n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , 
     n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , 
     n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , 
     n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , 
     n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , 
     n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , 
     n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , 
     n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , 
     n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , 
     n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , 
     n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , 
     n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , 
     n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , 
     n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , 
     n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , 
     n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , 
     n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , 
     n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , 
     n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , 
     n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , 
     n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , 
     n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , 
     n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , 
     n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , 
     n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , 
     n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , 
     n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , 
     n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , 
     n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , 
     n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , 
     n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , 
     n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , 
     n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , 
     n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , 
     n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , 
     n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , 
     n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , 
     n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , 
     n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , 
     n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , 
     n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , 
     n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , 
     n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , 
     n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , 
     n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , 
     n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , 
     n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , 
     n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , 
     n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , 
     n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , 
     n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , 
     n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , 
     n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , 
     n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , 
     n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , 
     n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , 
     n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , 
     n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , 
     n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , 
     n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , 
     n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , 
     n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , 
     n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , 
     n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , 
     n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , 
     n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , 
     n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , 
     n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , 
     n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , 
     n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , 
     n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , 
     n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , 
     n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , 
     n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , 
     n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , 
     n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , 
     n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , 
     n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , 
     n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , 
     n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , 
     n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , 
     n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , 
     n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , 
     n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , 
     n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , 
     n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , 
     n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , 
     n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , 
     n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , 
     n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , 
     n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , 
     n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , 
     n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , 
     n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , 
     n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , 
     n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , 
     n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , 
     n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , 
     n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , 
     n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , 
     n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , 
     n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , 
     n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , 
     n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , 
     n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , 
     n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , 
     n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , 
     n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , 
     n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , 
     n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , 
     n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , 
     n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , 
     n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , 
     n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , 
     n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , 
     n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , 
     n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , 
     n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , 
     n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , 
     n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , 
     n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , 
     n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , 
     n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , 
     n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , 
     n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , 
     n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , 
     n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , 
     n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , 
     n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , 
     n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , 
     n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , 
     n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , 
     n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , 
     n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , 
     n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , 
     n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , 
     n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , 
     n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , 
     n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , 
     n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , 
     n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , 
     n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , 
     n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , 
     n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , 
     n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , 
     n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , 
     n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , 
     n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , 
     n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , 
     n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , 
     n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , 
     n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , 
     n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , 
     n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , 
     n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , 
     n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , 
     n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , 
     n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , 
     n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , 
     n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , 
     n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , 
     n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , 
     n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , 
     n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , 
     n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , 
     n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , 
     n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , 
     n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , 
     n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , 
     n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , 
     n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , 
     n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , 
     n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , 
     n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , 
     n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , 
     n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , 
     n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , 
     n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , 
     n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , 
     n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , 
     n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , 
     n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , 
     n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , 
     n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , 
     n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , 
     n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , 
     n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , 
     n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , 
     n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , 
     n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , 
     n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , 
     n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , 
     n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , 
     n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , 
     n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , 
     n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , 
     n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , 
     n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , 
     n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , 
     n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , 
     n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , 
     n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , 
     n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , 
     n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , 
     n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , 
     n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , 
     n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , 
     n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , 
     n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , 
     n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , 
     n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , 
     n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , 
     n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , 
     n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , 
     n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , 
     n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , 
     n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , 
     n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , 
     n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , 
     n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , 
     n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , 
     n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , 
     n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , 
     n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , 
     n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , 
     n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , 
     n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , 
     n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , 
     n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , 
     n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , 
     n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , 
     n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , 
     n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , 
     n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , 
     n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , 
     n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , 
     n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , 
     n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , 
     n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , 
     n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , 
     n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , 
     n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , 
     n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , 
     n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , 
     n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , 
     n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , 
     n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , 
     n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , 
     n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , 
     n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , 
     n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , 
     n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , 
     n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , 
     n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , 
     n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , 
     n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , 
     n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , 
     n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , 
     n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , 
     n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , 
     n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , 
     n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , 
     n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , 
     n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , 
     n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , 
     n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , 
     n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , 
     n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , 
     n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , 
     n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , 
     n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , 
     n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , 
     n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , 
     n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , 
     n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , 
     n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , 
     n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , 
     n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , 
     n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , 
     n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , 
     n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , 
     n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , 
     n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , 
     n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , 
     n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , 
     n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , 
     n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , 
     n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , 
     n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , 
     n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , 
     n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , 
     n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , 
     n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , 
     n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , 
     n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , 
     n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , 
     n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , 
     n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , 
     n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , 
     n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , 
     n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , 
     n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , 
     n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , 
     n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , 
     n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , 
     n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , 
     n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , 
     n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , 
     n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , 
     n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , 
     n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , 
     n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , 
     n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , 
     n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , 
     n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , 
     n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , 
     n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , 
     n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , 
     n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , 
     n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , 
     n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , 
     n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , 
     n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , 
     n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , 
     n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , 
     n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , 
     n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , 
     n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , 
     n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , 
     n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , 
     n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , 
     n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , 
     n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , 
     n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , 
     n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , 
     n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , 
     n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , 
     n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , 
     n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , 
     n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , 
     n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , 
     n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , 
     n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , 
     n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , 
     n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , 
     n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , 
     n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , 
     n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , 
     n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , 
     n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , 
     n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , 
     n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , 
     n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , 
     n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , 
     n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , 
     n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , 
     n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , 
     n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , 
     n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , 
     n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , 
     n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , 
     n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , 
     n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , 
     n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , 
     n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , 
     n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , 
     n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , 
     n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , 
     n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , 
     n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , 
     n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , 
     n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , 
     n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , 
     n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , 
     n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , 
     n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , 
     n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , 
     n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , 
     n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , 
     n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , 
     n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , 
     n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , 
     n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , 
     n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , 
     n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , 
     n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , 
     n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , 
     n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , 
     n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , 
     n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , 
     n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , 
     n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , 
     n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , 
     n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , 
     n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , 
     n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , 
     n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , 
     n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , 
     n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , 
     n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , 
     n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , 
     n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , 
     n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , 
     n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , 
     n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , 
     n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , 
     n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , 
     n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , 
     n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , 
     n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , 
     n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , 
     n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , 
     n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , 
     n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , 
     n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , 
     n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , 
     n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , 
     n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , 
     n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , 
     n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , 
     n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , 
     n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , 
     n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , 
     n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , 
     n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , 
     n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , 
     n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , 
     n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , 
     n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , 
     n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , 
     n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , 
     n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , 
     n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , 
     n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , 
     n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , 
     n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , 
     n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , 
     n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , 
     n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , 
     n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , 
     n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , 
     n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , 
     n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , 
     n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , 
     n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , 
     n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , 
     n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , 
     n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , 
     n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , 
     n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , 
     n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , 
     n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , 
     n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , 
     n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , 
     n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , 
     n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , 
     n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , 
     n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , 
     n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , 
     n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , 
     n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , 
     n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , 
     n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , 
     n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , 
     n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , 
     n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , 
     n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , 
     n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , 
     n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , 
     n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , 
     n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , 
     n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , 
     n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , 
     n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , 
     n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , 
     n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , 
     n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , 
     n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , 
     n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , 
     n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , 
     n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , 
     n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , 
     n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , 
     n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , 
     n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , 
     n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , 
     n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , 
     n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , 
     n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , 
     n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , 
     n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , 
     n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , 
     n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , 
     n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , 
     n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , 
     n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , 
     n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , 
     n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , 
     n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , 
     n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , 
     n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , 
     n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , 
     n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , 
     n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , 
     n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , 
     n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , 
     n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , 
     n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , 
     n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , 
     n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , 
     n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , 
     n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , 
     n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , 
     n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , 
     n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , 
     n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , 
     n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , 
     n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , 
     n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , 
     n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , 
     n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , 
     n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , 
     n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , 
     n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , 
     n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , 
     n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , 
     n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , 
     n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , 
     n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , 
     n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , 
     n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , 
     n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , 
     n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , 
     n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , 
     n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , 
     n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , 
     n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , 
     n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , 
     n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , 
     n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , 
     n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , 
     n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , 
     n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , 
     n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , 
     n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , 
     n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , 
     n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , 
     n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , 
     n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , 
     n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , 
     n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , 
     n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , 
     n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , 
     n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , 
     n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , 
     n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , 
     n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , 
     n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , 
     n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , 
     n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , 
     n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , 
     n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , 
     n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , 
     n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , 
     n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , 
     n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , 
     n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , 
     n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , 
     n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , 
     n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , 
     n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , 
     n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , 
     n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , 
     n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , 
     n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , 
     n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , 
     n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , 
     n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , 
     n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , 
     n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , 
     n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , 
     n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , 
     n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , 
     n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , 
     n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , 
     n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , 
     n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , 
     n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , 
     n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , 
     n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , 
     n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , 
     n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , 
     n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , 
     n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , 
     n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , 
     n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , 
     n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , 
     n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , 
     n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , 
     n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , 
     n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , 
     n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , 
     n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , 
     n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , 
     n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , 
     n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , 
     n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , 
     n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , 
     n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , 
     n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , 
     n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , 
     n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , 
     n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , 
     n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , 
     n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , 
     n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , 
     n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , 
     n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , 
     n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , 
     n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , 
     n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , 
     n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , 
     n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , 
     n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , 
     n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , 
     n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , 
     n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , 
     n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , 
     n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , 
     n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , 
     n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , 
     n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , 
     n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , 
     n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , 
     n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , 
     n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , 
     n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , 
     n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , 
     n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , 
     n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , 
     n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , 
     n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , 
     n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , 
     n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , 
     n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , 
     n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , 
     n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , 
     n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , 
     n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , 
     n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , 
     n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , 
     n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , 
     n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , 
     n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , 
     n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , 
     n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , 
     n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , 
     n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , 
     n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , 
     n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , 
     n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , 
     n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , 
     n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , 
     n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , 
     n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , 
     n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , 
     n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , 
     n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , 
     n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , 
     n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , 
     n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , 
     n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , 
     n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , 
     n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , 
     n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , 
     n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , 
     n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , 
     n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , 
     n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , 
     n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , 
     n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , 
     n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , 
     n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , 
     n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , 
     n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , 
     n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , 
     n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , 
     n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , 
     n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , 
     n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , 
     n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , 
     n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , 
     n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , 
     n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , 
     n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , 
     n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , 
     n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , 
     n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , 
     n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , 
     n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , 
     n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , 
     n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , 
     n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , 
     n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , 
     n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , 
     n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , 
     n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , 
     n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , 
     n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , 
     n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , 
     n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , 
     n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , 
     n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , 
     n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , 
     n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , 
     n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , 
     n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , 
     n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , 
     n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , 
     n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , 
     n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , 
     n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , 
     n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , 
     n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , 
     n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , 
     n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , 
     n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , 
     n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , 
     n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , 
     n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , 
     n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , 
     n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , 
     n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , 
     n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , 
     n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , 
     n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , 
     n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , 
     n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , 
     n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , 
     n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , 
     n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , 
     n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , 
     n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , 
     n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , 
     n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , 
     n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , 
     n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , 
     n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , 
     n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , 
     n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , 
     n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , 
     n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , 
     n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , 
     n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , 
     n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , 
     n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , 
     n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , 
     n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , 
     n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , 
     n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , 
     n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , 
     n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , 
     n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , 
     n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , 
     n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , 
     n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , 
     n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , 
     n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , 
     n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , 
     n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , 
     n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , 
     n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , 
     n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , 
     n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , 
     n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , 
     n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , 
     n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , 
     n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , 
     n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , 
     n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , 
     n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , 
     n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , 
     n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , 
     n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , 
     n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , 
     n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , 
     n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , 
     n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , 
     n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , 
     n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , 
     n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , 
     n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , 
     n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , 
     n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , 
     n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , 
     n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , 
     n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , 
     n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , 
     n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , 
     n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , 
     n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , 
     n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , 
     n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , 
     n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , 
     n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , 
     n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , 
     n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , 
     n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , 
     n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , 
     n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , 
     n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , 
     n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , 
     n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , 
     n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , 
     n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , 
     n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , 
     n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , 
     n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , 
     n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , 
     n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , 
     n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , 
     n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , 
     n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , 
     n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , 
     n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , 
     n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , 
     n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , 
     n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , 
     n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , 
     n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , 
     n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , 
     n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , 
     n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , 
     n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , 
     n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , 
     n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , 
     n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , 
     n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , 
     n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , 
     n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , 
     n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , 
     n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , 
     n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , 
     n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , 
     n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , 
     n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , 
     n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , 
     n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , 
     n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , 
     n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , 
     n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , 
     n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , 
     n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , 
     n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , 
     n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , 
     n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , 
     n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , 
     n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , 
     n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , 
     n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , 
     n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , 
     n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , 
     n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , 
     n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , 
     n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , 
     n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , 
     n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , 
     n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , 
     n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , 
     n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , 
     n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , 
     n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , 
     n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , 
     n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , 
     n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , 
     n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , 
     n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , 
     n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , 
     n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , 
     n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , 
     n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , 
     n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , 
     n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , 
     n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , 
     n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , 
     n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , 
     n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , 
     n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , 
     n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , 
     n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , 
     n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , 
     n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , 
     n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , 
     n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , 
     n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , 
     n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , 
     n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , 
     n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , 
     n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , 
     n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , 
     n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , 
     n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , 
     n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , 
     n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , 
     n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , 
     n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , 
     n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , 
     n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , 
     n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , 
     n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , 
     n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , 
     n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , 
     n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , 
     n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , 
     n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , 
     n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , 
     n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , 
     n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , 
     n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , 
     n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , 
     n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , 
     n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , 
     n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , 
     n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , 
     n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , 
     n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , 
     n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , 
     n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , 
     n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , 
     n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , 
     n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , 
     n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , 
     n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , 
     n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , 
     n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , 
     n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , 
     n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , 
     n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , 
     n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , 
     n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , 
     n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , 
     n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , 
     n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , 
     n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , 
     n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , 
     n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , 
     n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , 
     n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , 
     n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , 
     n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , 
     n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , 
     n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , 
     n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , 
     n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , 
     n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , 
     n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , 
     n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , 
     n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , 
     n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , 
     n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , 
     n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , 
     n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , 
     n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , 
     n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , 
     n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , 
     n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , 
     n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , 
     n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , 
     n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , 
     n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , 
     n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , 
     n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , 
     n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , 
     n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , 
     n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , 
     n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , 
     n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , 
     n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , 
     n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , 
     n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , 
     n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , 
     n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , 
     n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , 
     n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , 
     n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , 
     n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , 
     n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , 
     n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , 
     n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , 
     n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , 
     n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , 
     n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , 
     n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , 
     n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , 
     n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , 
     n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , 
     n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , 
     n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , 
     n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , 
     n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , 
     n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , 
     n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , 
     n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , 
     n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , 
     n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , 
     n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , 
     n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , 
     n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , 
     n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , 
     n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , 
     n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , 
     n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , 
     n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , 
     n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , 
     n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , 
     n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , 
     n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , 
     n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , 
     n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , 
     n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , 
     n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , 
     n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , 
     n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , 
     n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , 
     n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , 
     n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , 
     n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , 
     n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , 
     n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , 
     n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , 
     n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , 
     n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , 
     n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , 
     n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , 
     n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , 
     n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , 
     n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , 
     n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , 
     n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , 
     n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , 
     n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , 
     n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , 
     n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , 
     n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , 
     n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , 
     n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , 
     n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , 
     n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , 
     n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , 
     n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , 
     n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , 
     n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , 
     n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , 
     n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , 
     n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , 
     n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , 
     n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , 
     n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , 
     n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , 
     n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , 
     n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , 
     n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , 
     n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , 
     n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , 
     n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , 
     n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , 
     n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , 
     n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , 
     n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , 
     n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , 
     n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , 
     n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , 
     n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , 
     n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , 
     n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , 
     n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , 
     n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , 
     n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , 
     n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , 
     n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , 
     n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , 
     n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , 
     n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , 
     n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , 
     n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , 
     n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , 
     n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , 
     n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , 
     n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , 
     n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , 
     n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , 
     n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , 
     n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , 
     n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , 
     n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , 
     n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , 
     n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , 
     n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , 
     n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , 
     n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , 
     n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , 
     n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , 
     n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , 
     n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , 
     n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , 
     n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , 
     n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , 
     n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , 
     n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , 
     n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , 
     n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , 
     n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , 
     n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , 
     n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , 
     n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , 
     n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , 
     n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , 
     n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , 
     n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , 
     n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , 
     n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , 
     n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , 
     n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , 
     n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , 
     n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , 
     n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , 
     n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , 
     n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , 
     n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , 
     n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , 
     n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , 
     n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , 
     n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , 
     n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , 
     n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , 
     n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , 
     n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , 
     n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , 
     n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , 
     n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , 
     n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , 
     n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , 
     n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , 
     n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , 
     n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , 
     n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , 
     n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , 
     n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , 
     n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , 
     n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , 
     n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , 
     n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , 
     n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , 
     n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , 
     n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , 
     n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , 
     n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , 
     n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , 
     n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , 
     n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , 
     n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , 
     n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , 
     n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , 
     n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , 
     n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , 
     n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , 
     n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , 
     n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , 
     n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , 
     n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , 
     n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , 
     n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , 
     n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , 
     n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , 
     n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , 
     n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , 
     n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , 
     n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , 
     n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , 
     n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , 
     n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , 
     n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , 
     n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , 
     n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , 
     n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , 
     n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , 
     n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , 
     n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , 
     n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , 
     n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , 
     n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , 
     n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , 
     n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , 
     n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , 
     n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , 
     n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , 
     n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , 
     n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , 
     n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , 
     n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , 
     n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , 
     n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , 
     n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , 
     n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , 
     n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , 
     n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , 
     n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , 
     n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , 
     n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , 
     n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , 
     n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , 
     n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , 
     n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , 
     n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , 
     n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , 
     n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , 
     n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , 
     n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , 
     n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , 
     n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , 
     n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , 
     n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , 
     n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , 
     n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , 
     n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , 
     n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , 
     n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , 
     n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , 
     n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , 
     n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , 
     n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , 
     n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , 
     n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , 
     n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , 
     n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , 
     n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , 
     n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , 
     n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , 
     n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , 
     n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , 
     n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , 
     n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , 
     n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , 
     n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , 
     n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , 
     n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , 
     n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , 
     n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , 
     n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , 
     n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , 
     n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , 
     n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , 
     n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , 
     n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , 
     n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , 
     n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , 
     n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , 
     n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , 
     n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , 
     n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , 
     n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , 
     n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , 
     n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , 
     n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , 
     n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , 
     n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , 
     n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , 
     n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , 
     n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , 
     n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , 
     n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , 
     n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , 
     n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , 
     n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , 
     n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , 
     n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , 
     n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , 
     n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , 
     n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , 
     n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , 
     n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , 
     n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , 
     n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , 
     n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , 
     n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , 
     n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , 
     n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , 
     n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , 
     n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , 
     n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , 
     n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , 
     n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , 
     n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , 
     n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , 
     n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , 
     n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , 
     n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , 
     n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , 
     n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , 
     n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , 
     n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , 
     n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , 
     n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , 
     n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , 
     n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , 
     n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , 
     n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , 
     n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , 
     n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , 
     n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , 
     n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , 
     n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , 
     n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , 
     n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , 
     n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , 
     n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , 
     n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , 
     n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , 
     n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , 
     n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , 
     n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , 
     n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , 
     n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , 
     n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , 
     n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , 
     n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , 
     n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , 
     n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , 
     n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , 
     n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , 
     n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , 
     n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , 
     n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , 
     n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , 
     n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , 
     n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , 
     n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , 
     n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , 
     n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , 
     n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , 
     n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , 
     n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , 
     n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , 
     n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , 
     n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , 
     n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , 
     n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , 
     n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , 
     n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , 
     n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , 
     n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , 
     n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , 
     n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , 
     n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , 
     n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , 
     n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , 
     n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , 
     n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , 
     n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , 
     n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , 
     n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , 
     n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , 
     n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , 
     n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , 
     n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , 
     n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , 
     n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , 
     n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , 
     n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , 
     n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , 
     n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , 
     n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , 
     n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , 
     n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , 
     n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , 
     n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , 
     n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , 
     n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , 
     n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , 
     n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , 
     n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , 
     n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , 
     n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , 
     n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , 
     n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , 
     n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , 
     n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , 
     n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , 
     n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , 
     n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , 
     n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , 
     n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , 
     n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , 
     n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , 
     n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , 
     n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , 
     n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , 
     n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , 
     n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , 
     n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , 
     n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , 
     n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , 
     n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , 
     n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , 
     n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , 
     n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , 
     n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , 
     n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , 
     n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , 
     n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , 
     n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , 
     n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , 
     n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , 
     n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , 
     n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , 
     n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , 
     n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , 
     n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , 
     n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , 
     n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , 
     n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , 
     n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , 
     n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , 
     n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , 
     n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , 
     n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , 
     n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , 
     n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , 
     n26777 , n26778 , n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , 
     n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , 
     n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , 
     n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , 
     n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , 
     n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , 
     n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , 
     n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , 
     n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , 
     n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , 
     n26877 , n26878 , n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , 
     n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , 
     n26897 , n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , 
     n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , 
     n26917 , n26918 , n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , 
     n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , 
     n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , 
     n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , 
     n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , 
     n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , 
     n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , 
     n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , 
     n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , 
     n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , 
     n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , 
     n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , 
     n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , 
     n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , 
     n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , 
     n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , 
     n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , 
     n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , 
     n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , 
     n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , 
     n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , 
     n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , 
     n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , 
     n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , 
     n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , 
     n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , 
     n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , 
     n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , 
     n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , 
     n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , 
     n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , 
     n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , 
     n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , 
     n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , 
     n27257 , n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , 
     n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , 
     n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , 
     n27287 , n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , 
     n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , 
     n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , 
     n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , 
     n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , 
     n27337 , n27338 , n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , 
     n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , 
     n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , 
     n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , 
     n27377 , n27378 , n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , 
     n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , 
     n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , 
     n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , 
     n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , 
     n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , 
     n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , 
     n27447 , n27448 , n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , 
     n27457 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , 
     n27467 , n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , 
     n27477 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , 
     n27487 , n27488 , n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , 
     n27497 , n27498 , n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , 
     n27507 , n27508 , n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , 
     n27517 , n27518 , n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , 
     n27527 , n27528 , n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , 
     n27537 , n27538 , n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , 
     n27547 , n27548 , n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , 
     n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , 
     n27567 , n27568 , n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , 
     n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , 
     n27587 , n27588 , n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , 
     n27597 , n27598 , n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , 
     n27607 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , 
     n27617 , n27618 , n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , 
     n27627 , n27628 , n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , 
     n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , 
     n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , 
     n27657 , n27658 , n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , 
     n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , 
     n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , 
     n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , 
     n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , 
     n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , 
     n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , 
     n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , 
     n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , 
     n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , 
     n27757 , n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , 
     n27767 , n27768 , n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , 
     n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , 
     n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , 
     n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , 
     n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , 
     n27817 , n27818 , n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , 
     n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , 
     n27837 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , 
     n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , 
     n27857 , n27858 , n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , 
     n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , 
     n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , 
     n27887 , n27888 , n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , 
     n27897 , n27898 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , 
     n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , 
     n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , 
     n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , 
     n27937 , n27938 , n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , 
     n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , 
     n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , 
     n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , 
     n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , 
     n27987 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , 
     n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , 
     n28007 , n28008 , n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , 
     n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , 
     n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , 
     n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , 
     n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , 
     n28057 , n28058 , n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , 
     n28067 , n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , 
     n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , 
     n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , 
     n28097 , n28098 , n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , 
     n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , 
     n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , 
     n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , 
     n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , 
     n28147 , n28148 , n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , 
     n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , 
     n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , 
     n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , 
     n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , 
     n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , 
     n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , 
     n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , 
     n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , 
     n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , 
     n28247 , n28248 , n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , 
     n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , 
     n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , 
     n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , 
     n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , 
     n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , 
     n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , 
     n28317 , n28318 , n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , 
     n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , 
     n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , 
     n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , 
     n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , 
     n28367 , n28368 , n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , 
     n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , 
     n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , 
     n28397 , n28398 , n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , 
     n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , 
     n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , 
     n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , 
     n28437 , n28438 , n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , 
     n28447 , n28448 , n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , 
     n28457 , n28458 , n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , 
     n28467 , n28468 , n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , n28475 , n28476 , 
     n28477 , n28478 , n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , 
     n28487 , n28488 , n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , n28495 , n28496 , 
     n28497 , n28498 , n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , 
     n28507 , n28508 , n28509 , n28510 , n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , 
     n28517 , n28518 , n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , 
     n28527 , n28528 , n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , 
     n28537 , n28538 , n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , n28545 , n28546 , 
     n28547 , n28548 , n28549 , n28550 , n28551 , n28552 , n28553 , n28554 , n28555 , n28556 , 
     n28557 , n28558 , n28559 , n28560 , n28561 , n28562 , n28563 , n28564 , n28565 , n28566 , 
     n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , n28575 , n28576 , 
     n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , n28585 , n28586 , 
     n28587 , n28588 , n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , n28595 , n28596 , 
     n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , n28605 , n28606 , 
     n28607 , n28608 , n28609 , n28610 , n28611 , n28612 , n28613 , n28614 , n28615 , n28616 , 
     n28617 , n28618 , n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , 
     n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , n28635 , n28636 , 
     n28637 , n28638 , n28639 , n28640 , n28641 , n28642 , n28643 , n28644 , n28645 , n28646 , 
     n28647 , n28648 , n28649 , n28650 , n28651 , n28652 , n28653 , n28654 , n28655 , n28656 , 
     n28657 , n28658 , n28659 , n28660 , n28661 , n28662 , n28663 , n28664 , n28665 , n28666 , 
     n28667 , n28668 , n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , n28675 , n28676 , 
     n28677 , n28678 , n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , n28685 , n28686 , 
     n28687 , n28688 , n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , n28695 , n28696 , 
     n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , n28705 , n28706 , 
     n28707 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , n28715 , n28716 , 
     n28717 , n28718 , n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , n28725 , n28726 , 
     n28727 , n28728 , n28729 , n28730 , n28731 , n28732 , n28733 , n28734 , n28735 , n28736 , 
     n28737 , n28738 , n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , n28745 , n28746 , 
     n28747 , n28748 , n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , n28755 , n28756 , 
     n28757 , n28758 , n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , 
     n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , 
     n28777 , n28778 , n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , n28785 , n28786 , 
     n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , 
     n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , 
     n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , 
     n28817 , n28818 , n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , 
     n28827 , n28828 , n28829 , n28830 , n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , 
     n28837 , n28838 , n28839 , n28840 , n28841 , n28842 , n28843 , n28844 , n28845 , n28846 , 
     n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , n28855 , n28856 , 
     n28857 , n28858 , n28859 , n28860 , n28861 , n28862 , n28863 , n28864 , n28865 , n28866 , 
     n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , n28875 , n28876 , 
     n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , n28885 , n28886 , 
     n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , n28895 , n28896 , 
     n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , n28905 , n28906 , 
     n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , n28915 , n28916 , 
     n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , n28925 , n28926 , 
     n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , n28935 , n28936 , 
     n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , n28945 , n28946 , 
     n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , n28955 , n28956 , 
     n28957 , n28958 , n28959 , n28960 , n28961 , n28962 , n28963 , n28964 , n28965 , n28966 , 
     n28967 , n28968 , n28969 , n28970 , n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , 
     n28977 , n28978 , n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , n28985 , n28986 , 
     n28987 , n28988 , n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , n28995 , n28996 , 
     n28997 , n28998 , n28999 , n29000 , n29001 , n29002 , n29003 , n29004 , n29005 , n29006 , 
     n29007 , n29008 , n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , n29015 , n29016 , 
     n29017 , n29018 , n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , n29025 , n29026 , 
     n29027 , n29028 , n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , n29035 , n29036 , 
     n29037 , n29038 , n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , n29045 , n29046 , 
     n29047 , n29048 , n29049 , n29050 , n29051 , n29052 , n29053 , n29054 , n29055 , n29056 , 
     n29057 , n29058 , n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , n29065 , n29066 , 
     n29067 , n29068 , n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , 
     n29077 , n29078 , n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , 
     n29087 , n29088 , n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , n29095 , n29096 , 
     n29097 , n29098 , n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , n29105 , n29106 , 
     n29107 , n29108 , n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , n29115 , n29116 , 
     n29117 , n29118 , n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , 
     n29127 , n29128 , n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , n29135 , n29136 , 
     n29137 , n29138 , n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , 
     n29147 , n29148 , n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , n29155 , n29156 , 
     n29157 , n29158 , n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , 
     n29167 , n29168 , n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , 
     n29177 , n29178 , n29179 , n29180 , n29181 , n29182 , n29183 , n29184 , n29185 , n29186 , 
     n29187 , n29188 , n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , n29195 , n29196 , 
     n29197 , n29198 , n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , n29205 , n29206 , 
     n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , n29215 , n29216 , 
     n29217 , n29218 , n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , n29225 , n29226 , 
     n29227 , n29228 , n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , n29235 , n29236 , 
     n29237 , n29238 , n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , n29245 , n29246 , 
     n29247 , n29248 , n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , n29255 , n29256 , 
     n29257 , n29258 , n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , n29265 , n29266 , 
     n29267 , n29268 , n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , 
     n29277 , n29278 , n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , 
     n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , n29295 , n29296 , 
     n29297 , n29298 , n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , n29305 , n29306 , 
     n29307 , n29308 , n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , n29315 , n29316 , 
     n29317 , n29318 , n29319 , n29320 , n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , 
     n29327 , n29328 , n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , 
     n29337 , n29338 , n29339 , n29340 , n29341 , n29342 , n29343 , n29344 , n29345 , n29346 , 
     n29347 , n29348 , n29349 , n29350 , n29351 , n29352 , n29353 , n29354 , n29355 , n29356 , 
     n29357 , n29358 , n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , n29365 , n29366 , 
     n29367 , n29368 , n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , n29375 , n29376 , 
     n29377 , n29378 , n29379 , n29380 , n29381 , n29382 , n29383 , n29384 , n29385 , n29386 , 
     n29387 , n29388 , n29389 , n29390 , n29391 , n29392 , n29393 , n29394 , n29395 , n29396 , 
     n29397 , n29398 , n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , n29405 , n29406 , 
     n29407 , n29408 , n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , n29415 , n29416 , 
     n29417 , n29418 , n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , 
     n29427 , n29428 , n29429 , n29430 , n29431 , n29432 , n29433 , n29434 , n29435 , n29436 , 
     n29437 , n29438 , n29439 , n29440 , n29441 , n29442 , n29443 , n29444 , n29445 , n29446 , 
     n29447 , n29448 , n29449 , n29450 , n29451 , n29452 , n29453 , n29454 , n29455 , n29456 , 
     n29457 , n29458 , n29459 , n29460 , n29461 , n29462 , n29463 , n29464 , n29465 , n29466 , 
     n29467 , n29468 , n29469 , n29470 , n29471 , n29472 , n29473 , n29474 , n29475 , n29476 , 
     n29477 , n29478 , n29479 , n29480 , n29481 , n29482 , n29483 , n29484 , n29485 , n29486 , 
     n29487 , n29488 , n29489 , n29490 , n29491 , n29492 , n29493 , n29494 , n29495 , n29496 , 
     n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , n29505 , n29506 , 
     n29507 , n29508 , n29509 , n29510 , n29511 , n29512 , n29513 , n29514 , n29515 , n29516 , 
     n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , n29523 , n29524 , n29525 , n29526 , 
     n29527 , n29528 , n29529 , n29530 , n29531 , n29532 , n29533 , n29534 , n29535 , n29536 , 
     n29537 , n29538 , n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , n29545 , n29546 , 
     n29547 , n29548 , n29549 , n29550 , n29551 , n29552 , n29553 , n29554 , n29555 , n29556 , 
     n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , n29563 , n29564 , n29565 , n29566 , 
     n29567 , n29568 , n29569 , n29570 , n29571 , n29572 , n29573 , n29574 , n29575 , n29576 , 
     n29577 , n29578 , n29579 , n29580 , n29581 , n29582 , n29583 , n29584 , n29585 , n29586 , 
     n29587 , n29588 , n29589 , n29590 , n29591 , n29592 , n29593 , n29594 , n29595 , n29596 , 
     n29597 , n29598 , n29599 , n29600 , n29601 , n29602 , n29603 , n29604 , n29605 , n29606 , 
     n29607 , n29608 , n29609 , n29610 , n29611 , n29612 , n29613 , n29614 , n29615 , n29616 , 
     n29617 , n29618 , n29619 , n29620 , n29621 , n29622 , n29623 , n29624 , n29625 , n29626 , 
     n29627 , n29628 , n29629 , n29630 , n29631 , n29632 , n29633 , n29634 , n29635 , n29636 , 
     n29637 , n29638 , n29639 , n29640 , n29641 , n29642 , n29643 , n29644 , n29645 , n29646 , 
     n29647 , n29648 , n29649 , n29650 , n29651 , n29652 , n29653 , n29654 , n29655 , n29656 , 
     n29657 , n29658 , n29659 , n29660 , n29661 , n29662 , n29663 , n29664 , n29665 , n29666 , 
     n29667 , n29668 , n29669 , n29670 , n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , 
     n29677 , n29678 , n29679 , n29680 , n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , 
     n29687 , n29688 , n29689 , n29690 , n29691 , n29692 , n29693 , n29694 , n29695 , n29696 , 
     n29697 , n29698 , n29699 , n29700 , n29701 , n29702 , n29703 , n29704 , n29705 , n29706 , 
     n29707 , n29708 , n29709 , n29710 , n29711 , n29712 , n29713 , n29714 , n29715 , n29716 , 
     n29717 , n29718 , n29719 , n29720 , n29721 , n29722 , n29723 , n29724 , n29725 , n29726 , 
     n29727 , n29728 , n29729 , n29730 , n29731 , n29732 , n29733 , n29734 , n29735 , n29736 , 
     n29737 , n29738 , n29739 , n29740 , n29741 , n29742 , n29743 , n29744 , n29745 , n29746 , 
     n29747 , n29748 , n29749 , n29750 , n29751 , n29752 , n29753 , n29754 , n29755 , n29756 , 
     n29757 , n29758 , n29759 , n29760 , n29761 , n29762 , n29763 , n29764 , n29765 , n29766 , 
     n29767 , n29768 , n29769 , n29770 , n29771 , n29772 , n29773 , n29774 , n29775 , n29776 , 
     n29777 , n29778 , n29779 , n29780 , n29781 , n29782 , n29783 , n29784 , n29785 , n29786 , 
     n29787 , n29788 , n29789 , n29790 , n29791 , n29792 , n29793 , n29794 , n29795 , n29796 , 
     n29797 , n29798 , n29799 , n29800 , n29801 , n29802 , n29803 , n29804 , n29805 , n29806 , 
     n29807 , n29808 , n29809 , n29810 , n29811 , n29812 , n29813 , n29814 , n29815 , n29816 , 
     n29817 , n29818 , n29819 , n29820 , n29821 , n29822 , n29823 , n29824 , n29825 , n29826 , 
     n29827 , n29828 , n29829 , n29830 , n29831 , n29832 , n29833 , n29834 , n29835 , n29836 , 
     n29837 , n29838 , n29839 , n29840 , n29841 , n29842 , n29843 , n29844 , n29845 , n29846 , 
     n29847 , n29848 , n29849 , n29850 , n29851 , n29852 , n29853 , n29854 , n29855 , n29856 , 
     n29857 , n29858 , n29859 , n29860 , n29861 , n29862 , n29863 , n29864 , n29865 , n29866 , 
     n29867 , n29868 , n29869 , n29870 , n29871 , n29872 , n29873 , n29874 , n29875 , n29876 , 
     n29877 , n29878 , n29879 , n29880 , n29881 , n29882 , n29883 , n29884 , n29885 , n29886 , 
     n29887 , n29888 , n29889 , n29890 , n29891 , n29892 , n29893 , n29894 , n29895 , n29896 , 
     n29897 , n29898 , n29899 , n29900 , n29901 , n29902 , n29903 , n29904 , n29905 , n29906 , 
     n29907 , n29908 , n29909 , n29910 , n29911 , n29912 , n29913 , n29914 , n29915 , n29916 , 
     n29917 , n29918 , n29919 , n29920 , n29921 , n29922 , n29923 , n29924 , n29925 , n29926 , 
     n29927 , n29928 , n29929 , n29930 , n29931 , n29932 , n29933 , n29934 , n29935 , n29936 , 
     n29937 , n29938 , n29939 , n29940 , n29941 , n29942 , n29943 , n29944 , n29945 , n29946 , 
     n29947 , n29948 , n29949 , n29950 , n29951 , n29952 , n29953 , n29954 , n29955 , n29956 , 
     n29957 , n29958 , n29959 , n29960 , n29961 , n29962 , n29963 , n29964 , n29965 , n29966 , 
     n29967 , n29968 , n29969 , n29970 , n29971 , n29972 , n29973 , n29974 , n29975 , n29976 , 
     n29977 , n29978 , n29979 , n29980 , n29981 , n29982 , n29983 , n29984 , n29985 , n29986 , 
     n29987 , n29988 , n29989 , n29990 , n29991 , n29992 , n29993 , n29994 , n29995 , n29996 , 
     n29997 , n29998 , n29999 , n30000 , n30001 , n30002 , n30003 , n30004 , n30005 , n30006 , 
     n30007 , n30008 , n30009 , n30010 , n30011 , n30012 , n30013 , n30014 , n30015 , n30016 , 
     n30017 , n30018 , n30019 , n30020 , n30021 , n30022 , n30023 , n30024 , n30025 , n30026 , 
     n30027 , n30028 , n30029 , n30030 , n30031 , n30032 , n30033 , n30034 , n30035 , n30036 , 
     n30037 , n30038 , n30039 , n30040 , n30041 , n30042 , n30043 , n30044 , n30045 , n30046 , 
     n30047 , n30048 , n30049 , n30050 , n30051 , n30052 , n30053 , n30054 , n30055 , n30056 , 
     n30057 , n30058 , n30059 , n30060 , n30061 , n30062 , n30063 , n30064 , n30065 , n30066 , 
     n30067 , n30068 , n30069 , n30070 , n30071 , n30072 , n30073 , n30074 , n30075 , n30076 , 
     n30077 , n30078 , n30079 , n30080 , n30081 , n30082 , n30083 , n30084 , n30085 , n30086 , 
     n30087 , n30088 , n30089 , n30090 , n30091 , n30092 , n30093 , n30094 , n30095 , n30096 , 
     n30097 , n30098 , n30099 , n30100 , n30101 , n30102 , n30103 , n30104 , n30105 , n30106 , 
     n30107 , n30108 , n30109 , n30110 , n30111 , n30112 , n30113 , n30114 , n30115 , n30116 , 
     n30117 , n30118 , n30119 , n30120 , n30121 , n30122 , n30123 , n30124 , n30125 , n30126 , 
     n30127 , n30128 , n30129 , n30130 , n30131 , n30132 , n30133 , n30134 , n30135 , n30136 , 
     n30137 , n30138 , n30139 , n30140 , n30141 , n30142 , n30143 , n30144 , n30145 , n30146 , 
     n30147 , n30148 , n30149 , n30150 , n30151 , n30152 , n30153 , n30154 , n30155 , n30156 , 
     n30157 , n30158 , n30159 , n30160 , n30161 , n30162 , n30163 , n30164 , n30165 , n30166 , 
     n30167 , n30168 , n30169 , n30170 , n30171 , n30172 , n30173 , n30174 , n30175 , n30176 , 
     n30177 , n30178 , n30179 , n30180 , n30181 , n30182 , n30183 , n30184 , n30185 , n30186 , 
     n30187 , n30188 , n30189 , n30190 , n30191 , n30192 , n30193 , n30194 , n30195 , n30196 , 
     n30197 , n30198 , n30199 , n30200 , n30201 , n30202 , n30203 , n30204 , n30205 , n30206 , 
     n30207 , n30208 , n30209 , n30210 , n30211 , n30212 , n30213 , n30214 , n30215 , n30216 , 
     n30217 , n30218 , n30219 , n30220 , n30221 , n30222 , n30223 , n30224 , n30225 , n30226 , 
     n30227 , n30228 , n30229 , n30230 , n30231 , n30232 , n30233 , n30234 , n30235 , n30236 , 
     n30237 , n30238 , n30239 , n30240 , n30241 , n30242 , n30243 , n30244 , n30245 , n30246 , 
     n30247 , n30248 , n30249 , n30250 , n30251 , n30252 , n30253 , n30254 , n30255 , n30256 , 
     n30257 , n30258 , n30259 , n30260 , n30261 , n30262 , n30263 , n30264 , n30265 , n30266 , 
     n30267 , n30268 , n30269 , n30270 , n30271 , n30272 , n30273 , n30274 , n30275 , n30276 , 
     n30277 , n30278 , n30279 , n30280 , n30281 , n30282 , n30283 , n30284 , n30285 , n30286 , 
     n30287 , n30288 , n30289 , n30290 , n30291 , n30292 , n30293 , n30294 , n30295 , n30296 , 
     n30297 , n30298 , n30299 , n30300 , n30301 , n30302 , n30303 , n30304 , n30305 , n30306 , 
     n30307 , n30308 , n30309 , n30310 , n30311 , n30312 , n30313 , n30314 , n30315 , n30316 , 
     n30317 , n30318 , n30319 , n30320 , n30321 , n30322 , n30323 , n30324 , n30325 , n30326 , 
     n30327 , n30328 , n30329 , n30330 , n30331 , n30332 , n30333 , n30334 , n30335 , n30336 , 
     n30337 , n30338 , n30339 , n30340 , n30341 , n30342 , n30343 , n30344 , n30345 , n30346 , 
     n30347 , n30348 , n30349 , n30350 , n30351 , n30352 , n30353 , n30354 , n30355 , n30356 , 
     n30357 , n30358 , n30359 , n30360 , n30361 , n30362 , n30363 , n30364 , n30365 , n30366 , 
     n30367 , n30368 , n30369 , n30370 , n30371 , n30372 , n30373 , n30374 , n30375 , n30376 , 
     n30377 , n30378 , n30379 , n30380 , n30381 , n30382 , n30383 , n30384 , n30385 , n30386 , 
     n30387 , n30388 , n30389 , n30390 , n30391 , n30392 , n30393 , n30394 , n30395 , n30396 , 
     n30397 , n30398 , n30399 , n30400 , n30401 , n30402 , n30403 , n30404 , n30405 , n30406 , 
     n30407 , n30408 , n30409 , n30410 , n30411 , n30412 , n30413 , n30414 , n30415 , n30416 , 
     n30417 , n30418 , n30419 , n30420 , n30421 , n30422 , n30423 , n30424 , n30425 , n30426 , 
     n30427 , n30428 , n30429 , n30430 , n30431 , n30432 , n30433 , n30434 , n30435 , n30436 , 
     n30437 , n30438 , n30439 , n30440 , n30441 , n30442 , n30443 , n30444 , n30445 , n30446 , 
     n30447 , n30448 , n30449 , n30450 , n30451 , n30452 , n30453 , n30454 , n30455 , n30456 , 
     n30457 , n30458 , n30459 , n30460 , n30461 , n30462 , n30463 , n30464 , n30465 , n30466 , 
     n30467 , n30468 , n30469 , n30470 , n30471 , n30472 , n30473 , n30474 , n30475 , n30476 , 
     n30477 , n30478 , n30479 , n30480 , n30481 , n30482 , n30483 , n30484 , n30485 , n30486 , 
     n30487 , n30488 , n30489 , n30490 , n30491 , n30492 , n30493 , n30494 , n30495 , n30496 , 
     n30497 , n30498 , n30499 , n30500 , n30501 , n30502 , n30503 , n30504 , n30505 , n30506 , 
     n30507 , n30508 , n30509 , n30510 , n30511 , n30512 , n30513 , n30514 , n30515 , n30516 , 
     n30517 , n30518 , n30519 , n30520 , n30521 , n30522 , n30523 , n30524 , n30525 , n30526 , 
     n30527 , n30528 , n30529 , n30530 , n30531 , n30532 , n30533 , n30534 , n30535 , n30536 , 
     n30537 , n30538 , n30539 , n30540 , n30541 , n30542 , n30543 , n30544 , n30545 , n30546 , 
     n30547 , n30548 , n30549 , n30550 , n30551 , n30552 , n30553 , n30554 , n30555 , n30556 , 
     n30557 , n30558 , n30559 , n30560 , n30561 , n30562 , n30563 , n30564 , n30565 , n30566 , 
     n30567 , n30568 , n30569 , n30570 , n30571 , n30572 , n30573 , n30574 , n30575 , n30576 , 
     n30577 , n30578 , n30579 , n30580 , n30581 , n30582 , n30583 , n30584 , n30585 , n30586 , 
     n30587 , n30588 , n30589 , n30590 , n30591 , n30592 , n30593 , n30594 , n30595 , n30596 , 
     n30597 , n30598 , n30599 , n30600 , n30601 , n30602 , n30603 , n30604 , n30605 , n30606 , 
     n30607 , n30608 , n30609 , n30610 , n30611 , n30612 , n30613 , n30614 , n30615 , n30616 , 
     n30617 , n30618 , n30619 , n30620 , n30621 , n30622 , n30623 , n30624 , n30625 , n30626 , 
     n30627 , n30628 , n30629 , n30630 , n30631 , n30632 , n30633 , n30634 , n30635 , n30636 , 
     n30637 , n30638 , n30639 , n30640 , n30641 , n30642 , n30643 , n30644 , n30645 , n30646 , 
     n30647 , n30648 , n30649 , n30650 , n30651 , n30652 , n30653 , n30654 , n30655 , n30656 , 
     n30657 , n30658 , n30659 , n30660 , n30661 , n30662 , n30663 , n30664 , n30665 , n30666 , 
     n30667 , n30668 , n30669 , n30670 , n30671 , n30672 , n30673 , n30674 , n30675 , n30676 , 
     n30677 , n30678 , n30679 , n30680 , n30681 , n30682 , n30683 , n30684 , n30685 , n30686 , 
     n30687 , n30688 , n30689 , n30690 , n30691 , n30692 , n30693 , n30694 , n30695 , n30696 , 
     n30697 , n30698 , n30699 , n30700 , n30701 , n30702 , n30703 , n30704 , n30705 , n30706 , 
     n30707 , n30708 , n30709 , n30710 , n30711 , n30712 , n30713 , n30714 , n30715 , n30716 , 
     n30717 , n30718 , n30719 , n30720 , n30721 , n30722 , n30723 , n30724 , n30725 , n30726 , 
     n30727 , n30728 , n30729 , n30730 , n30731 , n30732 , n30733 , n30734 , n30735 , n30736 , 
     n30737 , n30738 , n30739 , n30740 , n30741 , n30742 , n30743 , n30744 , n30745 , n30746 , 
     n30747 , n30748 , n30749 , n30750 , n30751 , n30752 , n30753 , n30754 , n30755 , n30756 , 
     n30757 , n30758 , n30759 , n30760 , n30761 , n30762 , n30763 , n30764 , n30765 , n30766 , 
     n30767 , n30768 , n30769 , n30770 , n30771 , n30772 , n30773 , n30774 , n30775 , n30776 , 
     n30777 , n30778 , n30779 , n30780 , n30781 , n30782 , n30783 , n30784 , n30785 , n30786 , 
     n30787 , n30788 , n30789 , n30790 , n30791 , n30792 , n30793 , n30794 , n30795 , n30796 , 
     n30797 , n30798 , n30799 , n30800 , n30801 , n30802 , n30803 , n30804 , n30805 , n30806 , 
     n30807 , n30808 , n30809 , n30810 , n30811 , n30812 , n30813 , n30814 , n30815 , n30816 , 
     n30817 , n30818 , n30819 , n30820 , n30821 , n30822 , n30823 , n30824 , n30825 , n30826 , 
     n30827 , n30828 , n30829 , n30830 , n30831 , n30832 , n30833 , n30834 , n30835 , n30836 , 
     n30837 , n30838 , n30839 , n30840 , n30841 , n30842 , n30843 , n30844 , n30845 , n30846 , 
     n30847 , n30848 , n30849 , n30850 , n30851 , n30852 , n30853 , n30854 , n30855 , n30856 , 
     n30857 , n30858 , n30859 , n30860 , n30861 , n30862 , n30863 , n30864 , n30865 , n30866 , 
     n30867 , n30868 , n30869 , n30870 , n30871 , n30872 , n30873 , n30874 , n30875 , n30876 , 
     n30877 , n30878 , n30879 , n30880 , n30881 , n30882 , n30883 , n30884 , n30885 , n30886 , 
     n30887 , n30888 , n30889 , n30890 , n30891 , n30892 , n30893 , n30894 , n30895 , n30896 , 
     n30897 , n30898 , n30899 , n30900 , n30901 , n30902 , n30903 , n30904 , n30905 , n30906 , 
     n30907 , n30908 , n30909 , n30910 , n30911 , n30912 , n30913 , n30914 , n30915 , n30916 , 
     n30917 , n30918 , n30919 , n30920 , n30921 , n30922 , n30923 , n30924 , n30925 , n30926 , 
     n30927 , n30928 , n30929 , n30930 , n30931 , n30932 , n30933 , n30934 , n30935 , n30936 , 
     n30937 , n30938 , n30939 , n30940 , n30941 , n30942 , n30943 , n30944 , n30945 , n30946 , 
     n30947 , n30948 , n30949 , n30950 , n30951 , n30952 , n30953 , n30954 , n30955 , n30956 , 
     n30957 , n30958 , n30959 , n30960 , n30961 , n30962 , n30963 , n30964 , n30965 , n30966 , 
     n30967 , n30968 , n30969 , n30970 , n30971 , n30972 , n30973 , n30974 , n30975 , n30976 , 
     n30977 , n30978 , n30979 , n30980 , n30981 , n30982 , n30983 , n30984 , n30985 , n30986 , 
     n30987 , n30988 , n30989 , n30990 , n30991 , n30992 , n30993 , n30994 , n30995 , n30996 , 
     n30997 , n30998 , n30999 , n31000 , n31001 , n31002 , n31003 , n31004 , n31005 , n31006 , 
     n31007 , n31008 , n31009 , n31010 , n31011 , n31012 , n31013 , n31014 , n31015 , n31016 , 
     n31017 , n31018 , n31019 , n31020 , n31021 , n31022 , n31023 , n31024 , n31025 , n31026 , 
     n31027 , n31028 , n31029 , n31030 , n31031 , n31032 , n31033 , n31034 , n31035 , n31036 , 
     n31037 , n31038 , n31039 , n31040 , n31041 , n31042 , n31043 , n31044 , n31045 , n31046 , 
     n31047 , n31048 , n31049 , n31050 , n31051 , n31052 , n31053 , n31054 , n31055 , n31056 , 
     n31057 , n31058 , n31059 , n31060 , n31061 , n31062 , n31063 , n31064 , n31065 , n31066 , 
     n31067 , n31068 , n31069 , n31070 , n31071 , n31072 , n31073 , n31074 , n31075 , n31076 , 
     n31077 , n31078 , n31079 , n31080 , n31081 , n31082 , n31083 , n31084 , n31085 , n31086 , 
     n31087 , n31088 , n31089 , n31090 , n31091 , n31092 , n31093 , n31094 , n31095 , n31096 , 
     n31097 , n31098 , n31099 , n31100 , n31101 , n31102 , n31103 , n31104 , n31105 , n31106 , 
     n31107 , n31108 , n31109 , n31110 , n31111 , n31112 , n31113 , n31114 , n31115 , n31116 , 
     n31117 , n31118 , n31119 , n31120 , n31121 , n31122 , n31123 , n31124 , n31125 , n31126 , 
     n31127 , n31128 , n31129 , n31130 , n31131 , n31132 , n31133 , n31134 , n31135 , n31136 , 
     n31137 , n31138 , n31139 , n31140 , n31141 , n31142 , n31143 , n31144 , n31145 , n31146 , 
     n31147 , n31148 , n31149 , n31150 , n31151 , n31152 , n31153 , n31154 , n31155 , n31156 , 
     n31157 , n31158 , n31159 , n31160 , n31161 , n31162 , n31163 , n31164 , n31165 , n31166 , 
     n31167 , n31168 , n31169 , n31170 , n31171 , n31172 , n31173 , n31174 , n31175 , n31176 , 
     n31177 , n31178 , n31179 , n31180 , n31181 , n31182 , n31183 , n31184 , n31185 , n31186 , 
     n31187 , n31188 , n31189 , n31190 , n31191 , n31192 , n31193 , n31194 , n31195 , n31196 , 
     n31197 , n31198 , n31199 , n31200 , n31201 , n31202 , n31203 , n31204 , n31205 , n31206 , 
     n31207 , n31208 , n31209 , n31210 , n31211 , n31212 , n31213 , n31214 , n31215 , n31216 , 
     n31217 , n31218 , n31219 , n31220 , n31221 , n31222 , n31223 , n31224 , n31225 , n31226 , 
     n31227 , n31228 , n31229 , n31230 , n31231 , n31232 , n31233 , n31234 , n31235 , n31236 , 
     n31237 , n31238 , n31239 , n31240 , n31241 , n31242 , n31243 , n31244 , n31245 , n31246 , 
     n31247 , n31248 , n31249 , n31250 , n31251 , n31252 , n31253 , n31254 , n31255 , n31256 , 
     n31257 , n31258 , n31259 , n31260 , n31261 , n31262 , n31263 , n31264 , n31265 , n31266 , 
     n31267 , n31268 , n31269 , n31270 , n31271 , n31272 , n31273 , n31274 , n31275 , n31276 , 
     n31277 , n31278 , n31279 , n31280 , n31281 , n31282 , n31283 , n31284 , n31285 , n31286 , 
     n31287 , n31288 , n31289 , n31290 , n31291 , n31292 , n31293 , n31294 , n31295 , n31296 , 
     n31297 , n31298 , n31299 , n31300 , n31301 , n31302 , n31303 , n31304 , n31305 , n31306 , 
     n31307 , n31308 , n31309 , n31310 , n31311 , n31312 , n31313 , n31314 , n31315 , n31316 , 
     n31317 , n31318 , n31319 , n31320 , n31321 , n31322 , n31323 , n31324 , n31325 , n31326 , 
     n31327 , n31328 , n31329 , n31330 , n31331 , n31332 , n31333 , n31334 , n31335 , n31336 , 
     n31337 , n31338 , n31339 , n31340 , n31341 , n31342 , n31343 , n31344 , n31345 , n31346 , 
     n31347 , n31348 , n31349 , n31350 , n31351 , n31352 , n31353 , n31354 , n31355 , n31356 , 
     n31357 , n31358 , n31359 , n31360 , n31361 , n31362 , n31363 , n31364 , n31365 , n31366 , 
     n31367 , n31368 , n31369 , n31370 , n31371 , n31372 , n31373 , n31374 , n31375 , n31376 , 
     n31377 , n31378 , n31379 , n31380 , n31381 , n31382 , n31383 , n31384 , n31385 , n31386 , 
     n31387 , n31388 , n31389 , n31390 , n31391 , n31392 , n31393 , n31394 , n31395 , n31396 , 
     n31397 , n31398 , n31399 , n31400 , n31401 , n31402 , n31403 , n31404 , n31405 , n31406 , 
     n31407 , n31408 , n31409 , n31410 , n31411 , n31412 , n31413 , n31414 , n31415 , n31416 , 
     n31417 , n31418 , n31419 , n31420 , n31421 , n31422 , n31423 , n31424 , n31425 , n31426 , 
     n31427 , n31428 , n31429 , n31430 , n31431 , n31432 , n31433 , n31434 , n31435 , n31436 , 
     n31437 , n31438 , n31439 , n31440 , n31441 , n31442 , n31443 , n31444 , n31445 , n31446 , 
     n31447 , n31448 , n31449 , n31450 , n31451 , n31452 , n31453 , n31454 , n31455 , n31456 , 
     n31457 , n31458 , n31459 , n31460 , n31461 , n31462 , n31463 , n31464 , n31465 , n31466 , 
     n31467 , n31468 , n31469 , n31470 , n31471 , n31472 , n31473 , n31474 , n31475 , n31476 , 
     n31477 , n31478 , n31479 , n31480 , n31481 , n31482 , n31483 , n31484 , n31485 , n31486 , 
     n31487 , n31488 , n31489 , n31490 , n31491 , n31492 , n31493 , n31494 , n31495 , n31496 , 
     n31497 , n31498 , n31499 , n31500 , n31501 , n31502 , n31503 , n31504 , n31505 , n31506 , 
     n31507 , n31508 , n31509 , n31510 , n31511 , n31512 , n31513 , n31514 , n31515 , n31516 , 
     n31517 , n31518 , n31519 , n31520 , n31521 , n31522 , n31523 , n31524 , n31525 , n31526 , 
     n31527 , n31528 , n31529 , n31530 , n31531 , n31532 , n31533 , n31534 , n31535 , n31536 , 
     n31537 , n31538 , n31539 , n31540 , n31541 , n31542 , n31543 , n31544 , n31545 , n31546 , 
     n31547 , n31548 , n31549 , n31550 , n31551 , n31552 , n31553 , n31554 , n31555 , n31556 , 
     n31557 , n31558 , n31559 , n31560 , n31561 , n31562 , n31563 , n31564 , n31565 , n31566 , 
     n31567 , n31568 , n31569 , n31570 , n31571 , n31572 , n31573 , n31574 , n31575 , n31576 , 
     n31577 , n31578 , n31579 , n31580 , n31581 , n31582 , n31583 , n31584 , n31585 , n31586 , 
     n31587 , n31588 , n31589 , n31590 , n31591 , n31592 , n31593 , n31594 , n31595 , n31596 , 
     n31597 , n31598 , n31599 , n31600 , n31601 , n31602 , n31603 , n31604 , n31605 , n31606 , 
     n31607 , n31608 , n31609 , n31610 , n31611 , n31612 , n31613 , n31614 , n31615 , n31616 , 
     n31617 , n31618 , n31619 , n31620 , n31621 , n31622 , n31623 , n31624 , n31625 , n31626 , 
     n31627 , n31628 , n31629 , n31630 , n31631 , n31632 , n31633 , n31634 , n31635 , n31636 , 
     n31637 , n31638 , n31639 , n31640 , n31641 , n31642 , n31643 , n31644 , n31645 , n31646 , 
     n31647 , n31648 , n31649 , n31650 , n31651 , n31652 , n31653 , n31654 , n31655 , n31656 , 
     n31657 , n31658 , n31659 , n31660 , n31661 , n31662 , n31663 , n31664 , n31665 , n31666 , 
     n31667 , n31668 , n31669 , n31670 , n31671 , n31672 , n31673 , n31674 , n31675 , n31676 , 
     n31677 , n31678 , n31679 , n31680 , n31681 , n31682 , n31683 , n31684 , n31685 , n31686 , 
     n31687 , n31688 , n31689 , n31690 , n31691 , n31692 , n31693 , n31694 , n31695 , n31696 , 
     n31697 , n31698 , n31699 , n31700 , n31701 , n31702 , n31703 , n31704 , n31705 , n31706 , 
     n31707 , n31708 , n31709 , n31710 , n31711 , n31712 , n31713 , n31714 , n31715 , n31716 , 
     n31717 , n31718 , n31719 , n31720 , n31721 , n31722 , n31723 , n31724 , n31725 , n31726 , 
     n31727 , n31728 , n31729 , n31730 , n31731 , n31732 , n31733 , n31734 , n31735 , n31736 , 
     n31737 , n31738 , n31739 , n31740 , n31741 , n31742 , n31743 , n31744 , n31745 , n31746 , 
     n31747 , n31748 , n31749 , n31750 , n31751 , n31752 , n31753 , n31754 , n31755 , n31756 , 
     n31757 , n31758 , n31759 , n31760 , n31761 , n31762 , n31763 , n31764 , n31765 , n31766 , 
     n31767 , n31768 , n31769 , n31770 , n31771 , n31772 , n31773 , n31774 , n31775 , n31776 , 
     n31777 , n31778 , n31779 , n31780 , n31781 , n31782 , n31783 , n31784 , n31785 , n31786 , 
     n31787 , n31788 , n31789 , n31790 , n31791 , n31792 , n31793 , n31794 , n31795 , n31796 , 
     n31797 , n31798 , n31799 , n31800 , n31801 , n31802 , n31803 , n31804 , n31805 , n31806 , 
     n31807 , n31808 , n31809 , n31810 , n31811 , n31812 , n31813 , n31814 , n31815 , n31816 , 
     n31817 , n31818 , n31819 , n31820 , n31821 , n31822 , n31823 , n31824 , n31825 , n31826 , 
     n31827 , n31828 , n31829 , n31830 , n31831 , n31832 , n31833 , n31834 , n31835 , n31836 , 
     n31837 , n31838 , n31839 , n31840 , n31841 , n31842 , n31843 , n31844 , n31845 , n31846 , 
     n31847 , n31848 , n31849 , n31850 , n31851 , n31852 , n31853 , n31854 , n31855 , n31856 , 
     n31857 , n31858 , n31859 , n31860 , n31861 , n31862 , n31863 , n31864 , n31865 , n31866 , 
     n31867 , n31868 , n31869 , n31870 , n31871 , n31872 , n31873 , n31874 , n31875 , n31876 , 
     n31877 , n31878 , n31879 , n31880 , n31881 , n31882 , n31883 , n31884 , n31885 , n31886 , 
     n31887 , n31888 , n31889 , n31890 , n31891 , n31892 , n31893 , n31894 , n31895 , n31896 , 
     n31897 , n31898 , n31899 , n31900 , n31901 , n31902 , n31903 , n31904 , n31905 , n31906 , 
     n31907 , n31908 , n31909 , n31910 , n31911 , n31912 , n31913 , n31914 , n31915 , n31916 , 
     n31917 , n31918 , n31919 , n31920 , n31921 , n31922 , n31923 , n31924 , n31925 , n31926 , 
     n31927 , n31928 , n31929 , n31930 , n31931 , n31932 , n31933 , n31934 , n31935 , n31936 , 
     n31937 , n31938 , n31939 , n31940 , n31941 , n31942 , n31943 , n31944 , n31945 , n31946 , 
     n31947 , n31948 , n31949 , n31950 , n31951 , n31952 , n31953 , n31954 , n31955 , n31956 , 
     n31957 , n31958 , n31959 , n31960 , n31961 , n31962 , n31963 , n31964 , n31965 , n31966 , 
     n31967 , n31968 , n31969 , n31970 , n31971 , n31972 , n31973 , n31974 , n31975 , n31976 , 
     n31977 , n31978 , n31979 , n31980 , n31981 , n31982 , n31983 , n31984 , n31985 , n31986 , 
     n31987 , n31988 , n31989 , n31990 , n31991 , n31992 , n31993 , n31994 , n31995 , n31996 , 
     n31997 , n31998 , n31999 , n32000 , n32001 , n32002 , n32003 , n32004 , n32005 , n32006 , 
     n32007 , n32008 , n32009 , n32010 , n32011 , n32012 , n32013 , n32014 , n32015 , n32016 , 
     n32017 , n32018 , n32019 , n32020 , n32021 , n32022 , n32023 , n32024 , n32025 , n32026 , 
     n32027 , n32028 , n32029 , n32030 , n32031 , n32032 , n32033 , n32034 , n32035 , n32036 , 
     n32037 , n32038 , n32039 , n32040 , n32041 , n32042 , n32043 , n32044 , n32045 , n32046 , 
     n32047 , n32048 , n32049 , n32050 , n32051 , n32052 , n32053 , n32054 , n32055 , n32056 , 
     n32057 , n32058 , n32059 , n32060 , n32061 , n32062 , n32063 , n32064 , n32065 , n32066 , 
     n32067 , n32068 , n32069 , n32070 , n32071 , n32072 , n32073 , n32074 , n32075 , n32076 , 
     n32077 , n32078 , n32079 , n32080 , n32081 , n32082 , n32083 , n32084 , n32085 , n32086 , 
     n32087 , n32088 , n32089 , n32090 , n32091 , n32092 , n32093 , n32094 , n32095 , n32096 , 
     n32097 , n32098 , n32099 , n32100 , n32101 , n32102 , n32103 , n32104 , n32105 , n32106 , 
     n32107 , n32108 , n32109 , n32110 , n32111 , n32112 , n32113 , n32114 , n32115 , n32116 , 
     n32117 , n32118 , n32119 , n32120 , n32121 , n32122 , n32123 , n32124 , n32125 , n32126 , 
     n32127 , n32128 , n32129 , n32130 , n32131 , n32132 , n32133 , n32134 , n32135 , n32136 , 
     n32137 , n32138 , n32139 , n32140 , n32141 , n32142 , n32143 , n32144 , n32145 , n32146 , 
     n32147 , n32148 , n32149 , n32150 , n32151 , n32152 , n32153 , n32154 , n32155 , n32156 , 
     n32157 , n32158 , n32159 , n32160 , n32161 , n32162 , n32163 , n32164 , n32165 , n32166 , 
     n32167 , n32168 , n32169 , n32170 , n32171 , n32172 , n32173 , n32174 , n32175 , n32176 , 
     n32177 , n32178 , n32179 , n32180 , n32181 , n32182 , n32183 , n32184 , n32185 , n32186 , 
     n32187 , n32188 , n32189 , n32190 , n32191 , n32192 , n32193 , n32194 , n32195 , n32196 , 
     n32197 , n32198 , n32199 , n32200 , n32201 , n32202 , n32203 , n32204 , n32205 , n32206 , 
     n32207 , n32208 , n32209 , n32210 , n32211 , n32212 , n32213 , n32214 , n32215 , n32216 , 
     n32217 , n32218 , n32219 , n32220 , n32221 , n32222 , n32223 , n32224 , n32225 , n32226 , 
     n32227 , n32228 , n32229 , n32230 , n32231 , n32232 , n32233 , n32234 , n32235 , n32236 , 
     n32237 , n32238 , n32239 , n32240 , n32241 , n32242 , n32243 , n32244 , n32245 , n32246 , 
     n32247 , n32248 , n32249 , n32250 , n32251 , n32252 , n32253 , n32254 , n32255 , n32256 , 
     n32257 , n32258 , n32259 , n32260 , n32261 , n32262 , n32263 , n32264 , n32265 , n32266 , 
     n32267 , n32268 , n32269 , n32270 , n32271 , n32272 , n32273 , n32274 , n32275 , n32276 , 
     n32277 , n32278 , n32279 , n32280 , n32281 , n32282 , n32283 , n32284 , n32285 , n32286 , 
     n32287 , n32288 , n32289 , n32290 , n32291 , n32292 , n32293 , n32294 , n32295 , n32296 , 
     n32297 , n32298 , n32299 , n32300 , n32301 , n32302 , n32303 , n32304 , n32305 , n32306 , 
     n32307 , n32308 , n32309 , n32310 , n32311 , n32312 , n32313 , n32314 , n32315 , n32316 , 
     n32317 , n32318 , n32319 , n32320 , n32321 , n32322 , n32323 , n32324 , n32325 , n32326 , 
     n32327 , n32328 , n32329 , n32330 , n32331 , n32332 , n32333 , n32334 , n32335 , n32336 , 
     n32337 , n32338 , n32339 , n32340 , n32341 , n32342 , n32343 , n32344 , n32345 , n32346 , 
     n32347 , n32348 , n32349 , n32350 , n32351 , n32352 , n32353 , n32354 , n32355 , n32356 , 
     n32357 , n32358 , n32359 , n32360 , n32361 , n32362 , n32363 , n32364 , n32365 , n32366 , 
     n32367 , n32368 , n32369 , n32370 , n32371 , n32372 , n32373 , n32374 , n32375 , n32376 , 
     n32377 , n32378 , n32379 , n32380 , n32381 , n32382 , n32383 , n32384 , n32385 , n32386 , 
     n32387 , n32388 , n32389 , n32390 , n32391 , n32392 , n32393 , n32394 , n32395 , n32396 , 
     n32397 , n32398 , n32399 , n32400 , n32401 , n32402 , n32403 , n32404 , n32405 , n32406 , 
     n32407 , n32408 , n32409 , n32410 , n32411 , n32412 , n32413 , n32414 , n32415 , n32416 , 
     n32417 , n32418 , n32419 , n32420 , n32421 , n32422 , n32423 , n32424 , n32425 , n32426 , 
     n32427 , n32428 , n32429 , n32430 , n32431 , n32432 , n32433 , n32434 , n32435 , n32436 , 
     n32437 , n32438 , n32439 , n32440 , n32441 , n32442 , n32443 , n32444 , n32445 , n32446 , 
     n32447 , n32448 , n32449 , n32450 , n32451 , n32452 , n32453 , n32454 , n32455 , n32456 , 
     n32457 , n32458 , n32459 , n32460 , n32461 , n32462 , n32463 , n32464 , n32465 , n32466 , 
     n32467 , n32468 , n32469 , n32470 , n32471 , n32472 , n32473 , n32474 , n32475 , n32476 , 
     n32477 , n32478 , n32479 , n32480 , n32481 , n32482 , n32483 , n32484 , n32485 , n32486 , 
     n32487 , n32488 , n32489 , n32490 , n32491 , n32492 , n32493 , n32494 , n32495 , n32496 , 
     n32497 , n32498 , n32499 , n32500 , n32501 , n32502 , n32503 , n32504 , n32505 , n32506 , 
     n32507 , n32508 , n32509 , n32510 , n32511 , n32512 , n32513 , n32514 , n32515 , n32516 , 
     n32517 , n32518 , n32519 , n32520 , n32521 , n32522 , n32523 , n32524 , n32525 , n32526 , 
     n32527 , n32528 , n32529 , n32530 , n32531 , n32532 , n32533 , n32534 , n32535 , n32536 , 
     n32537 , n32538 , n32539 , n32540 , n32541 , n32542 , n32543 , n32544 , n32545 , n32546 , 
     n32547 , n32548 , n32549 , n32550 , n32551 , n32552 , n32553 , n32554 , n32555 , n32556 , 
     n32557 , n32558 , n32559 , n32560 , n32561 , n32562 , n32563 , n32564 , n32565 , n32566 , 
     n32567 , n32568 , n32569 , n32570 , n32571 , n32572 , n32573 , n32574 , n32575 , n32576 , 
     n32577 , n32578 , n32579 , n32580 , n32581 , n32582 , n32583 , n32584 , n32585 , n32586 , 
     n32587 , n32588 , n32589 , n32590 , n32591 , n32592 , n32593 , n32594 , n32595 , n32596 , 
     n32597 , n32598 , n32599 , n32600 , n32601 , n32602 , n32603 , n32604 , n32605 , n32606 , 
     n32607 , n32608 , n32609 , n32610 , n32611 , n32612 , n32613 , n32614 , n32615 , n32616 , 
     n32617 , n32618 , n32619 , n32620 , n32621 , n32622 , n32623 , n32624 , n32625 , n32626 , 
     n32627 , n32628 , n32629 , n32630 , n32631 , n32632 , n32633 , n32634 , n32635 , n32636 , 
     n32637 , n32638 , n32639 , n32640 , n32641 , n32642 , n32643 , n32644 , n32645 , n32646 , 
     n32647 , n32648 , n32649 , n32650 , n32651 , n32652 , n32653 , n32654 , n32655 , n32656 , 
     n32657 , n32658 , n32659 , n32660 , n32661 , n32662 , n32663 , n32664 , n32665 , n32666 , 
     n32667 , n32668 , n32669 , n32670 , n32671 , n32672 , n32673 , n32674 , n32675 , n32676 , 
     n32677 , n32678 , n32679 , n32680 , n32681 , n32682 , n32683 , n32684 , n32685 , n32686 , 
     n32687 , n32688 , n32689 , n32690 , n32691 , n32692 , n32693 , n32694 , n32695 , n32696 , 
     n32697 , n32698 , n32699 , n32700 , n32701 , n32702 , n32703 , n32704 , n32705 , n32706 , 
     n32707 , n32708 , n32709 , n32710 , n32711 , n32712 , n32713 , n32714 , n32715 , n32716 , 
     n32717 , n32718 , n32719 , n32720 , n32721 , n32722 , n32723 , n32724 , n32725 , n32726 , 
     n32727 , n32728 , n32729 , n32730 , n32731 , n32732 , n32733 , n32734 , n32735 , n32736 , 
     n32737 , n32738 , n32739 , n32740 , n32741 , n32742 , n32743 , n32744 , n32745 , n32746 , 
     n32747 , n32748 , n32749 , n32750 , n32751 , n32752 , n32753 , n32754 , n32755 , n32756 , 
     n32757 , n32758 , n32759 , n32760 , n32761 , n32762 , n32763 , n32764 , n32765 , n32766 , 
     n32767 , n32768 , n32769 , n32770 , n32771 , n32772 , n32773 , n32774 , n32775 , n32776 , 
     n32777 , n32778 , n32779 , n32780 , n32781 , n32782 , n32783 , n32784 , n32785 , n32786 , 
     n32787 , n32788 , n32789 , n32790 , n32791 , n32792 , n32793 , n32794 , n32795 , n32796 , 
     n32797 , n32798 , n32799 , n32800 , n32801 , n32802 , n32803 , n32804 , n32805 , n32806 , 
     n32807 , n32808 , n32809 , n32810 , n32811 , n32812 , n32813 , n32814 , n32815 , n32816 , 
     n32817 , n32818 , n32819 , n32820 , n32821 , n32822 , n32823 , n32824 , n32825 , n32826 , 
     n32827 , n32828 , n32829 , n32830 , n32831 , n32832 , n32833 , n32834 , n32835 , n32836 , 
     n32837 , n32838 , n32839 , n32840 , n32841 , n32842 , n32843 , n32844 , n32845 , n32846 , 
     n32847 , n32848 , n32849 , n32850 , n32851 , n32852 , n32853 , n32854 , n32855 , n32856 , 
     n32857 , n32858 , n32859 , n32860 , n32861 , n32862 , n32863 , n32864 , n32865 , n32866 , 
     n32867 , n32868 , n32869 , n32870 , n32871 , n32872 , n32873 , n32874 , n32875 , n32876 , 
     n32877 , n32878 , n32879 , n32880 , n32881 , n32882 , n32883 , n32884 , n32885 , n32886 , 
     n32887 , n32888 , n32889 , n32890 , n32891 , n32892 , n32893 , n32894 , n32895 , n32896 , 
     n32897 , n32898 , n32899 , n32900 , n32901 , n32902 , n32903 , n32904 , n32905 , n32906 , 
     n32907 , n32908 , n32909 , n32910 , n32911 , n32912 , n32913 , n32914 , n32915 , n32916 , 
     n32917 , n32918 , n32919 , n32920 , n32921 , n32922 , n32923 , n32924 , n32925 , n32926 , 
     n32927 , n32928 , n32929 , n32930 , n32931 , n32932 , n32933 , n32934 , n32935 , n32936 , 
     n32937 , n32938 , n32939 , n32940 , n32941 , n32942 , n32943 , n32944 , n32945 , n32946 , 
     n32947 , n32948 , n32949 , n32950 , n32951 , n32952 , n32953 , n32954 , n32955 , n32956 , 
     n32957 , n32958 , n32959 , n32960 , n32961 , n32962 , n32963 , n32964 , n32965 , n32966 , 
     n32967 , n32968 , n32969 , n32970 , n32971 , n32972 , n32973 , n32974 , n32975 , n32976 , 
     n32977 , n32978 , n32979 , n32980 , n32981 , n32982 , n32983 , n32984 , n32985 , n32986 , 
     n32987 , n32988 , n32989 , n32990 , n32991 , n32992 , n32993 , n32994 , n32995 , n32996 , 
     n32997 , n32998 , n32999 , n33000 , n33001 , n33002 , n33003 , n33004 , n33005 , n33006 , 
     n33007 , n33008 , n33009 , n33010 , n33011 , n33012 , n33013 , n33014 , n33015 , n33016 , 
     n33017 , n33018 , n33019 , n33020 , n33021 , n33022 , n33023 , n33024 , n33025 , n33026 , 
     n33027 , n33028 , n33029 , n33030 , n33031 , n33032 , n33033 , n33034 , n33035 , n33036 , 
     n33037 , n33038 , n33039 , n33040 , n33041 , n33042 , n33043 , n33044 , n33045 , n33046 , 
     n33047 , n33048 , n33049 , n33050 , n33051 , n33052 , n33053 , n33054 , n33055 , n33056 , 
     n33057 , n33058 , n33059 , n33060 , n33061 , n33062 , n33063 , n33064 , n33065 , n33066 , 
     n33067 , n33068 , n33069 , n33070 , n33071 , n33072 , n33073 , n33074 , n33075 , n33076 , 
     n33077 , n33078 , n33079 , n33080 , n33081 , n33082 , n33083 , n33084 , n33085 , n33086 , 
     n33087 , n33088 , n33089 , n33090 , n33091 , n33092 , n33093 , n33094 , n33095 , n33096 , 
     n33097 , n33098 , n33099 , n33100 , n33101 , n33102 , n33103 , n33104 , n33105 , n33106 , 
     n33107 , n33108 , n33109 , n33110 , n33111 , n33112 , n33113 , n33114 , n33115 , n33116 , 
     n33117 , n33118 , n33119 , n33120 , n33121 , n33122 , n33123 , n33124 , n33125 , n33126 , 
     n33127 , n33128 , n33129 , n33130 , n33131 , n33132 , n33133 , n33134 , n33135 , n33136 , 
     n33137 , n33138 , n33139 , n33140 , n33141 , n33142 , n33143 , n33144 , n33145 , n33146 , 
     n33147 , n33148 , n33149 , n33150 , n33151 , n33152 , n33153 , n33154 , n33155 , n33156 , 
     n33157 , n33158 , n33159 , n33160 , n33161 , n33162 , n33163 , n33164 , n33165 , n33166 , 
     n33167 , n33168 , n33169 , n33170 , n33171 , n33172 , n33173 , n33174 , n33175 , n33176 , 
     n33177 , n33178 , n33179 , n33180 , n33181 , n33182 , n33183 , n33184 , n33185 , n33186 , 
     n33187 , n33188 , n33189 , n33190 , n33191 , n33192 , n33193 , n33194 , n33195 , n33196 , 
     n33197 , n33198 , n33199 , n33200 , n33201 , n33202 , n33203 , n33204 , n33205 , n33206 , 
     n33207 , n33208 , n33209 , n33210 , n33211 , n33212 , n33213 , n33214 , n33215 , n33216 , 
     n33217 , n33218 , n33219 , n33220 , n33221 , n33222 , n33223 , n33224 , n33225 , n33226 , 
     n33227 , n33228 , n33229 , n33230 , n33231 , n33232 , n33233 , n33234 , n33235 , n33236 , 
     n33237 , n33238 , n33239 , n33240 , n33241 , n33242 , n33243 , n33244 , n33245 , n33246 , 
     n33247 , n33248 , n33249 , n33250 , n33251 , n33252 , n33253 , n33254 , n33255 , n33256 , 
     n33257 , n33258 , n33259 , n33260 , n33261 , n33262 , n33263 , n33264 , n33265 , n33266 , 
     n33267 , n33268 , n33269 , n33270 , n33271 , n33272 , n33273 , n33274 , n33275 , n33276 , 
     n33277 , n33278 , n33279 , n33280 , n33281 , n33282 , n33283 , n33284 , n33285 , n33286 , 
     n33287 , n33288 , n33289 , n33290 , n33291 , n33292 , n33293 , n33294 , n33295 , n33296 , 
     n33297 , n33298 , n33299 , n33300 , n33301 , n33302 , n33303 , n33304 , n33305 , n33306 , 
     n33307 , n33308 , n33309 , n33310 , n33311 , n33312 , n33313 , n33314 , n33315 , n33316 , 
     n33317 , n33318 , n33319 , n33320 , n33321 , n33322 , n33323 , n33324 , n33325 , n33326 , 
     n33327 , n33328 , n33329 , n33330 , n33331 , n33332 , n33333 , n33334 , n33335 , n33336 , 
     n33337 , n33338 , n33339 , n33340 , n33341 , n33342 , n33343 , n33344 , n33345 , n33346 , 
     n33347 , n33348 , n33349 , n33350 , n33351 , n33352 , n33353 , n33354 , n33355 , n33356 , 
     n33357 , n33358 , n33359 , n33360 , n33361 , n33362 , n33363 , n33364 , n33365 , n33366 , 
     n33367 , n33368 , n33369 , n33370 , n33371 , n33372 , n33373 , n33374 , n33375 , n33376 , 
     n33377 , n33378 , n33379 , n33380 , n33381 , n33382 , n33383 , n33384 , n33385 , n33386 , 
     n33387 , n33388 , n33389 , n33390 , n33391 , n33392 , n33393 , n33394 , n33395 , n33396 , 
     n33397 , n33398 , n33399 , n33400 , n33401 , n33402 , n33403 , n33404 , n33405 , n33406 , 
     n33407 , n33408 , n33409 , n33410 , n33411 , n33412 , n33413 , n33414 , n33415 , n33416 , 
     n33417 , n33418 , n33419 , n33420 , n33421 , n33422 , n33423 , n33424 , n33425 , n33426 , 
     n33427 , n33428 , n33429 , n33430 , n33431 , n33432 , n33433 , n33434 , n33435 , n33436 , 
     n33437 , n33438 , n33439 , n33440 , n33441 , n33442 , n33443 , n33444 , n33445 , n33446 , 
     n33447 , n33448 , n33449 , n33450 , n33451 , n33452 , n33453 , n33454 , n33455 , n33456 , 
     n33457 , n33458 , n33459 , n33460 , n33461 , n33462 , n33463 , n33464 , n33465 , n33466 , 
     n33467 , n33468 , n33469 , n33470 , n33471 , n33472 , n33473 , n33474 , n33475 , n33476 , 
     n33477 , n33478 , n33479 , n33480 , n33481 , n33482 , n33483 , n33484 , n33485 , n33486 , 
     n33487 , n33488 , n33489 , n33490 , n33491 , n33492 , n33493 , n33494 , n33495 , n33496 , 
     n33497 , n33498 , n33499 , n33500 , n33501 , n33502 , n33503 , n33504 , n33505 , n33506 , 
     n33507 , n33508 , n33509 , n33510 , n33511 , n33512 , n33513 , n33514 , n33515 , n33516 , 
     n33517 , n33518 , n33519 , n33520 , n33521 , n33522 , n33523 , n33524 , n33525 , n33526 , 
     n33527 , n33528 , n33529 , n33530 , n33531 , n33532 , n33533 , n33534 , n33535 , n33536 , 
     n33537 , n33538 , n33539 , n33540 , n33541 , n33542 , n33543 , n33544 , n33545 , n33546 , 
     n33547 , n33548 , n33549 , n33550 , n33551 , n33552 , n33553 , n33554 , n33555 , n33556 , 
     n33557 , n33558 , n33559 , n33560 , n33561 , n33562 , n33563 , n33564 , n33565 , n33566 , 
     n33567 , n33568 , n33569 , n33570 , n33571 , n33572 , n33573 , n33574 , n33575 , n33576 , 
     n33577 , n33578 , n33579 , n33580 , n33581 , n33582 , n33583 , n33584 , n33585 , n33586 , 
     n33587 , n33588 , n33589 , n33590 , n33591 , n33592 , n33593 , n33594 , n33595 , n33596 , 
     n33597 , n33598 , n33599 , n33600 , n33601 , n33602 , n33603 , n33604 , n33605 , n33606 , 
     n33607 , n33608 , n33609 , n33610 , n33611 , n33612 , n33613 , n33614 , n33615 , n33616 , 
     n33617 , n33618 , n33619 , n33620 , n33621 , n33622 , n33623 , n33624 , n33625 , n33626 , 
     n33627 , n33628 , n33629 , n33630 , n33631 , n33632 , n33633 , n33634 , n33635 , n33636 , 
     n33637 , n33638 , n33639 , n33640 , n33641 , n33642 , n33643 , n33644 , n33645 , n33646 , 
     n33647 , n33648 , n33649 , n33650 , n33651 , n33652 , n33653 , n33654 , n33655 , n33656 , 
     n33657 , n33658 , n33659 , n33660 , n33661 , n33662 , n33663 , n33664 , n33665 , n33666 , 
     n33667 , n33668 , n33669 , n33670 , n33671 , n33672 , n33673 , n33674 , n33675 , n33676 , 
     n33677 , n33678 , n33679 , n33680 , n33681 , n33682 , n33683 , n33684 , n33685 , n33686 , 
     n33687 , n33688 , n33689 , n33690 , n33691 , n33692 , n33693 , n33694 , n33695 , n33696 , 
     n33697 , n33698 , n33699 , n33700 , n33701 , n33702 , n33703 , n33704 , n33705 , n33706 , 
     n33707 , n33708 , n33709 , n33710 , n33711 , n33712 , n33713 , n33714 , n33715 , n33716 , 
     n33717 , n33718 , n33719 , n33720 , n33721 , n33722 , n33723 , n33724 , n33725 , n33726 , 
     n33727 , n33728 , n33729 , n33730 , n33731 , n33732 , n33733 , n33734 , n33735 , n33736 , 
     n33737 , n33738 , n33739 , n33740 , n33741 , n33742 , n33743 , n33744 , n33745 , n33746 , 
     n33747 , n33748 , n33749 , n33750 , n33751 , n33752 , n33753 , n33754 , n33755 , n33756 , 
     n33757 , n33758 , n33759 , n33760 , n33761 , n33762 , n33763 , n33764 , n33765 , n33766 , 
     n33767 , n33768 , n33769 , n33770 , n33771 , n33772 , n33773 , n33774 , n33775 , n33776 , 
     n33777 , n33778 , n33779 , n33780 , n33781 , n33782 , n33783 , n33784 , n33785 , n33786 , 
     n33787 , n33788 , n33789 , n33790 , n33791 , n33792 , n33793 , n33794 , n33795 , n33796 , 
     n33797 , n33798 , n33799 , n33800 , n33801 , n33802 , n33803 , n33804 , n33805 , n33806 , 
     n33807 , n33808 , n33809 , n33810 , n33811 , n33812 , n33813 , n33814 , n33815 , n33816 , 
     n33817 , n33818 , n33819 , n33820 , n33821 , n33822 , n33823 , n33824 , n33825 , n33826 , 
     n33827 , n33828 , n33829 , n33830 , n33831 , n33832 , n33833 , n33834 , n33835 , n33836 , 
     n33837 , n33838 , n33839 , n33840 , n33841 , n33842 , n33843 , n33844 , n33845 , n33846 , 
     n33847 , n33848 , n33849 , n33850 , n33851 , n33852 , n33853 , n33854 , n33855 , n33856 , 
     n33857 , n33858 , n33859 , n33860 , n33861 , n33862 , n33863 , n33864 , n33865 , n33866 , 
     n33867 , n33868 , n33869 , n33870 , n33871 , n33872 , n33873 , n33874 , n33875 , n33876 , 
     n33877 , n33878 , n33879 , n33880 , n33881 , n33882 , n33883 , n33884 , n33885 , n33886 , 
     n33887 , n33888 , n33889 , n33890 , n33891 , n33892 , n33893 , n33894 , n33895 , n33896 , 
     n33897 , n33898 , n33899 , n33900 , n33901 , n33902 , n33903 , n33904 , n33905 , n33906 , 
     n33907 , n33908 , n33909 , n33910 , n33911 , n33912 , n33913 , n33914 , n33915 , n33916 , 
     n33917 , n33918 , n33919 , n33920 , n33921 , n33922 , n33923 , n33924 , n33925 , n33926 , 
     n33927 , n33928 , n33929 , n33930 , n33931 , n33932 , n33933 , n33934 , n33935 , n33936 , 
     n33937 , n33938 , n33939 , n33940 , n33941 , n33942 , n33943 , n33944 , n33945 , n33946 , 
     n33947 , n33948 , n33949 , n33950 , n33951 , n33952 , n33953 , n33954 , n33955 , n33956 , 
     n33957 , n33958 , n33959 , n33960 , n33961 , n33962 , n33963 , n33964 , n33965 , n33966 , 
     n33967 , n33968 , n33969 , n33970 , n33971 , n33972 , n33973 , n33974 , n33975 , n33976 , 
     n33977 , n33978 , n33979 , n33980 , n33981 , n33982 , n33983 , n33984 , n33985 , n33986 , 
     n33987 , n33988 , n33989 , n33990 , n33991 , n33992 , n33993 , n33994 , n33995 , n33996 , 
     n33997 , n33998 , n33999 , n34000 , n34001 , n34002 , n34003 , n34004 , n34005 , n34006 , 
     n34007 , n34008 , n34009 , n34010 , n34011 , n34012 , n34013 , n34014 , n34015 , n34016 , 
     n34017 , n34018 , n34019 , n34020 , n34021 , n34022 , n34023 , n34024 , n34025 , n34026 , 
     n34027 , n34028 , n34029 , n34030 , n34031 , n34032 , n34033 , n34034 , n34035 , n34036 , 
     n34037 , n34038 , n34039 , n34040 , n34041 , n34042 , n34043 , n34044 , n34045 , n34046 , 
     n34047 , n34048 , n34049 , n34050 , n34051 , n34052 , n34053 , n34054 , n34055 , n34056 , 
     n34057 , n34058 , n34059 , n34060 , n34061 , n34062 , n34063 , n34064 , n34065 , n34066 , 
     n34067 , n34068 , n34069 , n34070 , n34071 , n34072 , n34073 , n34074 , n34075 , n34076 , 
     n34077 , n34078 , n34079 , n34080 , n34081 , n34082 , n34083 , n34084 , n34085 , n34086 , 
     n34087 , n34088 , n34089 , n34090 , n34091 , n34092 , n34093 , n34094 , n34095 , n34096 , 
     n34097 , n34098 , n34099 , n34100 , n34101 , n34102 , n34103 , n34104 , n34105 , n34106 , 
     n34107 , n34108 , n34109 , n34110 , n34111 , n34112 , n34113 , n34114 , n34115 , n34116 , 
     n34117 , n34118 , n34119 , n34120 , n34121 , n34122 , n34123 , n34124 , n34125 , n34126 , 
     n34127 , n34128 , n34129 , n34130 , n34131 , n34132 , n34133 , n34134 , n34135 , n34136 , 
     n34137 , n34138 , n34139 , n34140 , n34141 , n34142 , n34143 , n34144 , n34145 , n34146 , 
     n34147 , n34148 , n34149 , n34150 , n34151 , n34152 , n34153 , n34154 , n34155 , n34156 , 
     n34157 , n34158 , n34159 , n34160 , n34161 , n34162 , n34163 , n34164 , n34165 , n34166 , 
     n34167 , n34168 , n34169 , n34170 , n34171 , n34172 , n34173 , n34174 , n34175 , n34176 , 
     n34177 , n34178 , n34179 , n34180 , n34181 , n34182 , n34183 , n34184 , n34185 , n34186 , 
     n34187 , n34188 , n34189 , n34190 , n34191 , n34192 , n34193 , n34194 , n34195 , n34196 , 
     n34197 , n34198 , n34199 , n34200 , n34201 , n34202 , n34203 , n34204 , n34205 , n34206 , 
     n34207 , n34208 , n34209 , n34210 , n34211 , n34212 , n34213 , n34214 , n34215 , n34216 , 
     n34217 , n34218 , n34219 , n34220 , n34221 , n34222 , n34223 , n34224 , n34225 , n34226 , 
     n34227 , n34228 , n34229 , n34230 , n34231 , n34232 , n34233 , n34234 , n34235 , n34236 , 
     n34237 , n34238 , n34239 , n34240 , n34241 , n34242 , n34243 , n34244 , n34245 , n34246 , 
     n34247 , n34248 , n34249 , n34250 , n34251 , n34252 , n34253 , n34254 , n34255 , n34256 , 
     n34257 , n34258 , n34259 , n34260 , n34261 , n34262 , n34263 , n34264 , n34265 , n34266 , 
     n34267 , n34268 , n34269 , n34270 , n34271 , n34272 , n34273 , n34274 , n34275 , n34276 , 
     n34277 , n34278 , n34279 , n34280 , n34281 , n34282 , n34283 , n34284 , n34285 , n34286 , 
     n34287 , n34288 , n34289 , n34290 , n34291 , n34292 , n34293 , n34294 , n34295 , n34296 , 
     n34297 , n34298 , n34299 , n34300 , n34301 , n34302 , n34303 , n34304 , n34305 , n34306 , 
     n34307 , n34308 , n34309 , n34310 , n34311 , n34312 , n34313 , n34314 , n34315 , n34316 , 
     n34317 , n34318 , n34319 , n34320 , n34321 , n34322 , n34323 , n34324 , n34325 , n34326 , 
     n34327 , n34328 , n34329 , n34330 , n34331 , n34332 , n34333 , n34334 , n34335 , n34336 , 
     n34337 , n34338 , n34339 , n34340 , n34341 , n34342 , n34343 , n34344 , n34345 , n34346 , 
     n34347 , n34348 , n34349 , n34350 , n34351 , n34352 , n34353 , n34354 , n34355 , n34356 , 
     n34357 , n34358 , n34359 , n34360 , n34361 , n34362 , n34363 , n34364 , n34365 , n34366 , 
     n34367 , n34368 , n34369 , n34370 , n34371 , n34372 , n34373 , n34374 , n34375 , n34376 , 
     n34377 , n34378 , n34379 , n34380 , n34381 , n34382 , n34383 , n34384 , n34385 , n34386 , 
     n34387 , n34388 , n34389 , n34390 , n34391 , n34392 , n34393 , n34394 , n34395 , n34396 , 
     n34397 , n34398 , n34399 , n34400 , n34401 , n34402 , n34403 , n34404 , n34405 , n34406 , 
     n34407 , n34408 , n34409 , n34410 , n34411 , n34412 , n34413 , n34414 , n34415 , n34416 , 
     n34417 , n34418 , n34419 , n34420 , n34421 , n34422 , n34423 , n34424 , n34425 , n34426 , 
     n34427 , n34428 , n34429 , n34430 , n34431 , n34432 , n34433 , n34434 , n34435 , n34436 , 
     n34437 , n34438 , n34439 , n34440 , n34441 , n34442 , n34443 , n34444 , n34445 , n34446 , 
     n34447 , n34448 , n34449 , n34450 , n34451 , n34452 , n34453 , n34454 , n34455 , n34456 , 
     n34457 , n34458 , n34459 , n34460 , n34461 , n34462 , n34463 , n34464 , n34465 , n34466 , 
     n34467 , n34468 , n34469 , n34470 , n34471 , n34472 , n34473 , n34474 , n34475 , n34476 , 
     n34477 , n34478 , n34479 , n34480 , n34481 , n34482 , n34483 , n34484 , n34485 , n34486 , 
     n34487 , n34488 , n34489 , n34490 , n34491 , n34492 , n34493 , n34494 , n34495 , n34496 , 
     n34497 , n34498 , n34499 , n34500 , n34501 , n34502 , n34503 , n34504 , n34505 , n34506 , 
     n34507 , n34508 , n34509 , n34510 , n34511 , n34512 , n34513 , n34514 , n34515 , n34516 , 
     n34517 , n34518 , n34519 , n34520 , n34521 , n34522 , n34523 , n34524 , n34525 , n34526 , 
     n34527 , n34528 , n34529 , n34530 , n34531 , n34532 , n34533 , n34534 , n34535 , n34536 , 
     n34537 , n34538 , n34539 , n34540 , n34541 , n34542 , n34543 , n34544 , n34545 , n34546 , 
     n34547 , n34548 , n34549 , n34550 , n34551 , n34552 , n34553 , n34554 , n34555 , n34556 , 
     n34557 , n34558 , n34559 , n34560 , n34561 , n34562 , n34563 , n34564 , n34565 , n34566 , 
     n34567 , n34568 , n34569 , n34570 , n34571 , n34572 , n34573 , n34574 , n34575 , n34576 , 
     n34577 , n34578 , n34579 , n34580 , n34581 , n34582 , n34583 , n34584 , n34585 , n34586 , 
     n34587 , n34588 , n34589 , n34590 , n34591 , n34592 , n34593 , n34594 , n34595 , n34596 , 
     n34597 , n34598 , n34599 , n34600 , n34601 , n34602 , n34603 , n34604 , n34605 , n34606 , 
     n34607 , n34608 , n34609 , n34610 , n34611 , n34612 , n34613 , n34614 , n34615 , n34616 , 
     n34617 , n34618 , n34619 , n34620 , n34621 , n34622 , n34623 , n34624 , n34625 , n34626 , 
     n34627 , n34628 , n34629 , n34630 , n34631 , n34632 , n34633 , n34634 , n34635 , n34636 , 
     n34637 , n34638 , n34639 , n34640 , n34641 , n34642 , n34643 , n34644 , n34645 , n34646 , 
     n34647 , n34648 , n34649 , n34650 , n34651 , n34652 , n34653 , n34654 , n34655 , n34656 , 
     n34657 , n34658 , n34659 , n34660 , n34661 , n34662 , n34663 , n34664 , n34665 , n34666 , 
     n34667 , n34668 , n34669 , n34670 , n34671 , n34672 , n34673 , n34674 , n34675 , n34676 , 
     n34677 , n34678 , n34679 , n34680 , n34681 , n34682 , n34683 , n34684 , n34685 , n34686 , 
     n34687 , n34688 , n34689 , n34690 , n34691 , n34692 , n34693 , n34694 , n34695 , n34696 , 
     n34697 , n34698 , n34699 , n34700 , n34701 , n34702 , n34703 , n34704 , n34705 , n34706 , 
     n34707 , n34708 , n34709 , n34710 , n34711 , n34712 , n34713 , n34714 , n34715 , n34716 , 
     n34717 , n34718 , n34719 , n34720 , n34721 , n34722 , n34723 , n34724 , n34725 , n34726 , 
     n34727 , n34728 , n34729 , n34730 , n34731 , n34732 , n34733 , n34734 , n34735 , n34736 , 
     n34737 , n34738 , n34739 , n34740 , n34741 , n34742 , n34743 , n34744 , n34745 , n34746 , 
     n34747 , n34748 , n34749 , n34750 , n34751 , n34752 , n34753 , n34754 , n34755 , n34756 , 
     n34757 , n34758 , n34759 , n34760 , n34761 , n34762 , n34763 , n34764 , n34765 , n34766 , 
     n34767 , n34768 , n34769 , n34770 , n34771 , n34772 , n34773 , n34774 , n34775 , n34776 , 
     n34777 , n34778 , n34779 , n34780 , n34781 , n34782 , n34783 , n34784 , n34785 , n34786 , 
     n34787 , n34788 , n34789 , n34790 , n34791 , n34792 , n34793 , n34794 , n34795 , n34796 , 
     n34797 , n34798 , n34799 , n34800 , n34801 , n34802 , n34803 , n34804 , n34805 , n34806 , 
     n34807 , n34808 , n34809 , n34810 , n34811 , n34812 , n34813 , n34814 , n34815 , n34816 , 
     n34817 , n34818 , n34819 , n34820 , n34821 , n34822 , n34823 , n34824 , n34825 , n34826 , 
     n34827 , n34828 , n34829 , n34830 , n34831 , n34832 , n34833 , n34834 , n34835 , n34836 , 
     n34837 , n34838 , n34839 , n34840 , n34841 , n34842 , n34843 , n34844 , n34845 , n34846 , 
     n34847 , n34848 , n34849 , n34850 , n34851 , n34852 , n34853 , n34854 , n34855 , n34856 , 
     n34857 , n34858 , n34859 , n34860 , n34861 , n34862 , n34863 , n34864 , n34865 , n34866 , 
     n34867 , n34868 , n34869 , n34870 , n34871 , n34872 , n34873 , n34874 , n34875 , n34876 , 
     n34877 , n34878 , n34879 , n34880 , n34881 , n34882 , n34883 , n34884 , n34885 , n34886 , 
     n34887 , n34888 , n34889 , n34890 , n34891 , n34892 , n34893 , n34894 , n34895 , n34896 , 
     n34897 , n34898 , n34899 , n34900 , n34901 , n34902 , n34903 , n34904 , n34905 , n34906 , 
     n34907 , n34908 , n34909 , n34910 , n34911 , n34912 , n34913 , n34914 , n34915 , n34916 , 
     n34917 , n34918 , n34919 , n34920 , n34921 , n34922 , n34923 , n34924 , n34925 , n34926 , 
     n34927 , n34928 , n34929 , n34930 , n34931 , n34932 , n34933 , n34934 , n34935 , n34936 , 
     n34937 , n34938 , n34939 , n34940 , n34941 , n34942 , n34943 , n34944 , n34945 , n34946 , 
     n34947 , n34948 , n34949 , n34950 , n34951 , n34952 , n34953 , n34954 , n34955 , n34956 , 
     n34957 , n34958 , n34959 , n34960 , n34961 , n34962 , n34963 , n34964 , n34965 , n34966 , 
     n34967 , n34968 , n34969 , n34970 , n34971 , n34972 , n34973 , n34974 , n34975 , n34976 , 
     n34977 , n34978 , n34979 , n34980 , n34981 , n34982 , n34983 , n34984 , n34985 , n34986 , 
     n34987 , n34988 , n34989 , n34990 , n34991 , n34992 , n34993 , n34994 , n34995 , n34996 , 
     n34997 , n34998 , n34999 , n35000 , n35001 , n35002 , n35003 , n35004 , n35005 , n35006 , 
     n35007 , n35008 , n35009 , n35010 , n35011 , n35012 , n35013 , n35014 , n35015 , n35016 , 
     n35017 , n35018 , n35019 , n35020 , n35021 , n35022 , n35023 , n35024 , n35025 , n35026 , 
     n35027 , n35028 , n35029 , n35030 , n35031 , n35032 , n35033 , n35034 , n35035 , n35036 , 
     n35037 , n35038 , n35039 , n35040 , n35041 , n35042 , n35043 , n35044 , n35045 , n35046 , 
     n35047 , n35048 , n35049 , n35050 , n35051 , n35052 , n35053 , n35054 , n35055 , n35056 , 
     n35057 , n35058 , n35059 , n35060 , n35061 , n35062 , n35063 , n35064 , n35065 , n35066 , 
     n35067 , n35068 , n35069 , n35070 , n35071 , n35072 , n35073 , n35074 , n35075 , n35076 , 
     n35077 , n35078 , n35079 , n35080 , n35081 , n35082 , n35083 , n35084 , n35085 , n35086 , 
     n35087 , n35088 , n35089 , n35090 , n35091 , n35092 , n35093 , n35094 , n35095 , n35096 , 
     n35097 , n35098 , n35099 , n35100 , n35101 , n35102 , n35103 , n35104 , n35105 , n35106 , 
     n35107 , n35108 , n35109 , n35110 , n35111 , n35112 , n35113 , n35114 , n35115 , n35116 , 
     n35117 , n35118 , n35119 , n35120 , n35121 , n35122 , n35123 , n35124 , n35125 , n35126 , 
     n35127 , n35128 , n35129 , n35130 , n35131 , n35132 , n35133 , n35134 , n35135 , n35136 , 
     n35137 , n35138 , n35139 , n35140 , n35141 , n35142 , n35143 , n35144 , n35145 , n35146 , 
     n35147 , n35148 , n35149 , n35150 , n35151 , n35152 , n35153 , n35154 , n35155 , n35156 , 
     n35157 , n35158 , n35159 , n35160 , n35161 , n35162 , n35163 , n35164 , n35165 , n35166 , 
     n35167 , n35168 , n35169 , n35170 , n35171 , n35172 , n35173 , n35174 , n35175 , n35176 , 
     n35177 , n35178 , n35179 , n35180 , n35181 , n35182 , n35183 , n35184 , n35185 , n35186 , 
     n35187 , n35188 , n35189 , n35190 , n35191 , n35192 , n35193 , n35194 , n35195 , n35196 , 
     n35197 , n35198 , n35199 , n35200 , n35201 , n35202 , n35203 , n35204 , n35205 , n35206 , 
     n35207 , n35208 , n35209 , n35210 , n35211 , n35212 , n35213 , n35214 , n35215 , n35216 , 
     n35217 , n35218 , n35219 , n35220 , n35221 , n35222 , n35223 , n35224 , n35225 , n35226 , 
     n35227 , n35228 , n35229 , n35230 , n35231 , n35232 , n35233 , n35234 , n35235 , n35236 , 
     n35237 , n35238 , n35239 , n35240 , n35241 , n35242 , n35243 , n35244 , n35245 , n35246 , 
     n35247 , n35248 , n35249 , n35250 , n35251 , n35252 , n35253 , n35254 , n35255 , n35256 , 
     n35257 , n35258 , n35259 , n35260 , n35261 , n35262 , n35263 , n35264 , n35265 , n35266 , 
     n35267 , n35268 , n35269 , n35270 , n35271 , n35272 , n35273 , n35274 , n35275 , n35276 , 
     n35277 , n35278 , n35279 , n35280 , n35281 , n35282 , n35283 , n35284 , n35285 , n35286 , 
     n35287 , n35288 , n35289 , n35290 , n35291 , n35292 , n35293 , n35294 , n35295 , n35296 , 
     n35297 , n35298 , n35299 , n35300 , n35301 , n35302 , n35303 , n35304 , n35305 , n35306 , 
     n35307 , n35308 , n35309 , n35310 , n35311 , n35312 , n35313 , n35314 , n35315 , n35316 , 
     n35317 , n35318 , n35319 , n35320 , n35321 , n35322 , n35323 , n35324 , n35325 , n35326 , 
     n35327 , n35328 , n35329 , n35330 , n35331 , n35332 , n35333 , n35334 , n35335 , n35336 , 
     n35337 , n35338 , n35339 , n35340 , n35341 , n35342 , n35343 , n35344 , n35345 , n35346 , 
     n35347 , n35348 , n35349 , n35350 , n35351 , n35352 , n35353 , n35354 , n35355 , n35356 , 
     n35357 , n35358 , n35359 , n35360 , n35361 , n35362 , n35363 , n35364 , n35365 , n35366 , 
     n35367 , n35368 , n35369 , n35370 , n35371 , n35372 , n35373 , n35374 , n35375 , n35376 , 
     n35377 , n35378 , n35379 , n35380 , n35381 , n35382 , n35383 , n35384 , n35385 , n35386 , 
     n35387 , n35388 , n35389 , n35390 , n35391 , n35392 , n35393 , n35394 , n35395 , n35396 , 
     n35397 , n35398 , n35399 , n35400 , n35401 , n35402 , n35403 , n35404 , n35405 , n35406 , 
     n35407 , n35408 , n35409 , n35410 , n35411 , n35412 , n35413 , n35414 , n35415 , n35416 , 
     n35417 , n35418 , n35419 , n35420 , n35421 , n35422 , n35423 , n35424 , n35425 , n35426 , 
     n35427 , n35428 , n35429 , n35430 , n35431 , n35432 , n35433 , n35434 , n35435 , n35436 , 
     n35437 , n35438 , n35439 , n35440 , n35441 , n35442 , n35443 , n35444 , n35445 , n35446 , 
     n35447 , n35448 , n35449 , n35450 , n35451 , n35452 , n35453 , n35454 , n35455 , n35456 , 
     n35457 , n35458 , n35459 , n35460 , n35461 , n35462 , n35463 , n35464 , n35465 , n35466 , 
     n35467 , n35468 , n35469 , n35470 , n35471 , n35472 , n35473 , n35474 , n35475 , n35476 , 
     n35477 , n35478 , n35479 , n35480 , n35481 , n35482 , n35483 , n35484 , n35485 , n35486 , 
     n35487 , n35488 , n35489 , n35490 , n35491 , n35492 , n35493 , n35494 , n35495 , n35496 , 
     n35497 , n35498 , n35499 , n35500 , n35501 , n35502 , n35503 , n35504 , n35505 , n35506 , 
     n35507 , n35508 , n35509 , n35510 , n35511 , n35512 , n35513 , n35514 , n35515 , n35516 , 
     n35517 , n35518 , n35519 , n35520 , n35521 , n35522 , n35523 , n35524 , n35525 , n35526 , 
     n35527 , n35528 , n35529 , n35530 , n35531 , n35532 , n35533 , n35534 , n35535 , n35536 , 
     n35537 , n35538 , n35539 , n35540 , n35541 , n35542 , n35543 , n35544 , n35545 , n35546 , 
     n35547 , n35548 , n35549 , n35550 , n35551 , n35552 , n35553 , n35554 , n35555 , n35556 , 
     n35557 , n35558 , n35559 , n35560 , n35561 , n35562 , n35563 , n35564 , n35565 , n35566 , 
     n35567 , n35568 , n35569 , n35570 , n35571 , n35572 , n35573 , n35574 , n35575 , n35576 , 
     n35577 , n35578 , n35579 , n35580 , n35581 , n35582 , n35583 , n35584 , n35585 , n35586 , 
     n35587 , n35588 , n35589 , n35590 , n35591 , n35592 , n35593 , n35594 , n35595 , n35596 , 
     n35597 , n35598 , n35599 , n35600 , n35601 , n35602 , n35603 , n35604 , n35605 , n35606 , 
     n35607 , n35608 , n35609 , n35610 , n35611 , n35612 , n35613 , n35614 , n35615 , n35616 , 
     n35617 , n35618 , n35619 , n35620 , n35621 , n35622 , n35623 , n35624 , n35625 , n35626 , 
     n35627 , n35628 , n35629 , n35630 , n35631 , n35632 , n35633 , n35634 , n35635 , n35636 , 
     n35637 , n35638 , n35639 , n35640 , n35641 , n35642 , n35643 , n35644 , n35645 , n35646 , 
     n35647 , n35648 , n35649 , n35650 , n35651 , n35652 , n35653 , n35654 , n35655 , n35656 , 
     n35657 , n35658 , n35659 , n35660 , n35661 , n35662 , n35663 , n35664 , n35665 , n35666 , 
     n35667 , n35668 , n35669 , n35670 , n35671 , n35672 , n35673 , n35674 , n35675 , n35676 , 
     n35677 , n35678 , n35679 , n35680 , n35681 , n35682 , n35683 , n35684 , n35685 , n35686 , 
     n35687 , n35688 , n35689 , n35690 , n35691 , n35692 , n35693 , n35694 , n35695 , n35696 , 
     n35697 , n35698 , n35699 , n35700 , n35701 , n35702 , n35703 , n35704 , n35705 , n35706 , 
     n35707 , n35708 , n35709 , n35710 , n35711 , n35712 , n35713 , n35714 , n35715 , n35716 , 
     n35717 , n35718 , n35719 , n35720 , n35721 , n35722 , n35723 , n35724 , n35725 , n35726 , 
     n35727 , n35728 , n35729 , n35730 , n35731 , n35732 , n35733 , n35734 , n35735 , n35736 , 
     n35737 , n35738 , n35739 , n35740 , n35741 , n35742 , n35743 , n35744 , n35745 , n35746 , 
     n35747 , n35748 , n35749 , n35750 , n35751 , n35752 , n35753 , n35754 , n35755 , n35756 , 
     n35757 , n35758 , n35759 , n35760 , n35761 , n35762 , n35763 , n35764 , n35765 , n35766 , 
     n35767 , n35768 , n35769 , n35770 , n35771 , n35772 , n35773 , n35774 , n35775 , n35776 , 
     n35777 , n35778 , n35779 , n35780 , n35781 , n35782 , n35783 , n35784 , n35785 , n35786 , 
     n35787 , n35788 , n35789 , n35790 , n35791 , n35792 , n35793 , n35794 , n35795 , n35796 , 
     n35797 , n35798 , n35799 , n35800 , n35801 , n35802 , n35803 , n35804 , n35805 , n35806 , 
     n35807 , n35808 , n35809 , n35810 , n35811 , n35812 , n35813 , n35814 , n35815 , n35816 , 
     n35817 , n35818 , n35819 , n35820 , n35821 , n35822 , n35823 , n35824 , n35825 , n35826 , 
     n35827 , n35828 , n35829 , n35830 , n35831 , n35832 , n35833 , n35834 , n35835 , n35836 , 
     n35837 , n35838 , n35839 , n35840 , n35841 , n35842 , n35843 , n35844 , n35845 , n35846 , 
     n35847 , n35848 , n35849 , n35850 , n35851 , n35852 , n35853 , n35854 , n35855 , n35856 , 
     n35857 , n35858 , n35859 , n35860 , n35861 , n35862 , n35863 , n35864 , n35865 , n35866 , 
     n35867 , n35868 , n35869 , n35870 , n35871 , n35872 , n35873 , n35874 , n35875 , n35876 , 
     n35877 , n35878 , n35879 , n35880 , n35881 , n35882 , n35883 , n35884 , n35885 , n35886 , 
     n35887 , n35888 , n35889 , n35890 , n35891 , n35892 , n35893 , n35894 , n35895 , n35896 , 
     n35897 , n35898 , n35899 , n35900 , n35901 , n35902 , n35903 , n35904 , n35905 , n35906 , 
     n35907 , n35908 , n35909 , n35910 , n35911 , n35912 , n35913 , n35914 , n35915 , n35916 , 
     n35917 , n35918 , n35919 , n35920 , n35921 , n35922 , n35923 , n35924 , n35925 , n35926 , 
     n35927 , n35928 , n35929 , n35930 , n35931 , n35932 , n35933 , n35934 , n35935 , n35936 , 
     n35937 , n35938 , n35939 , n35940 , n35941 , n35942 , n35943 , n35944 , n35945 , n35946 , 
     n35947 , n35948 , n35949 , n35950 , n35951 , n35952 , n35953 , n35954 , n35955 , n35956 , 
     n35957 , n35958 , n35959 , n35960 , n35961 , n35962 , n35963 , n35964 , n35965 , n35966 , 
     n35967 , n35968 , n35969 , n35970 , n35971 , n35972 , n35973 , n35974 , n35975 , n35976 , 
     n35977 , n35978 , n35979 , n35980 , n35981 , n35982 , n35983 , n35984 , n35985 , n35986 , 
     n35987 , n35988 , n35989 , n35990 , n35991 , n35992 , n35993 , n35994 , n35995 , n35996 , 
     n35997 , n35998 , n35999 , n36000 , n36001 , n36002 , n36003 , n36004 , n36005 , n36006 , 
     n36007 , n36008 , n36009 , n36010 , n36011 , n36012 , n36013 , n36014 , n36015 , n36016 , 
     n36017 , n36018 , n36019 , n36020 , n36021 , n36022 , n36023 , n36024 , n36025 , n36026 , 
     n36027 , n36028 , n36029 , n36030 , n36031 , n36032 , n36033 , n36034 , n36035 , n36036 , 
     n36037 , n36038 , n36039 , n36040 , n36041 , n36042 , n36043 , n36044 , n36045 , n36046 , 
     n36047 , n36048 , n36049 , n36050 , n36051 , n36052 , n36053 , n36054 , n36055 , n36056 , 
     n36057 , n36058 , n36059 , n36060 , n36061 , n36062 , n36063 , n36064 , n36065 , n36066 , 
     n36067 , n36068 , n36069 , n36070 , n36071 , n36072 , n36073 , n36074 , n36075 , n36076 , 
     n36077 , n36078 , n36079 , n36080 , n36081 , n36082 , n36083 , n36084 , n36085 , n36086 , 
     n36087 , n36088 , n36089 , n36090 , n36091 , n36092 , n36093 , n36094 , n36095 , n36096 , 
     n36097 , n36098 , n36099 , n36100 , n36101 , n36102 , n36103 , n36104 , n36105 , n36106 , 
     n36107 , n36108 , n36109 , n36110 , n36111 , n36112 , n36113 , n36114 , n36115 , n36116 , 
     n36117 , n36118 , n36119 , n36120 , n36121 , n36122 , n36123 , n36124 , n36125 , n36126 , 
     n36127 , n36128 , n36129 , n36130 , n36131 , n36132 , n36133 , n36134 , n36135 , n36136 , 
     n36137 , n36138 , n36139 , n36140 , n36141 , n36142 , n36143 , n36144 , n36145 , n36146 , 
     n36147 , n36148 , n36149 , n36150 , n36151 , n36152 , n36153 , n36154 , n36155 , n36156 , 
     n36157 , n36158 , n36159 , n36160 , n36161 , n36162 , n36163 , n36164 , n36165 , n36166 , 
     n36167 , n36168 , n36169 , n36170 , n36171 , n36172 , n36173 , n36174 , n36175 , n36176 , 
     n36177 , n36178 , n36179 , n36180 , n36181 , n36182 , n36183 , n36184 , n36185 , n36186 , 
     n36187 , n36188 , n36189 , n36190 , n36191 , n36192 , n36193 , n36194 , n36195 , n36196 , 
     n36197 , n36198 , n36199 , n36200 , n36201 , n36202 , n36203 , n36204 , n36205 , n36206 , 
     n36207 , n36208 , n36209 , n36210 , n36211 , n36212 , n36213 , n36214 , n36215 , n36216 , 
     n36217 , n36218 , n36219 , n36220 , n36221 , n36222 , n36223 , n36224 , n36225 , n36226 , 
     n36227 , n36228 , n36229 , n36230 , n36231 , n36232 , n36233 , n36234 , n36235 , n36236 , 
     n36237 , n36238 , n36239 , n36240 , n36241 , n36242 , n36243 , n36244 , n36245 , n36246 , 
     n36247 , n36248 , n36249 , n36250 , n36251 , n36252 , n36253 , n36254 , n36255 , n36256 , 
     n36257 , n36258 , n36259 , n36260 , n36261 , n36262 , n36263 , n36264 , n36265 , n36266 , 
     n36267 , n36268 , n36269 , n36270 , n36271 , n36272 , n36273 , n36274 , n36275 , n36276 , 
     n36277 , n36278 , n36279 , n36280 , n36281 , n36282 , n36283 , n36284 , n36285 , n36286 , 
     n36287 , n36288 , n36289 , n36290 , n36291 , n36292 , n36293 , n36294 , n36295 , n36296 , 
     n36297 , n36298 , n36299 , n36300 , n36301 , n36302 , n36303 , n36304 , n36305 , n36306 , 
     n36307 , n36308 , n36309 , n36310 , n36311 , n36312 , n36313 , n36314 , n36315 , n36316 , 
     n36317 , n36318 , n36319 , n36320 , n36321 , n36322 , n36323 , n36324 , n36325 , n36326 , 
     n36327 , n36328 , n36329 , n36330 , n36331 , n36332 , n36333 , n36334 , n36335 , n36336 , 
     n36337 , n36338 , n36339 , n36340 , n36341 , n36342 , n36343 , n36344 , n36345 , n36346 , 
     n36347 , n36348 , n36349 , n36350 , n36351 , n36352 , n36353 , n36354 , n36355 , n36356 , 
     n36357 , n36358 , n36359 , n36360 , n36361 , n36362 , n36363 , n36364 , n36365 , n36366 , 
     n36367 , n36368 , n36369 , n36370 , n36371 , n36372 , n36373 , n36374 , n36375 , n36376 , 
     n36377 , n36378 , n36379 , n36380 , n36381 , n36382 , n36383 , n36384 , n36385 , n36386 , 
     n36387 , n36388 , n36389 , n36390 , n36391 , n36392 , n36393 , n36394 , n36395 , n36396 , 
     n36397 , n36398 , n36399 , n36400 , n36401 , n36402 , n36403 , n36404 , n36405 , n36406 , 
     n36407 , n36408 , n36409 , n36410 , n36411 , n36412 , n36413 , n36414 , n36415 , n36416 , 
     n36417 , n36418 , n36419 , n36420 , n36421 , n36422 , n36423 , n36424 , n36425 , n36426 , 
     n36427 , n36428 , n36429 , n36430 , n36431 , n36432 , n36433 , n36434 , n36435 , n36436 , 
     n36437 , n36438 , n36439 , n36440 , n36441 , n36442 , n36443 , n36444 , n36445 , n36446 , 
     n36447 , n36448 , n36449 , n36450 , n36451 , n36452 , n36453 , n36454 , n36455 , n36456 , 
     n36457 , n36458 , n36459 , n36460 , n36461 , n36462 , n36463 , n36464 , n36465 , n36466 , 
     n36467 , n36468 , n36469 , n36470 , n36471 , n36472 , n36473 , n36474 , n36475 , n36476 , 
     n36477 , n36478 , n36479 , n36480 , n36481 , n36482 , n36483 , n36484 , n36485 , n36486 , 
     n36487 , n36488 , n36489 , n36490 , n36491 , n36492 , n36493 , n36494 , n36495 , n36496 , 
     n36497 , n36498 , n36499 , n36500 , n36501 , n36502 , n36503 , n36504 , n36505 , n36506 , 
     n36507 , n36508 , n36509 , n36510 , n36511 , n36512 , n36513 , n36514 , n36515 , n36516 , 
     n36517 , n36518 , n36519 , n36520 , n36521 , n36522 , n36523 , n36524 , n36525 , n36526 , 
     n36527 , n36528 , n36529 , n36530 , n36531 , n36532 , n36533 , n36534 , n36535 , n36536 , 
     n36537 , n36538 , n36539 , n36540 , n36541 , n36542 , n36543 , n36544 , n36545 , n36546 , 
     n36547 , n36548 , n36549 , n36550 , n36551 , n36552 , n36553 , n36554 , n36555 , n36556 , 
     n36557 , n36558 , n36559 , n36560 , n36561 , n36562 , n36563 , n36564 , n36565 , n36566 , 
     n36567 , n36568 , n36569 , n36570 , n36571 , n36572 , n36573 , n36574 , n36575 , n36576 , 
     n36577 , n36578 , n36579 , n36580 , n36581 , n36582 , n36583 , n36584 , n36585 , n36586 , 
     n36587 , n36588 , n36589 , n36590 , n36591 , n36592 , n36593 , n36594 , n36595 , n36596 , 
     n36597 , n36598 , n36599 , n36600 , n36601 , n36602 , n36603 , n36604 , n36605 , n36606 , 
     n36607 , n36608 , n36609 , n36610 , n36611 , n36612 , n36613 , n36614 , n36615 , n36616 , 
     n36617 , n36618 , n36619 , n36620 , n36621 , n36622 , n36623 , n36624 , n36625 , n36626 , 
     n36627 , n36628 , n36629 , n36630 , n36631 , n36632 , n36633 , n36634 , n36635 , n36636 , 
     n36637 , n36638 , n36639 , n36640 , n36641 , n36642 , n36643 , n36644 , n36645 , n36646 , 
     n36647 , n36648 , n36649 , n36650 , n36651 , n36652 , n36653 , n36654 , n36655 , n36656 , 
     n36657 , n36658 , n36659 , n36660 , n36661 , n36662 , n36663 , n36664 , n36665 , n36666 , 
     n36667 , n36668 , n36669 , n36670 , n36671 , n36672 , n36673 , n36674 , n36675 , n36676 , 
     n36677 , n36678 , n36679 , n36680 , n36681 , n36682 , n36683 , n36684 , n36685 , n36686 , 
     n36687 , n36688 , n36689 , n36690 , n36691 , n36692 , n36693 , n36694 , n36695 , n36696 , 
     n36697 , n36698 , n36699 , n36700 , n36701 , n36702 , n36703 , n36704 , n36705 , n36706 , 
     n36707 , n36708 , n36709 , n36710 , n36711 , n36712 , n36713 , n36714 , n36715 , n36716 , 
     n36717 , n36718 , n36719 , n36720 , n36721 , n36722 , n36723 , n36724 , n36725 , n36726 , 
     n36727 , n36728 , n36729 , n36730 , n36731 , n36732 , n36733 , n36734 , n36735 , n36736 , 
     n36737 , n36738 , n36739 , n36740 , n36741 , n36742 , n36743 , n36744 , n36745 , n36746 , 
     n36747 , n36748 , n36749 , n36750 , n36751 , n36752 , n36753 , n36754 , n36755 , n36756 , 
     n36757 , n36758 , n36759 , n36760 , n36761 , n36762 , n36763 , n36764 , n36765 , n36766 , 
     n36767 , n36768 , n36769 , n36770 , n36771 , n36772 , n36773 , n36774 , n36775 , n36776 , 
     n36777 , n36778 , n36779 , n36780 , n36781 , n36782 , n36783 , n36784 , n36785 , n36786 , 
     n36787 , n36788 , n36789 , n36790 , n36791 , n36792 , n36793 , n36794 , n36795 , n36796 , 
     n36797 , n36798 , n36799 , n36800 , n36801 , n36802 , n36803 , n36804 , n36805 , n36806 , 
     n36807 , n36808 , n36809 , n36810 , n36811 , n36812 , n36813 , n36814 , n36815 , n36816 , 
     n36817 , n36818 , n36819 , n36820 , n36821 , n36822 , n36823 , n36824 , n36825 , n36826 , 
     n36827 , n36828 , n36829 , n36830 , n36831 , n36832 , n36833 , n36834 , n36835 , n36836 , 
     n36837 , n36838 , n36839 , n36840 , n36841 , n36842 , n36843 , n36844 , n36845 , n36846 , 
     n36847 , n36848 , n36849 , n36850 , n36851 , n36852 , n36853 , n36854 , n36855 , n36856 , 
     n36857 , n36858 , n36859 , n36860 , n36861 , n36862 , n36863 , n36864 , n36865 , n36866 , 
     n36867 , n36868 , n36869 , n36870 , n36871 , n36872 , n36873 , n36874 , n36875 , n36876 , 
     n36877 , n36878 , n36879 , n36880 , n36881 , n36882 , n36883 , n36884 , n36885 , n36886 , 
     n36887 , n36888 , n36889 , n36890 , n36891 , n36892 , n36893 , n36894 , n36895 , n36896 , 
     n36897 , n36898 , n36899 , n36900 , n36901 , n36902 , n36903 , n36904 , n36905 , n36906 , 
     n36907 , n36908 , n36909 , n36910 , n36911 , n36912 , n36913 , n36914 , n36915 , n36916 , 
     n36917 , n36918 , n36919 , n36920 , n36921 , n36922 , n36923 , n36924 , n36925 , n36926 , 
     n36927 , n36928 , n36929 , n36930 , n36931 , n36932 , n36933 , n36934 , n36935 , n36936 , 
     n36937 , n36938 , n36939 , n36940 , n36941 , n36942 , n36943 , n36944 , n36945 , n36946 , 
     n36947 , n36948 , n36949 , n36950 , n36951 , n36952 , n36953 , n36954 , n36955 , n36956 , 
     n36957 , n36958 , n36959 , n36960 , n36961 , n36962 , n36963 , n36964 , n36965 , n36966 , 
     n36967 , n36968 , n36969 , n36970 , n36971 , n36972 , n36973 , n36974 , n36975 , n36976 , 
     n36977 , n36978 , n36979 , n36980 , n36981 , n36982 , n36983 , n36984 , n36985 , n36986 , 
     n36987 , n36988 , n36989 , n36990 , n36991 , n36992 , n36993 , n36994 , n36995 , n36996 , 
     n36997 , n36998 , n36999 , n37000 , n37001 , n37002 , n37003 , n37004 , n37005 , n37006 , 
     n37007 , n37008 , n37009 , n37010 , n37011 , n37012 , n37013 , n37014 , n37015 , n37016 , 
     n37017 , n37018 , n37019 , n37020 , n37021 , n37022 , n37023 , n37024 , n37025 , n37026 , 
     n37027 , n37028 , n37029 , n37030 , n37031 , n37032 , n37033 , n37034 , n37035 , n37036 , 
     n37037 , n37038 , n37039 , n37040 , n37041 , n37042 , n37043 , n37044 , n37045 , n37046 , 
     n37047 , n37048 , n37049 , n37050 , n37051 , n37052 , n37053 , n37054 , n37055 , n37056 , 
     n37057 , n37058 , n37059 , n37060 , n37061 , n37062 , n37063 , n37064 , n37065 , n37066 , 
     n37067 , n37068 , n37069 , n37070 , n37071 , n37072 , n37073 , n37074 , n37075 , n37076 , 
     n37077 , n37078 , n37079 , n37080 , n37081 , n37082 , n37083 , n37084 , n37085 , n37086 , 
     n37087 , n37088 , n37089 , n37090 , n37091 , n37092 , n37093 , n37094 , n37095 , n37096 , 
     n37097 , n37098 , n37099 , n37100 , n37101 , n37102 , n37103 , n37104 , n37105 , n37106 , 
     n37107 , n37108 , n37109 , n37110 , n37111 , n37112 , n37113 , n37114 , n37115 , n37116 , 
     n37117 , n37118 , n37119 , n37120 , n37121 , n37122 , n37123 , n37124 , n37125 , n37126 , 
     n37127 , n37128 , n37129 , n37130 , n37131 , n37132 , n37133 , n37134 , n37135 , n37136 , 
     n37137 , n37138 , n37139 , n37140 , n37141 , n37142 , n37143 , n37144 , n37145 , n37146 , 
     n37147 , n37148 , n37149 , n37150 , n37151 , n37152 , n37153 , n37154 , n37155 , n37156 , 
     n37157 , n37158 , n37159 , n37160 , n37161 , n37162 , n37163 , n37164 , n37165 , n37166 , 
     n37167 , n37168 , n37169 , n37170 , n37171 , n37172 , n37173 , n37174 , n37175 , n37176 , 
     n37177 , n37178 , n37179 , n37180 , n37181 , n37182 , n37183 , n37184 , n37185 , n37186 , 
     n37187 , n37188 , n37189 , n37190 , n37191 , n37192 , n37193 , n37194 , n37195 , n37196 , 
     n37197 , n37198 , n37199 , n37200 , n37201 , n37202 , n37203 , n37204 , n37205 , n37206 , 
     n37207 , n37208 , n37209 , n37210 , n37211 , n37212 , n37213 , n37214 , n37215 , n37216 , 
     n37217 , n37218 , n37219 , n37220 , n37221 , n37222 , n37223 , n37224 , n37225 , n37226 , 
     n37227 , n37228 , n37229 , n37230 , n37231 , n37232 , n37233 , n37234 , n37235 , n37236 , 
     n37237 , n37238 , n37239 , n37240 , n37241 , n37242 , n37243 , n37244 , n37245 , n37246 , 
     n37247 , n37248 , n37249 , n37250 , n37251 , n37252 , n37253 , n37254 , n37255 , n37256 , 
     n37257 , n37258 , n37259 , n37260 , n37261 , n37262 , n37263 , n37264 , n37265 , n37266 , 
     n37267 , n37268 , n37269 , n37270 , n37271 , n37272 , n37273 , n37274 , n37275 , n37276 , 
     n37277 , n37278 , n37279 , n37280 , n37281 , n37282 , n37283 , n37284 , n37285 , n37286 , 
     n37287 , n37288 , n37289 , n37290 , n37291 , n37292 , n37293 , n37294 , n37295 , n37296 , 
     n37297 , n37298 , n37299 , n37300 , n37301 , n37302 , n37303 , n37304 , n37305 , n37306 , 
     n37307 , n37308 , n37309 , n37310 , n37311 , n37312 , n37313 , n37314 , n37315 , n37316 , 
     n37317 , n37318 , n37319 , n37320 , n37321 , n37322 , n37323 , n37324 , n37325 , n37326 , 
     n37327 , n37328 , n37329 , n37330 , n37331 , n37332 , n37333 , n37334 , n37335 , n37336 , 
     n37337 , n37338 , n37339 , n37340 , n37341 , n37342 , n37343 , n37344 , n37345 , n37346 , 
     n37347 , n37348 , n37349 , n37350 , n37351 , n37352 , n37353 , n37354 , n37355 , n37356 , 
     n37357 , n37358 , n37359 , n37360 , n37361 , n37362 , n37363 , n37364 , n37365 , n37366 , 
     n37367 , n37368 , n37369 , n37370 , n37371 , n37372 , n37373 , n37374 , n37375 , n37376 , 
     n37377 , n37378 , n37379 , n37380 , n37381 , n37382 , n37383 , n37384 , n37385 , n37386 , 
     n37387 , n37388 , n37389 , n37390 , n37391 , n37392 , n37393 , n37394 , n37395 , n37396 , 
     n37397 , n37398 , n37399 , n37400 , n37401 , n37402 , n37403 , n37404 , n37405 , n37406 , 
     n37407 , n37408 , n37409 , n37410 , n37411 , n37412 , n37413 , n37414 , n37415 , n37416 , 
     n37417 , n37418 , n37419 , n37420 , n37421 , n37422 , n37423 , n37424 , n37425 , n37426 , 
     n37427 , n37428 , n37429 , n37430 , n37431 , n37432 , n37433 , n37434 , n37435 , n37436 , 
     n37437 , n37438 , n37439 , n37440 , n37441 , n37442 , n37443 , n37444 , n37445 , n37446 , 
     n37447 , n37448 , n37449 , n37450 , n37451 , n37452 , n37453 , n37454 , n37455 , n37456 , 
     n37457 , n37458 , n37459 , n37460 , n37461 , n37462 , n37463 , n37464 , n37465 , n37466 , 
     n37467 , n37468 , n37469 , n37470 , n37471 , n37472 , n37473 , n37474 , n37475 , n37476 , 
     n37477 , n37478 , n37479 , n37480 , n37481 , n37482 , n37483 , n37484 , n37485 , n37486 , 
     n37487 , n37488 , n37489 , n37490 , n37491 , n37492 , n37493 , n37494 , n37495 , n37496 , 
     n37497 , n37498 , n37499 , n37500 , n37501 , n37502 , n37503 , n37504 , n37505 , n37506 , 
     n37507 , n37508 , n37509 , n37510 , n37511 , n37512 , n37513 , n37514 , n37515 , n37516 , 
     n37517 , n37518 , n37519 , n37520 , n37521 , n37522 , n37523 , n37524 , n37525 , n37526 , 
     n37527 , n37528 , n37529 , n37530 , n37531 , n37532 , n37533 , n37534 , n37535 , n37536 , 
     n37537 , n37538 , n37539 , n37540 , n37541 , n37542 , n37543 , n37544 , n37545 , n37546 , 
     n37547 , n37548 , n37549 , n37550 , n37551 , n37552 , n37553 , n37554 , n37555 , n37556 , 
     n37557 , n37558 , n37559 , n37560 , n37561 , n37562 , n37563 , n37564 , n37565 , n37566 , 
     n37567 , n37568 , n37569 , n37570 , n37571 , n37572 , n37573 , n37574 , n37575 , n37576 , 
     n37577 , n37578 , n37579 , n37580 , n37581 , n37582 , n37583 , n37584 , n37585 , n37586 , 
     n37587 , n37588 , n37589 , n37590 , n37591 , n37592 , n37593 , n37594 , n37595 , n37596 , 
     n37597 , n37598 , n37599 , n37600 , n37601 , n37602 , n37603 , n37604 , n37605 , n37606 , 
     n37607 , n37608 , n37609 , n37610 , n37611 , n37612 , n37613 , n37614 , n37615 , n37616 , 
     n37617 , n37618 , n37619 , n37620 , n37621 , n37622 , n37623 , n37624 , n37625 , n37626 , 
     n37627 , n37628 , n37629 , n37630 , n37631 , n37632 , n37633 , n37634 , n37635 , n37636 , 
     n37637 , n37638 , n37639 , n37640 , n37641 , n37642 , n37643 , n37644 , n37645 , n37646 , 
     n37647 , n37648 , n37649 , n37650 , n37651 , n37652 , n37653 , n37654 , n37655 , n37656 , 
     n37657 , n37658 , n37659 , n37660 , n37661 , n37662 , n37663 , n37664 , n37665 , n37666 , 
     n37667 , n37668 , n37669 , n37670 , n37671 , n37672 , n37673 , n37674 , n37675 , n37676 , 
     n37677 , n37678 , n37679 , n37680 , n37681 , n37682 , n37683 , n37684 , n37685 , n37686 , 
     n37687 , n37688 , n37689 , n37690 , n37691 , n37692 , n37693 , n37694 , n37695 , n37696 , 
     n37697 , n37698 , n37699 , n37700 , n37701 , n37702 , n37703 , n37704 , n37705 , n37706 , 
     n37707 , n37708 , n37709 , n37710 , n37711 , n37712 , n37713 , n37714 , n37715 , n37716 , 
     n37717 , n37718 , n37719 , n37720 , n37721 , n37722 , n37723 , n37724 , n37725 , n37726 , 
     n37727 , n37728 , n37729 , n37730 , n37731 , n37732 , n37733 , n37734 , n37735 , n37736 , 
     n37737 , n37738 , n37739 , n37740 , n37741 , n37742 , n37743 , n37744 , n37745 , n37746 , 
     n37747 , n37748 , n37749 , n37750 , n37751 , n37752 , n37753 , n37754 , n37755 , n37756 , 
     n37757 , n37758 , n37759 , n37760 , n37761 , n37762 , n37763 , n37764 , n37765 , n37766 , 
     n37767 , n37768 , n37769 , n37770 , n37771 , n37772 , n37773 , n37774 , n37775 , n37776 , 
     n37777 , n37778 , n37779 , n37780 , n37781 , n37782 , n37783 , n37784 , n37785 , n37786 , 
     n37787 , n37788 , n37789 , n37790 , n37791 , n37792 , n37793 , n37794 , n37795 , n37796 , 
     n37797 , n37798 , n37799 , n37800 , n37801 , n37802 , n37803 , n37804 , n37805 , n37806 , 
     n37807 , n37808 , n37809 , n37810 , n37811 , n37812 , n37813 , n37814 , n37815 , n37816 , 
     n37817 , n37818 , n37819 , n37820 , n37821 , n37822 , n37823 , n37824 , n37825 , n37826 , 
     n37827 , n37828 , n37829 , n37830 , n37831 , n37832 , n37833 , n37834 , n37835 , n37836 , 
     n37837 , n37838 , n37839 , n37840 , n37841 , n37842 , n37843 , n37844 , n37845 , n37846 , 
     n37847 , n37848 , n37849 , n37850 , n37851 , n37852 , n37853 , n37854 , n37855 , n37856 , 
     n37857 , n37858 , n37859 , n37860 , n37861 , n37862 , n37863 , n37864 , n37865 , n37866 , 
     n37867 , n37868 , n37869 , n37870 , n37871 , n37872 , n37873 , n37874 , n37875 , n37876 , 
     n37877 , n37878 , n37879 , n37880 , n37881 , n37882 , n37883 , n37884 , n37885 , n37886 , 
     n37887 , n37888 , n37889 , n37890 , n37891 , n37892 , n37893 , n37894 , n37895 , n37896 , 
     n37897 , n37898 , n37899 , n37900 , n37901 , n37902 , n37903 , n37904 , n37905 , n37906 , 
     n37907 , n37908 , n37909 , n37910 , n37911 , n37912 , n37913 , n37914 , n37915 , n37916 , 
     n37917 , n37918 , n37919 , n37920 , n37921 , n37922 , n37923 , n37924 , n37925 , n37926 , 
     n37927 , n37928 , n37929 , n37930 , n37931 , n37932 , n37933 , n37934 , n37935 , n37936 , 
     n37937 , n37938 , n37939 , n37940 , n37941 , n37942 , n37943 , n37944 , n37945 , n37946 , 
     n37947 , n37948 , n37949 , n37950 , n37951 , n37952 , n37953 , n37954 , n37955 , n37956 , 
     n37957 , n37958 , n37959 , n37960 , n37961 , n37962 , n37963 , n37964 , n37965 , n37966 , 
     n37967 , n37968 , n37969 , n37970 , n37971 , n37972 , n37973 , n37974 , n37975 , n37976 , 
     n37977 , n37978 , n37979 , n37980 , n37981 , n37982 , n37983 , n37984 , n37985 , n37986 , 
     n37987 , n37988 , n37989 , n37990 , n37991 , n37992 , n37993 , n37994 , n37995 , n37996 , 
     n37997 , n37998 , n37999 , n38000 , n38001 , n38002 , n38003 , n38004 , n38005 , n38006 , 
     n38007 , n38008 , n38009 , n38010 , n38011 , n38012 , n38013 , n38014 , n38015 , n38016 , 
     n38017 , n38018 , n38019 , n38020 , n38021 , n38022 , n38023 , n38024 , n38025 , n38026 , 
     n38027 , n38028 , n38029 , n38030 , n38031 , n38032 , n38033 , n38034 , n38035 , n38036 , 
     n38037 , n38038 , n38039 , n38040 , n38041 , n38042 , n38043 , n38044 , n38045 , n38046 , 
     n38047 , n38048 , n38049 , n38050 , n38051 , n38052 , n38053 , n38054 , n38055 , n38056 , 
     n38057 , n38058 , n38059 , n38060 , n38061 , n38062 , n38063 , n38064 , n38065 , n38066 , 
     n38067 , n38068 , n38069 , n38070 , n38071 , n38072 , n38073 , n38074 , n38075 , n38076 , 
     n38077 , n38078 , n38079 , n38080 , n38081 , n38082 , n38083 , n38084 , n38085 , n38086 , 
     n38087 , n38088 , n38089 , n38090 , n38091 , n38092 , n38093 , n38094 , n38095 , n38096 , 
     n38097 , n38098 , n38099 , n38100 , n38101 , n38102 , n38103 , n38104 , n38105 , n38106 , 
     n38107 , n38108 , n38109 , n38110 , n38111 , n38112 , n38113 , n38114 , n38115 , n38116 , 
     n38117 , n38118 , n38119 , n38120 , n38121 , n38122 , n38123 , n38124 , n38125 , n38126 , 
     n38127 , n38128 , n38129 , n38130 , n38131 , n38132 , n38133 , n38134 , n38135 , n38136 , 
     n38137 , n38138 , n38139 , n38140 , n38141 , n38142 , n38143 , n38144 , n38145 , n38146 , 
     n38147 , n38148 , n38149 , n38150 , n38151 , n38152 , n38153 , n38154 , n38155 , n38156 , 
     n38157 , n38158 , n38159 , n38160 , n38161 , n38162 , n38163 , n38164 , n38165 , n38166 , 
     n38167 , n38168 , n38169 , n38170 , n38171 , n38172 , n38173 , n38174 , n38175 , n38176 , 
     n38177 , n38178 , n38179 , n38180 , n38181 , n38182 , n38183 , n38184 , n38185 , n38186 , 
     n38187 , n38188 , n38189 , n38190 , n38191 , n38192 , n38193 , n38194 , n38195 , n38196 , 
     n38197 , n38198 , n38199 , n38200 , n38201 , n38202 , n38203 , n38204 , n38205 , n38206 , 
     n38207 , n38208 , n38209 , n38210 , n38211 , n38212 , n38213 , n38214 , n38215 , n38216 , 
     n38217 , n38218 , n38219 , n38220 , n38221 , n38222 , n38223 , n38224 , n38225 , n38226 , 
     n38227 , n38228 , n38229 , n38230 , n38231 , n38232 , n38233 , n38234 , n38235 , n38236 , 
     n38237 , n38238 , n38239 , n38240 , n38241 , n38242 , n38243 , n38244 , n38245 , n38246 , 
     n38247 , n38248 , n38249 , n38250 , n38251 , n38252 , n38253 , n38254 , n38255 , n38256 , 
     n38257 , n38258 , n38259 , n38260 , n38261 , n38262 , n38263 , n38264 , n38265 , n38266 , 
     n38267 , n38268 , n38269 , n38270 , n38271 , n38272 , n38273 , n38274 , n38275 , n38276 , 
     n38277 , n38278 , n38279 , n38280 , n38281 , n38282 , n38283 , n38284 , n38285 , n38286 , 
     n38287 , n38288 , n38289 , n38290 , n38291 , n38292 , n38293 , n38294 , n38295 , n38296 , 
     n38297 , n38298 , n38299 , n38300 , n38301 , n38302 , n38303 , n38304 , n38305 , n38306 , 
     n38307 , n38308 , n38309 , n38310 , n38311 , n38312 , n38313 , n38314 , n38315 , n38316 , 
     n38317 , n38318 , n38319 , n38320 , n38321 , n38322 , n38323 , n38324 , n38325 , n38326 , 
     n38327 , n38328 , n38329 , n38330 , n38331 , n38332 , n38333 , n38334 , n38335 , n38336 , 
     n38337 , n38338 , n38339 , n38340 , n38341 , n38342 , n38343 , n38344 , n38345 , n38346 , 
     n38347 , n38348 , n38349 , n38350 , n38351 , n38352 , n38353 , n38354 , n38355 , n38356 , 
     n38357 , n38358 , n38359 , n38360 , n38361 , n38362 , n38363 , n38364 , n38365 , n38366 , 
     n38367 , n38368 , n38369 , n38370 , n38371 , n38372 , n38373 , n38374 , n38375 , n38376 , 
     n38377 , n38378 , n38379 , n38380 , n38381 , n38382 , n38383 , n38384 , n38385 , n38386 , 
     n38387 , n38388 , n38389 , n38390 , n38391 , n38392 , n38393 , n38394 , n38395 , n38396 , 
     n38397 , n38398 , n38399 , n38400 , n38401 , n38402 , n38403 , n38404 , n38405 , n38406 , 
     n38407 , n38408 , n38409 , n38410 , n38411 , n38412 , n38413 , n38414 , n38415 , n38416 , 
     n38417 , n38418 , n38419 , n38420 , n38421 , n38422 , n38423 , n38424 , n38425 , n38426 , 
     n38427 , n38428 , n38429 , n38430 , n38431 , n38432 , n38433 , n38434 , n38435 , n38436 , 
     n38437 , n38438 , n38439 , n38440 , n38441 , n38442 , n38443 , n38444 , n38445 , n38446 , 
     n38447 , n38448 , n38449 , n38450 , n38451 , n38452 , n38453 , n38454 , n38455 , n38456 , 
     n38457 , n38458 , n38459 , n38460 , n38461 , n38462 , n38463 , n38464 , n38465 , n38466 , 
     n38467 , n38468 , n38469 , n38470 , n38471 , n38472 , n38473 , n38474 , n38475 , n38476 , 
     n38477 , n38478 , n38479 , n38480 , n38481 , n38482 , n38483 , n38484 , n38485 , n38486 , 
     n38487 , n38488 , n38489 , n38490 , n38491 , n38492 , n38493 , n38494 , n38495 , n38496 , 
     n38497 , n38498 , n38499 , n38500 , n38501 , n38502 , n38503 , n38504 , n38505 , n38506 , 
     n38507 , n38508 , n38509 , n38510 , n38511 , n38512 , n38513 , n38514 , n38515 , n38516 , 
     n38517 , n38518 , n38519 , n38520 , n38521 , n38522 , n38523 , n38524 , n38525 , n38526 , 
     n38527 , n38528 , n38529 , n38530 , n38531 , n38532 , n38533 , n38534 , n38535 , n38536 , 
     n38537 , n38538 , n38539 , n38540 , n38541 , n38542 , n38543 , n38544 , n38545 , n38546 , 
     n38547 , n38548 , n38549 , n38550 , n38551 , n38552 , n38553 , n38554 , n38555 , n38556 , 
     n38557 , n38558 , n38559 , n38560 , n38561 , n38562 , n38563 , n38564 , n38565 , n38566 , 
     n38567 , n38568 , n38569 , n38570 , n38571 , n38572 , n38573 , n38574 , n38575 , n38576 , 
     n38577 , n38578 , n38579 , n38580 , n38581 , n38582 , n38583 , n38584 , n38585 , n38586 , 
     n38587 , n38588 , n38589 , n38590 , n38591 , n38592 , n38593 , n38594 , n38595 , n38596 , 
     n38597 , n38598 , n38599 , n38600 , n38601 , n38602 , n38603 , n38604 , n38605 , n38606 , 
     n38607 , n38608 , n38609 , n38610 , n38611 , n38612 , n38613 , n38614 , n38615 , n38616 , 
     n38617 , n38618 , n38619 , n38620 , n38621 , n38622 , n38623 , n38624 , n38625 , n38626 , 
     n38627 , n38628 , n38629 , n38630 , n38631 , n38632 , n38633 , n38634 , n38635 , n38636 , 
     n38637 , n38638 , n38639 , n38640 , n38641 , n38642 , n38643 , n38644 , n38645 , n38646 , 
     n38647 , n38648 , n38649 , n38650 , n38651 , n38652 , n38653 , n38654 , n38655 , n38656 , 
     n38657 , n38658 , n38659 , n38660 , n38661 , n38662 , n38663 , n38664 , n38665 , n38666 , 
     n38667 , n38668 , n38669 , n38670 , n38671 , n38672 , n38673 , n38674 , n38675 , n38676 , 
     n38677 , n38678 , n38679 , n38680 , n38681 , n38682 , n38683 , n38684 , n38685 , n38686 , 
     n38687 , n38688 , n38689 , n38690 , n38691 , n38692 , n38693 , n38694 , n38695 , n38696 , 
     n38697 , n38698 , n38699 , n38700 , n38701 , n38702 , n38703 , n38704 , n38705 , n38706 , 
     n38707 , n38708 , n38709 , n38710 , n38711 , n38712 , n38713 , n38714 , n38715 , n38716 , 
     n38717 , n38718 , n38719 , n38720 , n38721 , n38722 , n38723 , n38724 , n38725 , n38726 , 
     n38727 , n38728 , n38729 , n38730 , n38731 , n38732 , n38733 , n38734 , n38735 , n38736 , 
     n38737 , n38738 , n38739 , n38740 , n38741 , n38742 , n38743 , n38744 , n38745 , n38746 , 
     n38747 , n38748 , n38749 , n38750 , n38751 , n38752 , n38753 , n38754 , n38755 , n38756 , 
     n38757 , n38758 , n38759 , n38760 , n38761 , n38762 , n38763 , n38764 , n38765 , n38766 , 
     n38767 , n38768 , n38769 , n38770 , n38771 , n38772 , n38773 , n38774 , n38775 , n38776 , 
     n38777 , n38778 , n38779 , n38780 , n38781 , n38782 , n38783 , n38784 , n38785 , n38786 , 
     n38787 , n38788 , n38789 , n38790 , n38791 , n38792 , n38793 , n38794 , n38795 , n38796 , 
     n38797 , n38798 , n38799 , n38800 , n38801 , n38802 , n38803 , n38804 , n38805 , n38806 , 
     n38807 , n38808 , n38809 , n38810 , n38811 , n38812 , n38813 , n38814 , n38815 , n38816 , 
     n38817 , n38818 , n38819 , n38820 , n38821 , n38822 , n38823 , n38824 , n38825 , n38826 , 
     n38827 , n38828 , n38829 , n38830 , n38831 , n38832 , n38833 , n38834 , n38835 , n38836 , 
     n38837 , n38838 , n38839 , n38840 , n38841 , n38842 , n38843 , n38844 , n38845 , n38846 , 
     n38847 , n38848 , n38849 , n38850 , n38851 , n38852 , n38853 , n38854 , n38855 , n38856 , 
     n38857 , n38858 , n38859 , n38860 , n38861 , n38862 , n38863 , n38864 , n38865 , n38866 , 
     n38867 , n38868 , n38869 , n38870 , n38871 , n38872 , n38873 , n38874 , n38875 , n38876 , 
     n38877 , n38878 , n38879 , n38880 , n38881 , n38882 , n38883 , n38884 , n38885 , n38886 , 
     n38887 , n38888 , n38889 , n38890 , n38891 , n38892 , n38893 , n38894 , n38895 , n38896 , 
     n38897 , n38898 , n38899 , n38900 , n38901 , n38902 , n38903 , n38904 , n38905 , n38906 , 
     n38907 , n38908 , n38909 , n38910 , n38911 , n38912 , n38913 , n38914 , n38915 , n38916 , 
     n38917 , n38918 , n38919 , n38920 , n38921 , n38922 , n38923 , n38924 , n38925 , n38926 , 
     n38927 , n38928 , n38929 , n38930 , n38931 , n38932 , n38933 , n38934 , n38935 , n38936 , 
     n38937 , n38938 , n38939 , n38940 , n38941 , n38942 , n38943 , n38944 , n38945 , n38946 , 
     n38947 , n38948 , n38949 , n38950 , n38951 , n38952 , n38953 , n38954 , n38955 , n38956 , 
     n38957 , n38958 , n38959 , n38960 , n38961 , n38962 , n38963 , n38964 , n38965 , n38966 , 
     n38967 , n38968 , n38969 , n38970 , n38971 , n38972 , n38973 , n38974 , n38975 , n38976 , 
     n38977 , n38978 , n38979 , n38980 , n38981 , n38982 , n38983 , n38984 , n38985 , n38986 , 
     n38987 , n38988 , n38989 , n38990 , n38991 , n38992 , n38993 , n38994 , n38995 , n38996 , 
     n38997 , n38998 , n38999 , n39000 , n39001 , n39002 , n39003 , n39004 , n39005 , n39006 , 
     n39007 , n39008 , n39009 , n39010 , n39011 , n39012 , n39013 , n39014 , n39015 , n39016 , 
     n39017 , n39018 , n39019 , n39020 , n39021 , n39022 , n39023 , n39024 , n39025 , n39026 , 
     n39027 , n39028 , n39029 , n39030 , n39031 , n39032 , n39033 , n39034 , n39035 , n39036 , 
     n39037 , n39038 , n39039 , n39040 , n39041 , n39042 , n39043 , n39044 , n39045 , n39046 , 
     n39047 , n39048 , n39049 , n39050 , n39051 , n39052 , n39053 , n39054 , n39055 , n39056 , 
     n39057 , n39058 , n39059 , n39060 , n39061 , n39062 , n39063 , n39064 , n39065 , n39066 , 
     n39067 , n39068 , n39069 , n39070 , n39071 , n39072 , n39073 , n39074 , n39075 , n39076 , 
     n39077 , n39078 , n39079 , n39080 , n39081 , n39082 , n39083 , n39084 , n39085 , n39086 , 
     n39087 , n39088 , n39089 , n39090 , n39091 , n39092 , n39093 , n39094 , n39095 , n39096 , 
     n39097 , n39098 , n39099 , n39100 , n39101 , n39102 , n39103 , n39104 , n39105 , n39106 , 
     n39107 , n39108 , n39109 , n39110 , n39111 , n39112 , n39113 , n39114 , n39115 , n39116 , 
     n39117 , n39118 , n39119 , n39120 , n39121 , n39122 , n39123 , n39124 , n39125 , n39126 , 
     n39127 , n39128 , n39129 , n39130 , n39131 , n39132 , n39133 , n39134 , n39135 , n39136 , 
     n39137 , n39138 , n39139 , n39140 , n39141 , n39142 , n39143 , n39144 , n39145 , n39146 , 
     n39147 , n39148 , n39149 , n39150 , n39151 , n39152 , n39153 , n39154 , n39155 , n39156 , 
     n39157 , n39158 , n39159 , n39160 , n39161 , n39162 , n39163 , n39164 , n39165 , n39166 , 
     n39167 , n39168 , n39169 , n39170 , n39171 , n39172 , n39173 , n39174 , n39175 , n39176 , 
     n39177 , n39178 , n39179 , n39180 , n39181 , n39182 , n39183 , n39184 , n39185 , n39186 , 
     n39187 , n39188 , n39189 , n39190 , n39191 , n39192 , n39193 , n39194 , n39195 , n39196 , 
     n39197 , n39198 , n39199 , n39200 , n39201 , n39202 , n39203 , n39204 , n39205 , n39206 , 
     n39207 , n39208 , n39209 , n39210 , n39211 , n39212 , n39213 , n39214 , n39215 , n39216 , 
     n39217 , n39218 , n39219 , n39220 , n39221 , n39222 , n39223 , n39224 , n39225 , n39226 , 
     n39227 , n39228 , n39229 , n39230 , n39231 , n39232 , n39233 , n39234 , n39235 , n39236 , 
     n39237 , n39238 , n39239 , n39240 , n39241 , n39242 , n39243 , n39244 , n39245 , n39246 , 
     n39247 , n39248 , n39249 , n39250 , n39251 , n39252 , n39253 , n39254 , n39255 , n39256 , 
     n39257 , n39258 , n39259 , n39260 , n39261 , n39262 , n39263 , n39264 , n39265 , n39266 , 
     n39267 , n39268 , n39269 , n39270 , n39271 , n39272 , n39273 , n39274 , n39275 , n39276 , 
     n39277 , n39278 , n39279 , n39280 , n39281 , n39282 , n39283 , n39284 , n39285 , n39286 , 
     n39287 , n39288 , n39289 , n39290 , n39291 , n39292 , n39293 , n39294 , n39295 , n39296 , 
     n39297 , n39298 , n39299 , n39300 , n39301 , n39302 , n39303 , n39304 , n39305 , n39306 , 
     n39307 , n39308 , n39309 , n39310 , n39311 , n39312 , n39313 , n39314 , n39315 , n39316 , 
     n39317 , n39318 , n39319 , n39320 , n39321 , n39322 , n39323 , n39324 , n39325 , n39326 , 
     n39327 , n39328 , n39329 , n39330 , n39331 , n39332 , n39333 , n39334 , n39335 , n39336 , 
     n39337 , n39338 , n39339 , n39340 , n39341 , n39342 , n39343 , n39344 , n39345 , n39346 , 
     n39347 , n39348 , n39349 , n39350 , n39351 , n39352 , n39353 , n39354 , n39355 , n39356 , 
     n39357 , n39358 , n39359 , n39360 , n39361 , n39362 , n39363 , n39364 , n39365 , n39366 , 
     n39367 , n39368 , n39369 , n39370 , n39371 , n39372 , n39373 , n39374 , n39375 , n39376 , 
     n39377 , n39378 , n39379 , n39380 , n39381 , n39382 , n39383 , n39384 , n39385 , n39386 , 
     n39387 , n39388 , n39389 , n39390 , n39391 , n39392 , n39393 , n39394 , n39395 , n39396 , 
     n39397 , n39398 , n39399 , n39400 , n39401 , n39402 , n39403 , n39404 , n39405 , n39406 , 
     n39407 , n39408 , n39409 , n39410 , n39411 , n39412 , n39413 , n39414 , n39415 , n39416 , 
     n39417 , n39418 , n39419 , n39420 , n39421 , n39422 , n39423 , n39424 , n39425 , n39426 , 
     n39427 , n39428 , n39429 , n39430 , n39431 , n39432 , n39433 , n39434 , n39435 , n39436 , 
     n39437 , n39438 , n39439 , n39440 , n39441 , n39442 , n39443 , n39444 , n39445 , n39446 , 
     n39447 , n39448 , n39449 , n39450 , n39451 , n39452 , n39453 , n39454 , n39455 , n39456 , 
     n39457 , n39458 , n39459 , n39460 , n39461 , n39462 , n39463 , n39464 , n39465 , n39466 , 
     n39467 , n39468 , n39469 , n39470 , n39471 , n39472 , n39473 , n39474 , n39475 , n39476 , 
     n39477 , n39478 , n39479 , n39480 , n39481 , n39482 , n39483 , n39484 , n39485 , n39486 , 
     n39487 , n39488 , n39489 , n39490 , n39491 , n39492 , n39493 , n39494 , n39495 , n39496 , 
     n39497 , n39498 , n39499 , n39500 , n39501 , n39502 , n39503 , n39504 , n39505 , n39506 , 
     n39507 , n39508 , n39509 , n39510 , n39511 , n39512 , n39513 , n39514 , n39515 , n39516 , 
     n39517 , n39518 , n39519 , n39520 , n39521 , n39522 , n39523 , n39524 , n39525 , n39526 , 
     n39527 , n39528 , n39529 , n39530 , n39531 , n39532 , n39533 , n39534 , n39535 , n39536 , 
     n39537 , n39538 , n39539 , n39540 , n39541 , n39542 , n39543 , n39544 , n39545 , n39546 , 
     n39547 , n39548 , n39549 , n39550 , n39551 , n39552 , n39553 , n39554 , n39555 , n39556 , 
     n39557 , n39558 , n39559 , n39560 , n39561 , n39562 , n39563 , n39564 , n39565 , n39566 , 
     n39567 , n39568 , n39569 , n39570 , n39571 , n39572 , n39573 , n39574 , n39575 , n39576 , 
     n39577 , n39578 , n39579 , n39580 , n39581 , n39582 , n39583 , n39584 , n39585 , n39586 , 
     n39587 , n39588 , n39589 , n39590 , n39591 , n39592 , n39593 , n39594 , n39595 , n39596 , 
     n39597 , n39598 , n39599 , n39600 , n39601 , n39602 , n39603 , n39604 , n39605 , n39606 , 
     n39607 , n39608 , n39609 , n39610 , n39611 , n39612 , n39613 , n39614 , n39615 , n39616 , 
     n39617 , n39618 , n39619 , n39620 , n39621 , n39622 , n39623 , n39624 , n39625 , n39626 , 
     n39627 , n39628 , n39629 , n39630 , n39631 , n39632 , n39633 , n39634 , n39635 , n39636 , 
     n39637 , n39638 , n39639 , n39640 , n39641 , n39642 , n39643 , n39644 , n39645 , n39646 , 
     n39647 , n39648 , n39649 , n39650 , n39651 , n39652 , n39653 , n39654 , n39655 , n39656 , 
     n39657 , n39658 , n39659 , n39660 , n39661 , n39662 , n39663 , n39664 , n39665 , n39666 , 
     n39667 , n39668 , n39669 , n39670 , n39671 , n39672 , n39673 , n39674 , n39675 , n39676 , 
     n39677 , n39678 , n39679 , n39680 , n39681 , n39682 , n39683 , n39684 , n39685 , n39686 , 
     n39687 , n39688 , n39689 , n39690 , n39691 , n39692 , n39693 , n39694 , n39695 , n39696 , 
     n39697 , n39698 , n39699 , n39700 , n39701 , n39702 , n39703 , n39704 , n39705 , n39706 , 
     n39707 , n39708 , n39709 , n39710 , n39711 , n39712 , n39713 , n39714 , n39715 , n39716 , 
     n39717 , n39718 , n39719 , n39720 , n39721 , n39722 , n39723 , n39724 , n39725 , n39726 , 
     n39727 , n39728 , n39729 , n39730 , n39731 , n39732 , n39733 , n39734 , n39735 , n39736 , 
     n39737 , n39738 , n39739 , n39740 , n39741 , n39742 , n39743 , n39744 , n39745 , n39746 , 
     n39747 , n39748 , n39749 , n39750 , n39751 , n39752 , n39753 , n39754 , n39755 , n39756 , 
     n39757 , n39758 , n39759 , n39760 , n39761 , n39762 , n39763 , n39764 , n39765 , n39766 , 
     n39767 , n39768 , n39769 , n39770 , n39771 , n39772 , n39773 , n39774 , n39775 , n39776 , 
     n39777 , n39778 , n39779 , n39780 , n39781 , n39782 , n39783 , n39784 , n39785 , n39786 , 
     n39787 , n39788 , n39789 , n39790 , n39791 , n39792 , n39793 , n39794 , n39795 , n39796 , 
     n39797 , n39798 , n39799 , n39800 , n39801 , n39802 , n39803 , n39804 , n39805 , n39806 , 
     n39807 , n39808 , n39809 , n39810 , n39811 , n39812 , n39813 , n39814 , n39815 , n39816 , 
     n39817 , n39818 , n39819 , n39820 , n39821 , n39822 , n39823 , n39824 , n39825 , n39826 , 
     n39827 , n39828 , n39829 , n39830 , n39831 , n39832 , n39833 , n39834 , n39835 , n39836 , 
     n39837 , n39838 , n39839 , n39840 , n39841 , n39842 , n39843 , n39844 , n39845 , n39846 , 
     n39847 , n39848 , n39849 , n39850 , n39851 , n39852 , n39853 , n39854 , n39855 , n39856 , 
     n39857 , n39858 , n39859 , n39860 , n39861 , n39862 , n39863 , n39864 , n39865 , n39866 , 
     n39867 , n39868 , n39869 , n39870 , n39871 , n39872 , n39873 , n39874 , n39875 , n39876 , 
     n39877 , n39878 , n39879 , n39880 , n39881 , n39882 , n39883 , n39884 , n39885 , n39886 , 
     n39887 , n39888 , n39889 , n39890 , n39891 , n39892 , n39893 , n39894 , n39895 , n39896 , 
     n39897 , n39898 , n39899 , n39900 , n39901 , n39902 , n39903 , n39904 , n39905 , n39906 , 
     n39907 , n39908 , n39909 , n39910 , n39911 , n39912 , n39913 , n39914 , n39915 , n39916 , 
     n39917 , n39918 , n39919 , n39920 , n39921 , n39922 , n39923 , n39924 , n39925 , n39926 , 
     n39927 , n39928 , n39929 , n39930 , n39931 , n39932 , n39933 , n39934 , n39935 , n39936 , 
     n39937 , n39938 , n39939 , n39940 , n39941 , n39942 , n39943 , n39944 , n39945 , n39946 , 
     n39947 , n39948 , n39949 , n39950 , n39951 , n39952 , n39953 , n39954 , n39955 , n39956 , 
     n39957 , n39958 , n39959 , n39960 , n39961 , n39962 , n39963 , n39964 , n39965 , n39966 , 
     n39967 , n39968 , n39969 , n39970 , n39971 , n39972 , n39973 , n39974 , n39975 , n39976 , 
     n39977 , n39978 , n39979 , n39980 , n39981 , n39982 , n39983 , n39984 , n39985 , n39986 , 
     n39987 , n39988 , n39989 , n39990 , n39991 , n39992 , n39993 , n39994 , n39995 , n39996 , 
     n39997 , n39998 , n39999 , n40000 , n40001 , n40002 , n40003 , n40004 , n40005 , n40006 , 
     n40007 , n40008 , n40009 , n40010 , n40011 , n40012 , n40013 , n40014 , n40015 , n40016 , 
     n40017 , n40018 , n40019 , n40020 , n40021 , n40022 , n40023 , n40024 , n40025 , n40026 , 
     n40027 , n40028 , n40029 , n40030 , n40031 , n40032 , n40033 , n40034 , n40035 , n40036 , 
     n40037 , n40038 , n40039 , n40040 , n40041 , n40042 , n40043 , n40044 , n40045 , n40046 , 
     n40047 , n40048 , n40049 , n40050 , n40051 , n40052 , n40053 , n40054 , n40055 , n40056 , 
     n40057 , n40058 , n40059 , n40060 , n40061 , n40062 , n40063 , n40064 , n40065 , n40066 , 
     n40067 , n40068 , n40069 , n40070 , n40071 , n40072 , n40073 , n40074 , n40075 , n40076 , 
     n40077 , n40078 , n40079 , n40080 , n40081 , n40082 , n40083 , n40084 , n40085 , n40086 , 
     n40087 , n40088 , n40089 , n40090 , n40091 , n40092 , n40093 , n40094 , n40095 , n40096 , 
     n40097 , n40098 , n40099 , n40100 , n40101 , n40102 , n40103 , n40104 , n40105 , n40106 , 
     n40107 , n40108 , n40109 , n40110 , n40111 , n40112 , n40113 , n40114 , n40115 , n40116 , 
     n40117 , n40118 , n40119 , n40120 , n40121 , n40122 , n40123 , n40124 , n40125 , n40126 , 
     n40127 , n40128 , n40129 , n40130 , n40131 , n40132 , n40133 , n40134 , n40135 , n40136 , 
     n40137 , n40138 , n40139 , n40140 , n40141 , n40142 , n40143 , n40144 , n40145 , n40146 , 
     n40147 , n40148 , n40149 , n40150 , n40151 , n40152 , n40153 , n40154 , n40155 , n40156 , 
     n40157 , n40158 , n40159 , n40160 , n40161 , n40162 , n40163 , n40164 , n40165 , n40166 , 
     n40167 , n40168 , n40169 , n40170 , n40171 , n40172 , n40173 , n40174 , n40175 , n40176 , 
     n40177 , n40178 , n40179 , n40180 , n40181 , n40182 , n40183 , n40184 , n40185 , n40186 , 
     n40187 , n40188 , n40189 , n40190 , n40191 , n40192 , n40193 , n40194 , n40195 , n40196 , 
     n40197 , n40198 , n40199 , n40200 , n40201 , n40202 , n40203 , n40204 , n40205 , n40206 , 
     n40207 , n40208 , n40209 , n40210 , n40211 , n40212 , n40213 , n40214 , n40215 , n40216 , 
     n40217 , n40218 , n40219 , n40220 , n40221 , n40222 , n40223 , n40224 , n40225 , n40226 , 
     n40227 , n40228 , n40229 , n40230 , n40231 , n40232 , n40233 , n40234 , n40235 , n40236 , 
     n40237 , n40238 , n40239 , n40240 , n40241 , n40242 , n40243 , n40244 , n40245 , n40246 , 
     n40247 , n40248 , n40249 , n40250 , n40251 , n40252 , n40253 , n40254 , n40255 , n40256 , 
     n40257 , n40258 , n40259 , n40260 , n40261 , n40262 , n40263 , n40264 , n40265 , n40266 , 
     n40267 , n40268 , n40269 , n40270 , n40271 , n40272 , n40273 , n40274 , n40275 , n40276 , 
     n40277 , n40278 , n40279 , n40280 , n40281 , n40282 , n40283 , n40284 , n40285 , n40286 , 
     n40287 , n40288 , n40289 , n40290 , n40291 , n40292 , n40293 , n40294 , n40295 , n40296 , 
     n40297 , n40298 , n40299 , n40300 , n40301 , n40302 , n40303 , n40304 , n40305 , n40306 , 
     n40307 , n40308 , n40309 , n40310 , n40311 , n40312 , n40313 , n40314 , n40315 , n40316 , 
     n40317 , n40318 , n40319 , n40320 , n40321 , n40322 , n40323 , n40324 , n40325 , n40326 , 
     n40327 , n40328 , n40329 , n40330 , n40331 , n40332 , n40333 , n40334 , n40335 , n40336 , 
     n40337 , n40338 , n40339 , n40340 , n40341 , n40342 , n40343 , n40344 , n40345 , n40346 , 
     n40347 , n40348 , n40349 , n40350 , n40351 , n40352 , n40353 , n40354 , n40355 , n40356 , 
     n40357 , n40358 , n40359 , n40360 , n40361 , n40362 , n40363 , n40364 , n40365 , n40366 , 
     n40367 , n40368 , n40369 , n40370 , n40371 , n40372 , n40373 , n40374 , n40375 , n40376 , 
     n40377 , n40378 , n40379 , n40380 , n40381 , n40382 , n40383 , n40384 , n40385 , n40386 , 
     n40387 , n40388 , n40389 , n40390 , n40391 , n40392 , n40393 , n40394 , n40395 , n40396 , 
     n40397 , n40398 , n40399 , n40400 , n40401 , n40402 , n40403 , n40404 , n40405 , n40406 , 
     n40407 , n40408 , n40409 , n40410 , n40411 , n40412 , n40413 , n40414 , n40415 , n40416 , 
     n40417 , n40418 , n40419 , n40420 , n40421 , n40422 , n40423 , n40424 , n40425 , n40426 , 
     n40427 , n40428 , n40429 , n40430 , n40431 , n40432 , n40433 , n40434 , n40435 , n40436 , 
     n40437 , n40438 , n40439 , n40440 , n40441 , n40442 , n40443 , n40444 , n40445 , n40446 , 
     n40447 , n40448 , n40449 , n40450 , n40451 , n40452 , n40453 , n40454 , n40455 , n40456 , 
     n40457 , n40458 , n40459 , n40460 , n40461 , n40462 , n40463 , n40464 , n40465 , n40466 , 
     n40467 , n40468 , n40469 , n40470 , n40471 , n40472 , n40473 , n40474 , n40475 , n40476 , 
     n40477 , n40478 , n40479 , n40480 , n40481 , n40482 , n40483 , n40484 , n40485 , n40486 , 
     n40487 , n40488 , n40489 , n40490 , n40491 , n40492 , n40493 , n40494 , n40495 , n40496 , 
     n40497 , n40498 , n40499 , n40500 , n40501 , n40502 , n40503 , n40504 , n40505 , n40506 , 
     n40507 , n40508 , n40509 , n40510 , n40511 , n40512 , n40513 , n40514 , n40515 , n40516 , 
     n40517 , n40518 , n40519 , n40520 , n40521 , n40522 , n40523 , n40524 , n40525 , n40526 , 
     n40527 , n40528 , n40529 , n40530 , n40531 , n40532 , n40533 , n40534 , n40535 , n40536 , 
     n40537 , n40538 , n40539 , n40540 , n40541 , n40542 , n40543 , n40544 , n40545 , n40546 , 
     n40547 , n40548 , n40549 , n40550 , n40551 , n40552 , n40553 , n40554 , n40555 , n40556 , 
     n40557 , n40558 , n40559 , n40560 , n40561 , n40562 , n40563 , n40564 , n40565 , n40566 , 
     n40567 , n40568 , n40569 , n40570 , n40571 , n40572 , n40573 , n40574 , n40575 , n40576 , 
     n40577 , n40578 , n40579 , n40580 , n40581 , n40582 , n40583 , n40584 , n40585 , n40586 , 
     n40587 , n40588 , n40589 , n40590 , n40591 , n40592 , n40593 , n40594 , n40595 , n40596 , 
     n40597 , n40598 , n40599 , n40600 , n40601 , n40602 , n40603 , n40604 , n40605 , n40606 , 
     n40607 , n40608 , n40609 , n40610 , n40611 , n40612 , n40613 , n40614 , n40615 , n40616 , 
     n40617 , n40618 , n40619 , n40620 , n40621 , n40622 , n40623 , n40624 , n40625 , n40626 , 
     n40627 , n40628 , n40629 , n40630 , n40631 , n40632 , n40633 , n40634 , n40635 , n40636 , 
     n40637 , n40638 , n40639 , n40640 , n40641 , n40642 , n40643 , n40644 , n40645 , n40646 , 
     n40647 , n40648 , n40649 , n40650 , n40651 , n40652 , n40653 , n40654 , n40655 , n40656 , 
     n40657 , n40658 , n40659 , n40660 , n40661 , n40662 , n40663 , n40664 , n40665 , n40666 , 
     n40667 , n40668 , n40669 , n40670 , n40671 , n40672 , n40673 , n40674 , n40675 , n40676 , 
     n40677 , n40678 , n40679 , n40680 , n40681 , n40682 , n40683 , n40684 , n40685 , n40686 , 
     n40687 , n40688 , n40689 , n40690 , n40691 , n40692 , n40693 , n40694 , n40695 , n40696 , 
     n40697 , n40698 , n40699 , n40700 , n40701 , n40702 , n40703 , n40704 , n40705 , n40706 , 
     n40707 , n40708 , n40709 , n40710 , n40711 , n40712 , n40713 , n40714 , n40715 , n40716 , 
     n40717 , n40718 , n40719 , n40720 , n40721 , n40722 , n40723 , n40724 , n40725 , n40726 , 
     n40727 , n40728 , n40729 , n40730 , n40731 , n40732 , n40733 , n40734 , n40735 , n40736 , 
     n40737 , n40738 , n40739 , n40740 , n40741 , n40742 , n40743 , n40744 , n40745 , n40746 , 
     n40747 , n40748 , n40749 , n40750 , n40751 , n40752 , n40753 , n40754 , n40755 , n40756 , 
     n40757 , n40758 , n40759 , n40760 , n40761 , n40762 , n40763 , n40764 , n40765 , n40766 , 
     n40767 , n40768 , n40769 , n40770 , n40771 , n40772 , n40773 , n40774 , n40775 , n40776 , 
     n40777 , n40778 , n40779 , n40780 , n40781 , n40782 , n40783 , n40784 , n40785 , n40786 , 
     n40787 , n40788 , n40789 , n40790 , n40791 , n40792 , n40793 , n40794 , n40795 , n40796 , 
     n40797 , n40798 , n40799 , n40800 , n40801 , n40802 , n40803 , n40804 , n40805 , n40806 , 
     n40807 , n40808 , n40809 , n40810 , n40811 , n40812 , n40813 , n40814 , n40815 , n40816 , 
     n40817 , n40818 , n40819 , n40820 , n40821 , n40822 , n40823 , n40824 , n40825 , n40826 , 
     n40827 , n40828 , n40829 , n40830 , n40831 , n40832 , n40833 , n40834 , n40835 , n40836 , 
     n40837 , n40838 , n40839 , n40840 , n40841 , n40842 , n40843 , n40844 , n40845 , n40846 , 
     n40847 , n40848 , n40849 , n40850 , n40851 , n40852 , n40853 , n40854 , n40855 , n40856 , 
     n40857 , n40858 , n40859 , n40860 , n40861 , n40862 , n40863 , n40864 , n40865 , n40866 , 
     n40867 , n40868 , n40869 , n40870 , n40871 , n40872 , n40873 , n40874 , n40875 , n40876 , 
     n40877 , n40878 , n40879 , n40880 , n40881 , n40882 , n40883 , n40884 , n40885 , n40886 , 
     n40887 , n40888 , n40889 , n40890 , n40891 , n40892 , n40893 , n40894 , n40895 , n40896 , 
     n40897 , n40898 , n40899 , n40900 , n40901 , n40902 , n40903 , n40904 , n40905 , n40906 , 
     n40907 , n40908 , n40909 , n40910 , n40911 , n40912 , n40913 , n40914 , n40915 , n40916 , 
     n40917 , n40918 , n40919 , n40920 , n40921 , n40922 , n40923 , n40924 , n40925 , n40926 , 
     n40927 , n40928 , n40929 , n40930 , n40931 , n40932 , n40933 , n40934 , n40935 , n40936 , 
     n40937 , n40938 , n40939 , n40940 , n40941 , n40942 , n40943 , n40944 , n40945 , n40946 , 
     n40947 , n40948 , n40949 , n40950 , n40951 , n40952 , n40953 , n40954 , n40955 , n40956 , 
     n40957 , n40958 , n40959 , n40960 , n40961 , n40962 , n40963 , n40964 , n40965 , n40966 , 
     n40967 , n40968 , n40969 , n40970 , n40971 , n40972 , n40973 , n40974 , n40975 , n40976 , 
     n40977 , n40978 , n40979 , n40980 , n40981 , n40982 , n40983 , n40984 , n40985 , n40986 , 
     n40987 , n40988 , n40989 , n40990 , n40991 , n40992 , n40993 , n40994 , n40995 , n40996 , 
     n40997 , n40998 , n40999 , n41000 , n41001 , n41002 , n41003 , n41004 , n41005 , n41006 , 
     n41007 , n41008 , n41009 , n41010 , n41011 , n41012 , n41013 , n41014 , n41015 , n41016 , 
     n41017 , n41018 , n41019 , n41020 , n41021 , n41022 , n41023 , n41024 , n41025 , n41026 , 
     n41027 , n41028 , n41029 , n41030 , n41031 , n41032 , n41033 , n41034 , n41035 , n41036 , 
     n41037 , n41038 , n41039 , n41040 , n41041 , n41042 , n41043 , n41044 , n41045 , n41046 , 
     n41047 , n41048 , n41049 , n41050 , n41051 , n41052 , n41053 , n41054 , n41055 , n41056 , 
     n41057 , n41058 , n41059 , n41060 , n41061 , n41062 , n41063 , n41064 , n41065 , n41066 , 
     n41067 , n41068 , n41069 , n41070 , n41071 , n41072 , n41073 , n41074 , n41075 , n41076 , 
     n41077 , n41078 , n41079 , n41080 , n41081 , n41082 , n41083 , n41084 , n41085 , n41086 , 
     n41087 , n41088 , n41089 , n41090 , n41091 , n41092 , n41093 , n41094 , n41095 , n41096 , 
     n41097 , n41098 , n41099 , n41100 , n41101 , n41102 , n41103 , n41104 , n41105 , n41106 , 
     n41107 , n41108 , n41109 , n41110 , n41111 , n41112 , n41113 , n41114 , n41115 , n41116 , 
     n41117 , n41118 , n41119 , n41120 , n41121 , n41122 , n41123 , n41124 , n41125 , n41126 , 
     n41127 , n41128 , n41129 , n41130 , n41131 , n41132 , n41133 , n41134 , n41135 , n41136 , 
     n41137 , n41138 , n41139 , n41140 , n41141 , n41142 , n41143 , n41144 , n41145 , n41146 , 
     n41147 , n41148 , n41149 , n41150 , n41151 , n41152 , n41153 , n41154 , n41155 , n41156 , 
     n41157 , n41158 , n41159 , n41160 , n41161 , n41162 , n41163 , n41164 , n41165 , n41166 , 
     n41167 , n41168 , n41169 , n41170 , n41171 , n41172 , n41173 , n41174 , n41175 , n41176 , 
     n41177 , n41178 , n41179 , n41180 , n41181 , n41182 , n41183 , n41184 , n41185 , n41186 , 
     n41187 , n41188 , n41189 , n41190 , n41191 , n41192 , n41193 , n41194 , n41195 , n41196 , 
     n41197 , n41198 , n41199 , n41200 , n41201 , n41202 , n41203 , n41204 , n41205 , n41206 , 
     n41207 , n41208 , n41209 , n41210 , n41211 , n41212 , n41213 , n41214 , n41215 , n41216 , 
     n41217 , n41218 , n41219 , n41220 , n41221 , n41222 , n41223 , n41224 , n41225 , n41226 , 
     n41227 , n41228 , n41229 , n41230 , n41231 , n41232 , n41233 , n41234 , n41235 , n41236 , 
     n41237 , n41238 , n41239 , n41240 , n41241 , n41242 , n41243 , n41244 , n41245 , n41246 , 
     n41247 , n41248 , n41249 , n41250 , n41251 , n41252 , n41253 , n41254 , n41255 , n41256 , 
     n41257 , n41258 , n41259 , n41260 , n41261 , n41262 , n41263 , n41264 , n41265 , n41266 , 
     n41267 , n41268 , n41269 , n41270 , n41271 , n41272 , n41273 , n41274 , n41275 , n41276 , 
     n41277 , n41278 , n41279 , n41280 , n41281 , n41282 , n41283 , n41284 , n41285 , n41286 , 
     n41287 , n41288 , n41289 , n41290 , n41291 , n41292 , n41293 , n41294 , n41295 , n41296 , 
     n41297 , n41298 , n41299 , n41300 , n41301 , n41302 , n41303 , n41304 , n41305 , n41306 , 
     n41307 , n41308 , n41309 , n41310 , n41311 , n41312 , n41313 , n41314 , n41315 , n41316 , 
     n41317 , n41318 , n41319 , n41320 , n41321 , n41322 , n41323 , n41324 , n41325 , n41326 , 
     n41327 , n41328 , n41329 , n41330 , n41331 , n41332 , n41333 , n41334 , n41335 , n41336 , 
     n41337 , n41338 , n41339 , n41340 , n41341 , n41342 , n41343 , n41344 , n41345 , n41346 , 
     n41347 , n41348 , n41349 , n41350 , n41351 , n41352 , n41353 , n41354 , n41355 , n41356 , 
     n41357 , n41358 , n41359 , n41360 , n41361 , n41362 , n41363 , n41364 , n41365 , n41366 , 
     n41367 , n41368 , n41369 , n41370 , n41371 , n41372 , n41373 , n41374 , n41375 , n41376 , 
     n41377 , n41378 , n41379 , n41380 , n41381 , n41382 , n41383 , n41384 , n41385 , n41386 , 
     n41387 , n41388 , n41389 , n41390 , n41391 , n41392 , n41393 , n41394 , n41395 , n41396 , 
     n41397 , n41398 , n41399 , n41400 , n41401 , n41402 , n41403 , n41404 , n41405 , n41406 , 
     n41407 , n41408 , n41409 , n41410 , n41411 , n41412 , n41413 , n41414 , n41415 , n41416 , 
     n41417 , n41418 , n41419 , n41420 , n41421 , n41422 , n41423 , n41424 , n41425 , n41426 , 
     n41427 , n41428 , n41429 , n41430 , n41431 , n41432 , n41433 , n41434 , n41435 , n41436 , 
     n41437 , n41438 , n41439 , n41440 , n41441 , n41442 , n41443 , n41444 , n41445 , n41446 , 
     n41447 , n41448 , n41449 , n41450 , n41451 , n41452 , n41453 , n41454 , n41455 , n41456 , 
     n41457 , n41458 , n41459 , n41460 , n41461 , n41462 , n41463 , n41464 , n41465 , n41466 , 
     n41467 , n41468 , n41469 , n41470 , n41471 , n41472 , n41473 , n41474 , n41475 , n41476 , 
     n41477 , n41478 , n41479 , n41480 , n41481 , n41482 , n41483 , n41484 , n41485 , n41486 , 
     n41487 , n41488 , n41489 , n41490 , n41491 , n41492 , n41493 , n41494 , n41495 , n41496 , 
     n41497 , n41498 , n41499 , n41500 , n41501 , n41502 , n41503 , n41504 , n41505 , n41506 , 
     n41507 , n41508 , n41509 , n41510 , n41511 , n41512 , n41513 , n41514 , n41515 , n41516 , 
     n41517 , n41518 , n41519 , n41520 , n41521 , n41522 , n41523 , n41524 , n41525 , n41526 , 
     n41527 , n41528 , n41529 , n41530 , n41531 , n41532 , n41533 , n41534 , n41535 , n41536 , 
     n41537 , n41538 , n41539 , n41540 , n41541 , n41542 , n41543 , n41544 , n41545 , n41546 , 
     n41547 , n41548 , n41549 , n41550 , n41551 , n41552 , n41553 , n41554 , n41555 , n41556 , 
     n41557 , n41558 , n41559 , n41560 , n41561 , n41562 , n41563 , n41564 , n41565 , n41566 , 
     n41567 , n41568 , n41569 , n41570 , n41571 , n41572 , n41573 , n41574 , n41575 , n41576 , 
     n41577 , n41578 , n41579 , n41580 , n41581 , n41582 , n41583 , n41584 , n41585 , n41586 , 
     n41587 , n41588 , n41589 , n41590 , n41591 , n41592 , n41593 , n41594 , n41595 , n41596 , 
     n41597 , n41598 , n41599 , n41600 , n41601 , n41602 , n41603 , n41604 , n41605 , n41606 , 
     n41607 , n41608 , n41609 , n41610 , n41611 , n41612 , n41613 , n41614 , n41615 , n41616 , 
     n41617 , n41618 , n41619 , n41620 , n41621 , n41622 , n41623 , n41624 , n41625 , n41626 , 
     n41627 , n41628 , n41629 , n41630 , n41631 , n41632 , n41633 , n41634 , n41635 , n41636 , 
     n41637 , n41638 , n41639 , n41640 , n41641 , n41642 , n41643 , n41644 , n41645 , n41646 , 
     n41647 , n41648 , n41649 , n41650 , n41651 , n41652 , n41653 , n41654 , n41655 , n41656 , 
     n41657 , n41658 , n41659 , n41660 , n41661 , n41662 , n41663 , n41664 , n41665 , n41666 , 
     n41667 , n41668 , n41669 , n41670 , n41671 , n41672 , n41673 , n41674 , n41675 , n41676 , 
     n41677 , n41678 , n41679 , n41680 , n41681 , n41682 , n41683 , n41684 , n41685 , n41686 , 
     n41687 , n41688 , n41689 , n41690 , n41691 , n41692 , n41693 , n41694 , n41695 , n41696 , 
     n41697 , n41698 , n41699 , n41700 , n41701 , n41702 , n41703 , n41704 , n41705 , n41706 , 
     n41707 , n41708 , n41709 , n41710 , n41711 , n41712 , n41713 , n41714 , n41715 , n41716 , 
     n41717 , n41718 , n41719 , n41720 , n41721 , n41722 , n41723 , n41724 , n41725 , n41726 , 
     n41727 , n41728 , n41729 , n41730 , n41731 , n41732 , n41733 , n41734 , n41735 , n41736 , 
     n41737 , n41738 , n41739 , n41740 , n41741 , n41742 , n41743 , n41744 , n41745 , n41746 , 
     n41747 , n41748 , n41749 , n41750 , n41751 , n41752 , n41753 , n41754 , n41755 , n41756 , 
     n41757 , n41758 , n41759 , n41760 , n41761 , n41762 , n41763 , n41764 , n41765 , n41766 , 
     n41767 , n41768 , n41769 , n41770 , n41771 , n41772 , n41773 , n41774 , n41775 , n41776 , 
     n41777 , n41778 , n41779 , n41780 , n41781 , n41782 , n41783 , n41784 , n41785 , n41786 , 
     n41787 , n41788 , n41789 , n41790 , n41791 , n41792 , n41793 , n41794 , n41795 , n41796 , 
     n41797 , n41798 , n41799 , n41800 , n41801 , n41802 , n41803 , n41804 , n41805 , n41806 , 
     n41807 , n41808 , n41809 , n41810 , n41811 , n41812 , n41813 , n41814 , n41815 , n41816 , 
     n41817 , n41818 , n41819 , n41820 , n41821 , n41822 , n41823 , n41824 , n41825 , n41826 , 
     n41827 , n41828 , n41829 , n41830 , n41831 , n41832 , n41833 , n41834 , n41835 , n41836 , 
     n41837 , n41838 , n41839 , n41840 , n41841 , n41842 , n41843 , n41844 , n41845 , n41846 , 
     n41847 , n41848 , n41849 , n41850 , n41851 , n41852 , n41853 , n41854 , n41855 , n41856 , 
     n41857 , n41858 , n41859 , n41860 , n41861 , n41862 , n41863 , n41864 , n41865 , n41866 , 
     n41867 , n41868 , n41869 , n41870 , n41871 , n41872 , n41873 , n41874 , n41875 , n41876 , 
     n41877 , n41878 , n41879 , n41880 , n41881 , n41882 , n41883 , n41884 , n41885 , n41886 , 
     n41887 , n41888 , n41889 , n41890 , n41891 , n41892 , n41893 , n41894 , n41895 , n41896 , 
     n41897 , n41898 , n41899 , n41900 , n41901 , n41902 , n41903 , n41904 , n41905 , n41906 , 
     n41907 , n41908 , n41909 , n41910 , n41911 , n41912 , n41913 , n41914 , n41915 , n41916 , 
     n41917 , n41918 , n41919 , n41920 , n41921 , n41922 , n41923 , n41924 , n41925 , n41926 , 
     n41927 , n41928 , n41929 , n41930 , n41931 , n41932 , n41933 , n41934 , n41935 , n41936 , 
     n41937 , n41938 , n41939 , n41940 , n41941 , n41942 , n41943 , n41944 , n41945 , n41946 , 
     n41947 , n41948 , n41949 , n41950 , n41951 , n41952 , n41953 , n41954 , n41955 , n41956 , 
     n41957 , n41958 , n41959 , n41960 , n41961 , n41962 , n41963 , n41964 , n41965 , n41966 , 
     n41967 , n41968 , n41969 , n41970 , n41971 , n41972 , n41973 , n41974 , n41975 , n41976 , 
     n41977 , n41978 , n41979 , n41980 , n41981 , n41982 , n41983 , n41984 , n41985 , n41986 , 
     n41987 , n41988 , n41989 , n41990 , n41991 , n41992 , n41993 , n41994 , n41995 , n41996 , 
     n41997 , n41998 , n41999 , n42000 , n42001 , n42002 , n42003 , n42004 , n42005 , n42006 , 
     n42007 , n42008 , n42009 , n42010 , n42011 , n42012 , n42013 , n42014 , n42015 , n42016 , 
     n42017 , n42018 , n42019 , n42020 , n42021 , n42022 , n42023 , n42024 , n42025 , n42026 , 
     n42027 , n42028 , n42029 , n42030 , n42031 , n42032 , n42033 , n42034 , n42035 , n42036 , 
     n42037 , n42038 , n42039 , n42040 , n42041 , n42042 , n42043 , n42044 , n42045 , n42046 , 
     n42047 , n42048 , n42049 , n42050 , n42051 , n42052 , n42053 , n42054 , n42055 , n42056 , 
     n42057 , n42058 , n42059 , n42060 , n42061 , n42062 , n42063 , n42064 , n42065 , n42066 , 
     n42067 , n42068 , n42069 , n42070 , n42071 , n42072 , n42073 , n42074 , n42075 , n42076 , 
     n42077 , n42078 , n42079 , n42080 , n42081 , n42082 , n42083 , n42084 , n42085 , n42086 , 
     n42087 , n42088 , n42089 , n42090 , n42091 , n42092 , n42093 , n42094 , n42095 , n42096 , 
     n42097 , n42098 , n42099 , n42100 , n42101 , n42102 , n42103 , n42104 , n42105 , n42106 , 
     n42107 , n42108 , n42109 , n42110 , n42111 , n42112 , n42113 , n42114 , n42115 , n42116 , 
     n42117 , n42118 , n42119 , n42120 , n42121 , n42122 , n42123 , n42124 , n42125 , n42126 , 
     n42127 , n42128 , n42129 , n42130 , n42131 , n42132 , n42133 , n42134 , n42135 , n42136 , 
     n42137 , n42138 , n42139 , n42140 , n42141 , n42142 , n42143 , n42144 , n42145 , n42146 , 
     n42147 , n42148 , n42149 , n42150 , n42151 , n42152 , n42153 , n42154 , n42155 , n42156 , 
     n42157 , n42158 , n42159 , n42160 , n42161 , n42162 , n42163 , n42164 , n42165 , n42166 , 
     n42167 , n42168 , n42169 , n42170 , n42171 , n42172 , n42173 , n42174 , n42175 , n42176 , 
     n42177 , n42178 , n42179 , n42180 , n42181 , n42182 , n42183 , n42184 , n42185 , n42186 , 
     n42187 , n42188 , n42189 , n42190 , n42191 , n42192 , n42193 , n42194 , n42195 , n42196 , 
     n42197 , n42198 , n42199 , n42200 , n42201 , n42202 , n42203 , n42204 , n42205 , n42206 , 
     n42207 , n42208 , n42209 , n42210 , n42211 , n42212 , n42213 , n42214 , n42215 , n42216 , 
     n42217 , n42218 , n42219 , n42220 , n42221 , n42222 , n42223 , n42224 , n42225 , n42226 , 
     n42227 , n42228 , n42229 , n42230 , n42231 , n42232 , n42233 , n42234 , n42235 , n42236 , 
     n42237 , n42238 , n42239 , n42240 , n42241 , n42242 , n42243 , n42244 , n42245 , n42246 , 
     n42247 , n42248 , n42249 , n42250 , n42251 , n42252 , n42253 , n42254 , n42255 , n42256 , 
     n42257 , n42258 , n42259 , n42260 , n42261 , n42262 , n42263 , n42264 , n42265 , n42266 , 
     n42267 , n42268 , n42269 , n42270 , n42271 , n42272 , n42273 , n42274 , n42275 , n42276 , 
     n42277 , n42278 , n42279 , n42280 , n42281 , n42282 , n42283 , n42284 , n42285 , n42286 , 
     n42287 , n42288 , n42289 , n42290 , n42291 , n42292 , n42293 , n42294 , n42295 , n42296 , 
     n42297 , n42298 , n42299 , n42300 , n42301 , n42302 , n42303 , n42304 , n42305 , n42306 , 
     n42307 , n42308 , n42309 , n42310 , n42311 , n42312 , n42313 , n42314 , n42315 , n42316 , 
     n42317 , n42318 , n42319 , n42320 , n42321 , n42322 , n42323 , n42324 , n42325 , n42326 , 
     n42327 , n42328 , n42329 , n42330 , n42331 , n42332 , n42333 , n42334 , n42335 , n42336 , 
     n42337 , n42338 , n42339 , n42340 , n42341 , n42342 , n42343 , n42344 , n42345 , n42346 , 
     n42347 , n42348 , n42349 , n42350 , n42351 , n42352 , n42353 , n42354 , n42355 , n42356 , 
     n42357 , n42358 , n42359 , n42360 , n42361 , n42362 , n42363 , n42364 , n42365 , n42366 , 
     n42367 , n42368 , n42369 , n42370 , n42371 , n42372 , n42373 , n42374 , n42375 , n42376 , 
     n42377 , n42378 , n42379 , n42380 , n42381 , n42382 , n42383 , n42384 , n42385 , n42386 , 
     n42387 , n42388 , n42389 , n42390 , n42391 , n42392 , n42393 , n42394 , n42395 , n42396 , 
     n42397 , n42398 , n42399 , n42400 , n42401 , n42402 , n42403 , n42404 , n42405 , n42406 , 
     n42407 , n42408 , n42409 , n42410 , n42411 , n42412 , n42413 , n42414 , n42415 , n42416 , 
     n42417 , n42418 , n42419 , n42420 , n42421 , n42422 , n42423 , n42424 , n42425 , n42426 , 
     n42427 , n42428 , n42429 , n42430 , n42431 , n42432 , n42433 , n42434 , n42435 , n42436 , 
     n42437 , n42438 , n42439 , n42440 , n42441 , n42442 , n42443 , n42444 , n42445 , n42446 , 
     n42447 , n42448 , n42449 , n42450 , n42451 , n42452 , n42453 , n42454 , n42455 , n42456 , 
     n42457 , n42458 , n42459 , n42460 , n42461 , n42462 , n42463 , n42464 , n42465 , n42466 , 
     n42467 , n42468 , n42469 , n42470 , n42471 , n42472 , n42473 , n42474 , n42475 , n42476 , 
     n42477 , n42478 , n42479 , n42480 , n42481 , n42482 , n42483 , n42484 , n42485 , n42486 , 
     n42487 , n42488 , n42489 , n42490 , n42491 , n42492 , n42493 , n42494 , n42495 , n42496 , 
     n42497 , n42498 , n42499 , n42500 , n42501 , n42502 , n42503 , n42504 , n42505 , n42506 , 
     n42507 , n42508 , n42509 , n42510 , n42511 , n42512 , n42513 , n42514 , n42515 , n42516 , 
     n42517 , n42518 , n42519 , n42520 , n42521 , n42522 , n42523 , n42524 , n42525 , n42526 , 
     n42527 , n42528 , n42529 , n42530 , n42531 , n42532 , n42533 , n42534 , n42535 , n42536 , 
     n42537 , n42538 , n42539 , n42540 , n42541 , n42542 , n42543 , n42544 , n42545 , n42546 , 
     n42547 , n42548 , n42549 , n42550 , n42551 , n42552 , n42553 , n42554 , n42555 , n42556 , 
     n42557 , n42558 , n42559 , n42560 , n42561 , n42562 , n42563 , n42564 , n42565 , n42566 , 
     n42567 , n42568 , n42569 , n42570 , n42571 , n42572 , n42573 , n42574 , n42575 , n42576 , 
     n42577 , n42578 , n42579 , n42580 , n42581 , n42582 , n42583 , n42584 , n42585 , n42586 , 
     n42587 , n42588 , n42589 , n42590 , n42591 , n42592 , n42593 , n42594 , n42595 , n42596 , 
     n42597 , n42598 , n42599 , n42600 , n42601 , n42602 , n42603 , n42604 , n42605 , n42606 , 
     n42607 , n42608 , n42609 , n42610 , n42611 , n42612 , n42613 , n42614 , n42615 , n42616 , 
     n42617 , n42618 , n42619 , n42620 , n42621 , n42622 , n42623 , n42624 , n42625 , n42626 , 
     n42627 , n42628 , n42629 , n42630 , n42631 , n42632 , n42633 , n42634 , n42635 , n42636 , 
     n42637 , n42638 , n42639 , n42640 , n42641 , n42642 , n42643 , n42644 , n42645 , n42646 , 
     n42647 , n42648 , n42649 , n42650 , n42651 , n42652 , n42653 , n42654 , n42655 , n42656 , 
     n42657 , n42658 , n42659 , n42660 , n42661 , n42662 , n42663 , n42664 , n42665 , n42666 , 
     n42667 , n42668 , n42669 , n42670 , n42671 , n42672 , n42673 , n42674 , n42675 , n42676 , 
     n42677 , n42678 , n42679 , n42680 , n42681 , n42682 , n42683 , n42684 , n42685 , n42686 , 
     n42687 , n42688 , n42689 , n42690 , n42691 , n42692 , n42693 , n42694 , n42695 , n42696 , 
     n42697 , n42698 , n42699 , n42700 , n42701 , n42702 , n42703 , n42704 , n42705 , n42706 , 
     n42707 , n42708 , n42709 , n42710 , n42711 , n42712 , n42713 , n42714 , n42715 , n42716 , 
     n42717 , n42718 , n42719 , n42720 , n42721 , n42722 , n42723 , n42724 , n42725 , n42726 , 
     n42727 , n42728 , n42729 , n42730 , n42731 , n42732 , n42733 , n42734 , n42735 , n42736 , 
     n42737 , n42738 , n42739 , n42740 , n42741 , n42742 , n42743 , n42744 , n42745 , n42746 , 
     n42747 , n42748 , n42749 , n42750 , n42751 , n42752 , n42753 , n42754 , n42755 , n42756 , 
     n42757 , n42758 , n42759 , n42760 , n42761 , n42762 , n42763 , n42764 , n42765 , n42766 , 
     n42767 , n42768 , n42769 , n42770 , n42771 , n42772 , n42773 , n42774 , n42775 , n42776 , 
     n42777 , n42778 , n42779 , n42780 , n42781 , n42782 , n42783 , n42784 , n42785 , n42786 , 
     n42787 , n42788 , n42789 , n42790 , n42791 , n42792 , n42793 , n42794 , n42795 , n42796 , 
     n42797 , n42798 , n42799 , n42800 , n42801 , n42802 , n42803 , n42804 , n42805 , n42806 , 
     n42807 , n42808 , n42809 , n42810 , n42811 , n42812 , n42813 , n42814 , n42815 , n42816 , 
     n42817 , n42818 , n42819 , n42820 , n42821 , n42822 , n42823 , n42824 , n42825 , n42826 , 
     n42827 , n42828 , n42829 , n42830 , n42831 , n42832 , n42833 , n42834 , n42835 , n42836 , 
     n42837 , n42838 , n42839 , n42840 , n42841 , n42842 , n42843 , n42844 , n42845 , n42846 , 
     n42847 , n42848 , n42849 , n42850 , n42851 , n42852 , n42853 , n42854 , n42855 , n42856 , 
     n42857 , n42858 , n42859 , n42860 , n42861 , n42862 , n42863 , n42864 , n42865 , n42866 , 
     n42867 , n42868 , n42869 , n42870 , n42871 , n42872 , n42873 , n42874 , n42875 , n42876 , 
     n42877 , n42878 , n42879 , n42880 , n42881 , n42882 , n42883 , n42884 , n42885 , n42886 , 
     n42887 , n42888 , n42889 , n42890 , n42891 , n42892 , n42893 , n42894 , n42895 , n42896 , 
     n42897 , n42898 , n42899 , n42900 , n42901 , n42902 , n42903 , n42904 , n42905 , n42906 , 
     n42907 , n42908 , n42909 , n42910 , n42911 , n42912 , n42913 , n42914 , n42915 , n42916 , 
     n42917 , n42918 , n42919 , n42920 , n42921 , n42922 , n42923 , n42924 , n42925 , n42926 , 
     n42927 , n42928 , n42929 , n42930 , n42931 , n42932 , n42933 , n42934 , n42935 , n42936 , 
     n42937 , n42938 , n42939 , n42940 , n42941 , n42942 , n42943 , n42944 , n42945 , n42946 , 
     n42947 , n42948 , n42949 , n42950 , n42951 , n42952 , n42953 , n42954 , n42955 , n42956 , 
     n42957 , n42958 , n42959 , n42960 , n42961 , n42962 , n42963 , n42964 , n42965 , n42966 , 
     n42967 , n42968 , n42969 , n42970 , n42971 , n42972 , n42973 , n42974 , n42975 , n42976 , 
     n42977 , n42978 , n42979 , n42980 , n42981 , n42982 , n42983 , n42984 , n42985 , n42986 , 
     n42987 , n42988 , n42989 , n42990 , n42991 , n42992 , n42993 , n42994 , n42995 , n42996 , 
     n42997 , n42998 , n42999 , n43000 , n43001 , n43002 , n43003 , n43004 , n43005 , n43006 , 
     n43007 , n43008 , n43009 , n43010 , n43011 , n43012 , n43013 , n43014 , n43015 , n43016 , 
     n43017 , n43018 , n43019 , n43020 , n43021 , n43022 , n43023 , n43024 , n43025 , n43026 , 
     n43027 , n43028 , n43029 , n43030 , n43031 , n43032 , n43033 , n43034 , n43035 , n43036 , 
     n43037 , n43038 , n43039 , n43040 , n43041 , n43042 , n43043 , n43044 , n43045 , n43046 , 
     n43047 , n43048 , n43049 , n43050 , n43051 , n43052 , n43053 , n43054 , n43055 , n43056 , 
     n43057 , n43058 , n43059 , n43060 , n43061 , n43062 , n43063 , n43064 , n43065 , n43066 , 
     n43067 , n43068 , n43069 , n43070 , n43071 , n43072 , n43073 , n43074 , n43075 , n43076 , 
     n43077 , n43078 , n43079 , n43080 , n43081 , n43082 , n43083 , n43084 , n43085 , n43086 , 
     n43087 , n43088 , n43089 , n43090 , n43091 , n43092 , n43093 , n43094 , n43095 , n43096 , 
     n43097 , n43098 , n43099 , n43100 , n43101 , n43102 , n43103 , n43104 , n43105 , n43106 , 
     n43107 , n43108 , n43109 , n43110 , n43111 , n43112 , n43113 , n43114 , n43115 , n43116 , 
     n43117 , n43118 , n43119 , n43120 , n43121 , n43122 , n43123 , n43124 , n43125 , n43126 , 
     n43127 , n43128 , n43129 , n43130 , n43131 , n43132 , n43133 , n43134 , n43135 , n43136 , 
     n43137 , n43138 , n43139 , n43140 , n43141 , n43142 , n43143 , n43144 , n43145 , n43146 , 
     n43147 , n43148 , n43149 , n43150 , n43151 , n43152 , n43153 , n43154 , n43155 , n43156 , 
     n43157 , n43158 , n43159 , n43160 , n43161 , n43162 , n43163 , n43164 , n43165 , n43166 , 
     n43167 , n43168 , n43169 , n43170 , n43171 , n43172 , n43173 , n43174 , n43175 , n43176 , 
     n43177 , n43178 , n43179 , n43180 , n43181 , n43182 , n43183 , n43184 , n43185 , n43186 , 
     n43187 , n43188 , n43189 , n43190 , n43191 , n43192 , n43193 , n43194 , n43195 , n43196 , 
     n43197 , n43198 , n43199 , n43200 , n43201 , n43202 , n43203 , n43204 , n43205 , n43206 , 
     n43207 , n43208 , n43209 , n43210 , n43211 , n43212 , n43213 , n43214 , n43215 , n43216 , 
     n43217 , n43218 , n43219 , n43220 , n43221 , n43222 , n43223 , n43224 , n43225 , n43226 , 
     n43227 , n43228 , n43229 , n43230 , n43231 , n43232 , n43233 , n43234 , n43235 , n43236 , 
     n43237 , n43238 , n43239 , n43240 , n43241 , n43242 , n43243 , n43244 , n43245 , n43246 , 
     n43247 , n43248 , n43249 , n43250 , n43251 , n43252 , n43253 , n43254 , n43255 , n43256 , 
     n43257 , n43258 , n43259 , n43260 , n43261 , n43262 , n43263 , n43264 , n43265 , n43266 , 
     n43267 , n43268 , n43269 , n43270 , n43271 , n43272 , n43273 , n43274 , n43275 , n43276 , 
     n43277 , n43278 , n43279 , n43280 , n43281 , n43282 , n43283 , n43284 , n43285 , n43286 , 
     n43287 , n43288 , n43289 , n43290 , n43291 , n43292 , n43293 , n43294 , n43295 , n43296 , 
     n43297 , n43298 , n43299 , n43300 , n43301 , n43302 , n43303 , n43304 , n43305 , n43306 , 
     n43307 , n43308 , n43309 , n43310 , n43311 , n43312 , n43313 , n43314 , n43315 , n43316 , 
     n43317 , n43318 , n43319 , n43320 , n43321 , n43322 , n43323 , n43324 , n43325 , n43326 , 
     n43327 , n43328 , n43329 , n43330 , n43331 , n43332 , n43333 , n43334 , n43335 , n43336 , 
     n43337 , n43338 , n43339 , n43340 , n43341 , n43342 , n43343 , n43344 , n43345 , n43346 , 
     n43347 , n43348 , n43349 , n43350 , n43351 , n43352 , n43353 , n43354 , n43355 , n43356 , 
     n43357 , n43358 , n43359 , n43360 , n43361 , n43362 , n43363 , n43364 , n43365 , n43366 , 
     n43367 , n43368 , n43369 , n43370 , n43371 , n43372 , n43373 , n43374 , n43375 , n43376 , 
     n43377 , n43378 , n43379 , n43380 , n43381 , n43382 , n43383 , n43384 , n43385 , n43386 , 
     n43387 , n43388 , n43389 , n43390 , n43391 , n43392 , n43393 , n43394 , n43395 , n43396 , 
     n43397 , n43398 , n43399 , n43400 , n43401 , n43402 , n43403 , n43404 , n43405 , n43406 , 
     n43407 , n43408 , n43409 , n43410 , n43411 , n43412 , n43413 , n43414 , n43415 , n43416 , 
     n43417 , n43418 , n43419 , n43420 , n43421 , n43422 , n43423 , n43424 , n43425 , n43426 , 
     n43427 , n43428 , n43429 , n43430 , n43431 , n43432 , n43433 , n43434 , n43435 , n43436 , 
     n43437 , n43438 , n43439 , n43440 , n43441 , n43442 , n43443 , n43444 , n43445 , n43446 , 
     n43447 , n43448 , n43449 , n43450 , n43451 , n43452 , n43453 , n43454 , n43455 , n43456 , 
     n43457 , n43458 , n43459 , n43460 , n43461 , n43462 , n43463 , n43464 , n43465 , n43466 , 
     n43467 , n43468 , n43469 , n43470 , n43471 , n43472 , n43473 , n43474 , n43475 , n43476 , 
     n43477 , n43478 , n43479 , n43480 , n43481 , n43482 , n43483 , n43484 , n43485 , n43486 , 
     n43487 , n43488 , n43489 , n43490 , n43491 , n43492 , n43493 , n43494 , n43495 , n43496 , 
     n43497 , n43498 , n43499 , n43500 , n43501 , n43502 , n43503 , n43504 , n43505 , n43506 , 
     n43507 , n43508 , n43509 , n43510 , n43511 , n43512 , n43513 , n43514 , n43515 , n43516 , 
     n43517 , n43518 , n43519 , n43520 , n43521 , n43522 , n43523 , n43524 , n43525 , n43526 , 
     n43527 , n43528 , n43529 , n43530 , n43531 , n43532 , n43533 , n43534 , n43535 , n43536 , 
     n43537 , n43538 , n43539 , n43540 , n43541 , n43542 , n43543 , n43544 , n43545 , n43546 , 
     n43547 , n43548 , n43549 , n43550 , n43551 , n43552 , n43553 , n43554 , n43555 , n43556 , 
     n43557 , n43558 , n43559 , n43560 , n43561 , n43562 , n43563 , n43564 , n43565 , n43566 , 
     n43567 , n43568 , n43569 , n43570 , n43571 , n43572 , n43573 , n43574 , n43575 , n43576 , 
     n43577 , n43578 , n43579 , n43580 , n43581 , n43582 , n43583 , n43584 , n43585 , n43586 , 
     n43587 , n43588 , n43589 , n43590 , n43591 , n43592 , n43593 , n43594 , n43595 , n43596 , 
     n43597 , n43598 , n43599 , n43600 , n43601 , n43602 , n43603 , n43604 , n43605 , n43606 , 
     n43607 , n43608 , n43609 , n43610 , n43611 , n43612 , n43613 , n43614 , n43615 , n43616 , 
     n43617 , n43618 , n43619 , n43620 , n43621 , n43622 , n43623 , n43624 , n43625 , n43626 , 
     n43627 , n43628 , n43629 , n43630 , n43631 , n43632 , n43633 , n43634 , n43635 , n43636 , 
     n43637 , n43638 , n43639 , n43640 , n43641 , n43642 , n43643 , n43644 , n43645 , n43646 , 
     n43647 , n43648 , n43649 , n43650 , n43651 , n43652 , n43653 , n43654 , n43655 , n43656 , 
     n43657 , n43658 , n43659 , n43660 , n43661 , n43662 , n43663 , n43664 , n43665 , n43666 , 
     n43667 , n43668 , n43669 , n43670 , n43671 , n43672 , n43673 , n43674 , n43675 , n43676 , 
     n43677 , n43678 , n43679 , n43680 , n43681 , n43682 , n43683 , n43684 , n43685 , n43686 , 
     n43687 , n43688 , n43689 , n43690 , n43691 , n43692 , n43693 , n43694 , n43695 , n43696 , 
     n43697 , n43698 , n43699 , n43700 , n43701 , n43702 , n43703 , n43704 , n43705 , n43706 , 
     n43707 , n43708 , n43709 , n43710 , n43711 , n43712 , n43713 , n43714 , n43715 , n43716 , 
     n43717 , n43718 , n43719 , n43720 , n43721 , n43722 , n43723 , n43724 , n43725 , n43726 , 
     n43727 , n43728 , n43729 , n43730 , n43731 , n43732 , n43733 , n43734 , n43735 , n43736 , 
     n43737 , n43738 , n43739 , n43740 , n43741 , n43742 , n43743 , n43744 , n43745 , n43746 , 
     n43747 , n43748 , n43749 , n43750 , n43751 , n43752 , n43753 , n43754 , n43755 , n43756 , 
     n43757 , n43758 , n43759 , n43760 , n43761 , n43762 , n43763 , n43764 , n43765 , n43766 , 
     n43767 , n43768 , n43769 , n43770 , n43771 , n43772 , n43773 , n43774 , n43775 , n43776 , 
     n43777 , n43778 , n43779 , n43780 , n43781 , n43782 , n43783 , n43784 , n43785 , n43786 , 
     n43787 , n43788 , n43789 , n43790 , n43791 , n43792 , n43793 , n43794 , n43795 , n43796 , 
     n43797 , n43798 , n43799 , n43800 , n43801 , n43802 , n43803 , n43804 , n43805 , n43806 , 
     n43807 , n43808 , n43809 , n43810 , n43811 , n43812 , n43813 , n43814 , n43815 , n43816 , 
     n43817 , n43818 , n43819 , n43820 , n43821 , n43822 , n43823 , n43824 , n43825 , n43826 , 
     n43827 , n43828 , n43829 , n43830 , n43831 , n43832 , n43833 , n43834 , n43835 , n43836 , 
     n43837 , n43838 , n43839 , n43840 , n43841 , n43842 , n43843 , n43844 , n43845 , n43846 , 
     n43847 , n43848 , n43849 , n43850 , n43851 , n43852 , n43853 , n43854 , n43855 , n43856 , 
     n43857 , n43858 , n43859 , n43860 , n43861 , n43862 , n43863 , n43864 , n43865 , n43866 , 
     n43867 , n43868 , n43869 , n43870 , n43871 , n43872 , n43873 , n43874 , n43875 , n43876 , 
     n43877 , n43878 , n43879 , n43880 , n43881 , n43882 , n43883 , n43884 , n43885 , n43886 , 
     n43887 , n43888 , n43889 , n43890 , n43891 , n43892 , n43893 , n43894 , n43895 , n43896 , 
     n43897 , n43898 , n43899 , n43900 , n43901 , n43902 , n43903 , n43904 , n43905 , n43906 , 
     n43907 , n43908 , n43909 , n43910 , n43911 , n43912 , n43913 , n43914 , n43915 , n43916 , 
     n43917 , n43918 , n43919 , n43920 , n43921 , n43922 , n43923 , n43924 , n43925 , n43926 , 
     n43927 , n43928 , n43929 , n43930 , n43931 , n43932 , n43933 , n43934 , n43935 , n43936 , 
     n43937 , n43938 , n43939 , n43940 , n43941 , n43942 , n43943 , n43944 , n43945 , n43946 , 
     n43947 , n43948 , n43949 , n43950 , n43951 , n43952 , n43953 , n43954 , n43955 , n43956 , 
     n43957 , n43958 , n43959 , n43960 , n43961 , n43962 , n43963 , n43964 , n43965 , n43966 , 
     n43967 , n43968 , n43969 , n43970 , n43971 , n43972 , n43973 , n43974 , n43975 , n43976 , 
     n43977 , n43978 , n43979 , n43980 , n43981 , n43982 , n43983 , n43984 , n43985 , n43986 , 
     n43987 , n43988 , n43989 , n43990 , n43991 , n43992 , n43993 , n43994 , n43995 , n43996 , 
     n43997 , n43998 , n43999 , n44000 , n44001 , n44002 , n44003 , n44004 , n44005 , n44006 , 
     n44007 , n44008 , n44009 , n44010 , n44011 , n44012 , n44013 , n44014 , n44015 , n44016 , 
     n44017 , n44018 , n44019 , n44020 , n44021 , n44022 , n44023 , n44024 , n44025 , n44026 , 
     n44027 , n44028 , n44029 , n44030 , n44031 , n44032 , n44033 , n44034 , n44035 , n44036 , 
     n44037 , n44038 , n44039 , n44040 , n44041 , n44042 , n44043 , n44044 , n44045 , n44046 , 
     n44047 , n44048 , n44049 , n44050 , n44051 , n44052 , n44053 , n44054 , n44055 , n44056 , 
     n44057 , n44058 , n44059 , n44060 , n44061 , n44062 , n44063 , n44064 , n44065 , n44066 , 
     n44067 , n44068 , n44069 , n44070 , n44071 , n44072 , n44073 , n44074 , n44075 , n44076 , 
     n44077 , n44078 , n44079 , n44080 , n44081 , n44082 , n44083 , n44084 , n44085 , n44086 , 
     n44087 , n44088 , n44089 , n44090 , n44091 , n44092 , n44093 , n44094 , n44095 , n44096 , 
     n44097 , n44098 , n44099 , n44100 , n44101 , n44102 , n44103 , n44104 , n44105 , n44106 , 
     n44107 , n44108 , n44109 , n44110 , n44111 , n44112 , n44113 , n44114 , n44115 , n44116 , 
     n44117 , n44118 , n44119 , n44120 , n44121 , n44122 , n44123 , n44124 , n44125 , n44126 , 
     n44127 , n44128 , n44129 , n44130 , n44131 , n44132 , n44133 , n44134 , n44135 , n44136 , 
     n44137 , n44138 , n44139 , n44140 , n44141 , n44142 , n44143 , n44144 , n44145 , n44146 , 
     n44147 , n44148 , n44149 , n44150 , n44151 , n44152 , n44153 , n44154 , n44155 , n44156 , 
     n44157 , n44158 , n44159 , n44160 , n44161 , n44162 , n44163 , n44164 , n44165 , n44166 , 
     n44167 , n44168 , n44169 , n44170 , n44171 , n44172 , n44173 , n44174 , n44175 , n44176 , 
     n44177 , n44178 , n44179 , n44180 , n44181 , n44182 , n44183 , n44184 , n44185 , n44186 , 
     n44187 , n44188 , n44189 , n44190 , n44191 , n44192 , n44193 , n44194 , n44195 , n44196 , 
     n44197 , n44198 , n44199 , n44200 , n44201 , n44202 , n44203 , n44204 , n44205 , n44206 , 
     n44207 , n44208 , n44209 , n44210 , n44211 , n44212 , n44213 , n44214 , n44215 , n44216 , 
     n44217 , n44218 , n44219 , n44220 , n44221 , n44222 , n44223 , n44224 , n44225 , n44226 , 
     n44227 , n44228 , n44229 , n44230 , n44231 , n44232 , n44233 , n44234 , n44235 , n44236 , 
     n44237 , n44238 , n44239 , n44240 , n44241 , n44242 , n44243 , n44244 , n44245 , n44246 , 
     n44247 , n44248 , n44249 , n44250 , n44251 , n44252 , n44253 , n44254 , n44255 , n44256 , 
     n44257 , n44258 , n44259 , n44260 , n44261 , n44262 , n44263 , n44264 , n44265 , n44266 , 
     n44267 , n44268 , n44269 , n44270 , n44271 , n44272 , n44273 , n44274 , n44275 , n44276 , 
     n44277 , n44278 , n44279 , n44280 , n44281 , n44282 , n44283 , n44284 , n44285 , n44286 , 
     n44287 , n44288 , n44289 , n44290 , n44291 , n44292 , n44293 , n44294 , n44295 , n44296 , 
     n44297 , n44298 , n44299 , n44300 , n44301 , n44302 , n44303 , n44304 , n44305 , n44306 , 
     n44307 , n44308 , n44309 , n44310 , n44311 , n44312 , n44313 , n44314 , n44315 , n44316 , 
     n44317 , n44318 , n44319 , n44320 , n44321 , n44322 , n44323 , n44324 , n44325 , n44326 , 
     n44327 , n44328 , n44329 , n44330 , n44331 , n44332 , n44333 , n44334 , n44335 , n44336 , 
     n44337 , n44338 , n44339 , n44340 , n44341 , n44342 , n44343 , n44344 , n44345 , n44346 , 
     n44347 , n44348 , n44349 , n44350 , n44351 , n44352 , n44353 , n44354 , n44355 , n44356 , 
     n44357 , n44358 , n44359 , n44360 , n44361 , n44362 , n44363 , n44364 , n44365 , n44366 , 
     n44367 , n44368 , n44369 , n44370 , n44371 , n44372 , n44373 , n44374 , n44375 , n44376 , 
     n44377 , n44378 , n44379 , n44380 , n44381 , n44382 , n44383 , n44384 , n44385 , n44386 , 
     n44387 , n44388 , n44389 , n44390 , n44391 , n44392 , n44393 , n44394 , n44395 , n44396 , 
     n44397 , n44398 , n44399 , n44400 , n44401 , n44402 , n44403 , n44404 , n44405 , n44406 , 
     n44407 , n44408 , n44409 , n44410 , n44411 , n44412 , n44413 , n44414 , n44415 , n44416 , 
     n44417 , n44418 , n44419 , n44420 , n44421 , n44422 , n44423 , n44424 , n44425 , n44426 , 
     n44427 , n44428 , n44429 , n44430 , n44431 , n44432 , n44433 , n44434 , n44435 , n44436 , 
     n44437 , n44438 , n44439 , n44440 , n44441 , n44442 , n44443 , n44444 , n44445 , n44446 , 
     n44447 , n44448 , n44449 , n44450 , n44451 , n44452 , n44453 , n44454 , n44455 , n44456 , 
     n44457 , n44458 , n44459 , n44460 , n44461 , n44462 , n44463 , n44464 , n44465 , n44466 , 
     n44467 , n44468 , n44469 , n44470 , n44471 , n44472 , n44473 , n44474 , n44475 , n44476 , 
     n44477 , n44478 , n44479 , n44480 , n44481 , n44482 , n44483 , n44484 , n44485 , n44486 , 
     n44487 , n44488 , n44489 , n44490 , n44491 , n44492 , n44493 , n44494 , n44495 , n44496 , 
     n44497 , n44498 , n44499 , n44500 , n44501 , n44502 , n44503 , n44504 , n44505 , n44506 , 
     n44507 , n44508 , n44509 , n44510 , n44511 , n44512 , n44513 , n44514 , n44515 , n44516 , 
     n44517 , n44518 , n44519 , n44520 , n44521 , n44522 , n44523 , n44524 , n44525 , n44526 , 
     n44527 , n44528 , n44529 , n44530 , n44531 , n44532 , n44533 , n44534 , n44535 , n44536 , 
     n44537 , n44538 , n44539 , n44540 , n44541 , n44542 , n44543 , n44544 , n44545 , n44546 , 
     n44547 , n44548 , n44549 , n44550 , n44551 , n44552 , n44553 , n44554 , n44555 , n44556 , 
     n44557 , n44558 , n44559 , n44560 , n44561 , n44562 , n44563 , n44564 , n44565 , n44566 , 
     n44567 , n44568 , n44569 , n44570 , n44571 , n44572 , n44573 , n44574 , n44575 , n44576 , 
     n44577 , n44578 , n44579 , n44580 , n44581 , n44582 , n44583 , n44584 , n44585 , n44586 , 
     n44587 , n44588 , n44589 , n44590 , n44591 , n44592 , n44593 , n44594 , n44595 , n44596 , 
     n44597 , n44598 , n44599 , n44600 , n44601 , n44602 , n44603 , n44604 , n44605 , n44606 , 
     n44607 , n44608 , n44609 , n44610 , n44611 , n44612 , n44613 , n44614 , n44615 , n44616 , 
     n44617 , n44618 , n44619 , n44620 , n44621 , n44622 , n44623 , n44624 , n44625 , n44626 , 
     n44627 , n44628 , n44629 , n44630 , n44631 , n44632 , n44633 , n44634 , n44635 , n44636 , 
     n44637 , n44638 , n44639 , n44640 , n44641 , n44642 , n44643 , n44644 , n44645 , n44646 , 
     n44647 , n44648 , n44649 , n44650 , n44651 , n44652 , n44653 , n44654 , n44655 , n44656 , 
     n44657 , n44658 , n44659 , n44660 , n44661 , n44662 , n44663 , n44664 , n44665 , n44666 , 
     n44667 , n44668 , n44669 , n44670 , n44671 , n44672 , n44673 , n44674 , n44675 , n44676 , 
     n44677 , n44678 , n44679 , n44680 , n44681 , n44682 , n44683 , n44684 , n44685 , n44686 , 
     n44687 , n44688 , n44689 , n44690 , n44691 , n44692 , n44693 , n44694 , n44695 , n44696 , 
     n44697 , n44698 , n44699 , n44700 , n44701 , n44702 , n44703 , n44704 , n44705 , n44706 , 
     n44707 , n44708 , n44709 , n44710 , n44711 , n44712 , n44713 , n44714 , n44715 , n44716 , 
     n44717 , n44718 , n44719 , n44720 , n44721 , n44722 , n44723 , n44724 , n44725 , n44726 , 
     n44727 , n44728 , n44729 , n44730 , n44731 , n44732 , n44733 , n44734 , n44735 , n44736 , 
     n44737 , n44738 , n44739 , n44740 , n44741 , n44742 , n44743 , n44744 , n44745 , n44746 , 
     n44747 , n44748 , n44749 , n44750 , n44751 , n44752 , n44753 , n44754 , n44755 , n44756 , 
     n44757 , n44758 , n44759 , n44760 , n44761 , n44762 , n44763 , n44764 , n44765 , n44766 , 
     n44767 , n44768 , n44769 , n44770 , n44771 , n44772 , n44773 , n44774 , n44775 , n44776 , 
     n44777 , n44778 , n44779 , n44780 , n44781 , n44782 , n44783 , n44784 , n44785 , n44786 , 
     n44787 , n44788 , n44789 , n44790 , n44791 , n44792 , n44793 , n44794 , n44795 , n44796 , 
     n44797 , n44798 , n44799 , n44800 , n44801 , n44802 , n44803 , n44804 , n44805 , n44806 , 
     n44807 , n44808 , n44809 , n44810 , n44811 , n44812 , n44813 , n44814 , n44815 , n44816 , 
     n44817 , n44818 , n44819 , n44820 , n44821 , n44822 , n44823 , n44824 , n44825 , n44826 , 
     n44827 , n44828 , n44829 , n44830 , n44831 , n44832 , n44833 , n44834 , n44835 , n44836 , 
     n44837 , n44838 , n44839 , n44840 , n44841 , n44842 , n44843 , n44844 , n44845 , n44846 , 
     n44847 , n44848 , n44849 , n44850 , n44851 , n44852 , n44853 , n44854 , n44855 , n44856 , 
     n44857 , n44858 , n44859 , n44860 , n44861 , n44862 , n44863 , n44864 , n44865 , n44866 , 
     n44867 , n44868 , n44869 , n44870 , n44871 , n44872 , n44873 , n44874 , n44875 , n44876 , 
     n44877 , n44878 , n44879 , n44880 , n44881 , n44882 , n44883 , n44884 , n44885 , n44886 , 
     n44887 , n44888 , n44889 , n44890 , n44891 , n44892 , n44893 , n44894 , n44895 , n44896 , 
     n44897 , n44898 , n44899 , n44900 , n44901 , n44902 , n44903 , n44904 , n44905 , n44906 , 
     n44907 , n44908 , n44909 , n44910 , n44911 , n44912 , n44913 , n44914 , n44915 , n44916 , 
     n44917 , n44918 , n44919 , n44920 , n44921 , n44922 , n44923 , n44924 , n44925 , n44926 , 
     n44927 , n44928 , n44929 , n44930 , n44931 , n44932 , n44933 , n44934 , n44935 , n44936 , 
     n44937 , n44938 , n44939 , n44940 , n44941 , n44942 , n44943 , n44944 , n44945 , n44946 , 
     n44947 , n44948 , n44949 , n44950 , n44951 , n44952 , n44953 , n44954 , n44955 , n44956 , 
     n44957 , n44958 , n44959 , n44960 , n44961 , n44962 , n44963 , n44964 , n44965 , n44966 , 
     n44967 , n44968 , n44969 , n44970 , n44971 , n44972 , n44973 , n44974 , n44975 , n44976 , 
     n44977 , n44978 , n44979 , n44980 , n44981 , n44982 , n44983 , n44984 , n44985 , n44986 , 
     n44987 , n44988 , n44989 , n44990 , n44991 , n44992 , n44993 , n44994 , n44995 , n44996 , 
     n44997 , n44998 , n44999 , n45000 , n45001 , n45002 , n45003 , n45004 , n45005 , n45006 , 
     n45007 , n45008 , n45009 , n45010 , n45011 , n45012 , n45013 , n45014 , n45015 , n45016 , 
     n45017 , n45018 , n45019 , n45020 , n45021 , n45022 , n45023 , n45024 , n45025 , n45026 , 
     n45027 , n45028 , n45029 , n45030 , n45031 , n45032 , n45033 , n45034 , n45035 , n45036 , 
     n45037 , n45038 , n45039 , n45040 , n45041 , n45042 , n45043 , n45044 , n45045 , n45046 , 
     n45047 , n45048 , n45049 , n45050 , n45051 , n45052 , n45053 , n45054 , n45055 , n45056 , 
     n45057 , n45058 , n45059 , n45060 , n45061 , n45062 , n45063 , n45064 , n45065 , n45066 , 
     n45067 , n45068 , n45069 , n45070 , n45071 , n45072 , n45073 , n45074 , n45075 , n45076 , 
     n45077 , n45078 , n45079 , n45080 , n45081 , n45082 , n45083 , n45084 , n45085 , n45086 , 
     n45087 , n45088 , n45089 , n45090 , n45091 , n45092 , n45093 , n45094 , n45095 , n45096 , 
     n45097 , n45098 , n45099 , n45100 , n45101 , n45102 , n45103 , n45104 , n45105 , n45106 , 
     n45107 , n45108 , n45109 , n45110 , n45111 , n45112 , n45113 , n45114 , n45115 , n45116 , 
     n45117 , n45118 , n45119 , n45120 , n45121 , n45122 , n45123 , n45124 , n45125 , n45126 , 
     n45127 , n45128 , n45129 , n45130 , n45131 , n45132 , n45133 , n45134 , n45135 , n45136 , 
     n45137 , n45138 , n45139 , n45140 , n45141 , n45142 , n45143 , n45144 , n45145 , n45146 , 
     n45147 , n45148 , n45149 , n45150 , n45151 , n45152 , n45153 , n45154 , n45155 , n45156 , 
     n45157 , n45158 , n45159 , n45160 , n45161 , n45162 , n45163 , n45164 , n45165 , n45166 , 
     n45167 , n45168 , n45169 , n45170 , n45171 , n45172 , n45173 , n45174 , n45175 , n45176 , 
     n45177 , n45178 , n45179 , n45180 , n45181 , n45182 , n45183 , n45184 , n45185 , n45186 , 
     n45187 , n45188 , n45189 , n45190 , n45191 , n45192 , n45193 , n45194 , n45195 , n45196 , 
     n45197 , n45198 , n45199 , n45200 , n45201 , n45202 , n45203 , n45204 , n45205 , n45206 , 
     n45207 , n45208 , n45209 , n45210 , n45211 , n45212 , n45213 , n45214 , n45215 , n45216 , 
     n45217 , n45218 , n45219 , n45220 , n45221 , n45222 , n45223 , n45224 , n45225 , n45226 , 
     n45227 , n45228 , n45229 , n45230 , n45231 , n45232 , n45233 , n45234 , n45235 , n45236 , 
     n45237 , n45238 , n45239 , n45240 , n45241 , n45242 , n45243 , n45244 , n45245 , n45246 , 
     n45247 , n45248 , n45249 , n45250 , n45251 , n45252 , n45253 , n45254 , n45255 , n45256 , 
     n45257 , n45258 , n45259 , n45260 , n45261 , n45262 , n45263 , n45264 , n45265 , n45266 , 
     n45267 , n45268 , n45269 , n45270 , n45271 , n45272 , n45273 , n45274 , n45275 , n45276 , 
     n45277 , n45278 , n45279 , n45280 , n45281 , n45282 , n45283 , n45284 , n45285 , n45286 , 
     n45287 , n45288 , n45289 , n45290 , n45291 , n45292 , n45293 , n45294 , n45295 , n45296 , 
     n45297 , n45298 , n45299 , n45300 , n45301 , n45302 , n45303 , n45304 , n45305 , n45306 , 
     n45307 , n45308 , n45309 , n45310 , n45311 , n45312 , n45313 , n45314 , n45315 , n45316 , 
     n45317 , n45318 , n45319 , n45320 , n45321 , n45322 , n45323 , n45324 , n45325 , n45326 , 
     n45327 , n45328 , n45329 , n45330 , n45331 , n45332 , n45333 , n45334 , n45335 , n45336 , 
     n45337 , n45338 , n45339 , n45340 , n45341 , n45342 , n45343 , n45344 , n45345 , n45346 , 
     n45347 , n45348 , n45349 , n45350 , n45351 , n45352 , n45353 , n45354 , n45355 , n45356 , 
     n45357 , n45358 , n45359 , n45360 , n45361 , n45362 , n45363 , n45364 , n45365 , n45366 , 
     n45367 , n45368 , n45369 , n45370 , n45371 , n45372 , n45373 , n45374 , n45375 , n45376 , 
     n45377 , n45378 , n45379 , n45380 , n45381 , n45382 , n45383 , n45384 , n45385 , n45386 , 
     n45387 , n45388 , n45389 , n45390 , n45391 , n45392 , n45393 , n45394 , n45395 , n45396 , 
     n45397 , n45398 , n45399 , n45400 , n45401 , n45402 , n45403 , n45404 , n45405 , n45406 , 
     n45407 , n45408 , n45409 , n45410 , n45411 , n45412 , n45413 , n45414 , n45415 , n45416 , 
     n45417 , n45418 , n45419 , n45420 , n45421 , n45422 , n45423 , n45424 , n45425 , n45426 , 
     n45427 , n45428 , n45429 , n45430 , n45431 , n45432 , n45433 , n45434 , n45435 , n45436 , 
     n45437 , n45438 , n45439 , n45440 , n45441 , n45442 , n45443 , n45444 , n45445 , n45446 , 
     n45447 , n45448 , n45449 , n45450 , n45451 , n45452 , n45453 , n45454 , n45455 , n45456 , 
     n45457 , n45458 , n45459 , n45460 , n45461 , n45462 , n45463 , n45464 , n45465 , n45466 , 
     n45467 , n45468 , n45469 , n45470 , n45471 , n45472 , n45473 , n45474 , n45475 , n45476 , 
     n45477 , n45478 , n45479 , n45480 , n45481 , n45482 , n45483 , n45484 , n45485 , n45486 , 
     n45487 , n45488 , n45489 , n45490 , n45491 , n45492 , n45493 , n45494 , n45495 , n45496 , 
     n45497 , n45498 , n45499 , n45500 , n45501 , n45502 , n45503 , n45504 , n45505 , n45506 , 
     n45507 , n45508 , n45509 , n45510 , n45511 , n45512 , n45513 , n45514 , n45515 , n45516 , 
     n45517 , n45518 , n45519 , n45520 , n45521 , n45522 , n45523 , n45524 , n45525 , n45526 , 
     n45527 , n45528 , n45529 , n45530 , n45531 , n45532 , n45533 , n45534 , n45535 , n45536 , 
     n45537 , n45538 , n45539 , n45540 , n45541 , n45542 , n45543 , n45544 , n45545 , n45546 , 
     n45547 , n45548 , n45549 , n45550 , n45551 , n45552 , n45553 , n45554 , n45555 , n45556 , 
     n45557 , n45558 , n45559 , n45560 , n45561 , n45562 , n45563 , n45564 , n45565 , n45566 , 
     n45567 , n45568 , n45569 , n45570 , n45571 , n45572 , n45573 , n45574 , n45575 , n45576 , 
     n45577 , n45578 , n45579 , n45580 , n45581 , n45582 , n45583 , n45584 , n45585 , n45586 , 
     n45587 , n45588 , n45589 , n45590 , n45591 , n45592 , n45593 , n45594 , n45595 , n45596 , 
     n45597 , n45598 , n45599 , n45600 , n45601 , n45602 , n45603 , n45604 , n45605 , n45606 , 
     n45607 , n45608 , n45609 , n45610 , n45611 , n45612 , n45613 , n45614 , n45615 , n45616 , 
     n45617 , n45618 , n45619 , n45620 , n45621 , n45622 , n45623 , n45624 , n45625 , n45626 , 
     n45627 , n45628 , n45629 , n45630 , n45631 , n45632 , n45633 , n45634 , n45635 , n45636 , 
     n45637 , n45638 , n45639 , n45640 , n45641 , n45642 , n45643 , n45644 , n45645 , n45646 , 
     n45647 , n45648 , n45649 , n45650 , n45651 , n45652 , n45653 , n45654 , n45655 , n45656 , 
     n45657 , n45658 , n45659 , n45660 , n45661 , n45662 , n45663 , n45664 , n45665 , n45666 , 
     n45667 , n45668 , n45669 , n45670 , n45671 , n45672 , n45673 , n45674 , n45675 , n45676 , 
     n45677 , n45678 , n45679 , n45680 , n45681 , n45682 , n45683 , n45684 , n45685 , n45686 , 
     n45687 , n45688 , n45689 , n45690 , n45691 , n45692 , n45693 , n45694 , n45695 , n45696 , 
     n45697 , n45698 , n45699 , n45700 , n45701 , n45702 , n45703 , n45704 , n45705 , n45706 , 
     n45707 , n45708 , n45709 , n45710 , n45711 , n45712 , n45713 , n45714 , n45715 , n45716 , 
     n45717 , n45718 , n45719 , n45720 , n45721 , n45722 , n45723 , n45724 , n45725 , n45726 , 
     n45727 , n45728 , n45729 , n45730 , n45731 , n45732 , n45733 , n45734 , n45735 , n45736 , 
     n45737 , n45738 , n45739 , n45740 , n45741 , n45742 , n45743 , n45744 , n45745 , n45746 , 
     n45747 , n45748 , n45749 , n45750 , n45751 , n45752 , n45753 , n45754 , n45755 , n45756 , 
     n45757 , n45758 , n45759 , n45760 , n45761 , n45762 , n45763 , n45764 , n45765 , n45766 , 
     n45767 , n45768 , n45769 , n45770 , n45771 , n45772 , n45773 , n45774 , n45775 , n45776 , 
     n45777 , n45778 , n45779 , n45780 , n45781 , n45782 , n45783 , n45784 , n45785 , n45786 , 
     n45787 , n45788 , n45789 , n45790 , n45791 , n45792 , n45793 , n45794 , n45795 , n45796 , 
     n45797 , n45798 , n45799 , n45800 , n45801 , n45802 , n45803 , n45804 , n45805 , n45806 , 
     n45807 , n45808 , n45809 , n45810 , n45811 , n45812 , n45813 , n45814 , n45815 , n45816 , 
     n45817 , n45818 , n45819 , n45820 , n45821 , n45822 , n45823 , n45824 , n45825 , n45826 , 
     n45827 , n45828 , n45829 , n45830 , n45831 , n45832 , n45833 , n45834 , n45835 , n45836 , 
     n45837 , n45838 , n45839 , n45840 , n45841 , n45842 , n45843 , n45844 , n45845 , n45846 , 
     n45847 , n45848 , n45849 , n45850 , n45851 , n45852 , n45853 , n45854 , n45855 , n45856 , 
     n45857 , n45858 , n45859 , n45860 , n45861 , n45862 , n45863 , n45864 , n45865 , n45866 , 
     n45867 , n45868 , n45869 , n45870 , n45871 , n45872 , n45873 , n45874 , n45875 , n45876 , 
     n45877 , n45878 , n45879 , n45880 , n45881 , n45882 , n45883 , n45884 , n45885 , n45886 , 
     n45887 , n45888 , n45889 , n45890 , n45891 , n45892 , n45893 , n45894 , n45895 , n45896 , 
     n45897 , n45898 , n45899 , n45900 , n45901 , n45902 , n45903 , n45904 , n45905 , n45906 , 
     n45907 , n45908 , n45909 , n45910 , n45911 , n45912 , n45913 , n45914 , n45915 , n45916 , 
     n45917 , n45918 , n45919 , n45920 , n45921 , n45922 , n45923 , n45924 , n45925 , n45926 , 
     n45927 , n45928 , n45929 , n45930 , n45931 , n45932 , n45933 , n45934 , n45935 , n45936 , 
     n45937 , n45938 , n45939 , n45940 , n45941 , n45942 , n45943 , n45944 , n45945 , n45946 , 
     n45947 , n45948 , n45949 , n45950 , n45951 , n45952 , n45953 , n45954 , n45955 , n45956 , 
     n45957 , n45958 , n45959 , n45960 , n45961 , n45962 , n45963 , n45964 , n45965 , n45966 , 
     n45967 , n45968 , n45969 , n45970 , n45971 , n45972 , n45973 , n45974 , n45975 , n45976 , 
     n45977 , n45978 , n45979 , n45980 , n45981 , n45982 , n45983 , n45984 , n45985 , n45986 , 
     n45987 , n45988 , n45989 , n45990 , n45991 , n45992 , n45993 , n45994 , n45995 , n45996 , 
     n45997 , n45998 , n45999 , n46000 , n46001 , n46002 , n46003 , n46004 , n46005 , n46006 , 
     n46007 , n46008 , n46009 , n46010 , n46011 , n46012 , n46013 , n46014 , n46015 , n46016 , 
     n46017 , n46018 , n46019 , n46020 , n46021 , n46022 , n46023 , n46024 , n46025 , n46026 , 
     n46027 , n46028 , n46029 , n46030 , n46031 , n46032 , n46033 , n46034 , n46035 , n46036 , 
     n46037 , n46038 , n46039 , n46040 , n46041 , n46042 , n46043 , n46044 , n46045 , n46046 , 
     n46047 , n46048 , n46049 , n46050 , n46051 , n46052 , n46053 , n46054 , n46055 , n46056 , 
     n46057 , n46058 , n46059 , n46060 , n46061 , n46062 , n46063 , n46064 , n46065 , n46066 , 
     n46067 , n46068 , n46069 , n46070 , n46071 , n46072 , n46073 , n46074 , n46075 , n46076 , 
     n46077 , n46078 , n46079 , n46080 , n46081 , n46082 , n46083 , n46084 , n46085 , n46086 , 
     n46087 , n46088 , n46089 , n46090 , n46091 , n46092 , n46093 , n46094 , n46095 , n46096 , 
     n46097 , n46098 , n46099 , n46100 , n46101 , n46102 , n46103 , n46104 , n46105 , n46106 , 
     n46107 , n46108 , n46109 , n46110 , n46111 , n46112 , n46113 , n46114 , n46115 , n46116 , 
     n46117 , n46118 , n46119 , n46120 , n46121 , n46122 , n46123 , n46124 , n46125 , n46126 , 
     n46127 , n46128 , n46129 , n46130 , n46131 , n46132 , n46133 , n46134 , n46135 , n46136 , 
     n46137 , n46138 , n46139 , n46140 , n46141 , n46142 , n46143 , n46144 , n46145 , n46146 , 
     n46147 , n46148 , n46149 , n46150 , n46151 , n46152 , n46153 , n46154 , n46155 , n46156 , 
     n46157 , n46158 , n46159 , n46160 , n46161 , n46162 , n46163 , n46164 , n46165 , n46166 , 
     n46167 , n46168 , n46169 , n46170 , n46171 , n46172 , n46173 , n46174 , n46175 , n46176 , 
     n46177 , n46178 , n46179 , n46180 , n46181 , n46182 , n46183 , n46184 , n46185 , n46186 , 
     n46187 , n46188 , n46189 , n46190 , n46191 , n46192 , n46193 , n46194 , n46195 , n46196 , 
     n46197 , n46198 , n46199 , n46200 , n46201 , n46202 , n46203 , n46204 , n46205 , n46206 , 
     n46207 , n46208 , n46209 , n46210 , n46211 , n46212 , n46213 , n46214 , n46215 , n46216 , 
     n46217 , n46218 , n46219 , n46220 , n46221 , n46222 , n46223 , n46224 , n46225 , n46226 , 
     n46227 , n46228 , n46229 , n46230 , n46231 , n46232 , n46233 , n46234 , n46235 , n46236 , 
     n46237 , n46238 , n46239 , n46240 , n46241 , n46242 , n46243 , n46244 , n46245 , n46246 , 
     n46247 , n46248 , n46249 , n46250 , n46251 , n46252 , n46253 , n46254 , n46255 , n46256 , 
     n46257 , n46258 , n46259 , n46260 , n46261 , n46262 , n46263 , n46264 , n46265 , n46266 , 
     n46267 , n46268 , n46269 , n46270 , n46271 , n46272 , n46273 , n46274 , n46275 , n46276 , 
     n46277 , n46278 , n46279 , n46280 , n46281 , n46282 , n46283 , n46284 , n46285 , n46286 , 
     n46287 , n46288 , n46289 , n46290 , n46291 , n46292 , n46293 , n46294 , n46295 , n46296 , 
     n46297 , n46298 , n46299 , n46300 , n46301 , n46302 , n46303 , n46304 , n46305 , n46306 , 
     n46307 , n46308 , n46309 , n46310 , n46311 , n46312 , n46313 , n46314 , n46315 , n46316 , 
     n46317 , n46318 , n46319 , n46320 , n46321 , n46322 , n46323 , n46324 , n46325 , n46326 , 
     n46327 , n46328 , n46329 , n46330 , n46331 , n46332 , n46333 , n46334 , n46335 , n46336 , 
     n46337 , n46338 , n46339 , n46340 , n46341 , n46342 , n46343 , n46344 , n46345 , n46346 , 
     n46347 , n46348 , n46349 , n46350 , n46351 , n46352 , n46353 , n46354 , n46355 , n46356 , 
     n46357 , n46358 , n46359 , n46360 , n46361 , n46362 , n46363 , n46364 , n46365 , n46366 , 
     n46367 , n46368 , n46369 , n46370 , n46371 , n46372 , n46373 , n46374 , n46375 , n46376 , 
     n46377 , n46378 , n46379 , n46380 , n46381 , n46382 , n46383 , n46384 , n46385 , n46386 , 
     n46387 , n46388 , n46389 , n46390 , n46391 , n46392 , n46393 , n46394 , n46395 , n46396 , 
     n46397 , n46398 , n46399 , n46400 , n46401 , n46402 , n46403 , n46404 , n46405 , n46406 , 
     n46407 , n46408 , n46409 , n46410 , n46411 , n46412 , n46413 , n46414 , n46415 , n46416 , 
     n46417 , n46418 , n46419 , n46420 , n46421 , n46422 , n46423 , n46424 , n46425 , n46426 , 
     n46427 , n46428 , n46429 , n46430 , n46431 , n46432 , n46433 , n46434 , n46435 , n46436 , 
     n46437 , n46438 , n46439 , n46440 , n46441 , n46442 , n46443 , n46444 , n46445 , n46446 , 
     n46447 , n46448 , n46449 , n46450 , n46451 , n46452 , n46453 , n46454 , n46455 , n46456 , 
     n46457 , n46458 , n46459 , n46460 , n46461 , n46462 , n46463 , n46464 , n46465 , n46466 , 
     n46467 , n46468 , n46469 , n46470 , n46471 , n46472 , n46473 , n46474 , n46475 , n46476 , 
     n46477 , n46478 , n46479 , n46480 , n46481 , n46482 , n46483 , n46484 , n46485 , n46486 , 
     n46487 , n46488 , n46489 , n46490 , n46491 , n46492 , n46493 , n46494 , n46495 , n46496 , 
     n46497 , n46498 , n46499 , n46500 , n46501 , n46502 , n46503 , n46504 , n46505 , n46506 , 
     n46507 , n46508 , n46509 , n46510 , n46511 , n46512 , n46513 , n46514 , n46515 , n46516 , 
     n46517 , n46518 , n46519 , n46520 , n46521 , n46522 , n46523 , n46524 , n46525 , n46526 , 
     n46527 , n46528 , n46529 , n46530 , n46531 , n46532 , n46533 , n46534 , n46535 , n46536 , 
     n46537 , n46538 , n46539 , n46540 , n46541 , n46542 , n46543 , n46544 , n46545 , n46546 , 
     n46547 , n46548 , n46549 , n46550 , n46551 , n46552 , n46553 , n46554 , n46555 , n46556 , 
     n46557 , n46558 , n46559 , n46560 , n46561 , n46562 , n46563 , n46564 , n46565 , n46566 , 
     n46567 , n46568 , n46569 , n46570 , n46571 , n46572 , n46573 , n46574 , n46575 , n46576 , 
     n46577 , n46578 , n46579 , n46580 , n46581 , n46582 , n46583 , n46584 , n46585 , n46586 , 
     n46587 , n46588 , n46589 , n46590 , n46591 , n46592 , n46593 , n46594 , n46595 , n46596 , 
     n46597 , n46598 , n46599 , n46600 , n46601 , n46602 , n46603 , n46604 , n46605 , n46606 , 
     n46607 , n46608 , n46609 , n46610 , n46611 , n46612 , n46613 , n46614 , n46615 , n46616 , 
     n46617 , n46618 , n46619 , n46620 , n46621 , n46622 , n46623 , n46624 , n46625 , n46626 , 
     n46627 , n46628 , n46629 , n46630 , n46631 , n46632 , n46633 , n46634 , n46635 , n46636 , 
     n46637 , n46638 , n46639 , n46640 , n46641 , n46642 , n46643 , n46644 , n46645 , n46646 , 
     n46647 , n46648 , n46649 , n46650 , n46651 , n46652 , n46653 , n46654 , n46655 , n46656 , 
     n46657 , n46658 , n46659 , n46660 , n46661 , n46662 , n46663 , n46664 , n46665 , n46666 , 
     n46667 , n46668 , n46669 , n46670 , n46671 , n46672 , n46673 , n46674 , n46675 , n46676 , 
     n46677 , n46678 , n46679 , n46680 , n46681 , n46682 , n46683 , n46684 , n46685 , n46686 , 
     n46687 , n46688 , n46689 , n46690 , n46691 , n46692 , n46693 , n46694 , n46695 , n46696 , 
     n46697 , n46698 , n46699 , n46700 , n46701 , n46702 , n46703 , n46704 , n46705 , n46706 , 
     n46707 , n46708 , n46709 , n46710 , n46711 , n46712 , n46713 , n46714 , n46715 , n46716 , 
     n46717 , n46718 , n46719 , n46720 , n46721 , n46722 , n46723 , n46724 , n46725 , n46726 , 
     n46727 , n46728 , n46729 , n46730 , n46731 , n46732 , n46733 , n46734 , n46735 , n46736 , 
     n46737 , n46738 , n46739 , n46740 , n46741 , n46742 , n46743 , n46744 , n46745 , n46746 , 
     n46747 , n46748 , n46749 , n46750 , n46751 , n46752 , n46753 , n46754 , n46755 , n46756 , 
     n46757 , n46758 , n46759 , n46760 , n46761 , n46762 , n46763 , n46764 , n46765 , n46766 , 
     n46767 , n46768 , n46769 , n46770 , n46771 , n46772 , n46773 , n46774 , n46775 , n46776 , 
     n46777 , n46778 , n46779 , n46780 , n46781 , n46782 , n46783 , n46784 , n46785 , n46786 , 
     n46787 , n46788 , n46789 , n46790 , n46791 , n46792 , n46793 , n46794 , n46795 , n46796 , 
     n46797 , n46798 , n46799 , n46800 , n46801 , n46802 , n46803 , n46804 , n46805 , n46806 , 
     n46807 , n46808 , n46809 , n46810 , n46811 , n46812 , n46813 , n46814 , n46815 , n46816 , 
     n46817 , n46818 , n46819 , n46820 , n46821 , n46822 , n46823 , n46824 , n46825 , n46826 , 
     n46827 , n46828 , n46829 , n46830 , n46831 , n46832 , n46833 , n46834 , n46835 , n46836 , 
     n46837 , n46838 , n46839 , n46840 , n46841 , n46842 , n46843 , n46844 , n46845 , n46846 , 
     n46847 , n46848 , n46849 , n46850 , n46851 , n46852 , n46853 , n46854 , n46855 , n46856 , 
     n46857 , n46858 , n46859 , n46860 , n46861 , n46862 , n46863 , n46864 , n46865 , n46866 , 
     n46867 , n46868 , n46869 , n46870 , n46871 , n46872 , n46873 , n46874 , n46875 , n46876 , 
     n46877 , n46878 , n46879 , n46880 , n46881 , n46882 , n46883 , n46884 , n46885 , n46886 , 
     n46887 , n46888 , n46889 , n46890 , n46891 , n46892 , n46893 , n46894 , n46895 , n46896 , 
     n46897 , n46898 , n46899 , n46900 , n46901 , n46902 , n46903 , n46904 , n46905 , n46906 , 
     n46907 , n46908 , n46909 , n46910 , n46911 , n46912 , n46913 , n46914 , n46915 , n46916 , 
     n46917 , n46918 , n46919 , n46920 , n46921 , n46922 , n46923 , n46924 , n46925 , n46926 , 
     n46927 , n46928 , n46929 , n46930 , n46931 , n46932 , n46933 , n46934 , n46935 , n46936 , 
     n46937 , n46938 , n46939 , n46940 , n46941 , n46942 , n46943 , n46944 , n46945 , n46946 , 
     n46947 , n46948 , n46949 , n46950 , n46951 , n46952 , n46953 , n46954 , n46955 , n46956 , 
     n46957 , n46958 , n46959 , n46960 , n46961 , n46962 , n46963 , n46964 , n46965 , n46966 , 
     n46967 , n46968 , n46969 , n46970 , n46971 , n46972 , n46973 , n46974 , n46975 , n46976 , 
     n46977 , n46978 , n46979 , n46980 , n46981 , n46982 , n46983 , n46984 , n46985 , n46986 , 
     n46987 , n46988 , n46989 , n46990 , n46991 , n46992 , n46993 , n46994 , n46995 , n46996 , 
     n46997 , n46998 , n46999 , n47000 , n47001 , n47002 , n47003 , n47004 , n47005 , n47006 , 
     n47007 , n47008 , n47009 , n47010 , n47011 , n47012 , n47013 , n47014 , n47015 , n47016 , 
     n47017 , n47018 , n47019 , n47020 , n47021 , n47022 , n47023 , n47024 , n47025 , n47026 , 
     n47027 , n47028 , n47029 , n47030 , n47031 , n47032 , n47033 , n47034 , n47035 , n47036 , 
     n47037 , n47038 , n47039 , n47040 , n47041 , n47042 , n47043 , n47044 , n47045 , n47046 , 
     n47047 , n47048 , n47049 , n47050 , n47051 , n47052 , n47053 , n47054 , n47055 , n47056 , 
     n47057 , n47058 , n47059 , n47060 , n47061 , n47062 , n47063 , n47064 , n47065 , n47066 , 
     n47067 , n47068 , n47069 , n47070 , n47071 , n47072 , n47073 , n47074 , n47075 , n47076 , 
     n47077 , n47078 , n47079 , n47080 , n47081 , n47082 , n47083 , n47084 , n47085 , n47086 , 
     n47087 , n47088 , n47089 , n47090 , n47091 , n47092 , n47093 , n47094 , n47095 , n47096 , 
     n47097 , n47098 , n47099 , n47100 , n47101 , n47102 , n47103 , n47104 , n47105 , n47106 , 
     n47107 , n47108 , n47109 , n47110 , n47111 , n47112 , n47113 , n47114 , n47115 , n47116 , 
     n47117 , n47118 , n47119 , n47120 , n47121 , n47122 , n47123 , n47124 , n47125 , n47126 , 
     n47127 , n47128 , n47129 , n47130 , n47131 , n47132 , n47133 , n47134 , n47135 , n47136 , 
     n47137 , n47138 , n47139 , n47140 , n47141 , n47142 , n47143 , n47144 , n47145 , n47146 , 
     n47147 , n47148 , n47149 , n47150 , n47151 , n47152 , n47153 , n47154 , n47155 , n47156 , 
     n47157 , n47158 , n47159 , n47160 , n47161 , n47162 , n47163 , n47164 , n47165 , n47166 , 
     n47167 , n47168 , n47169 , n47170 , n47171 , n47172 , n47173 , n47174 , n47175 , n47176 , 
     n47177 , n47178 , n47179 , n47180 , n47181 , n47182 , n47183 , n47184 , n47185 , n47186 , 
     n47187 , n47188 , n47189 , n47190 , n47191 , n47192 , n47193 , n47194 , n47195 , n47196 , 
     n47197 , n47198 , n47199 , n47200 , n47201 , n47202 , n47203 , n47204 , n47205 , n47206 , 
     n47207 , n47208 , n47209 , n47210 , n47211 , n47212 , n47213 , n47214 , n47215 , n47216 , 
     n47217 , n47218 , n47219 , n47220 , n47221 , n47222 , n47223 , n47224 , n47225 , n47226 , 
     n47227 , n47228 , n47229 , n47230 , n47231 , n47232 , n47233 , n47234 , n47235 , n47236 , 
     n47237 , n47238 , n47239 , n47240 , n47241 , n47242 , n47243 , n47244 , n47245 , n47246 , 
     n47247 , n47248 , n47249 , n47250 , n47251 , n47252 , n47253 , n47254 , n47255 , n47256 , 
     n47257 , n47258 , n47259 , n47260 , n47261 , n47262 , n47263 , n47264 , n47265 , n47266 , 
     n47267 , n47268 , n47269 , n47270 , n47271 , n47272 , n47273 , n47274 , n47275 , n47276 , 
     n47277 , n47278 , n47279 , n47280 , n47281 , n47282 , n47283 , n47284 , n47285 , n47286 , 
     n47287 , n47288 , n47289 , n47290 , n47291 , n47292 , n47293 , n47294 , n47295 , n47296 , 
     n47297 , n47298 , n47299 , n47300 , n47301 , n47302 , n47303 , n47304 , n47305 , n47306 , 
     n47307 , n47308 , n47309 , n47310 , n47311 , n47312 , n47313 , n47314 , n47315 , n47316 , 
     n47317 , n47318 , n47319 , n47320 , n47321 , n47322 , n47323 , n47324 , n47325 , n47326 , 
     n47327 , n47328 , n47329 , n47330 , n47331 , n47332 , n47333 , n47334 , n47335 , n47336 , 
     n47337 , n47338 , n47339 , n47340 , n47341 , n47342 , n47343 , n47344 , n47345 , n47346 , 
     n47347 , n47348 , n47349 , n47350 , n47351 , n47352 , n47353 , n47354 , n47355 , n47356 , 
     n47357 , n47358 , n47359 , n47360 , n47361 , n47362 , n47363 , n47364 , n47365 , n47366 , 
     n47367 , n47368 , n47369 , n47370 , n47371 , n47372 , n47373 , n47374 , n47375 , n47376 , 
     n47377 , n47378 , n47379 , n47380 , n47381 , n47382 , n47383 , n47384 , n47385 , n47386 , 
     n47387 , n47388 , n47389 , n47390 , n47391 , n47392 , n47393 , n47394 , n47395 , n47396 , 
     n47397 , n47398 , n47399 , n47400 , n47401 , n47402 , n47403 , n47404 , n47405 , n47406 , 
     n47407 , n47408 , n47409 , n47410 , n47411 , n47412 , n47413 , n47414 , n47415 , n47416 , 
     n47417 , n47418 , n47419 , n47420 , n47421 , n47422 , n47423 , n47424 , n47425 , n47426 , 
     n47427 , n47428 , n47429 , n47430 , n47431 , n47432 , n47433 , n47434 , n47435 , n47436 , 
     n47437 , n47438 , n47439 , n47440 , n47441 , n47442 , n47443 , n47444 , n47445 , n47446 , 
     n47447 , n47448 , n47449 , n47450 , n47451 , n47452 , n47453 , n47454 , n47455 , n47456 , 
     n47457 , n47458 , n47459 , n47460 , n47461 , n47462 , n47463 , n47464 , n47465 , n47466 , 
     n47467 , n47468 , n47469 , n47470 , n47471 , n47472 , n47473 , n47474 , n47475 , n47476 , 
     n47477 , n47478 , n47479 , n47480 , n47481 , n47482 , n47483 , n47484 , n47485 , n47486 , 
     n47487 , n47488 , n47489 , n47490 , n47491 , n47492 , n47493 , n47494 , n47495 , n47496 , 
     n47497 , n47498 , n47499 , n47500 , n47501 , n47502 , n47503 , n47504 , n47505 , n47506 , 
     n47507 , n47508 , n47509 , n47510 , n47511 , n47512 , n47513 , n47514 , n47515 , n47516 , 
     n47517 , n47518 , n47519 , n47520 , n47521 , n47522 , n47523 , n47524 , n47525 , n47526 , 
     n47527 , n47528 , n47529 , n47530 , n47531 , n47532 , n47533 , n47534 , n47535 , n47536 , 
     n47537 , n47538 , n47539 , n47540 , n47541 , n47542 , n47543 , n47544 , n47545 , n47546 , 
     n47547 , n47548 , n47549 , n47550 , n47551 , n47552 , n47553 , n47554 , n47555 , n47556 , 
     n47557 , n47558 , n47559 , n47560 , n47561 , n47562 , n47563 , n47564 , n47565 , n47566 , 
     n47567 , n47568 , n47569 , n47570 , n47571 , n47572 , n47573 , n47574 , n47575 , n47576 , 
     n47577 , n47578 , n47579 , n47580 , n47581 , n47582 , n47583 , n47584 , n47585 , n47586 , 
     n47587 , n47588 , n47589 , n47590 , n47591 , n47592 , n47593 , n47594 , n47595 , n47596 , 
     n47597 , n47598 , n47599 , n47600 , n47601 , n47602 , n47603 , n47604 , n47605 , n47606 , 
     n47607 , n47608 , n47609 , n47610 , n47611 , n47612 , n47613 , n47614 , n47615 , n47616 , 
     n47617 , n47618 , n47619 , n47620 , n47621 , n47622 , n47623 , n47624 , n47625 , n47626 , 
     n47627 , n47628 , n47629 , n47630 , n47631 , n47632 , n47633 , n47634 , n47635 , n47636 , 
     n47637 , n47638 , n47639 , n47640 , n47641 , n47642 , n47643 , n47644 , n47645 , n47646 , 
     n47647 , n47648 , n47649 , n47650 , n47651 , n47652 , n47653 , n47654 , n47655 , n47656 , 
     n47657 , n47658 , n47659 , n47660 , n47661 , n47662 , n47663 , n47664 , n47665 , n47666 , 
     n47667 , n47668 , n47669 , n47670 , n47671 , n47672 , n47673 , n47674 , n47675 , n47676 , 
     n47677 , n47678 , n47679 , n47680 , n47681 , n47682 , n47683 , n47684 , n47685 , n47686 , 
     n47687 , n47688 , n47689 , n47690 , n47691 , n47692 , n47693 , n47694 , n47695 , n47696 , 
     n47697 , n47698 , n47699 , n47700 , n47701 , n47702 , n47703 , n47704 , n47705 , n47706 , 
     n47707 , n47708 , n47709 , n47710 , n47711 , n47712 , n47713 , n47714 , n47715 , n47716 , 
     n47717 , n47718 , n47719 , n47720 , n47721 , n47722 , n47723 , n47724 , n47725 , n47726 , 
     n47727 , n47728 , n47729 , n47730 , n47731 , n47732 , n47733 , n47734 , n47735 , n47736 , 
     n47737 , n47738 , n47739 , n47740 , n47741 , n47742 , n47743 , n47744 , n47745 , n47746 , 
     n47747 , n47748 , n47749 , n47750 , n47751 , n47752 , n47753 , n47754 , n47755 , n47756 , 
     n47757 , n47758 , n47759 , n47760 , n47761 , n47762 , n47763 , n47764 , n47765 , n47766 , 
     n47767 , n47768 , n47769 , n47770 , n47771 , n47772 , n47773 , n47774 , n47775 , n47776 , 
     n47777 , n47778 , n47779 , n47780 , n47781 , n47782 , n47783 , n47784 , n47785 , n47786 , 
     n47787 , n47788 , n47789 , n47790 , n47791 , n47792 , n47793 , n47794 , n47795 , n47796 , 
     n47797 , n47798 , n47799 , n47800 , n47801 , n47802 , n47803 , n47804 , n47805 , n47806 , 
     n47807 , n47808 , n47809 , n47810 , n47811 , n47812 , n47813 , n47814 , n47815 , n47816 , 
     n47817 , n47818 , n47819 , n47820 , n47821 , n47822 , n47823 , n47824 , n47825 , n47826 , 
     n47827 , n47828 , n47829 , n47830 , n47831 , n47832 , n47833 , n47834 , n47835 , n47836 , 
     n47837 , n47838 , n47839 , n47840 , n47841 , n47842 , n47843 , n47844 , n47845 , n47846 , 
     n47847 , n47848 , n47849 , n47850 , n47851 , n47852 , n47853 , n47854 , n47855 , n47856 , 
     n47857 , n47858 , n47859 , n47860 , n47861 , n47862 , n47863 , n47864 , n47865 , n47866 , 
     n47867 , n47868 , n47869 , n47870 , n47871 , n47872 , n47873 , n47874 , n47875 , n47876 , 
     n47877 , n47878 , n47879 , n47880 , n47881 , n47882 , n47883 , n47884 , n47885 , n47886 , 
     n47887 , n47888 , n47889 , n47890 , n47891 , n47892 , n47893 , n47894 , n47895 , n47896 , 
     n47897 , n47898 , n47899 , n47900 , n47901 , n47902 , n47903 , n47904 , n47905 , n47906 , 
     n47907 , n47908 , n47909 , n47910 , n47911 , n47912 , n47913 , n47914 , n47915 , n47916 , 
     n47917 , n47918 , n47919 , n47920 , n47921 , n47922 , n47923 , n47924 , n47925 , n47926 , 
     n47927 , n47928 , n47929 , n47930 , n47931 , n47932 , n47933 , n47934 , n47935 , n47936 , 
     n47937 , n47938 , n47939 , n47940 , n47941 , n47942 , n47943 , n47944 , n47945 , n47946 , 
     n47947 , n47948 , n47949 , n47950 , n47951 , n47952 , n47953 , n47954 , n47955 , n47956 , 
     n47957 , n47958 , n47959 , n47960 , n47961 , n47962 , n47963 , n47964 , n47965 , n47966 , 
     n47967 , n47968 , n47969 , n47970 , n47971 , n47972 , n47973 , n47974 , n47975 , n47976 , 
     n47977 , n47978 , n47979 , n47980 , n47981 , n47982 , n47983 , n47984 , n47985 , n47986 , 
     n47987 , n47988 , n47989 , n47990 , n47991 , n47992 , n47993 , n47994 , n47995 , n47996 , 
     n47997 , n47998 , n47999 , n48000 , n48001 , n48002 , n48003 , n48004 , n48005 , n48006 , 
     n48007 , n48008 , n48009 , n48010 , n48011 , n48012 , n48013 , n48014 , n48015 , n48016 , 
     n48017 , n48018 , n48019 , n48020 , n48021 , n48022 , n48023 , n48024 , n48025 , n48026 , 
     n48027 , n48028 , n48029 , n48030 , n48031 , n48032 , n48033 , n48034 , n48035 , n48036 , 
     n48037 , n48038 , n48039 , n48040 , n48041 , n48042 , n48043 , n48044 , n48045 , n48046 , 
     n48047 , n48048 , n48049 , n48050 , n48051 , n48052 , n48053 , n48054 , n48055 , n48056 , 
     n48057 , n48058 , n48059 , n48060 , n48061 , n48062 , n48063 , n48064 , n48065 , n48066 , 
     n48067 , n48068 , n48069 , n48070 , n48071 , n48072 , n48073 , n48074 , n48075 , n48076 , 
     n48077 , n48078 , n48079 , n48080 , n48081 , n48082 , n48083 , n48084 , n48085 , n48086 , 
     n48087 , n48088 , n48089 , n48090 , n48091 , n48092 , n48093 , n48094 , n48095 , n48096 , 
     n48097 , n48098 , n48099 , n48100 , n48101 , n48102 , n48103 , n48104 , n48105 , n48106 , 
     n48107 , n48108 , n48109 , n48110 , n48111 , n48112 , n48113 , n48114 , n48115 , n48116 , 
     n48117 , n48118 , n48119 , n48120 , n48121 , n48122 , n48123 , n48124 , n48125 , n48126 , 
     n48127 , n48128 , n48129 , n48130 , n48131 , n48132 , n48133 , n48134 , n48135 , n48136 , 
     n48137 , n48138 , n48139 , n48140 , n48141 , n48142 , n48143 , n48144 , n48145 , n48146 , 
     n48147 , n48148 , n48149 , n48150 , n48151 , n48152 , n48153 , n48154 , n48155 , n48156 , 
     n48157 , n48158 , n48159 , n48160 , n48161 , n48162 , n48163 , n48164 , n48165 , n48166 , 
     n48167 , n48168 , n48169 , n48170 , n48171 , n48172 , n48173 , n48174 , n48175 , n48176 , 
     n48177 , n48178 , n48179 , n48180 , n48181 , n48182 , n48183 , n48184 , n48185 , n48186 , 
     n48187 , n48188 , n48189 , n48190 , n48191 , n48192 , n48193 , n48194 , n48195 , n48196 , 
     n48197 , n48198 , n48199 , n48200 , n48201 , n48202 , n48203 , n48204 , n48205 , n48206 , 
     n48207 , n48208 , n48209 , n48210 , n48211 , n48212 , n48213 , n48214 , n48215 , n48216 , 
     n48217 , n48218 , n48219 , n48220 , n48221 , n48222 , n48223 , n48224 , n48225 , n48226 , 
     n48227 , n48228 , n48229 , n48230 , n48231 , n48232 , n48233 , n48234 , n48235 , n48236 , 
     n48237 , n48238 , n48239 , n48240 , n48241 , n48242 , n48243 , n48244 , n48245 , n48246 , 
     n48247 , n48248 , n48249 , n48250 , n48251 , n48252 , n48253 , n48254 , n48255 , n48256 , 
     n48257 , n48258 , n48259 , n48260 , n48261 , n48262 , n48263 , n48264 , n48265 , n48266 , 
     n48267 , n48268 , n48269 , n48270 , n48271 , n48272 , n48273 , n48274 , n48275 , n48276 , 
     n48277 , n48278 , n48279 , n48280 , n48281 , n48282 , n48283 , n48284 , n48285 , n48286 , 
     n48287 , n48288 , n48289 , n48290 , n48291 , n48292 , n48293 , n48294 , n48295 , n48296 , 
     n48297 , n48298 , n48299 , n48300 , n48301 , n48302 , n48303 , n48304 , n48305 , n48306 , 
     n48307 , n48308 , n48309 , n48310 , n48311 , n48312 , n48313 , n48314 , n48315 , n48316 , 
     n48317 , n48318 , n48319 , n48320 , n48321 , n48322 , n48323 , n48324 , n48325 , n48326 , 
     n48327 , n48328 , n48329 , n48330 , n48331 , n48332 , n48333 , n48334 , n48335 , n48336 , 
     n48337 , n48338 , n48339 , n48340 , n48341 , n48342 , n48343 , n48344 , n48345 , n48346 , 
     n48347 , n48348 , n48349 , n48350 , n48351 , n48352 , n48353 , n48354 , n48355 , n48356 , 
     n48357 , n48358 , n48359 , n48360 , n48361 , n48362 , n48363 , n48364 , n48365 , n48366 , 
     n48367 , n48368 , n48369 , n48370 , n48371 , n48372 , n48373 , n48374 , n48375 , n48376 , 
     n48377 , n48378 , n48379 , n48380 , n48381 , n48382 , n48383 , n48384 , n48385 , n48386 , 
     n48387 , n48388 , n48389 , n48390 , n48391 , n48392 , n48393 , n48394 , n48395 , n48396 , 
     n48397 , n48398 , n48399 , n48400 , n48401 , n48402 , n48403 , n48404 , n48405 , n48406 , 
     n48407 , n48408 , n48409 , n48410 , n48411 , n48412 , n48413 , n48414 , n48415 , n48416 , 
     n48417 , n48418 , n48419 , n48420 , n48421 , n48422 , n48423 , n48424 , n48425 , n48426 , 
     n48427 , n48428 , n48429 , n48430 , n48431 , n48432 , n48433 , n48434 , n48435 , n48436 , 
     n48437 , n48438 , n48439 , n48440 , n48441 , n48442 , n48443 , n48444 , n48445 , n48446 , 
     n48447 , n48448 , n48449 , n48450 , n48451 , n48452 , n48453 , n48454 , n48455 , n48456 , 
     n48457 , n48458 , n48459 , n48460 , n48461 , n48462 , n48463 , n48464 , n48465 , n48466 , 
     n48467 , n48468 , n48469 , n48470 , n48471 , n48472 , n48473 , n48474 , n48475 , n48476 , 
     n48477 , n48478 , n48479 , n48480 , n48481 , n48482 , n48483 , n48484 , n48485 , n48486 , 
     n48487 , n48488 , n48489 , n48490 , n48491 , n48492 , n48493 , n48494 , n48495 , n48496 , 
     n48497 , n48498 , n48499 , n48500 , n48501 , n48502 , n48503 , n48504 , n48505 , n48506 , 
     n48507 , n48508 , n48509 , n48510 , n48511 , n48512 , n48513 , n48514 , n48515 , n48516 , 
     n48517 , n48518 , n48519 , n48520 , n48521 , n48522 , n48523 , n48524 , n48525 , n48526 , 
     n48527 , n48528 , n48529 , n48530 , n48531 , n48532 , n48533 , n48534 , n48535 , n48536 , 
     n48537 , n48538 , n48539 , n48540 , n48541 , n48542 , n48543 , n48544 , n48545 , n48546 , 
     n48547 , n48548 , n48549 , n48550 , n48551 , n48552 , n48553 , n48554 , n48555 , n48556 , 
     n48557 , n48558 , n48559 , n48560 , n48561 , n48562 , n48563 , n48564 , n48565 , n48566 , 
     n48567 , n48568 , n48569 , n48570 , n48571 , n48572 , n48573 , n48574 , n48575 , n48576 , 
     n48577 , n48578 , n48579 , n48580 , n48581 , n48582 , n48583 , n48584 , n48585 , n48586 , 
     n48587 , n48588 , n48589 , n48590 , n48591 , n48592 , n48593 , n48594 , n48595 , n48596 , 
     n48597 , n48598 , n48599 , n48600 , n48601 , n48602 , n48603 , n48604 , n48605 , n48606 , 
     n48607 , n48608 , n48609 , n48610 , n48611 , n48612 , n48613 , n48614 , n48615 , n48616 , 
     n48617 , n48618 , n48619 , n48620 , n48621 , n48622 , n48623 , n48624 , n48625 , n48626 , 
     n48627 , n48628 , n48629 , n48630 , n48631 , n48632 , n48633 , n48634 , n48635 , n48636 , 
     n48637 , n48638 , n48639 , n48640 , n48641 , n48642 , n48643 , n48644 , n48645 , n48646 , 
     n48647 , n48648 , n48649 , n48650 , n48651 , n48652 , n48653 , n48654 , n48655 , n48656 , 
     n48657 , n48658 , n48659 , n48660 , n48661 , n48662 , n48663 , n48664 , n48665 , n48666 , 
     n48667 , n48668 , n48669 , n48670 , n48671 , n48672 , n48673 , n48674 , n48675 , n48676 , 
     n48677 , n48678 , n48679 , n48680 , n48681 , n48682 , n48683 , n48684 , n48685 , n48686 , 
     n48687 , n48688 , n48689 , n48690 , n48691 , n48692 , n48693 , n48694 , n48695 , n48696 , 
     n48697 , n48698 , n48699 , n48700 , n48701 , n48702 , n48703 , n48704 , n48705 , n48706 , 
     n48707 , n48708 , n48709 , n48710 , n48711 , n48712 , n48713 , n48714 , n48715 , n48716 , 
     n48717 , n48718 , n48719 , n48720 , n48721 , n48722 , n48723 , n48724 , n48725 , n48726 , 
     n48727 , n48728 , n48729 , n48730 , n48731 , n48732 , n48733 , n48734 , n48735 , n48736 , 
     n48737 , n48738 , n48739 , n48740 , n48741 , n48742 , n48743 , n48744 , n48745 , n48746 , 
     n48747 , n48748 , n48749 , n48750 , n48751 , n48752 , n48753 , n48754 , n48755 , n48756 , 
     n48757 , n48758 , n48759 , n48760 , n48761 , n48762 , n48763 , n48764 , n48765 , n48766 , 
     n48767 , n48768 , n48769 , n48770 , n48771 , n48772 , n48773 , n48774 , n48775 , n48776 , 
     n48777 , n48778 , n48779 , n48780 , n48781 , n48782 , n48783 , n48784 , n48785 , n48786 , 
     n48787 , n48788 , n48789 , n48790 , n48791 , n48792 , n48793 , n48794 , n48795 , n48796 , 
     n48797 , n48798 , n48799 , n48800 , n48801 , n48802 , n48803 , n48804 , n48805 , n48806 , 
     n48807 , n48808 , n48809 , n48810 , n48811 , n48812 , n48813 , n48814 , n48815 , n48816 , 
     n48817 , n48818 , n48819 , n48820 , n48821 , n48822 , n48823 , n48824 , n48825 , n48826 , 
     n48827 , n48828 , n48829 , n48830 , n48831 , n48832 , n48833 , n48834 , n48835 , n48836 , 
     n48837 , n48838 , n48839 , n48840 , n48841 , n48842 , n48843 , n48844 , n48845 , n48846 , 
     n48847 , n48848 , n48849 , n48850 , n48851 , n48852 , n48853 , n48854 , n48855 , n48856 , 
     n48857 , n48858 , n48859 , n48860 , n48861 , n48862 , n48863 , n48864 , n48865 , n48866 , 
     n48867 , n48868 , n48869 , n48870 , n48871 , n48872 , n48873 , n48874 , n48875 , n48876 , 
     n48877 , n48878 , n48879 , n48880 , n48881 , n48882 , n48883 , n48884 , n48885 , n48886 , 
     n48887 , n48888 , n48889 , n48890 , n48891 , n48892 , n48893 , n48894 , n48895 , n48896 , 
     n48897 , n48898 , n48899 , n48900 , n48901 , n48902 , n48903 , n48904 , n48905 , n48906 , 
     n48907 , n48908 , n48909 , n48910 , n48911 , n48912 , n48913 , n48914 , n48915 , n48916 , 
     n48917 , n48918 , n48919 , n48920 , n48921 , n48922 , n48923 , n48924 , n48925 , n48926 , 
     n48927 , n48928 , n48929 , n48930 , n48931 , n48932 , n48933 , n48934 , n48935 , n48936 , 
     n48937 , n48938 , n48939 , n48940 , n48941 , n48942 , n48943 , n48944 , n48945 , n48946 , 
     n48947 , n48948 , n48949 , n48950 , n48951 , n48952 , n48953 , n48954 , n48955 , n48956 , 
     n48957 , n48958 , n48959 , n48960 , n48961 , n48962 , n48963 , n48964 , n48965 , n48966 , 
     n48967 , n48968 , n48969 , n48970 , n48971 , n48972 , n48973 , n48974 , n48975 , n48976 , 
     n48977 , n48978 , n48979 , n48980 , n48981 , n48982 , n48983 , n48984 , n48985 , n48986 , 
     n48987 , n48988 , n48989 , n48990 , n48991 , n48992 , n48993 , n48994 , n48995 , n48996 , 
     n48997 , n48998 , n48999 , n49000 , n49001 , n49002 , n49003 , n49004 , n49005 , n49006 , 
     n49007 , n49008 , n49009 , n49010 , n49011 , n49012 , n49013 , n49014 , n49015 , n49016 , 
     n49017 , n49018 , n49019 , n49020 , n49021 , n49022 , n49023 , n49024 , n49025 , n49026 , 
     n49027 , n49028 , n49029 , n49030 , n49031 , n49032 , n49033 , n49034 , n49035 , n49036 , 
     n49037 , n49038 , n49039 , n49040 , n49041 , n49042 , n49043 , n49044 , n49045 , n49046 , 
     n49047 , n49048 , n49049 , n49050 , n49051 , n49052 , n49053 , n49054 , n49055 , n49056 , 
     n49057 , n49058 , n49059 , n49060 , n49061 , n49062 , n49063 , n49064 , n49065 , n49066 , 
     n49067 , n49068 , n49069 , n49070 , n49071 , n49072 , n49073 , n49074 , n49075 , n49076 , 
     n49077 , n49078 , n49079 , n49080 , n49081 , n49082 , n49083 , n49084 , n49085 , n49086 , 
     n49087 , n49088 , n49089 , n49090 , n49091 , n49092 , n49093 , n49094 , n49095 , n49096 , 
     n49097 , n49098 , n49099 , n49100 , n49101 , n49102 , n49103 , n49104 , n49105 , n49106 , 
     n49107 , n49108 , n49109 , n49110 , n49111 , n49112 , n49113 , n49114 , n49115 , n49116 , 
     n49117 , n49118 , n49119 , n49120 , n49121 , n49122 , n49123 , n49124 , n49125 , n49126 , 
     n49127 , n49128 , n49129 , n49130 , n49131 , n49132 , n49133 , n49134 , n49135 , n49136 , 
     n49137 , n49138 , n49139 , n49140 , n49141 , n49142 , n49143 , n49144 , n49145 , n49146 , 
     n49147 , n49148 , n49149 , n49150 , n49151 , n49152 , n49153 , n49154 , n49155 , n49156 , 
     n49157 , n49158 , n49159 , n49160 , n49161 , n49162 , n49163 , n49164 , n49165 , n49166 , 
     n49167 , n49168 , n49169 , n49170 , n49171 , n49172 , n49173 , n49174 , n49175 , n49176 , 
     n49177 , n49178 , n49179 , n49180 , n49181 , n49182 , n49183 , n49184 , n49185 , n49186 , 
     n49187 , n49188 , n49189 , n49190 , n49191 , n49192 , n49193 , n49194 , n49195 , n49196 , 
     n49197 , n49198 , n49199 , n49200 , n49201 , n49202 , n49203 , n49204 , n49205 , n49206 , 
     n49207 , n49208 , n49209 , n49210 , n49211 , n49212 , n49213 , n49214 , n49215 , n49216 , 
     n49217 , n49218 , n49219 , n49220 , n49221 , n49222 , n49223 , n49224 , n49225 , n49226 , 
     n49227 , n49228 , n49229 , n49230 , n49231 , n49232 , n49233 , n49234 , n49235 , n49236 , 
     n49237 , n49238 , n49239 , n49240 , n49241 , n49242 , n49243 , n49244 , n49245 , n49246 , 
     n49247 , n49248 , n49249 , n49250 , n49251 , n49252 , n49253 , n49254 , n49255 , n49256 , 
     n49257 , n49258 , n49259 , n49260 , n49261 , n49262 , n49263 , n49264 , n49265 , n49266 , 
     n49267 , n49268 , n49269 , n49270 , n49271 , n49272 , n49273 , n49274 , n49275 , n49276 , 
     n49277 , n49278 , n49279 , n49280 , n49281 , n49282 , n49283 , n49284 , n49285 , n49286 , 
     n49287 , n49288 , n49289 , n49290 , n49291 , n49292 , n49293 , n49294 , n49295 , n49296 , 
     n49297 , n49298 , n49299 , n49300 , n49301 , n49302 , n49303 , n49304 , n49305 , n49306 , 
     n49307 , n49308 , n49309 , n49310 , n49311 , n49312 , n49313 , n49314 , n49315 , n49316 , 
     n49317 , n49318 , n49319 , n49320 , n49321 , n49322 , n49323 , n49324 , n49325 , n49326 , 
     n49327 , n49328 , n49329 , n49330 , n49331 , n49332 , n49333 , n49334 , n49335 , n49336 , 
     n49337 , n49338 , n49339 , n49340 , n49341 , n49342 , n49343 , n49344 , n49345 , n49346 , 
     n49347 , n49348 , n49349 , n49350 , n49351 , n49352 , n49353 , n49354 , n49355 , n49356 , 
     n49357 , n49358 , n49359 , n49360 , n49361 , n49362 , n49363 , n49364 , n49365 , n49366 , 
     n49367 , n49368 , n49369 , n49370 , n49371 , n49372 , n49373 , n49374 , n49375 , n49376 , 
     n49377 , n49378 , n49379 , n49380 , n49381 , n49382 , n49383 , n49384 , n49385 , n49386 , 
     n49387 , n49388 , n49389 , n49390 , n49391 , n49392 , n49393 , n49394 , n49395 , n49396 , 
     n49397 , n49398 , n49399 , n49400 , n49401 , n49402 , n49403 , n49404 , n49405 , n49406 , 
     n49407 , n49408 , n49409 , n49410 , n49411 , n49412 , n49413 , n49414 , n49415 , n49416 , 
     n49417 , n49418 , n49419 , n49420 , n49421 , n49422 , n49423 , n49424 , n49425 , n49426 , 
     n49427 , n49428 , n49429 , n49430 , n49431 , n49432 , n49433 , n49434 , n49435 , n49436 , 
     n49437 , n49438 , n49439 , n49440 , n49441 , n49442 , n49443 , n49444 , n49445 , n49446 , 
     n49447 , n49448 , n49449 , n49450 , n49451 , n49452 , n49453 , n49454 , n49455 , n49456 , 
     n49457 , n49458 , n49459 , n49460 , n49461 , n49462 , n49463 , n49464 , n49465 , n49466 , 
     n49467 , n49468 , n49469 , n49470 , n49471 , n49472 , n49473 , n49474 , n49475 , n49476 , 
     n49477 , n49478 , n49479 , n49480 , n49481 , n49482 , n49483 , n49484 , n49485 , n49486 , 
     n49487 , n49488 , n49489 , n49490 , n49491 , n49492 , n49493 , n49494 , n49495 , n49496 , 
     n49497 , n49498 , n49499 , n49500 , n49501 , n49502 , n49503 , n49504 , n49505 , n49506 , 
     n49507 , n49508 , n49509 , n49510 , n49511 , n49512 , n49513 , n49514 , n49515 , n49516 , 
     n49517 , n49518 , n49519 , n49520 , n49521 , n49522 , n49523 , n49524 , n49525 , n49526 , 
     n49527 , n49528 , n49529 , n49530 , n49531 , n49532 , n49533 , n49534 , n49535 , n49536 , 
     n49537 , n49538 , n49539 , n49540 , n49541 , n49542 , n49543 , n49544 , n49545 , n49546 , 
     n49547 , n49548 , n49549 , n49550 , n49551 , n49552 , n49553 , n49554 , n49555 , n49556 , 
     n49557 , n49558 , n49559 , n49560 , n49561 , n49562 , n49563 , n49564 , n49565 , n49566 , 
     n49567 , n49568 , n49569 , n49570 , n49571 , n49572 , n49573 , n49574 , n49575 , n49576 , 
     n49577 , n49578 , n49579 , n49580 , n49581 , n49582 , n49583 , n49584 , n49585 , n49586 , 
     n49587 , n49588 , n49589 , n49590 , n49591 , n49592 , n49593 , n49594 , n49595 , n49596 , 
     n49597 , n49598 , n49599 , n49600 , n49601 , n49602 , n49603 , n49604 , n49605 , n49606 , 
     n49607 , n49608 , n49609 , n49610 , n49611 , n49612 , n49613 , n49614 , n49615 , n49616 , 
     n49617 , n49618 , n49619 , n49620 , n49621 , n49622 , n49623 , n49624 , n49625 , n49626 , 
     n49627 , n49628 , n49629 , n49630 , n49631 , n49632 , n49633 , n49634 , n49635 , n49636 , 
     n49637 , n49638 , n49639 , n49640 , n49641 , n49642 , n49643 , n49644 , n49645 , n49646 , 
     n49647 , n49648 , n49649 , n49650 , n49651 , n49652 , n49653 , n49654 , n49655 , n49656 , 
     n49657 , n49658 , n49659 , n49660 , n49661 , n49662 , n49663 , n49664 , n49665 , n49666 , 
     n49667 , n49668 , n49669 , n49670 , n49671 , n49672 , n49673 , n49674 , n49675 , n49676 , 
     n49677 , n49678 , n49679 , n49680 , n49681 , n49682 , n49683 , n49684 , n49685 , n49686 , 
     n49687 , n49688 , n49689 , n49690 , n49691 , n49692 , n49693 , n49694 , n49695 , n49696 , 
     n49697 , n49698 , n49699 , n49700 , n49701 , n49702 , n49703 , n49704 , n49705 , n49706 , 
     n49707 , n49708 , n49709 , n49710 , n49711 , n49712 , n49713 , n49714 , n49715 , n49716 , 
     n49717 , n49718 , n49719 , n49720 , n49721 , n49722 , n49723 , n49724 , n49725 , n49726 , 
     n49727 , n49728 , n49729 , n49730 , n49731 , n49732 , n49733 , n49734 , n49735 , n49736 , 
     n49737 , n49738 , n49739 , n49740 , n49741 , n49742 , n49743 , n49744 , n49745 , n49746 , 
     n49747 , n49748 , n49749 , n49750 , n49751 , n49752 , n49753 , n49754 , n49755 , n49756 , 
     n49757 , n49758 , n49759 , n49760 , n49761 , n49762 , n49763 , n49764 , n49765 , n49766 , 
     n49767 , n49768 , n49769 , n49770 , n49771 , n49772 , n49773 , n49774 , n49775 , n49776 , 
     n49777 , n49778 , n49779 , n49780 , n49781 , n49782 , n49783 , n49784 , n49785 , n49786 , 
     n49787 , n49788 , n49789 , n49790 , n49791 , n49792 , n49793 , n49794 , n49795 , n49796 , 
     n49797 , n49798 , n49799 , n49800 , n49801 , n49802 , n49803 , n49804 , n49805 , n49806 , 
     n49807 , n49808 , n49809 , n49810 , n49811 , n49812 , n49813 , n49814 , n49815 , n49816 , 
     n49817 , n49818 , n49819 , n49820 , n49821 , n49822 , n49823 , n49824 , n49825 , n49826 , 
     n49827 , n49828 , n49829 , n49830 , n49831 , n49832 , n49833 , n49834 , n49835 , n49836 , 
     n49837 , n49838 , n49839 , n49840 , n49841 , n49842 , n49843 , n49844 , n49845 , n49846 , 
     n49847 , n49848 , n49849 , n49850 , n49851 , n49852 , n49853 , n49854 , n49855 , n49856 , 
     n49857 , n49858 , n49859 , n49860 , n49861 , n49862 , n49863 , n49864 , n49865 , n49866 , 
     n49867 , n49868 , n49869 , n49870 , n49871 , n49872 , n49873 , n49874 , n49875 , n49876 , 
     n49877 , n49878 , n49879 , n49880 , n49881 , n49882 , n49883 , n49884 , n49885 , n49886 , 
     n49887 , n49888 , n49889 , n49890 , n49891 , n49892 , n49893 , n49894 , n49895 , n49896 , 
     n49897 , n49898 , n49899 , n49900 , n49901 , n49902 , n49903 , n49904 , n49905 , n49906 , 
     n49907 , n49908 , n49909 , n49910 , n49911 , n49912 , n49913 , n49914 , n49915 , n49916 , 
     n49917 , n49918 , n49919 , n49920 , n49921 , n49922 , n49923 , n49924 , n49925 , n49926 , 
     n49927 , n49928 , n49929 , n49930 , n49931 , n49932 , n49933 , n49934 , n49935 , n49936 , 
     n49937 , n49938 , n49939 , n49940 , n49941 , n49942 , n49943 , n49944 , n49945 , n49946 , 
     n49947 , n49948 , n49949 , n49950 , n49951 , n49952 , n49953 , n49954 , n49955 , n49956 , 
     n49957 , n49958 , n49959 , n49960 , n49961 , n49962 , n49963 , n49964 , n49965 , n49966 , 
     n49967 , n49968 , n49969 , n49970 , n49971 , n49972 , n49973 , n49974 , n49975 , n49976 , 
     n49977 , n49978 , n49979 , n49980 , n49981 , n49982 , n49983 , n49984 , n49985 , n49986 , 
     n49987 , n49988 , n49989 , n49990 , n49991 , n49992 , n49993 , n49994 , n49995 , n49996 , 
     n49997 , n49998 , n49999 , n50000 , n50001 , n50002 , n50003 , n50004 , n50005 , n50006 , 
     n50007 , n50008 , n50009 , n50010 , n50011 , n50012 , n50013 , n50014 , n50015 , n50016 , 
     n50017 , n50018 , n50019 , n50020 , n50021 , n50022 , n50023 , n50024 , n50025 , n50026 , 
     n50027 , n50028 , n50029 , n50030 , n50031 , n50032 , n50033 , n50034 , n50035 , n50036 , 
     n50037 , n50038 , n50039 , n50040 , n50041 , n50042 , n50043 , n50044 , n50045 , n50046 , 
     n50047 , n50048 , n50049 , n50050 , n50051 , n50052 , n50053 , n50054 , n50055 , n50056 , 
     n50057 , n50058 , n50059 , n50060 , n50061 , n50062 , n50063 , n50064 , n50065 , n50066 , 
     n50067 , n50068 , n50069 , n50070 , n50071 , n50072 , n50073 , n50074 , n50075 , n50076 , 
     n50077 , n50078 , n50079 , n50080 , n50081 , n50082 , n50083 , n50084 , n50085 , n50086 , 
     n50087 , n50088 , n50089 , n50090 , n50091 , n50092 , n50093 , n50094 , n50095 , n50096 , 
     n50097 , n50098 , n50099 , n50100 , n50101 , n50102 , n50103 , n50104 , n50105 , n50106 , 
     n50107 , n50108 , n50109 , n50110 , n50111 , n50112 , n50113 , n50114 , n50115 , n50116 , 
     n50117 , n50118 , n50119 , n50120 , n50121 , n50122 , n50123 , n50124 , n50125 , n50126 , 
     n50127 , n50128 , n50129 , n50130 , n50131 , n50132 , n50133 , n50134 , n50135 , n50136 , 
     n50137 , n50138 , n50139 , n50140 , n50141 , n50142 , n50143 , n50144 , n50145 , n50146 , 
     n50147 , n50148 , n50149 , n50150 , n50151 , n50152 , n50153 , n50154 , n50155 , n50156 , 
     n50157 , n50158 , n50159 , n50160 , n50161 , n50162 , n50163 , n50164 , n50165 , n50166 , 
     n50167 , n50168 , n50169 , n50170 , n50171 , n50172 , n50173 , n50174 , n50175 , n50176 , 
     n50177 , n50178 , n50179 , n50180 , n50181 , n50182 , n50183 , n50184 , n50185 , n50186 , 
     n50187 , n50188 , n50189 , n50190 , n50191 , n50192 , n50193 , n50194 , n50195 , n50196 , 
     n50197 , n50198 , n50199 , n50200 , n50201 , n50202 , n50203 , n50204 , n50205 , n50206 , 
     n50207 , n50208 , n50209 , n50210 , n50211 , n50212 , n50213 , n50214 , n50215 , n50216 , 
     n50217 , n50218 , n50219 , n50220 , n50221 , n50222 , n50223 , n50224 , n50225 , n50226 , 
     n50227 , n50228 , n50229 , n50230 , n50231 , n50232 , n50233 , n50234 , n50235 , n50236 , 
     n50237 , n50238 , n50239 , n50240 , n50241 , n50242 , n50243 , n50244 , n50245 , n50246 , 
     n50247 , n50248 , n50249 , n50250 , n50251 , n50252 , n50253 , n50254 , n50255 , n50256 , 
     n50257 , n50258 , n50259 , n50260 , n50261 , n50262 , n50263 , n50264 , n50265 , n50266 , 
     n50267 , n50268 , n50269 , n50270 , n50271 , n50272 , n50273 , n50274 , n50275 , n50276 , 
     n50277 , n50278 , n50279 , n50280 , n50281 , n50282 , n50283 , n50284 , n50285 , n50286 , 
     n50287 , n50288 , n50289 , n50290 , n50291 , n50292 , n50293 , n50294 , n50295 , n50296 , 
     n50297 , n50298 , n50299 , n50300 , n50301 , n50302 , n50303 , n50304 , n50305 , n50306 , 
     n50307 , n50308 , n50309 , n50310 , n50311 , n50312 , n50313 , n50314 , n50315 , n50316 , 
     n50317 , n50318 , n50319 , n50320 , n50321 , n50322 , n50323 , n50324 , n50325 , n50326 , 
     n50327 , n50328 , n50329 , n50330 , n50331 , n50332 , n50333 , n50334 , n50335 , n50336 , 
     n50337 , n50338 , n50339 , n50340 , n50341 , n50342 , n50343 , n50344 , n50345 , n50346 , 
     n50347 , n50348 , n50349 , n50350 , n50351 , n50352 , n50353 , n50354 , n50355 , n50356 , 
     n50357 , n50358 , n50359 , n50360 , n50361 , n50362 , n50363 , n50364 , n50365 , n50366 , 
     n50367 , n50368 , n50369 , n50370 , n50371 , n50372 , n50373 , n50374 , n50375 , n50376 , 
     n50377 , n50378 , n50379 , n50380 , n50381 , n50382 , n50383 , n50384 , n50385 , n50386 , 
     n50387 , n50388 , n50389 , n50390 , n50391 , n50392 , n50393 , n50394 , n50395 , n50396 , 
     n50397 , n50398 , n50399 , n50400 , n50401 , n50402 , n50403 , n50404 , n50405 , n50406 , 
     n50407 , n50408 , n50409 , n50410 , n50411 , n50412 , n50413 , n50414 , n50415 , n50416 , 
     n50417 , n50418 , n50419 , n50420 , n50421 , n50422 , n50423 , n50424 , n50425 , n50426 , 
     n50427 , n50428 , n50429 , n50430 , n50431 , n50432 , n50433 , n50434 , n50435 , n50436 , 
     n50437 , n50438 , n50439 , n50440 , n50441 , n50442 , n50443 , n50444 , n50445 , n50446 , 
     n50447 , n50448 , n50449 , n50450 , n50451 , n50452 , n50453 , n50454 , n50455 , n50456 , 
     n50457 , n50458 , n50459 , n50460 , n50461 , n50462 , n50463 , n50464 , n50465 , n50466 , 
     n50467 , n50468 , n50469 , n50470 , n50471 , n50472 , n50473 , n50474 , n50475 , n50476 , 
     n50477 , n50478 , n50479 , n50480 , n50481 , n50482 , n50483 , n50484 , n50485 , n50486 , 
     n50487 , n50488 , n50489 , n50490 , n50491 , n50492 , n50493 , n50494 , n50495 , n50496 , 
     n50497 , n50498 , n50499 , n50500 , n50501 , n50502 , n50503 , n50504 , n50505 , n50506 , 
     n50507 , n50508 , n50509 , n50510 , n50511 , n50512 , n50513 , n50514 , n50515 , n50516 , 
     n50517 , n50518 , n50519 , n50520 , n50521 , n50522 , n50523 , n50524 , n50525 , n50526 , 
     n50527 , n50528 , n50529 , n50530 , n50531 , n50532 , n50533 , n50534 , n50535 , n50536 , 
     n50537 , n50538 , n50539 , n50540 , n50541 , n50542 , n50543 , n50544 , n50545 , n50546 , 
     n50547 , n50548 , n50549 , n50550 , n50551 , n50552 , n50553 , n50554 , n50555 , n50556 , 
     n50557 , n50558 , n50559 , n50560 , n50561 , n50562 , n50563 , n50564 , n50565 , n50566 , 
     n50567 , n50568 , n50569 , n50570 , n50571 , n50572 , n50573 , n50574 , n50575 , n50576 , 
     n50577 , n50578 , n50579 , n50580 , n50581 , n50582 , n50583 , n50584 , n50585 , n50586 , 
     n50587 , n50588 , n50589 , n50590 , n50591 , n50592 , n50593 , n50594 , n50595 , n50596 , 
     n50597 , n50598 , n50599 , n50600 , n50601 , n50602 , n50603 , n50604 , n50605 , n50606 , 
     n50607 , n50608 , n50609 , n50610 , n50611 , n50612 , n50613 , n50614 , n50615 , n50616 , 
     n50617 , n50618 , n50619 , n50620 , n50621 , n50622 , n50623 , n50624 , n50625 , n50626 , 
     n50627 , n50628 , n50629 , n50630 , n50631 , n50632 , n50633 , n50634 , n50635 , n50636 , 
     n50637 , n50638 , n50639 , n50640 , n50641 , n50642 , n50643 , n50644 , n50645 , n50646 , 
     n50647 , n50648 , n50649 , n50650 , n50651 , n50652 , n50653 , n50654 , n50655 , n50656 , 
     n50657 , n50658 , n50659 , n50660 , n50661 , n50662 , n50663 , n50664 , n50665 , n50666 , 
     n50667 , n50668 , n50669 , n50670 , n50671 , n50672 , n50673 , n50674 , n50675 , n50676 , 
     n50677 , n50678 , n50679 , n50680 , n50681 , n50682 , n50683 , n50684 , n50685 , n50686 , 
     n50687 , n50688 , n50689 , n50690 , n50691 , n50692 , n50693 , n50694 , n50695 , n50696 , 
     n50697 , n50698 , n50699 , n50700 , n50701 , n50702 , n50703 , n50704 , n50705 , n50706 , 
     n50707 , n50708 , n50709 , n50710 , n50711 , n50712 , n50713 , n50714 , n50715 , n50716 , 
     n50717 , n50718 , n50719 , n50720 , n50721 , n50722 , n50723 , n50724 , n50725 , n50726 , 
     n50727 , n50728 , n50729 , n50730 , n50731 , n50732 , n50733 , n50734 , n50735 , n50736 , 
     n50737 , n50738 , n50739 , n50740 , n50741 , n50742 , n50743 , n50744 , n50745 , n50746 , 
     n50747 , n50748 , n50749 , n50750 , n50751 , n50752 , n50753 , n50754 , n50755 , n50756 , 
     n50757 , n50758 , n50759 , n50760 , n50761 , n50762 , n50763 , n50764 , n50765 , n50766 , 
     n50767 , n50768 , n50769 , n50770 , n50771 , n50772 , n50773 , n50774 , n50775 , n50776 , 
     n50777 , n50778 , n50779 , n50780 , n50781 , n50782 , n50783 , n50784 , n50785 , n50786 , 
     n50787 , n50788 , n50789 , n50790 , n50791 , n50792 , n50793 , n50794 , n50795 , n50796 , 
     n50797 , n50798 , n50799 , n50800 , n50801 , n50802 , n50803 , n50804 , n50805 , n50806 , 
     n50807 , n50808 , n50809 , n50810 , n50811 , n50812 , n50813 , n50814 , n50815 , n50816 , 
     n50817 , n50818 , n50819 , n50820 , n50821 , n50822 , n50823 , n50824 , n50825 , n50826 , 
     n50827 , n50828 , n50829 , n50830 , n50831 , n50832 , n50833 , n50834 , n50835 , n50836 , 
     n50837 , n50838 , n50839 , n50840 , n50841 , n50842 , n50843 , n50844 , n50845 , n50846 , 
     n50847 , n50848 , n50849 , n50850 , n50851 , n50852 , n50853 , n50854 , n50855 , n50856 , 
     n50857 , n50858 , n50859 , n50860 , n50861 , n50862 , n50863 , n50864 , n50865 , n50866 , 
     n50867 , n50868 , n50869 , n50870 , n50871 , n50872 , n50873 , n50874 , n50875 , n50876 , 
     n50877 , n50878 , n50879 , n50880 , n50881 , n50882 , n50883 , n50884 , n50885 , n50886 , 
     n50887 , n50888 , n50889 , n50890 , n50891 , n50892 , n50893 , n50894 , n50895 , n50896 , 
     n50897 , n50898 , n50899 , n50900 , n50901 , n50902 , n50903 , n50904 , n50905 , n50906 , 
     n50907 , n50908 , n50909 , n50910 , n50911 , n50912 , n50913 , n50914 , n50915 , n50916 , 
     n50917 , n50918 , n50919 , n50920 , n50921 , n50922 , n50923 , n50924 , n50925 , n50926 , 
     n50927 , n50928 , n50929 , n50930 , n50931 , n50932 , n50933 , n50934 , n50935 , n50936 , 
     n50937 , n50938 , n50939 , n50940 , n50941 , n50942 , n50943 , n50944 , n50945 , n50946 , 
     n50947 , n50948 , n50949 , n50950 , n50951 , n50952 , n50953 , n50954 , n50955 , n50956 , 
     n50957 , n50958 , n50959 , n50960 , n50961 , n50962 , n50963 , n50964 , n50965 , n50966 , 
     n50967 , n50968 , n50969 , n50970 , n50971 , n50972 , n50973 , n50974 , n50975 , n50976 , 
     n50977 , n50978 , n50979 , n50980 , n50981 , n50982 , n50983 , n50984 , n50985 , n50986 , 
     n50987 , n50988 , n50989 , n50990 , n50991 , n50992 , n50993 , n50994 , n50995 , n50996 , 
     n50997 , n50998 , n50999 , n51000 , n51001 , n51002 , n51003 , n51004 , n51005 , n51006 , 
     n51007 , n51008 , n51009 , n51010 , n51011 , n51012 , n51013 , n51014 , n51015 , n51016 , 
     n51017 , n51018 , n51019 , n51020 , n51021 , n51022 , n51023 , n51024 , n51025 , n51026 , 
     n51027 , n51028 , n51029 , n51030 , n51031 , n51032 , n51033 , n51034 , n51035 , n51036 , 
     n51037 , n51038 , n51039 , n51040 , n51041 , n51042 , n51043 , n51044 , n51045 , n51046 , 
     n51047 , n51048 , n51049 , n51050 , n51051 , n51052 , n51053 , n51054 , n51055 , n51056 , 
     n51057 , n51058 , n51059 , n51060 , n51061 , n51062 , n51063 , n51064 , n51065 , n51066 , 
     n51067 , n51068 , n51069 , n51070 , n51071 , n51072 , n51073 , n51074 , n51075 , n51076 , 
     n51077 , n51078 , n51079 , n51080 , n51081 , n51082 , n51083 , n51084 , n51085 , n51086 , 
     n51087 , n51088 , n51089 , n51090 , n51091 , n51092 , n51093 , n51094 , n51095 , n51096 , 
     n51097 , n51098 , n51099 , n51100 , n51101 , n51102 , n51103 , n51104 , n51105 , n51106 , 
     n51107 , n51108 , n51109 , n51110 , n51111 , n51112 , n51113 , n51114 , n51115 , n51116 , 
     n51117 , n51118 , n51119 , n51120 , n51121 , n51122 , n51123 , n51124 , n51125 , n51126 , 
     n51127 , n51128 , n51129 , n51130 , n51131 , n51132 , n51133 , n51134 , n51135 , n51136 , 
     n51137 , n51138 , n51139 , n51140 , n51141 , n51142 , n51143 , n51144 , n51145 , n51146 , 
     n51147 , n51148 , n51149 , n51150 , n51151 , n51152 , n51153 , n51154 , n51155 , n51156 , 
     n51157 , n51158 , n51159 , n51160 , n51161 , n51162 , n51163 , n51164 , n51165 , n51166 , 
     n51167 , n51168 , n51169 , n51170 , n51171 , n51172 , n51173 , n51174 , n51175 , n51176 , 
     n51177 , n51178 , n51179 , n51180 , n51181 , n51182 , n51183 , n51184 , n51185 , n51186 , 
     n51187 , n51188 , n51189 , n51190 , n51191 , n51192 , n51193 , n51194 , n51195 , n51196 , 
     n51197 , n51198 , n51199 , n51200 , n51201 , n51202 , n51203 , n51204 , n51205 , n51206 , 
     n51207 , n51208 , n51209 , n51210 , n51211 , n51212 , n51213 , n51214 , n51215 , n51216 , 
     n51217 , n51218 , n51219 , n51220 , n51221 , n51222 , n51223 , n51224 , n51225 , n51226 , 
     n51227 , n51228 , n51229 , n51230 , n51231 , n51232 , n51233 , n51234 , n51235 , n51236 , 
     n51237 , n51238 , n51239 , n51240 , n51241 , n51242 , n51243 , n51244 , n51245 , n51246 , 
     n51247 , n51248 , n51249 , n51250 , n51251 , n51252 , n51253 , n51254 , n51255 , n51256 , 
     n51257 , n51258 , n51259 , n51260 , n51261 , n51262 , n51263 , n51264 , n51265 , n51266 , 
     n51267 , n51268 , n51269 , n51270 , n51271 , n51272 , n51273 , n51274 , n51275 , n51276 , 
     n51277 , n51278 , n51279 , n51280 , n51281 , n51282 , n51283 , n51284 , n51285 , n51286 , 
     n51287 , n51288 , n51289 , n51290 , n51291 , n51292 , n51293 , n51294 , n51295 , n51296 , 
     n51297 , n51298 , n51299 , n51300 , n51301 , n51302 , n51303 , n51304 , n51305 , n51306 , 
     n51307 , n51308 , n51309 , n51310 , n51311 , n51312 , n51313 , n51314 , n51315 , n51316 , 
     n51317 , n51318 , n51319 , n51320 , n51321 , n51322 , n51323 , n51324 , n51325 , n51326 , 
     n51327 , n51328 , n51329 , n51330 , n51331 , n51332 , n51333 , n51334 , n51335 , n51336 , 
     n51337 , n51338 , n51339 , n51340 , n51341 , n51342 , n51343 , n51344 , n51345 , n51346 , 
     n51347 , n51348 , n51349 , n51350 , n51351 , n51352 , n51353 , n51354 , n51355 , n51356 , 
     n51357 , n51358 , n51359 , n51360 , n51361 , n51362 , n51363 , n51364 , n51365 , n51366 , 
     n51367 , n51368 , n51369 , n51370 , n51371 , n51372 , n51373 , n51374 , n51375 , n51376 , 
     n51377 , n51378 , n51379 , n51380 , n51381 , n51382 , n51383 , n51384 , n51385 , n51386 , 
     n51387 , n51388 , n51389 , n51390 , n51391 , n51392 , n51393 , n51394 , n51395 , n51396 , 
     n51397 , n51398 , n51399 , n51400 , n51401 , n51402 , n51403 , n51404 , n51405 , n51406 , 
     n51407 , n51408 , n51409 , n51410 , n51411 , n51412 , n51413 , n51414 , n51415 , n51416 , 
     n51417 , n51418 , n51419 , n51420 , n51421 , n51422 , n51423 , n51424 , n51425 , n51426 , 
     n51427 , n51428 , n51429 , n51430 , n51431 , n51432 , n51433 , n51434 , n51435 , n51436 , 
     n51437 , n51438 , n51439 , n51440 , n51441 , n51442 , n51443 , n51444 , n51445 , n51446 , 
     n51447 , n51448 , n51449 , n51450 , n51451 , n51452 , n51453 , n51454 , n51455 , n51456 , 
     n51457 , n51458 , n51459 , n51460 , n51461 , n51462 , n51463 , n51464 , n51465 , n51466 , 
     n51467 , n51468 , n51469 , n51470 , n51471 , n51472 , n51473 , n51474 , n51475 , n51476 , 
     n51477 , n51478 , n51479 , n51480 , n51481 , n51482 , n51483 , n51484 , n51485 , n51486 , 
     n51487 , n51488 , n51489 , n51490 , n51491 , n51492 , n51493 , n51494 , n51495 , n51496 , 
     n51497 , n51498 , n51499 , n51500 , n51501 , n51502 , n51503 , n51504 , n51505 , n51506 , 
     n51507 , n51508 , n51509 , n51510 , n51511 , n51512 , n51513 , n51514 , n51515 , n51516 , 
     n51517 , n51518 , n51519 , n51520 , n51521 , n51522 , n51523 , n51524 , n51525 , n51526 , 
     n51527 , n51528 , n51529 , n51530 , n51531 , n51532 , n51533 , n51534 , n51535 , n51536 , 
     n51537 , n51538 , n51539 , n51540 , n51541 , n51542 , n51543 , n51544 , n51545 , n51546 , 
     n51547 , n51548 , n51549 , n51550 , n51551 , n51552 , n51553 , n51554 , n51555 , n51556 , 
     n51557 , n51558 , n51559 , n51560 , n51561 , n51562 , n51563 , n51564 , n51565 , n51566 , 
     n51567 , n51568 , n51569 , n51570 , n51571 , n51572 , n51573 , n51574 , n51575 , n51576 , 
     n51577 , n51578 , n51579 , n51580 , n51581 , n51582 , n51583 , n51584 , n51585 , n51586 , 
     n51587 , n51588 , n51589 , n51590 , n51591 , n51592 , n51593 , n51594 , n51595 , n51596 , 
     n51597 , n51598 , n51599 , n51600 , n51601 , n51602 , n51603 , n51604 , n51605 , n51606 , 
     n51607 , n51608 , n51609 , n51610 , n51611 , n51612 , n51613 , n51614 , n51615 , n51616 , 
     n51617 , n51618 , n51619 , n51620 , n51621 , n51622 , n51623 , n51624 , n51625 , n51626 , 
     n51627 , n51628 , n51629 , n51630 , n51631 , n51632 , n51633 , n51634 , n51635 , n51636 , 
     n51637 , n51638 , n51639 , n51640 , n51641 , n51642 , n51643 , n51644 , n51645 , n51646 , 
     n51647 , n51648 , n51649 , n51650 , n51651 , n51652 , n51653 , n51654 , n51655 , n51656 , 
     n51657 , n51658 , n51659 , n51660 , n51661 , n51662 , n51663 , n51664 , n51665 , n51666 , 
     n51667 , n51668 , n51669 , n51670 , n51671 , n51672 , n51673 , n51674 , n51675 , n51676 , 
     n51677 , n51678 , n51679 , n51680 , n51681 , n51682 , n51683 , n51684 , n51685 , n51686 , 
     n51687 , n51688 , n51689 , n51690 , n51691 , n51692 , n51693 , n51694 , n51695 , n51696 , 
     n51697 , n51698 , n51699 , n51700 , n51701 , n51702 , n51703 , n51704 , n51705 , n51706 , 
     n51707 , n51708 , n51709 , n51710 , n51711 , n51712 , n51713 , n51714 , n51715 , n51716 , 
     n51717 , n51718 , n51719 , n51720 , n51721 , n51722 , n51723 , n51724 , n51725 , n51726 , 
     n51727 , n51728 , n51729 , n51730 , n51731 , n51732 , n51733 , n51734 , n51735 , n51736 , 
     n51737 , n51738 , n51739 , n51740 , n51741 , n51742 , n51743 , n51744 , n51745 , n51746 , 
     n51747 , n51748 , n51749 , n51750 , n51751 , n51752 , n51753 , n51754 , n51755 , n51756 , 
     n51757 , n51758 , n51759 , n51760 , n51761 , n51762 , n51763 , n51764 , n51765 , n51766 , 
     n51767 , n51768 , n51769 , n51770 , n51771 , n51772 , n51773 , n51774 , n51775 , n51776 , 
     n51777 , n51778 , n51779 , n51780 , n51781 , n51782 , n51783 , n51784 , n51785 , n51786 , 
     n51787 , n51788 , n51789 , n51790 , n51791 , n51792 , n51793 , n51794 , n51795 , n51796 , 
     n51797 , n51798 , n51799 , n51800 , n51801 , n51802 , n51803 , n51804 , n51805 , n51806 , 
     n51807 , n51808 , n51809 , n51810 , n51811 , n51812 , n51813 , n51814 , n51815 , n51816 , 
     n51817 , n51818 , n51819 , n51820 , n51821 , n51822 , n51823 , n51824 , n51825 , n51826 , 
     n51827 , n51828 , n51829 , n51830 , n51831 , n51832 , n51833 , n51834 , n51835 , n51836 , 
     n51837 , n51838 , n51839 , n51840 , n51841 , n51842 , n51843 , n51844 , n51845 , n51846 , 
     n51847 , n51848 , n51849 , n51850 , n51851 , n51852 , n51853 , n51854 , n51855 , n51856 , 
     n51857 , n51858 , n51859 , n51860 , n51861 , n51862 , n51863 , n51864 , n51865 , n51866 , 
     n51867 , n51868 , n51869 , n51870 , n51871 , n51872 , n51873 , n51874 , n51875 , n51876 , 
     n51877 , n51878 , n51879 , n51880 , n51881 , n51882 , n51883 , n51884 , n51885 , n51886 , 
     n51887 , n51888 , n51889 , n51890 , n51891 , n51892 , n51893 , n51894 , n51895 , n51896 , 
     n51897 , n51898 , n51899 , n51900 , n51901 , n51902 , n51903 , n51904 , n51905 , n51906 , 
     n51907 , n51908 , n51909 , n51910 , n51911 , n51912 , n51913 , n51914 , n51915 , n51916 , 
     n51917 , n51918 , n51919 , n51920 , n51921 , n51922 , n51923 , n51924 , n51925 , n51926 , 
     n51927 , n51928 , n51929 , n51930 , n51931 , n51932 , n51933 , n51934 , n51935 , n51936 , 
     n51937 , n51938 , n51939 , n51940 , n51941 , n51942 , n51943 , n51944 , n51945 , n51946 , 
     n51947 , n51948 , n51949 , n51950 , n51951 , n51952 , n51953 , n51954 , n51955 , n51956 , 
     n51957 , n51958 , n51959 , n51960 , n51961 , n51962 , n51963 , n51964 , n51965 , n51966 , 
     n51967 , n51968 , n51969 , n51970 , n51971 , n51972 , n51973 , n51974 , n51975 , n51976 , 
     n51977 , n51978 , n51979 , n51980 , n51981 , n51982 , n51983 , n51984 , n51985 , n51986 , 
     n51987 , n51988 , n51989 , n51990 , n51991 , n51992 , n51993 , n51994 , n51995 , n51996 , 
     n51997 , n51998 , n51999 , n52000 , n52001 , n52002 , n52003 , n52004 , n52005 , n52006 , 
     n52007 , n52008 , n52009 , n52010 , n52011 , n52012 , n52013 , n52014 , n52015 , n52016 , 
     n52017 , n52018 , n52019 , n52020 , n52021 , n52022 , n52023 , n52024 , n52025 , n52026 , 
     n52027 , n52028 , n52029 , n52030 , n52031 , n52032 , n52033 , n52034 , n52035 , n52036 , 
     n52037 , n52038 , n52039 , n52040 , n52041 , n52042 , n52043 , n52044 , n52045 , n52046 , 
     n52047 , n52048 , n52049 , n52050 , n52051 , n52052 , n52053 , n52054 , n52055 , n52056 , 
     n52057 , n52058 , n52059 , n52060 , n52061 , n52062 , n52063 , n52064 , n52065 , n52066 , 
     n52067 , n52068 , n52069 , n52070 , n52071 , n52072 , n52073 , n52074 , n52075 , n52076 , 
     n52077 , n52078 , n52079 , n52080 , n52081 , n52082 , n52083 , n52084 , n52085 , n52086 , 
     n52087 , n52088 , n52089 , n52090 , n52091 , n52092 , n52093 , n52094 , n52095 , n52096 , 
     n52097 , n52098 , n52099 , n52100 , n52101 , n52102 , n52103 , n52104 , n52105 , n52106 , 
     n52107 , n52108 , n52109 , n52110 , n52111 , n52112 , n52113 , n52114 , n52115 , n52116 , 
     n52117 , n52118 , n52119 , n52120 , n52121 , n52122 , n52123 , n52124 , n52125 , n52126 , 
     n52127 , n52128 , n52129 , n52130 , n52131 , n52132 , n52133 , n52134 , n52135 , n52136 , 
     n52137 , n52138 , n52139 , n52140 , n52141 , n52142 , n52143 , n52144 , n52145 , n52146 , 
     n52147 , n52148 , n52149 , n52150 , n52151 , n52152 , n52153 , n52154 , n52155 , n52156 , 
     n52157 , n52158 , n52159 , n52160 , n52161 , n52162 , n52163 , n52164 , n52165 , n52166 , 
     n52167 , n52168 , n52169 , n52170 , n52171 , n52172 , n52173 , n52174 , n52175 , n52176 , 
     n52177 , n52178 , n52179 , n52180 , n52181 , n52182 , n52183 , n52184 , n52185 , n52186 , 
     n52187 , n52188 , n52189 , n52190 , n52191 , n52192 , n52193 , n52194 , n52195 , n52196 , 
     n52197 , n52198 , n52199 , n52200 , n52201 , n52202 , n52203 , n52204 , n52205 , n52206 , 
     n52207 , n52208 , n52209 , n52210 , n52211 , n52212 , n52213 , n52214 , n52215 , n52216 , 
     n52217 , n52218 , n52219 , n52220 , n52221 , n52222 , n52223 , n52224 , n52225 , n52226 , 
     n52227 , n52228 , n52229 , n52230 , n52231 , n52232 , n52233 , n52234 , n52235 , n52236 , 
     n52237 , n52238 , n52239 , n52240 , n52241 , n52242 , n52243 , n52244 , n52245 , n52246 , 
     n52247 , n52248 , n52249 , n52250 , n52251 , n52252 , n52253 , n52254 , n52255 , n52256 , 
     n52257 , n52258 , n52259 , n52260 , n52261 , n52262 , n52263 , n52264 , n52265 , n52266 , 
     n52267 , n52268 , n52269 , n52270 , n52271 , n52272 , n52273 , n52274 , n52275 , n52276 , 
     n52277 , n52278 , n52279 , n52280 , n52281 , n52282 , n52283 , n52284 , n52285 , n52286 , 
     n52287 , n52288 , n52289 , n52290 , n52291 , n52292 , n52293 , n52294 , n52295 , n52296 , 
     n52297 , n52298 , n52299 , n52300 , n52301 , n52302 , n52303 , n52304 , n52305 , n52306 , 
     n52307 , n52308 , n52309 , n52310 , n52311 , n52312 , n52313 , n52314 , n52315 , n52316 , 
     n52317 , n52318 , n52319 , n52320 , n52321 , n52322 , n52323 , n52324 , n52325 , n52326 , 
     n52327 , n52328 , n52329 , n52330 , n52331 , n52332 , n52333 , n52334 , n52335 , n52336 , 
     n52337 , n52338 , n52339 , n52340 , n52341 , n52342 , n52343 , n52344 , n52345 , n52346 , 
     n52347 , n52348 , n52349 , n52350 , n52351 , n52352 , n52353 , n52354 , n52355 , n52356 , 
     n52357 , n52358 , n52359 , n52360 , n52361 , n52362 , n52363 , n52364 , n52365 , n52366 , 
     n52367 , n52368 , n52369 , n52370 , n52371 , n52372 , n52373 , n52374 , n52375 , n52376 , 
     n52377 , n52378 , n52379 , n52380 , n52381 , n52382 , n52383 , n52384 , n52385 , n52386 , 
     n52387 , n52388 , n52389 , n52390 , n52391 , n52392 , n52393 , n52394 , n52395 , n52396 , 
     n52397 , n52398 , n52399 , n52400 , n52401 , n52402 , n52403 , n52404 , n52405 , n52406 , 
     n52407 , n52408 , n52409 , n52410 , n52411 , n52412 , n52413 , n52414 , n52415 , n52416 , 
     n52417 , n52418 , n52419 , n52420 , n52421 , n52422 , n52423 , n52424 , n52425 , n52426 , 
     n52427 , n52428 , n52429 , n52430 , n52431 , n52432 , n52433 , n52434 , n52435 , n52436 , 
     n52437 , n52438 , n52439 , n52440 , n52441 , n52442 , n52443 , n52444 , n52445 , n52446 , 
     n52447 , n52448 , n52449 , n52450 , n52451 , n52452 , n52453 , n52454 , n52455 , n52456 , 
     n52457 , n52458 , n52459 , n52460 , n52461 , n52462 , n52463 , n52464 , n52465 , n52466 , 
     n52467 , n52468 , n52469 , n52470 , n52471 , n52472 , n52473 , n52474 , n52475 , n52476 , 
     n52477 , n52478 , n52479 , n52480 , n52481 , n52482 , n52483 , n52484 , n52485 , n52486 , 
     n52487 , n52488 , n52489 , n52490 , n52491 , n52492 , n52493 , n52494 , n52495 , n52496 , 
     n52497 , n52498 , n52499 , n52500 , n52501 , n52502 , n52503 , n52504 , n52505 , n52506 , 
     n52507 , n52508 , n52509 , n52510 , n52511 , n52512 , n52513 , n52514 , n52515 , n52516 , 
     n52517 , n52518 , n52519 , n52520 , n52521 , n52522 , n52523 , n52524 , n52525 , n52526 , 
     n52527 , n52528 , n52529 , n52530 , n52531 , n52532 , n52533 , n52534 , n52535 , n52536 , 
     n52537 , n52538 , n52539 , n52540 , n52541 , n52542 , n52543 , n52544 , n52545 , n52546 , 
     n52547 , n52548 , n52549 , n52550 , n52551 , n52552 , n52553 , n52554 , n52555 , n52556 , 
     n52557 , n52558 , n52559 , n52560 , n52561 , n52562 , n52563 , n52564 , n52565 , n52566 , 
     n52567 , n52568 , n52569 , n52570 , n52571 , n52572 , n52573 , n52574 , n52575 , n52576 , 
     n52577 , n52578 , n52579 , n52580 , n52581 , n52582 , n52583 , n52584 , n52585 , n52586 , 
     n52587 , n52588 , n52589 , n52590 , n52591 , n52592 , n52593 , n52594 , n52595 , n52596 , 
     n52597 , n52598 , n52599 , n52600 , n52601 , n52602 , n52603 , n52604 , n52605 , n52606 , 
     n52607 , n52608 , n52609 , n52610 , n52611 , n52612 , n52613 , n52614 , n52615 , n52616 , 
     n52617 , n52618 , n52619 , n52620 , n52621 , n52622 , n52623 , n52624 , n52625 , n52626 , 
     n52627 , n52628 , n52629 , n52630 , n52631 , n52632 , n52633 , n52634 , n52635 , n52636 , 
     n52637 , n52638 , n52639 , n52640 , n52641 , n52642 , n52643 , n52644 , n52645 , n52646 , 
     n52647 , n52648 , n52649 , n52650 , n52651 , n52652 , n52653 , n52654 , n52655 , n52656 , 
     n52657 , n52658 , n52659 , n52660 , n52661 , n52662 , n52663 , n52664 , n52665 , n52666 , 
     n52667 , n52668 , n52669 , n52670 , n52671 , n52672 , n52673 , n52674 , n52675 , n52676 , 
     n52677 , n52678 , n52679 , n52680 , n52681 , n52682 , n52683 , n52684 , n52685 , n52686 , 
     n52687 , n52688 , n52689 , n52690 , n52691 , n52692 , n52693 , n52694 , n52695 , n52696 , 
     n52697 , n52698 , n52699 , n52700 , n52701 , n52702 , n52703 , n52704 , n52705 , n52706 , 
     n52707 , n52708 , n52709 , n52710 , n52711 , n52712 , n52713 , n52714 , n52715 , n52716 , 
     n52717 , n52718 , n52719 , n52720 , n52721 , n52722 , n52723 , n52724 , n52725 , n52726 , 
     n52727 , n52728 , n52729 , n52730 , n52731 , n52732 , n52733 , n52734 , n52735 , n52736 , 
     n52737 , n52738 , n52739 , n52740 , n52741 , n52742 , n52743 , n52744 , n52745 , n52746 , 
     n52747 , n52748 , n52749 , n52750 , n52751 , n52752 , n52753 , n52754 , n52755 , n52756 , 
     n52757 , n52758 , n52759 , n52760 , n52761 , n52762 , n52763 , n52764 , n52765 , n52766 , 
     n52767 , n52768 , n52769 , n52770 , n52771 , n52772 , n52773 , n52774 , n52775 , n52776 , 
     n52777 , n52778 , n52779 , n52780 , n52781 , n52782 , n52783 , n52784 , n52785 , n52786 , 
     n52787 , n52788 , n52789 , n52790 , n52791 , n52792 , n52793 , n52794 , n52795 , n52796 , 
     n52797 , n52798 , n52799 , n52800 , n52801 , n52802 , n52803 , n52804 , n52805 , n52806 , 
     n52807 , n52808 , n52809 , n52810 , n52811 , n52812 , n52813 , n52814 , n52815 , n52816 , 
     n52817 , n52818 , n52819 , n52820 , n52821 , n52822 , n52823 , n52824 , n52825 , n52826 , 
     n52827 , n52828 , n52829 , n52830 , n52831 , n52832 , n52833 , n52834 , n52835 , n52836 , 
     n52837 , n52838 , n52839 , n52840 , n52841 , n52842 , n52843 , n52844 , n52845 , n52846 , 
     n52847 , n52848 , n52849 , n52850 , n52851 , n52852 , n52853 , n52854 , n52855 , n52856 , 
     n52857 , n52858 , n52859 , n52860 , n52861 , n52862 , n52863 , n52864 , n52865 , n52866 , 
     n52867 , n52868 , n52869 , n52870 , n52871 , n52872 , n52873 , n52874 , n52875 , n52876 , 
     n52877 , n52878 , n52879 , n52880 , n52881 , n52882 , n52883 , n52884 , n52885 , n52886 , 
     n52887 , n52888 , n52889 , n52890 , n52891 , n52892 , n52893 , n52894 , n52895 , n52896 , 
     n52897 , n52898 , n52899 , n52900 , n52901 , n52902 , n52903 , n52904 , n52905 , n52906 , 
     n52907 , n52908 , n52909 , n52910 , n52911 , n52912 , n52913 , n52914 , n52915 , n52916 , 
     n52917 , n52918 , n52919 , n52920 , n52921 , n52922 , n52923 , n52924 , n52925 , n52926 , 
     n52927 , n52928 , n52929 , n52930 , n52931 , n52932 , n52933 , n52934 , n52935 , n52936 , 
     n52937 , n52938 , n52939 , n52940 , n52941 , n52942 , n52943 , n52944 , n52945 , n52946 , 
     n52947 , n52948 , n52949 , n52950 , n52951 , n52952 , n52953 , n52954 , n52955 , n52956 , 
     n52957 , n52958 , n52959 , n52960 , n52961 , n52962 , n52963 , n52964 , n52965 , n52966 , 
     n52967 , n52968 , n52969 , n52970 , n52971 , n52972 , n52973 , n52974 , n52975 , n52976 , 
     n52977 , n52978 , n52979 , n52980 , n52981 , n52982 , n52983 , n52984 , n52985 , n52986 , 
     n52987 , n52988 , n52989 , n52990 , n52991 , n52992 , n52993 , n52994 , n52995 , n52996 , 
     n52997 , n52998 , n52999 , n53000 , n53001 , n53002 , n53003 , n53004 , n53005 , n53006 , 
     n53007 , n53008 , n53009 , n53010 , n53011 , n53012 , n53013 , n53014 , n53015 , n53016 , 
     n53017 , n53018 , n53019 , n53020 , n53021 , n53022 , n53023 , n53024 , n53025 , n53026 , 
     n53027 , n53028 , n53029 , n53030 , n53031 , n53032 , n53033 , n53034 , n53035 , n53036 , 
     n53037 , n53038 , n53039 , n53040 , n53041 , n53042 , n53043 , n53044 , n53045 , n53046 , 
     n53047 , n53048 , n53049 , n53050 , n53051 , n53052 , n53053 , n53054 , n53055 , n53056 , 
     n53057 , n53058 , n53059 , n53060 , n53061 , n53062 , n53063 , n53064 , n53065 , n53066 , 
     n53067 , n53068 , n53069 , n53070 , n53071 , n53072 , n53073 , n53074 , n53075 , n53076 , 
     n53077 , n53078 , n53079 , n53080 , n53081 , n53082 , n53083 , n53084 , n53085 , n53086 , 
     n53087 , n53088 , n53089 , n53090 , n53091 , n53092 , n53093 , n53094 , n53095 , n53096 , 
     n53097 , n53098 , n53099 , n53100 , n53101 , n53102 , n53103 , n53104 , n53105 , n53106 , 
     n53107 , n53108 , n53109 , n53110 , n53111 , n53112 , n53113 , n53114 , n53115 , n53116 , 
     n53117 , n53118 , n53119 , n53120 , n53121 , n53122 , n53123 , n53124 , n53125 , n53126 , 
     n53127 , n53128 , n53129 , n53130 , n53131 , n53132 , n53133 , n53134 , n53135 , n53136 , 
     n53137 , n53138 , n53139 , n53140 , n53141 , n53142 , n53143 , n53144 , n53145 , n53146 , 
     n53147 , n53148 , n53149 , n53150 , n53151 , n53152 , n53153 , n53154 , n53155 , n53156 , 
     n53157 , n53158 , n53159 , n53160 , n53161 , n53162 , n53163 , n53164 , n53165 , n53166 , 
     n53167 , n53168 , n53169 , n53170 , n53171 , n53172 , n53173 , n53174 , n53175 , n53176 , 
     n53177 , n53178 , n53179 , n53180 , n53181 , n53182 , n53183 , n53184 , n53185 , n53186 , 
     n53187 , n53188 , n53189 , n53190 , n53191 , n53192 , n53193 , n53194 , n53195 , n53196 , 
     n53197 , n53198 , n53199 , n53200 , n53201 , n53202 , n53203 , n53204 , n53205 , n53206 , 
     n53207 , n53208 , n53209 , n53210 , n53211 , n53212 , n53213 , n53214 , n53215 , n53216 , 
     n53217 , n53218 , n53219 , n53220 , n53221 , n53222 , n53223 , n53224 , n53225 , n53226 , 
     n53227 , n53228 , n53229 , n53230 , n53231 , n53232 , n53233 , n53234 , n53235 , n53236 , 
     n53237 , n53238 , n53239 , n53240 , n53241 , n53242 , n53243 , n53244 , n53245 , n53246 , 
     n53247 , n53248 , n53249 , n53250 , n53251 , n53252 , n53253 , n53254 , n53255 , n53256 , 
     n53257 , n53258 , n53259 , n53260 , n53261 , n53262 , n53263 , n53264 , n53265 , n53266 , 
     n53267 , n53268 , n53269 , n53270 , n53271 , n53272 , n53273 , n53274 , n53275 , n53276 , 
     n53277 , n53278 , n53279 , n53280 , n53281 , n53282 , n53283 , n53284 , n53285 , n53286 , 
     n53287 , n53288 , n53289 , n53290 , n53291 , n53292 , n53293 , n53294 , n53295 , n53296 , 
     n53297 , n53298 , n53299 , n53300 , n53301 , n53302 , n53303 , n53304 , n53305 , n53306 , 
     n53307 , n53308 , n53309 , n53310 , n53311 , n53312 , n53313 , n53314 , n53315 , n53316 , 
     n53317 , n53318 , n53319 , n53320 , n53321 , n53322 , n53323 , n53324 , n53325 , n53326 , 
     n53327 , n53328 , n53329 , n53330 , n53331 , n53332 , n53333 , n53334 , n53335 , n53336 , 
     n53337 , n53338 , n53339 , n53340 , n53341 , n53342 , n53343 , n53344 , n53345 , n53346 , 
     n53347 , n53348 , n53349 , n53350 , n53351 , n53352 , n53353 , n53354 , n53355 , n53356 , 
     n53357 , n53358 , n53359 , n53360 , n53361 , n53362 , n53363 , n53364 , n53365 , n53366 , 
     n53367 , n53368 , n53369 , n53370 , n53371 , n53372 , n53373 , n53374 , n53375 , n53376 , 
     n53377 , n53378 , n53379 , n53380 , n53381 , n53382 , n53383 , n53384 , n53385 , n53386 , 
     n53387 , n53388 , n53389 , n53390 , n53391 , n53392 , n53393 , n53394 , n53395 , n53396 , 
     n53397 , n53398 , n53399 , n53400 , n53401 , n53402 , n53403 , n53404 , n53405 , n53406 , 
     n53407 , n53408 , n53409 , n53410 , n53411 , n53412 , n53413 , n53414 , n53415 , n53416 , 
     n53417 , n53418 , n53419 , n53420 , n53421 , n53422 , n53423 , n53424 , n53425 , n53426 , 
     n53427 , n53428 , n53429 , n53430 , n53431 , n53432 , n53433 , n53434 , n53435 , n53436 , 
     n53437 , n53438 , n53439 , n53440 , n53441 , n53442 , n53443 , n53444 , n53445 , n53446 , 
     n53447 , n53448 , n53449 , n53450 , n53451 , n53452 , n53453 , n53454 , n53455 , n53456 , 
     n53457 , n53458 , n53459 , n53460 , n53461 , n53462 , n53463 , n53464 , n53465 , n53466 , 
     n53467 , n53468 , n53469 , n53470 , n53471 , n53472 , n53473 , n53474 , n53475 , n53476 , 
     n53477 , n53478 , n53479 , n53480 , n53481 , n53482 , n53483 , n53484 , n53485 , n53486 , 
     n53487 , n53488 , n53489 , n53490 , n53491 , n53492 , n53493 , n53494 , n53495 , n53496 , 
     n53497 , n53498 , n53499 , n53500 , n53501 , n53502 , n53503 , n53504 , n53505 , n53506 , 
     n53507 , n53508 , n53509 , n53510 , n53511 , n53512 , n53513 , n53514 , n53515 , n53516 , 
     n53517 , n53518 , n53519 , n53520 , n53521 , n53522 , n53523 , n53524 , n53525 , n53526 , 
     n53527 , n53528 , n53529 , n53530 , n53531 , n53532 , n53533 , n53534 , n53535 , n53536 , 
     n53537 , n53538 , n53539 , n53540 , n53541 , n53542 , n53543 , n53544 , n53545 , n53546 , 
     n53547 , n53548 , n53549 , n53550 , n53551 , n53552 , n53553 , n53554 , n53555 , n53556 , 
     n53557 , n53558 , n53559 , n53560 , n53561 , n53562 , n53563 , n53564 , n53565 , n53566 , 
     n53567 , n53568 , n53569 , n53570 , n53571 , n53572 , n53573 , n53574 , n53575 , n53576 , 
     n53577 , n53578 , n53579 , n53580 , n53581 , n53582 , n53583 , n53584 , n53585 , n53586 , 
     n53587 , n53588 , n53589 , n53590 , n53591 , n53592 , n53593 , n53594 , n53595 , n53596 , 
     n53597 , n53598 , n53599 , n53600 , n53601 , n53602 , n53603 , n53604 , n53605 , n53606 , 
     n53607 , n53608 , n53609 , n53610 , n53611 , n53612 , n53613 , n53614 , n53615 , n53616 , 
     n53617 , n53618 , n53619 , n53620 , n53621 , n53622 , n53623 , n53624 , n53625 , n53626 , 
     n53627 , n53628 , n53629 , n53630 , n53631 , n53632 , n53633 , n53634 , n53635 , n53636 , 
     n53637 , n53638 , n53639 , n53640 , n53641 , n53642 , n53643 , n53644 , n53645 , n53646 , 
     n53647 , n53648 , n53649 , n53650 , n53651 , n53652 , n53653 , n53654 , n53655 , n53656 , 
     n53657 , n53658 , n53659 , n53660 , n53661 , n53662 , n53663 , n53664 , n53665 , n53666 , 
     n53667 , n53668 , n53669 , n53670 , n53671 , n53672 , n53673 , n53674 , n53675 , n53676 , 
     n53677 , n53678 , n53679 , n53680 , n53681 , n53682 , n53683 , n53684 , n53685 , n53686 , 
     n53687 , n53688 , n53689 , n53690 , n53691 , n53692 , n53693 , n53694 , n53695 , n53696 , 
     n53697 , n53698 , n53699 , n53700 , n53701 , n53702 , n53703 , n53704 , n53705 , n53706 , 
     n53707 , n53708 , n53709 , n53710 , n53711 , n53712 , n53713 , n53714 , n53715 , n53716 , 
     n53717 , n53718 , n53719 , n53720 , n53721 , n53722 , n53723 , n53724 , n53725 , n53726 , 
     n53727 , n53728 , n53729 , n53730 , n53731 , n53732 , n53733 , n53734 , n53735 , n53736 , 
     n53737 , n53738 , n53739 , n53740 , n53741 , n53742 , n53743 , n53744 , n53745 , n53746 , 
     n53747 , n53748 , n53749 , n53750 , n53751 , n53752 , n53753 , n53754 , n53755 , n53756 , 
     n53757 , n53758 , n53759 , n53760 , n53761 , n53762 , n53763 , n53764 , n53765 , n53766 , 
     n53767 , n53768 , n53769 , n53770 , n53771 , n53772 , n53773 , n53774 , n53775 , n53776 , 
     n53777 , n53778 , n53779 , n53780 , n53781 , n53782 , n53783 , n53784 , n53785 , n53786 , 
     n53787 , n53788 , n53789 , n53790 , n53791 , n53792 , n53793 , n53794 , n53795 , n53796 , 
     n53797 , n53798 , n53799 , n53800 , n53801 , n53802 , n53803 , n53804 , n53805 , n53806 , 
     n53807 , n53808 , n53809 , n53810 , n53811 , n53812 , n53813 , n53814 , n53815 , n53816 , 
     n53817 , n53818 , n53819 , n53820 , n53821 , n53822 , n53823 , n53824 , n53825 , n53826 , 
     n53827 , n53828 , n53829 , n53830 , n53831 , n53832 , n53833 , n53834 , n53835 , n53836 , 
     n53837 , n53838 , n53839 , n53840 , n53841 , n53842 , n53843 , n53844 , n53845 , n53846 , 
     n53847 , n53848 , n53849 , n53850 , n53851 , n53852 , n53853 , n53854 , n53855 , n53856 , 
     n53857 , n53858 , n53859 , n53860 , n53861 , n53862 , n53863 , n53864 , n53865 , n53866 , 
     n53867 , n53868 , n53869 , n53870 , n53871 , n53872 , n53873 , n53874 , n53875 , n53876 , 
     n53877 , n53878 , n53879 , n53880 , n53881 , n53882 , n53883 , n53884 , n53885 , n53886 , 
     n53887 , n53888 , n53889 , n53890 , n53891 , n53892 , n53893 , n53894 , n53895 , n53896 , 
     n53897 , n53898 , n53899 , n53900 , n53901 , n53902 , n53903 , n53904 , n53905 , n53906 , 
     n53907 , n53908 , n53909 , n53910 , n53911 , n53912 , n53913 , n53914 , n53915 , n53916 , 
     n53917 , n53918 , n53919 , n53920 , n53921 , n53922 , n53923 , n53924 , n53925 , n53926 , 
     n53927 , n53928 , n53929 , n53930 , n53931 , n53932 , n53933 , n53934 , n53935 , n53936 , 
     n53937 , n53938 , n53939 , n53940 , n53941 , n53942 , n53943 , n53944 , n53945 , n53946 , 
     n53947 , n53948 , n53949 , n53950 , n53951 , n53952 , n53953 , n53954 , n53955 , n53956 , 
     n53957 , n53958 , n53959 , n53960 , n53961 , n53962 , n53963 , n53964 , n53965 , n53966 , 
     n53967 , n53968 , n53969 , n53970 , n53971 , n53972 , n53973 , n53974 , n53975 , n53976 , 
     n53977 , n53978 , n53979 , n53980 , n53981 , n53982 , n53983 , n53984 , n53985 , n53986 , 
     n53987 , n53988 , n53989 , n53990 , n53991 , n53992 , n53993 , n53994 , n53995 , n53996 , 
     n53997 , n53998 , n53999 , n54000 , n54001 , n54002 , n54003 , n54004 , n54005 , n54006 , 
     n54007 , n54008 , n54009 , n54010 , n54011 , n54012 , n54013 , n54014 , n54015 , n54016 , 
     n54017 , n54018 , n54019 , n54020 , n54021 , n54022 , n54023 , n54024 , n54025 , n54026 , 
     n54027 , n54028 , n54029 , n54030 , n54031 , n54032 , n54033 , n54034 , n54035 , n54036 , 
     n54037 , n54038 , n54039 , n54040 , n54041 , n54042 , n54043 , n54044 , n54045 , n54046 , 
     n54047 , n54048 , n54049 , n54050 , n54051 , n54052 , n54053 , n54054 , n54055 , n54056 , 
     n54057 , n54058 , n54059 , n54060 , n54061 , n54062 , n54063 , n54064 , n54065 , n54066 , 
     n54067 , n54068 , n54069 , n54070 , n54071 , n54072 , n54073 , n54074 , n54075 , n54076 , 
     n54077 , n54078 , n54079 , n54080 , n54081 , n54082 , n54083 , n54084 , n54085 , n54086 , 
     n54087 , n54088 , n54089 , n54090 , n54091 , n54092 , n54093 , n54094 , n54095 , n54096 , 
     n54097 , n54098 , n54099 , n54100 , n54101 , n54102 , n54103 , n54104 , n54105 , n54106 , 
     n54107 , n54108 , n54109 , n54110 , n54111 , n54112 , n54113 , n54114 , n54115 , n54116 , 
     n54117 , n54118 , n54119 , n54120 , n54121 , n54122 , n54123 , n54124 , n54125 , n54126 , 
     n54127 , n54128 , n54129 , n54130 , n54131 , n54132 , n54133 , n54134 , n54135 , n54136 , 
     n54137 , n54138 , n54139 , n54140 , n54141 , n54142 , n54143 , n54144 , n54145 , n54146 , 
     n54147 , n54148 , n54149 , n54150 , n54151 , n54152 , n54153 , n54154 , n54155 , n54156 , 
     n54157 , n54158 , n54159 , n54160 , n54161 , n54162 , n54163 , n54164 , n54165 , n54166 , 
     n54167 , n54168 , n54169 , n54170 , n54171 , n54172 , n54173 , n54174 , n54175 , n54176 , 
     n54177 , n54178 , n54179 , n54180 , n54181 , n54182 , n54183 , n54184 , n54185 , n54186 , 
     n54187 , n54188 , n54189 , n54190 , n54191 , n54192 , n54193 , n54194 , n54195 , n54196 , 
     n54197 , n54198 , n54199 , n54200 , n54201 , n54202 , n54203 , n54204 , n54205 , n54206 , 
     n54207 , n54208 , n54209 , n54210 , n54211 , n54212 , n54213 , n54214 , n54215 , n54216 , 
     n54217 , n54218 , n54219 , n54220 , n54221 , n54222 , n54223 , n54224 , n54225 , n54226 , 
     n54227 , n54228 , n54229 , n54230 , n54231 , n54232 , n54233 , n54234 , n54235 , n54236 , 
     n54237 , n54238 , n54239 , n54240 , n54241 , n54242 , n54243 , n54244 , n54245 , n54246 , 
     n54247 , n54248 , n54249 , n54250 , n54251 , n54252 , n54253 , n54254 , n54255 , n54256 , 
     n54257 , n54258 , n54259 , n54260 , n54261 , n54262 , n54263 , n54264 , n54265 , n54266 , 
     n54267 , n54268 , n54269 , n54270 , n54271 , n54272 , n54273 , n54274 , n54275 , n54276 , 
     n54277 , n54278 , n54279 , n54280 , n54281 , n54282 , n54283 , n54284 , n54285 , n54286 , 
     n54287 , n54288 , n54289 , n54290 , n54291 , n54292 , n54293 , n54294 , n54295 , n54296 , 
     n54297 , n54298 , n54299 , n54300 , n54301 , n54302 , n54303 , n54304 , n54305 , n54306 , 
     n54307 , n54308 , n54309 , n54310 , n54311 , n54312 , n54313 , n54314 , n54315 , n54316 , 
     n54317 , n54318 , n54319 , n54320 , n54321 , n54322 , n54323 , n54324 , n54325 , n54326 , 
     n54327 , n54328 , n54329 , n54330 , n54331 , n54332 , n54333 , n54334 , n54335 , n54336 , 
     n54337 , n54338 , n54339 , n54340 , n54341 , n54342 , n54343 , n54344 , n54345 , n54346 , 
     n54347 , n54348 , n54349 , n54350 , n54351 , n54352 , n54353 , n54354 , n54355 , n54356 , 
     n54357 , n54358 , n54359 , n54360 , n54361 , n54362 , n54363 , n54364 , n54365 , n54366 , 
     n54367 , n54368 , n54369 , n54370 , n54371 , n54372 , n54373 , n54374 , n54375 , n54376 , 
     n54377 , n54378 , n54379 , n54380 , n54381 , n54382 , n54383 , n54384 , n54385 , n54386 , 
     n54387 , n54388 , n54389 , n54390 , n54391 , n54392 , n54393 , n54394 , n54395 , n54396 , 
     n54397 , n54398 , n54399 , n54400 , n54401 , n54402 , n54403 , n54404 , n54405 , n54406 , 
     n54407 , n54408 , n54409 , n54410 , n54411 , n54412 , n54413 , n54414 , n54415 , n54416 , 
     n54417 , n54418 , n54419 , n54420 , n54421 , n54422 , n54423 , n54424 , n54425 , n54426 , 
     n54427 , n54428 , n54429 , n54430 , n54431 , n54432 , n54433 , n54434 , n54435 , n54436 , 
     n54437 , n54438 , n54439 , n54440 , n54441 , n54442 , n54443 , n54444 , n54445 , n54446 , 
     n54447 , n54448 , n54449 , n54450 , n54451 , n54452 , n54453 , n54454 , n54455 , n54456 , 
     n54457 , n54458 , n54459 , n54460 , n54461 , n54462 , n54463 , n54464 , n54465 , n54466 , 
     n54467 , n54468 , n54469 , n54470 , n54471 , n54472 , n54473 , n54474 , n54475 , n54476 , 
     n54477 , n54478 , n54479 , n54480 , n54481 , n54482 , n54483 , n54484 , n54485 , n54486 , 
     n54487 , n54488 , n54489 , n54490 , n54491 , n54492 , n54493 , n54494 , n54495 , n54496 , 
     n54497 , n54498 , n54499 , n54500 , n54501 , n54502 , n54503 , n54504 , n54505 , n54506 , 
     n54507 , n54508 , n54509 , n54510 , n54511 , n54512 , n54513 , n54514 , n54515 , n54516 , 
     n54517 , n54518 , n54519 , n54520 , n54521 , n54522 , n54523 , n54524 , n54525 , n54526 , 
     n54527 , n54528 , n54529 , n54530 , n54531 , n54532 , n54533 , n54534 , n54535 , n54536 , 
     n54537 , n54538 , n54539 , n54540 , n54541 , n54542 , n54543 , n54544 , n54545 , n54546 , 
     n54547 , n54548 , n54549 , n54550 , n54551 , n54552 , n54553 , n54554 , n54555 , n54556 , 
     n54557 , n54558 , n54559 , n54560 , n54561 , n54562 , n54563 , n54564 , n54565 , n54566 , 
     n54567 , n54568 , n54569 , n54570 , n54571 , n54572 , n54573 , n54574 , n54575 , n54576 , 
     n54577 , n54578 , n54579 , n54580 , n54581 , n54582 , n54583 , n54584 , n54585 , n54586 , 
     n54587 , n54588 , n54589 , n54590 , n54591 , n54592 , n54593 , n54594 , n54595 , n54596 , 
     n54597 , n54598 , n54599 , n54600 , n54601 , n54602 , n54603 , n54604 , n54605 , n54606 , 
     n54607 , n54608 , n54609 , n54610 , n54611 , n54612 , n54613 , n54614 , n54615 , n54616 , 
     n54617 , n54618 , n54619 , n54620 , n54621 , n54622 , n54623 , n54624 , n54625 , n54626 , 
     n54627 , n54628 , n54629 , n54630 , n54631 , n54632 , n54633 , n54634 , n54635 , n54636 , 
     n54637 , n54638 , n54639 , n54640 , n54641 , n54642 , n54643 , n54644 , n54645 , n54646 , 
     n54647 , n54648 , n54649 , n54650 , n54651 , n54652 , n54653 , n54654 , n54655 , n54656 , 
     n54657 , n54658 , n54659 , n54660 , n54661 , n54662 , n54663 , n54664 , n54665 , n54666 , 
     n54667 , n54668 , n54669 , n54670 , n54671 , n54672 , n54673 , n54674 , n54675 , n54676 , 
     n54677 , n54678 , n54679 , n54680 , n54681 , n54682 , n54683 , n54684 , n54685 , n54686 , 
     n54687 , n54688 , n54689 , n54690 , n54691 , n54692 , n54693 , n54694 , n54695 , n54696 , 
     n54697 , n54698 , n54699 , n54700 , n54701 , n54702 , n54703 , n54704 , n54705 , n54706 , 
     n54707 , n54708 , n54709 , n54710 , n54711 , n54712 , n54713 , n54714 , n54715 , n54716 , 
     n54717 , n54718 , n54719 , n54720 , n54721 , n54722 , n54723 , n54724 , n54725 , n54726 , 
     n54727 , n54728 , n54729 , n54730 , n54731 , n54732 , n54733 , n54734 , n54735 , n54736 , 
     n54737 , n54738 , n54739 , n54740 , n54741 , n54742 , n54743 , n54744 , n54745 , n54746 , 
     n54747 , n54748 , n54749 , n54750 , n54751 , n54752 , n54753 , n54754 , n54755 , n54756 , 
     n54757 , n54758 , n54759 , n54760 , n54761 , n54762 , n54763 , n54764 , n54765 , n54766 , 
     n54767 , n54768 , n54769 , n54770 , n54771 , n54772 , n54773 , n54774 , n54775 , n54776 , 
     n54777 , n54778 , n54779 , n54780 , n54781 , n54782 , n54783 , n54784 , n54785 , n54786 , 
     n54787 , n54788 , n54789 , n54790 , n54791 , n54792 , n54793 , n54794 , n54795 , n54796 , 
     n54797 , n54798 , n54799 , n54800 , n54801 , n54802 , n54803 , n54804 , n54805 , n54806 , 
     n54807 , n54808 , n54809 , n54810 , n54811 , n54812 , n54813 , n54814 , n54815 , n54816 , 
     n54817 , n54818 , n54819 , n54820 , n54821 , n54822 , n54823 , n54824 , n54825 , n54826 , 
     n54827 , n54828 , n54829 , n54830 , n54831 , n54832 , n54833 , n54834 , n54835 , n54836 , 
     n54837 , n54838 , n54839 , n54840 , n54841 , n54842 , n54843 , n54844 , n54845 , n54846 , 
     n54847 , n54848 , n54849 , n54850 , n54851 , n54852 , n54853 , n54854 , n54855 , n54856 , 
     n54857 , n54858 , n54859 , n54860 , n54861 , n54862 , n54863 , n54864 , n54865 , n54866 , 
     n54867 , n54868 , n54869 , n54870 , n54871 , n54872 , n54873 , n54874 , n54875 , n54876 , 
     n54877 , n54878 , n54879 , n54880 , n54881 , n54882 , n54883 , n54884 , n54885 , n54886 , 
     n54887 , n54888 , n54889 , n54890 , n54891 , n54892 , n54893 , n54894 , n54895 , n54896 , 
     n54897 , n54898 , n54899 , n54900 , n54901 , n54902 , n54903 , n54904 , n54905 , n54906 , 
     n54907 , n54908 , n54909 , n54910 , n54911 , n54912 , n54913 , n54914 , n54915 , n54916 , 
     n54917 , n54918 , n54919 , n54920 , n54921 , n54922 , n54923 , n54924 , n54925 , n54926 , 
     n54927 , n54928 , n54929 , n54930 , n54931 , n54932 , n54933 , n54934 , n54935 , n54936 , 
     n54937 , n54938 , n54939 , n54940 , n54941 , n54942 , n54943 , n54944 , n54945 , n54946 , 
     n54947 , n54948 , n54949 , n54950 , n54951 , n54952 , n54953 , n54954 , n54955 , n54956 , 
     n54957 , n54958 , n54959 , n54960 , n54961 , n54962 , n54963 , n54964 , n54965 , n54966 , 
     n54967 , n54968 , n54969 , n54970 , n54971 , n54972 , n54973 , n54974 , n54975 , n54976 , 
     n54977 , n54978 , n54979 , n54980 , n54981 , n54982 , n54983 , n54984 , n54985 , n54986 , 
     n54987 , n54988 , n54989 , n54990 , n54991 , n54992 , n54993 , n54994 , n54995 , n54996 , 
     n54997 , n54998 , n54999 , n55000 , n55001 , n55002 , n55003 , n55004 , n55005 , n55006 , 
     n55007 , n55008 , n55009 , n55010 , n55011 , n55012 , n55013 , n55014 , n55015 , n55016 , 
     n55017 , n55018 , n55019 , n55020 , n55021 , n55022 , n55023 , n55024 , n55025 , n55026 , 
     n55027 , n55028 , n55029 , n55030 , n55031 , n55032 , n55033 , n55034 , n55035 , n55036 , 
     n55037 , n55038 , n55039 , n55040 , n55041 , n55042 , n55043 , n55044 , n55045 , n55046 , 
     n55047 , n55048 , n55049 , n55050 , n55051 , n55052 , n55053 , n55054 , n55055 , n55056 , 
     n55057 , n55058 , n55059 , n55060 , n55061 , n55062 , n55063 , n55064 , n55065 , n55066 , 
     n55067 , n55068 , n55069 , n55070 , n55071 , n55072 , n55073 , n55074 , n55075 , n55076 , 
     n55077 , n55078 , n55079 , n55080 , n55081 , n55082 , n55083 , n55084 , n55085 , n55086 , 
     n55087 , n55088 , n55089 , n55090 , n55091 , n55092 , n55093 , n55094 , n55095 , n55096 , 
     n55097 , n55098 , n55099 , n55100 , n55101 , n55102 , n55103 , n55104 , n55105 , n55106 , 
     n55107 , n55108 , n55109 , n55110 , n55111 , n55112 , n55113 , n55114 , n55115 , n55116 , 
     n55117 , n55118 , n55119 , n55120 , n55121 , n55122 , n55123 , n55124 , n55125 , n55126 , 
     n55127 , n55128 , n55129 , n55130 , n55131 , n55132 , n55133 , n55134 , n55135 , n55136 , 
     n55137 , n55138 , n55139 , n55140 , n55141 , n55142 , n55143 , n55144 , n55145 , n55146 , 
     n55147 , n55148 , n55149 , n55150 , n55151 , n55152 , n55153 , n55154 , n55155 , n55156 , 
     n55157 , n55158 , n55159 , n55160 , n55161 , n55162 , n55163 , n55164 , n55165 , n55166 , 
     n55167 , n55168 , n55169 , n55170 , n55171 , n55172 , n55173 , n55174 , n55175 , n55176 , 
     n55177 , n55178 , n55179 , n55180 , n55181 , n55182 , n55183 , n55184 , n55185 , n55186 , 
     n55187 , n55188 , n55189 , n55190 , n55191 , n55192 , n55193 , n55194 , n55195 , n55196 , 
     n55197 , n55198 , n55199 , n55200 , n55201 , n55202 , n55203 , n55204 , n55205 , n55206 , 
     n55207 , n55208 , n55209 , n55210 , n55211 , n55212 , n55213 , n55214 , n55215 , n55216 , 
     n55217 , n55218 , n55219 , n55220 , n55221 , n55222 , n55223 , n55224 , n55225 , n55226 , 
     n55227 , n55228 , n55229 , n55230 , n55231 , n55232 , n55233 , n55234 , n55235 , n55236 , 
     n55237 , n55238 , n55239 , n55240 , n55241 , n55242 , n55243 , n55244 , n55245 , n55246 , 
     n55247 , n55248 , n55249 , n55250 , n55251 , n55252 , n55253 , n55254 , n55255 , n55256 , 
     n55257 , n55258 , n55259 , n55260 , n55261 , n55262 , n55263 , n55264 , n55265 , n55266 , 
     n55267 , n55268 , n55269 , n55270 , n55271 , n55272 , n55273 , n55274 , n55275 , n55276 , 
     n55277 , n55278 , n55279 , n55280 , n55281 , n55282 , n55283 , n55284 , n55285 , n55286 , 
     n55287 , n55288 , n55289 , n55290 , n55291 , n55292 , n55293 , n55294 , n55295 , n55296 , 
     n55297 , n55298 , n55299 , n55300 , n55301 , n55302 , n55303 , n55304 , n55305 , n55306 , 
     n55307 , n55308 , n55309 , n55310 , n55311 , n55312 , n55313 , n55314 , n55315 , n55316 , 
     n55317 , n55318 , n55319 , n55320 , n55321 , n55322 , n55323 , n55324 , n55325 , n55326 , 
     n55327 , n55328 , n55329 , n55330 , n55331 , n55332 , n55333 , n55334 , n55335 , n55336 , 
     n55337 , n55338 , n55339 , n55340 , n55341 , n55342 , n55343 , n55344 , n55345 , n55346 , 
     n55347 , n55348 , n55349 , n55350 , n55351 , n55352 , n55353 , n55354 , n55355 , n55356 , 
     n55357 , n55358 , n55359 , n55360 , n55361 , n55362 , n55363 , n55364 , n55365 , n55366 , 
     n55367 , n55368 , n55369 , n55370 , n55371 , n55372 , n55373 , n55374 , n55375 , n55376 , 
     n55377 , n55378 , n55379 , n55380 , n55381 , n55382 , n55383 , n55384 , n55385 , n55386 , 
     n55387 , n55388 , n55389 , n55390 , n55391 , n55392 , n55393 , n55394 , n55395 , n55396 , 
     n55397 , n55398 , n55399 , n55400 , n55401 , n55402 , n55403 , n55404 , n55405 , n55406 , 
     n55407 , n55408 , n55409 , n55410 , n55411 , n55412 , n55413 , n55414 , n55415 , n55416 , 
     n55417 , n55418 , n55419 , n55420 , n55421 , n55422 , n55423 , n55424 , n55425 , n55426 , 
     n55427 , n55428 , n55429 , n55430 , n55431 , n55432 , n55433 , n55434 , n55435 , n55436 , 
     n55437 , n55438 , n55439 , n55440 , n55441 , n55442 , n55443 , n55444 , n55445 , n55446 , 
     n55447 , n55448 , n55449 , n55450 , n55451 , n55452 , n55453 , n55454 , n55455 , n55456 , 
     n55457 , n55458 , n55459 , n55460 , n55461 , n55462 , n55463 , n55464 , n55465 , n55466 , 
     n55467 , n55468 , n55469 , n55470 , n55471 , n55472 , n55473 , n55474 , n55475 , n55476 , 
     n55477 , n55478 , n55479 , n55480 , n55481 , n55482 , n55483 , n55484 , n55485 , n55486 , 
     n55487 , n55488 , n55489 , n55490 , n55491 , n55492 , n55493 , n55494 , n55495 , n55496 , 
     n55497 , n55498 , n55499 , n55500 , n55501 , n55502 , n55503 , n55504 , n55505 , n55506 , 
     n55507 , n55508 , n55509 , n55510 , n55511 , n55512 , n55513 , n55514 , n55515 , n55516 , 
     n55517 , n55518 , n55519 , n55520 , n55521 , n55522 , n55523 , n55524 , n55525 , n55526 , 
     n55527 , n55528 , n55529 , n55530 , n55531 , n55532 , n55533 , n55534 , n55535 , n55536 , 
     n55537 , n55538 , n55539 , n55540 , n55541 , n55542 , n55543 , n55544 , n55545 , n55546 , 
     n55547 , n55548 , n55549 , n55550 , n55551 , n55552 , n55553 , n55554 , n55555 , n55556 , 
     n55557 , n55558 , n55559 , n55560 , n55561 , n55562 , n55563 , n55564 , n55565 , n55566 , 
     n55567 , n55568 , n55569 , n55570 , n55571 , n55572 , n55573 , n55574 , n55575 , n55576 , 
     n55577 , n55578 , n55579 , n55580 , n55581 , n55582 , n55583 , n55584 , n55585 , n55586 , 
     n55587 , n55588 , n55589 , n55590 , n55591 , n55592 , n55593 , n55594 , n55595 , n55596 , 
     n55597 , n55598 , n55599 , n55600 , n55601 , n55602 , n55603 , n55604 , n55605 , n55606 , 
     n55607 , n55608 , n55609 , n55610 , n55611 , n55612 , n55613 , n55614 , n55615 , n55616 , 
     n55617 , n55618 , n55619 , n55620 , n55621 , n55622 , n55623 , n55624 , n55625 , n55626 , 
     n55627 , n55628 , n55629 , n55630 , n55631 , n55632 , n55633 , n55634 , n55635 , n55636 , 
     n55637 , n55638 , n55639 , n55640 , n55641 , n55642 , n55643 , n55644 , n55645 , n55646 , 
     n55647 , n55648 , n55649 , n55650 , n55651 , n55652 , n55653 , n55654 , n55655 , n55656 , 
     n55657 , n55658 , n55659 , n55660 , n55661 , n55662 , n55663 , n55664 , n55665 , n55666 , 
     n55667 , n55668 , n55669 , n55670 , n55671 , n55672 , n55673 , n55674 , n55675 , n55676 , 
     n55677 , n55678 , n55679 , n55680 , n55681 , n55682 , n55683 , n55684 , n55685 , n55686 , 
     n55687 , n55688 , n55689 , n55690 , n55691 , n55692 , n55693 , n55694 , n55695 , n55696 , 
     n55697 , n55698 , n55699 , n55700 , n55701 , n55702 , n55703 , n55704 , n55705 , n55706 , 
     n55707 , n55708 , n55709 , n55710 , n55711 , n55712 , n55713 , n55714 , n55715 , n55716 , 
     n55717 , n55718 , n55719 , n55720 , n55721 , n55722 , n55723 , n55724 , n55725 , n55726 , 
     n55727 , n55728 , n55729 , n55730 , n55731 , n55732 , n55733 , n55734 , n55735 , n55736 , 
     n55737 , n55738 , n55739 , n55740 , n55741 , n55742 , n55743 , n55744 , n55745 , n55746 , 
     n55747 , n55748 , n55749 , n55750 , n55751 , n55752 , n55753 , n55754 , n55755 , n55756 , 
     n55757 , n55758 , n55759 , n55760 , n55761 , n55762 , n55763 , n55764 , n55765 , n55766 , 
     n55767 , n55768 , n55769 , n55770 , n55771 , n55772 , n55773 , n55774 , n55775 , n55776 , 
     n55777 , n55778 , n55779 , n55780 , n55781 , n55782 , n55783 , n55784 , n55785 , n55786 , 
     n55787 , n55788 , n55789 , n55790 , n55791 , n55792 , n55793 , n55794 , n55795 , n55796 , 
     n55797 , n55798 , n55799 , n55800 , n55801 , n55802 , n55803 , n55804 , n55805 , n55806 , 
     n55807 , n55808 , n55809 , n55810 , n55811 , n55812 , n55813 , n55814 , n55815 , n55816 , 
     n55817 , n55818 , n55819 , n55820 , n55821 , n55822 , n55823 , n55824 , n55825 , n55826 , 
     n55827 , n55828 , n55829 , n55830 , n55831 , n55832 , n55833 , n55834 , n55835 , n55836 , 
     n55837 , n55838 , n55839 , n55840 , n55841 , n55842 , n55843 , n55844 , n55845 , n55846 , 
     n55847 , n55848 , n55849 , n55850 , n55851 , n55852 , n55853 , n55854 , n55855 , n55856 , 
     n55857 , n55858 , n55859 , n55860 , n55861 , n55862 , n55863 , n55864 , n55865 , n55866 , 
     n55867 , n55868 , n55869 , n55870 , n55871 , n55872 , n55873 , n55874 , n55875 , n55876 , 
     n55877 , n55878 , n55879 , n55880 , n55881 , n55882 , n55883 , n55884 , n55885 , n55886 , 
     n55887 , n55888 , n55889 , n55890 , n55891 , n55892 , n55893 , n55894 , n55895 , n55896 , 
     n55897 , n55898 , n55899 , n55900 , n55901 , n55902 , n55903 , n55904 , n55905 , n55906 , 
     n55907 , n55908 , n55909 , n55910 , n55911 , n55912 , n55913 , n55914 , n55915 , n55916 , 
     n55917 , n55918 , n55919 , n55920 , n55921 , n55922 , n55923 , n55924 , n55925 , n55926 , 
     n55927 , n55928 , n55929 , n55930 , n55931 , n55932 , n55933 , n55934 , n55935 , n55936 , 
     n55937 , n55938 , n55939 , n55940 , n55941 , n55942 , n55943 , n55944 , n55945 , n55946 , 
     n55947 , n55948 , n55949 , n55950 , n55951 , n55952 , n55953 , n55954 , n55955 , n55956 , 
     n55957 , n55958 , n55959 , n55960 , n55961 , n55962 , n55963 , n55964 , n55965 , n55966 , 
     n55967 , n55968 , n55969 , n55970 , n55971 , n55972 , n55973 , n55974 , n55975 , n55976 , 
     n55977 , n55978 , n55979 , n55980 , n55981 , n55982 , n55983 , n55984 , n55985 , n55986 , 
     n55987 , n55988 , n55989 , n55990 , n55991 , n55992 , n55993 , n55994 , n55995 , n55996 , 
     n55997 , n55998 , n55999 , n56000 , n56001 , n56002 , n56003 , n56004 , n56005 , n56006 , 
     n56007 , n56008 , n56009 , n56010 , n56011 , n56012 , n56013 , n56014 , n56015 , n56016 , 
     n56017 , n56018 , n56019 , n56020 , n56021 , n56022 , n56023 , n56024 , n56025 , n56026 , 
     n56027 , n56028 , n56029 , n56030 , n56031 , n56032 , n56033 , n56034 , n56035 , n56036 , 
     n56037 , n56038 , n56039 , n56040 , n56041 , n56042 , n56043 , n56044 , n56045 , n56046 , 
     n56047 , n56048 , n56049 , n56050 , n56051 , n56052 , n56053 , n56054 , n56055 , n56056 , 
     n56057 , n56058 , n56059 , n56060 , n56061 , n56062 , n56063 , n56064 , n56065 , n56066 , 
     n56067 , n56068 , n56069 , n56070 , n56071 , n56072 , n56073 , n56074 , n56075 , n56076 , 
     n56077 , n56078 , n56079 , n56080 , n56081 , n56082 , n56083 , n56084 , n56085 , n56086 , 
     n56087 , n56088 , n56089 , n56090 , n56091 , n56092 , n56093 , n56094 , n56095 , n56096 , 
     n56097 , n56098 , n56099 , n56100 , n56101 , n56102 , n56103 , n56104 , n56105 , n56106 , 
     n56107 , n56108 , n56109 , n56110 , n56111 , n56112 , n56113 , n56114 , n56115 , n56116 , 
     n56117 , n56118 , n56119 , n56120 , n56121 , n56122 , n56123 , n56124 , n56125 , n56126 , 
     n56127 , n56128 , n56129 , n56130 , n56131 , n56132 , n56133 , n56134 , n56135 , n56136 , 
     n56137 , n56138 , n56139 , n56140 , n56141 , n56142 , n56143 , n56144 , n56145 , n56146 , 
     n56147 , n56148 , n56149 , n56150 , n56151 , n56152 , n56153 , n56154 , n56155 , n56156 , 
     n56157 , n56158 , n56159 , n56160 , n56161 , n56162 , n56163 , n56164 , n56165 , n56166 , 
     n56167 , n56168 , n56169 , n56170 , n56171 , n56172 , n56173 , n56174 , n56175 , n56176 , 
     n56177 , n56178 , n56179 , n56180 , n56181 , n56182 , n56183 , n56184 , n56185 , n56186 , 
     n56187 , n56188 , n56189 , n56190 , n56191 , n56192 , n56193 , n56194 , n56195 , n56196 , 
     n56197 , n56198 , n56199 , n56200 , n56201 , n56202 , n56203 , n56204 , n56205 , n56206 , 
     n56207 , n56208 , n56209 , n56210 , n56211 , n56212 , n56213 , n56214 , n56215 , n56216 , 
     n56217 , n56218 , n56219 , n56220 , n56221 , n56222 , n56223 , n56224 , n56225 , n56226 , 
     n56227 , n56228 , n56229 , n56230 , n56231 , n56232 , n56233 , n56234 , n56235 , n56236 , 
     n56237 , n56238 , n56239 , n56240 , n56241 , n56242 , n56243 , n56244 , n56245 , n56246 , 
     n56247 , n56248 , n56249 , n56250 , n56251 , n56252 , n56253 , n56254 , n56255 , n56256 , 
     n56257 , n56258 , n56259 , n56260 , n56261 , n56262 , n56263 , n56264 , n56265 , n56266 , 
     n56267 , n56268 , n56269 , n56270 , n56271 , n56272 , n56273 , n56274 , n56275 , n56276 , 
     n56277 , n56278 , n56279 , n56280 , n56281 , n56282 , n56283 , n56284 , n56285 , n56286 , 
     n56287 , n56288 , n56289 , n56290 , n56291 , n56292 , n56293 , n56294 , n56295 , n56296 , 
     n56297 , n56298 , n56299 , n56300 , n56301 , n56302 , n56303 , n56304 , n56305 , n56306 , 
     n56307 , n56308 , n56309 , n56310 , n56311 , n56312 , n56313 , n56314 , n56315 , n56316 , 
     n56317 , n56318 , n56319 , n56320 , n56321 , n56322 , n56323 , n56324 , n56325 , n56326 , 
     n56327 , n56328 , n56329 , n56330 , n56331 , n56332 , n56333 , n56334 , n56335 , n56336 , 
     n56337 , n56338 , n56339 , n56340 , n56341 , n56342 , n56343 , n56344 , n56345 , n56346 , 
     n56347 , n56348 , n56349 , n56350 , n56351 , n56352 , n56353 , n56354 , n56355 , n56356 , 
     n56357 , n56358 , n56359 , n56360 , n56361 , n56362 , n56363 , n56364 , n56365 , n56366 , 
     n56367 , n56368 , n56369 , n56370 , n56371 , n56372 , n56373 , n56374 , n56375 , n56376 , 
     n56377 , n56378 , n56379 , n56380 , n56381 , n56382 , n56383 , n56384 , n56385 , n56386 , 
     n56387 , n56388 , n56389 , n56390 , n56391 , n56392 , n56393 , n56394 , n56395 , n56396 , 
     n56397 , n56398 , n56399 , n56400 , n56401 , n56402 , n56403 , n56404 , n56405 , n56406 , 
     n56407 , n56408 , n56409 , n56410 , n56411 , n56412 , n56413 , n56414 , n56415 , n56416 , 
     n56417 , n56418 , n56419 , n56420 , n56421 , n56422 , n56423 , n56424 , n56425 , n56426 , 
     n56427 , n56428 , n56429 , n56430 , n56431 , n56432 , n56433 , n56434 , n56435 , n56436 , 
     n56437 , n56438 , n56439 , n56440 , n56441 , n56442 , n56443 , n56444 , n56445 , n56446 , 
     n56447 , n56448 , n56449 , n56450 , n56451 , n56452 , n56453 , n56454 , n56455 , n56456 , 
     n56457 , n56458 , n56459 , n56460 , n56461 , n56462 , n56463 , n56464 , n56465 , n56466 , 
     n56467 , n56468 , n56469 , n56470 , n56471 , n56472 , n56473 , n56474 , n56475 , n56476 , 
     n56477 , n56478 , n56479 , n56480 , n56481 , n56482 , n56483 , n56484 , n56485 , n56486 , 
     n56487 , n56488 , n56489 , n56490 , n56491 , n56492 , n56493 , n56494 , n56495 , n56496 , 
     n56497 , n56498 , n56499 , n56500 , n56501 , n56502 , n56503 , n56504 , n56505 , n56506 , 
     n56507 , n56508 , n56509 , n56510 , n56511 , n56512 , n56513 , n56514 , n56515 , n56516 , 
     n56517 , n56518 , n56519 , n56520 , n56521 , n56522 , n56523 , n56524 , n56525 , n56526 , 
     n56527 , n56528 , n56529 , n56530 , n56531 , n56532 , n56533 , n56534 , n56535 , n56536 , 
     n56537 , n56538 , n56539 , n56540 , n56541 , n56542 , n56543 , n56544 , n56545 , n56546 , 
     n56547 , n56548 , n56549 , n56550 , n56551 , n56552 , n56553 , n56554 , n56555 , n56556 , 
     n56557 , n56558 , n56559 , n56560 , n56561 , n56562 , n56563 , n56564 , n56565 , n56566 , 
     n56567 , n56568 , n56569 , n56570 , n56571 , n56572 , n56573 , n56574 , n56575 , n56576 , 
     n56577 , n56578 , n56579 , n56580 , n56581 , n56582 , n56583 , n56584 , n56585 , n56586 , 
     n56587 , n56588 , n56589 , n56590 , n56591 , n56592 , n56593 , n56594 , n56595 , n56596 , 
     n56597 , n56598 , n56599 , n56600 , n56601 , n56602 , n56603 , n56604 , n56605 , n56606 , 
     n56607 , n56608 , n56609 , n56610 , n56611 , n56612 , n56613 , n56614 , n56615 , n56616 , 
     n56617 , n56618 , n56619 , n56620 , n56621 , n56622 , n56623 , n56624 , n56625 , n56626 , 
     n56627 , n56628 , n56629 , n56630 , n56631 , n56632 , n56633 , n56634 , n56635 , n56636 , 
     n56637 , n56638 , n56639 , n56640 , n56641 , n56642 , n56643 , n56644 , n56645 , n56646 , 
     n56647 , n56648 , n56649 , n56650 , n56651 , n56652 , n56653 , n56654 , n56655 , n56656 , 
     n56657 , n56658 , n56659 , n56660 , n56661 , n56662 , n56663 , n56664 , n56665 , n56666 , 
     n56667 , n56668 , n56669 , n56670 , n56671 , n56672 , n56673 , n56674 , n56675 , n56676 , 
     n56677 , n56678 , n56679 , n56680 , n56681 , n56682 , n56683 , n56684 , n56685 , n56686 , 
     n56687 , n56688 , n56689 , n56690 , n56691 , n56692 , n56693 , n56694 , n56695 , n56696 , 
     n56697 , n56698 , n56699 , n56700 , n56701 , n56702 , n56703 , n56704 , n56705 , n56706 , 
     n56707 , n56708 , n56709 , n56710 , n56711 , n56712 , n56713 , n56714 , n56715 , n56716 , 
     n56717 , n56718 , n56719 , n56720 , n56721 , n56722 , n56723 , n56724 , n56725 , n56726 , 
     n56727 , n56728 , n56729 , n56730 , n56731 , n56732 , n56733 , n56734 , n56735 , n56736 , 
     n56737 , n56738 , n56739 , n56740 , n56741 , n56742 , n56743 , n56744 , n56745 , n56746 , 
     n56747 , n56748 , n56749 , n56750 , n56751 , n56752 , n56753 , n56754 , n56755 , n56756 , 
     n56757 , n56758 , n56759 , n56760 , n56761 , n56762 , n56763 , n56764 , n56765 , n56766 , 
     n56767 , n56768 , n56769 , n56770 , n56771 , n56772 , n56773 , n56774 , n56775 , n56776 , 
     n56777 , n56778 , n56779 , n56780 , n56781 , n56782 , n56783 , n56784 , n56785 , n56786 , 
     n56787 , n56788 , n56789 , n56790 , n56791 , n56792 , n56793 , n56794 , n56795 , n56796 , 
     n56797 , n56798 , n56799 , n56800 , n56801 , n56802 , n56803 , n56804 , n56805 , n56806 , 
     n56807 , n56808 , n56809 , n56810 , n56811 , n56812 , n56813 , n56814 , n56815 , n56816 , 
     n56817 , n56818 , n56819 , n56820 , n56821 , n56822 , n56823 , n56824 , n56825 , n56826 , 
     n56827 , n56828 , n56829 , n56830 , n56831 , n56832 , n56833 , n56834 , n56835 , n56836 , 
     n56837 , n56838 , n56839 , n56840 , n56841 , n56842 , n56843 , n56844 , n56845 , n56846 , 
     n56847 , n56848 , n56849 , n56850 , n56851 , n56852 , n56853 , n56854 , n56855 , n56856 , 
     n56857 , n56858 , n56859 , n56860 , n56861 , n56862 , n56863 , n56864 , n56865 , n56866 , 
     n56867 , n56868 , n56869 , n56870 , n56871 , n56872 , n56873 , n56874 , n56875 , n56876 , 
     n56877 , n56878 , n56879 , n56880 , n56881 , n56882 , n56883 , n56884 , n56885 , n56886 , 
     n56887 , n56888 , n56889 , n56890 , n56891 , n56892 , n56893 , n56894 , n56895 , n56896 , 
     n56897 , n56898 , n56899 , n56900 , n56901 , n56902 , n56903 , n56904 , n56905 , n56906 , 
     n56907 , n56908 , n56909 , n56910 , n56911 , n56912 , n56913 , n56914 , n56915 , n56916 , 
     n56917 , n56918 , n56919 , n56920 , n56921 , n56922 , n56923 , n56924 , n56925 , n56926 , 
     n56927 , n56928 , n56929 , n56930 , n56931 , n56932 , n56933 , n56934 , n56935 , n56936 , 
     n56937 , n56938 , n56939 , n56940 , n56941 , n56942 , n56943 , n56944 , n56945 , n56946 , 
     n56947 , n56948 , n56949 , n56950 , n56951 , n56952 , n56953 , n56954 , n56955 , n56956 , 
     n56957 , n56958 , n56959 , n56960 , n56961 , n56962 , n56963 , n56964 , n56965 , n56966 , 
     n56967 , n56968 , n56969 , n56970 , n56971 , n56972 , n56973 , n56974 , n56975 , n56976 , 
     n56977 , n56978 , n56979 , n56980 , n56981 , n56982 , n56983 , n56984 , n56985 , n56986 , 
     n56987 , n56988 , n56989 , n56990 , n56991 , n56992 , n56993 , n56994 , n56995 , n56996 , 
     n56997 , n56998 , n56999 , n57000 , n57001 , n57002 , n57003 , n57004 , n57005 , n57006 , 
     n57007 , n57008 , n57009 , n57010 , n57011 , n57012 , n57013 , n57014 , n57015 , n57016 , 
     n57017 , n57018 , n57019 , n57020 , n57021 , n57022 , n57023 , n57024 , n57025 , n57026 , 
     n57027 , n57028 , n57029 , n57030 , n57031 , n57032 , n57033 , n57034 , n57035 , n57036 , 
     n57037 , n57038 , n57039 , n57040 , n57041 , n57042 , n57043 , n57044 , n57045 , n57046 , 
     n57047 , n57048 , n57049 , n57050 , n57051 , n57052 , n57053 , n57054 , n57055 , n57056 , 
     n57057 , n57058 , n57059 , n57060 , n57061 , n57062 , n57063 , n57064 , n57065 , n57066 , 
     n57067 , n57068 , n57069 , n57070 , n57071 , n57072 , n57073 , n57074 , n57075 , n57076 , 
     n57077 , n57078 , n57079 , n57080 , n57081 , n57082 , n57083 , n57084 , n57085 , n57086 , 
     n57087 , n57088 , n57089 , n57090 , n57091 , n57092 , n57093 , n57094 , n57095 , n57096 , 
     n57097 , n57098 , n57099 , n57100 , n57101 , n57102 , n57103 , n57104 , n57105 , n57106 , 
     n57107 , n57108 , n57109 , n57110 , n57111 , n57112 , n57113 , n57114 , n57115 , n57116 , 
     n57117 , n57118 , n57119 , n57120 , n57121 , n57122 , n57123 , n57124 , n57125 , n57126 , 
     n57127 , n57128 , n57129 , n57130 , n57131 , n57132 , n57133 , n57134 , n57135 , n57136 , 
     n57137 , n57138 , n57139 , n57140 , n57141 , n57142 , n57143 , n57144 , n57145 , n57146 , 
     n57147 , n57148 , n57149 , n57150 , n57151 , n57152 , n57153 , n57154 , n57155 , n57156 , 
     n57157 , n57158 , n57159 , n57160 , n57161 , n57162 , n57163 , n57164 , n57165 , n57166 , 
     n57167 , n57168 , n57169 , n57170 , n57171 , n57172 , n57173 , n57174 , n57175 , n57176 , 
     n57177 , n57178 , n57179 , n57180 , n57181 , n57182 , n57183 , n57184 , n57185 , n57186 , 
     n57187 , n57188 , n57189 , n57190 , n57191 , n57192 , n57193 , n57194 , n57195 , n57196 , 
     n57197 , n57198 , n57199 , n57200 , n57201 , n57202 , n57203 , n57204 , n57205 , n57206 , 
     n57207 , n57208 , n57209 , n57210 , n57211 , n57212 , n57213 , n57214 , n57215 , n57216 , 
     n57217 , n57218 , n57219 , n57220 , n57221 , n57222 , n57223 , n57224 , n57225 , n57226 , 
     n57227 , n57228 , n57229 , n57230 , n57231 , n57232 , n57233 , n57234 , n57235 , n57236 , 
     n57237 , n57238 , n57239 , n57240 , n57241 , n57242 , n57243 , n57244 , n57245 , n57246 , 
     n57247 , n57248 , n57249 , n57250 , n57251 , n57252 , n57253 , n57254 , n57255 , n57256 , 
     n57257 , n57258 , n57259 , n57260 , n57261 , n57262 , n57263 , n57264 , n57265 , n57266 , 
     n57267 , n57268 , n57269 , n57270 , n57271 , n57272 , n57273 , n57274 , n57275 , n57276 , 
     n57277 , n57278 , n57279 , n57280 , n57281 , n57282 , n57283 , n57284 , n57285 , n57286 , 
     n57287 , n57288 , n57289 , n57290 , n57291 , n57292 , n57293 , n57294 , n57295 , n57296 , 
     n57297 , n57298 , n57299 , n57300 , n57301 , n57302 , n57303 , n57304 , n57305 , n57306 , 
     n57307 , n57308 , n57309 , n57310 , n57311 , n57312 , n57313 , n57314 , n57315 , n57316 , 
     n57317 , n57318 , n57319 , n57320 , n57321 , n57322 , n57323 , n57324 , n57325 , n57326 , 
     n57327 , n57328 , n57329 , n57330 , n57331 , n57332 , n57333 , n57334 , n57335 , n57336 , 
     n57337 , n57338 , n57339 , n57340 , n57341 , n57342 , n57343 , n57344 , n57345 , n57346 , 
     n57347 , n57348 , n57349 , n57350 , n57351 , n57352 , n57353 , n57354 , n57355 , n57356 , 
     n57357 , n57358 , n57359 , n57360 , n57361 , n57362 , n57363 , n57364 , n57365 , n57366 , 
     n57367 , n57368 , n57369 , n57370 , n57371 , n57372 , n57373 , n57374 , n57375 , n57376 , 
     n57377 , n57378 , n57379 , n57380 , n57381 , n57382 , n57383 , n57384 , n57385 , n57386 , 
     n57387 , n57388 , n57389 , n57390 , n57391 , n57392 , n57393 , n57394 , n57395 , n57396 , 
     n57397 , n57398 , n57399 , n57400 , n57401 , n57402 , n57403 , n57404 , n57405 , n57406 , 
     n57407 , n57408 , n57409 , n57410 , n57411 , n57412 , n57413 , n57414 , n57415 , n57416 , 
     n57417 , n57418 , n57419 , n57420 , n57421 , n57422 , n57423 , n57424 , n57425 , n57426 , 
     n57427 , n57428 , n57429 , n57430 , n57431 , n57432 , n57433 , n57434 , n57435 , n57436 , 
     n57437 , n57438 , n57439 , n57440 , n57441 , n57442 , n57443 , n57444 , n57445 , n57446 , 
     n57447 , n57448 , n57449 , n57450 , n57451 , n57452 , n57453 , n57454 , n57455 , n57456 , 
     n57457 , n57458 , n57459 , n57460 , n57461 , n57462 , n57463 , n57464 , n57465 , n57466 , 
     n57467 , n57468 , n57469 , n57470 , n57471 , n57472 , n57473 , n57474 , n57475 , n57476 , 
     n57477 , n57478 , n57479 , n57480 , n57481 , n57482 , n57483 , n57484 , n57485 , n57486 , 
     n57487 , n57488 , n57489 , n57490 , n57491 , n57492 , n57493 , n57494 , n57495 , n57496 , 
     n57497 , n57498 , n57499 , n57500 , n57501 , n57502 , n57503 , n57504 , n57505 , n57506 , 
     n57507 , n57508 , n57509 , n57510 , n57511 , n57512 , n57513 , n57514 , n57515 , n57516 , 
     n57517 , n57518 , n57519 , n57520 , n57521 , n57522 , n57523 , n57524 , n57525 , n57526 , 
     n57527 , n57528 , n57529 , n57530 , n57531 , n57532 , n57533 , n57534 , n57535 , n57536 , 
     n57537 , n57538 , n57539 , n57540 , n57541 , n57542 , n57543 , n57544 , n57545 , n57546 , 
     n57547 , n57548 , n57549 , n57550 , n57551 , n57552 , n57553 , n57554 , n57555 , n57556 , 
     n57557 , n57558 , n57559 , n57560 , n57561 , n57562 , n57563 , n57564 , n57565 , n57566 , 
     n57567 , n57568 , n57569 , n57570 , n57571 , n57572 , n57573 , n57574 , n57575 , n57576 , 
     n57577 , n57578 , n57579 , n57580 , n57581 , n57582 , n57583 , n57584 , n57585 , n57586 , 
     n57587 , n57588 , n57589 , n57590 , n57591 , n57592 , n57593 , n57594 , n57595 , n57596 , 
     n57597 , n57598 , n57599 , n57600 , n57601 , n57602 , n57603 , n57604 , n57605 , n57606 , 
     n57607 , n57608 , n57609 , n57610 , n57611 , n57612 , n57613 , n57614 , n57615 , n57616 , 
     n57617 , n57618 , n57619 , n57620 , n57621 , n57622 , n57623 , n57624 , n57625 , n57626 , 
     n57627 , n57628 , n57629 , n57630 , n57631 , n57632 , n57633 , n57634 , n57635 , n57636 , 
     n57637 , n57638 , n57639 , n57640 , n57641 , n57642 , n57643 , n57644 , n57645 , n57646 , 
     n57647 , n57648 , n57649 , n57650 , n57651 , n57652 , n57653 , n57654 , n57655 , n57656 , 
     n57657 , n57658 , n57659 , n57660 , n57661 , n57662 , n57663 , n57664 , n57665 , n57666 , 
     n57667 , n57668 , n57669 , n57670 , n57671 , n57672 , n57673 , n57674 , n57675 , n57676 , 
     n57677 , n57678 , n57679 , n57680 , n57681 , n57682 , n57683 , n57684 , n57685 , n57686 , 
     n57687 , n57688 , n57689 , n57690 , n57691 , n57692 , n57693 , n57694 , n57695 , n57696 , 
     n57697 , n57698 , n57699 , n57700 , n57701 , n57702 , n57703 , n57704 , n57705 , n57706 , 
     n57707 , n57708 , n57709 , n57710 , n57711 , n57712 , n57713 , n57714 , n57715 , n57716 , 
     n57717 , n57718 , n57719 , n57720 , n57721 , n57722 , n57723 , n57724 , n57725 , n57726 , 
     n57727 , n57728 , n57729 , n57730 , n57731 , n57732 , n57733 , n57734 , n57735 , n57736 , 
     n57737 , n57738 , n57739 , n57740 , n57741 , n57742 , n57743 , n57744 , n57745 , n57746 , 
     n57747 , n57748 , n57749 , n57750 , n57751 , n57752 , n57753 , n57754 , n57755 , n57756 , 
     n57757 , n57758 , n57759 , n57760 , n57761 , n57762 , n57763 , n57764 , n57765 , n57766 , 
     n57767 , n57768 , n57769 , n57770 , n57771 , n57772 , n57773 , n57774 , n57775 , n57776 , 
     n57777 , n57778 , n57779 , n57780 , n57781 , n57782 , n57783 , n57784 , n57785 , n57786 , 
     n57787 , n57788 , n57789 , n57790 , n57791 , n57792 , n57793 , n57794 , n57795 , n57796 , 
     n57797 , n57798 , n57799 , n57800 , n57801 , n57802 , n57803 , n57804 , n57805 , n57806 , 
     n57807 , n57808 , n57809 , n57810 , n57811 , n57812 , n57813 , n57814 , n57815 , n57816 , 
     n57817 , n57818 , n57819 , n57820 , n57821 , n57822 , n57823 , n57824 , n57825 , n57826 , 
     n57827 , n57828 , n57829 , n57830 , n57831 , n57832 , n57833 , n57834 , n57835 , n57836 , 
     n57837 , n57838 , n57839 , n57840 , n57841 , n57842 , n57843 , n57844 , n57845 , n57846 , 
     n57847 , n57848 , n57849 , n57850 , n57851 , n57852 , n57853 , n57854 , n57855 , n57856 , 
     n57857 , n57858 , n57859 , n57860 , n57861 , n57862 , n57863 , n57864 , n57865 , n57866 , 
     n57867 , n57868 , n57869 , n57870 , n57871 , n57872 , n57873 , n57874 , n57875 , n57876 , 
     n57877 , n57878 , n57879 , n57880 , n57881 , n57882 , n57883 , n57884 , n57885 , n57886 , 
     n57887 , n57888 , n57889 , n57890 , n57891 , n57892 , n57893 , n57894 , n57895 , n57896 , 
     n57897 , n57898 , n57899 , n57900 , n57901 , n57902 , n57903 , n57904 , n57905 , n57906 , 
     n57907 , n57908 , n57909 , n57910 , n57911 , n57912 , n57913 , n57914 , n57915 , n57916 , 
     n57917 , n57918 , n57919 , n57920 , n57921 , n57922 , n57923 , n57924 , n57925 , n57926 , 
     n57927 , n57928 , n57929 , n57930 , n57931 , n57932 , n57933 , n57934 , n57935 , n57936 , 
     n57937 , n57938 , n57939 , n57940 , n57941 , n57942 , n57943 , n57944 , n57945 , n57946 , 
     n57947 , n57948 , n57949 , n57950 , n57951 , n57952 , n57953 , n57954 , n57955 , n57956 , 
     n57957 , n57958 , n57959 , n57960 , n57961 , n57962 , n57963 , n57964 , n57965 , n57966 , 
     n57967 , n57968 , n57969 , n57970 , n57971 , n57972 , n57973 , n57974 , n57975 , n57976 , 
     n57977 , n57978 , n57979 , n57980 , n57981 , n57982 , n57983 , n57984 , n57985 , n57986 , 
     n57987 , n57988 , n57989 , n57990 , n57991 , n57992 , n57993 , n57994 , n57995 , n57996 , 
     n57997 , n57998 , n57999 , n58000 , n58001 , n58002 , n58003 , n58004 , n58005 , n58006 , 
     n58007 , n58008 , n58009 , n58010 , n58011 , n58012 , n58013 , n58014 , n58015 , n58016 , 
     n58017 , n58018 , n58019 , n58020 , n58021 , n58022 , n58023 , n58024 , n58025 , n58026 , 
     n58027 , n58028 , n58029 , n58030 , n58031 , n58032 , n58033 , n58034 , n58035 , n58036 , 
     n58037 , n58038 , n58039 , n58040 , n58041 , n58042 , n58043 , n58044 , n58045 , n58046 , 
     n58047 , n58048 , n58049 , n58050 , n58051 , n58052 , n58053 , n58054 , n58055 , n58056 , 
     n58057 , n58058 , n58059 , n58060 , n58061 , n58062 , n58063 , n58064 , n58065 , n58066 , 
     n58067 , n58068 , n58069 , n58070 , n58071 , n58072 , n58073 , n58074 , n58075 , n58076 , 
     n58077 , n58078 , n58079 , n58080 , n58081 , n58082 , n58083 , n58084 , n58085 , n58086 , 
     n58087 , n58088 , n58089 , n58090 , n58091 , n58092 , n58093 , n58094 , n58095 , n58096 , 
     n58097 , n58098 , n58099 , n58100 , n58101 , n58102 , n58103 , n58104 , n58105 , n58106 , 
     n58107 , n58108 , n58109 , n58110 , n58111 , n58112 , n58113 , n58114 , n58115 , n58116 , 
     n58117 , n58118 , n58119 , n58120 , n58121 , n58122 , n58123 , n58124 , n58125 , n58126 , 
     n58127 , n58128 , n58129 , n58130 , n58131 , n58132 , n58133 , n58134 , n58135 , n58136 , 
     n58137 , n58138 , n58139 , n58140 , n58141 , n58142 , n58143 , n58144 , n58145 , n58146 , 
     n58147 , n58148 , n58149 , n58150 , n58151 , n58152 , n58153 , n58154 , n58155 , n58156 , 
     n58157 , n58158 , n58159 , n58160 , n58161 , n58162 , n58163 , n58164 , n58165 , n58166 , 
     n58167 , n58168 , n58169 , n58170 , n58171 , n58172 , n58173 , n58174 , n58175 , n58176 , 
     n58177 , n58178 , n58179 , n58180 , n58181 , n58182 , n58183 , n58184 , n58185 , n58186 , 
     n58187 , n58188 , n58189 , n58190 , n58191 , n58192 , n58193 , n58194 , n58195 , n58196 , 
     n58197 , n58198 , n58199 , n58200 , n58201 , n58202 , n58203 , n58204 , n58205 , n58206 , 
     n58207 , n58208 , n58209 , n58210 , n58211 , n58212 , n58213 , n58214 , n58215 , n58216 , 
     n58217 , n58218 , n58219 , n58220 , n58221 , n58222 , n58223 , n58224 , n58225 , n58226 , 
     n58227 , n58228 , n58229 , n58230 , n58231 , n58232 , n58233 , n58234 , n58235 , n58236 , 
     n58237 , n58238 , n58239 , n58240 , n58241 , n58242 , n58243 , n58244 , n58245 , n58246 , 
     n58247 , n58248 , n58249 , n58250 , n58251 , n58252 , n58253 , n58254 , n58255 , n58256 , 
     n58257 , n58258 , n58259 , n58260 , n58261 , n58262 , n58263 , n58264 , n58265 , n58266 , 
     n58267 , n58268 , n58269 , n58270 , n58271 , n58272 , n58273 , n58274 , n58275 , n58276 , 
     n58277 , n58278 , n58279 , n58280 , n58281 , n58282 , n58283 , n58284 , n58285 , n58286 , 
     n58287 , n58288 , n58289 , n58290 , n58291 , n58292 , n58293 , n58294 , n58295 , n58296 , 
     n58297 , n58298 , n58299 , n58300 , n58301 , n58302 , n58303 , n58304 , n58305 , n58306 , 
     n58307 , n58308 , n58309 , n58310 , n58311 , n58312 , n58313 , n58314 , n58315 , n58316 , 
     n58317 , n58318 , n58319 , n58320 , n58321 , n58322 , n58323 , n58324 , n58325 , n58326 , 
     n58327 , n58328 , n58329 , n58330 , n58331 , n58332 , n58333 , n58334 , n58335 , n58336 , 
     n58337 , n58338 , n58339 , n58340 , n58341 , n58342 , n58343 , n58344 , n58345 , n58346 , 
     n58347 , n58348 , n58349 , n58350 , n58351 , n58352 , n58353 , n58354 , n58355 , n58356 , 
     n58357 , n58358 , n58359 , n58360 , n58361 , n58362 , n58363 , n58364 , n58365 , n58366 , 
     n58367 , n58368 , n58369 , n58370 , n58371 , n58372 , n58373 , n58374 , n58375 , n58376 , 
     n58377 , n58378 , n58379 , n58380 , n58381 , n58382 , n58383 , n58384 , n58385 , n58386 , 
     n58387 , n58388 , n58389 , n58390 , n58391 , n58392 , n58393 , n58394 , n58395 , n58396 , 
     n58397 , n58398 , n58399 , n58400 , n58401 , n58402 , n58403 , n58404 , n58405 , n58406 , 
     n58407 , n58408 , n58409 , n58410 , n58411 , n58412 , n58413 , n58414 , n58415 , n58416 , 
     n58417 , n58418 , n58419 , n58420 , n58421 , n58422 , n58423 , n58424 , n58425 , n58426 , 
     n58427 , n58428 , n58429 , n58430 , n58431 , n58432 , n58433 , n58434 , n58435 , n58436 , 
     n58437 , n58438 , n58439 , n58440 , n58441 , n58442 , n58443 , n58444 , n58445 , n58446 , 
     n58447 , n58448 , n58449 , n58450 , n58451 , n58452 , n58453 , n58454 , n58455 , n58456 , 
     n58457 , n58458 , n58459 , n58460 , n58461 , n58462 , n58463 , n58464 , n58465 , n58466 , 
     n58467 , n58468 , n58469 , n58470 , n58471 , n58472 , n58473 , n58474 , n58475 , n58476 , 
     n58477 , n58478 , n58479 , n58480 , n58481 , n58482 , n58483 , n58484 , n58485 , n58486 , 
     n58487 , n58488 , n58489 , n58490 , n58491 , n58492 , n58493 , n58494 , n58495 , n58496 , 
     n58497 , n58498 , n58499 , n58500 , n58501 , n58502 , n58503 , n58504 , n58505 , n58506 , 
     n58507 , n58508 , n58509 , n58510 , n58511 , n58512 , n58513 , n58514 , n58515 , n58516 , 
     n58517 , n58518 , n58519 , n58520 , n58521 , n58522 , n58523 , n58524 , n58525 , n58526 , 
     n58527 , n58528 , n58529 , n58530 , n58531 , n58532 , n58533 , n58534 , n58535 , n58536 , 
     n58537 , n58538 , n58539 , n58540 , n58541 , n58542 , n58543 , n58544 , n58545 , n58546 , 
     n58547 , n58548 , n58549 , n58550 , n58551 , n58552 , n58553 , n58554 , n58555 , n58556 , 
     n58557 , n58558 , n58559 , n58560 , n58561 , n58562 , n58563 , n58564 , n58565 , n58566 , 
     n58567 , n58568 , n58569 , n58570 , n58571 , n58572 , n58573 , n58574 , n58575 , n58576 , 
     n58577 , n58578 , n58579 , n58580 , n58581 , n58582 , n58583 , n58584 , n58585 , n58586 , 
     n58587 , n58588 , n58589 , n58590 , n58591 , n58592 , n58593 , n58594 , n58595 , n58596 , 
     n58597 , n58598 , n58599 , n58600 , n58601 , n58602 , n58603 , n58604 , n58605 , n58606 , 
     n58607 , n58608 , n58609 , n58610 , n58611 , n58612 , n58613 , n58614 , n58615 , n58616 , 
     n58617 , n58618 , n58619 , n58620 , n58621 , n58622 , n58623 , n58624 , n58625 , n58626 , 
     n58627 , n58628 , n58629 , n58630 , n58631 , n58632 , n58633 , n58634 , n58635 , n58636 , 
     n58637 , n58638 , n58639 , n58640 , n58641 , n58642 , n58643 , n58644 , n58645 , n58646 , 
     n58647 , n58648 , n58649 , n58650 , n58651 , n58652 , n58653 , n58654 , n58655 , n58656 , 
     n58657 , n58658 , n58659 , n58660 , n58661 , n58662 , n58663 , n58664 , n58665 , n58666 , 
     n58667 , n58668 , n58669 , n58670 , n58671 , n58672 , n58673 , n58674 , n58675 , n58676 , 
     n58677 , n58678 , n58679 , n58680 , n58681 , n58682 , n58683 , n58684 , n58685 , n58686 , 
     n58687 , n58688 , n58689 , n58690 , n58691 , n58692 , n58693 , n58694 , n58695 , n58696 , 
     n58697 , n58698 , n58699 , n58700 , n58701 , n58702 , n58703 , n58704 , n58705 , n58706 , 
     n58707 , n58708 , n58709 , n58710 , n58711 , n58712 , n58713 , n58714 , n58715 , n58716 , 
     n58717 , n58718 , n58719 , n58720 , n58721 , n58722 , n58723 , n58724 , n58725 , n58726 , 
     n58727 , n58728 , n58729 , n58730 , n58731 , n58732 , n58733 , n58734 , n58735 , n58736 , 
     n58737 , n58738 , n58739 , n58740 , n58741 , n58742 , n58743 , n58744 , n58745 , n58746 , 
     n58747 , n58748 , n58749 , n58750 , n58751 , n58752 , n58753 , n58754 , n58755 , n58756 , 
     n58757 , n58758 , n58759 , n58760 , n58761 , n58762 , n58763 , n58764 , n58765 , n58766 , 
     n58767 , n58768 , n58769 , n58770 , n58771 , n58772 , n58773 , n58774 , n58775 , n58776 , 
     n58777 , n58778 , n58779 , n58780 , n58781 , n58782 , n58783 , n58784 , n58785 , n58786 , 
     n58787 , n58788 , n58789 , n58790 , n58791 , n58792 , n58793 , n58794 , n58795 , n58796 , 
     n58797 , n58798 , n58799 , n58800 , n58801 , n58802 , n58803 , n58804 , n58805 , n58806 , 
     n58807 , n58808 , n58809 , n58810 , n58811 , n58812 , n58813 , n58814 , n58815 , n58816 , 
     n58817 , n58818 , n58819 , n58820 , n58821 , n58822 , n58823 , n58824 , n58825 , n58826 , 
     n58827 , n58828 , n58829 , n58830 , n58831 , n58832 , n58833 , n58834 , n58835 , n58836 , 
     n58837 , n58838 , n58839 , n58840 , n58841 , n58842 , n58843 , n58844 , n58845 , n58846 , 
     n58847 , n58848 , n58849 , n58850 , n58851 , n58852 , n58853 , n58854 , n58855 , n58856 , 
     n58857 , n58858 , n58859 , n58860 , n58861 , n58862 , n58863 , n58864 , n58865 , n58866 , 
     n58867 , n58868 , n58869 , n58870 , n58871 , n58872 , n58873 , n58874 , n58875 , n58876 , 
     n58877 , n58878 , n58879 , n58880 , n58881 , n58882 , n58883 , n58884 , n58885 , n58886 , 
     n58887 , n58888 , n58889 , n58890 , n58891 , n58892 , n58893 , n58894 , n58895 , n58896 , 
     n58897 , n58898 , n58899 , n58900 , n58901 , n58902 , n58903 , n58904 , n58905 , n58906 , 
     n58907 , n58908 , n58909 , n58910 , n58911 , n58912 , n58913 , n58914 , n58915 , n58916 , 
     n58917 , n58918 , n58919 , n58920 , n58921 , n58922 , n58923 , n58924 , n58925 , n58926 , 
     n58927 , n58928 , n58929 , n58930 , n58931 , n58932 , n58933 , n58934 , n58935 , n58936 , 
     n58937 , n58938 , n58939 , n58940 , n58941 , n58942 , n58943 , n58944 , n58945 , n58946 , 
     n58947 , n58948 , n58949 , n58950 , n58951 , n58952 , n58953 , n58954 , n58955 , n58956 , 
     n58957 , n58958 , n58959 , n58960 , n58961 , n58962 , n58963 , n58964 , n58965 , n58966 , 
     n58967 , n58968 , n58969 , n58970 , n58971 , n58972 , n58973 , n58974 , n58975 , n58976 , 
     n58977 , n58978 , n58979 , n58980 , n58981 , n58982 , n58983 , n58984 , n58985 , n58986 , 
     n58987 , n58988 , n58989 , n58990 , n58991 , n58992 , n58993 , n58994 , n58995 , n58996 , 
     n58997 , n58998 , n58999 , n59000 , n59001 , n59002 , n59003 , n59004 , n59005 , n59006 , 
     n59007 , n59008 , n59009 , n59010 , n59011 , n59012 , n59013 , n59014 , n59015 , n59016 , 
     n59017 , n59018 , n59019 , n59020 , n59021 , n59022 , n59023 , n59024 , n59025 , n59026 , 
     n59027 , n59028 , n59029 , n59030 , n59031 , n59032 , n59033 , n59034 , n59035 , n59036 , 
     n59037 , n59038 , n59039 , n59040 , n59041 , n59042 , n59043 , n59044 , n59045 , n59046 , 
     n59047 , n59048 , n59049 , n59050 , n59051 , n59052 , n59053 , n59054 , n59055 , n59056 , 
     n59057 , n59058 , n59059 , n59060 , n59061 , n59062 , n59063 , n59064 , n59065 , n59066 , 
     n59067 , n59068 , n59069 , n59070 , n59071 , n59072 , n59073 , n59074 , n59075 , n59076 , 
     n59077 , n59078 , n59079 , n59080 , n59081 , n59082 , n59083 , n59084 , n59085 , n59086 , 
     n59087 , n59088 , n59089 , n59090 , n59091 , n59092 , n59093 , n59094 , n59095 , n59096 , 
     n59097 , n59098 , n59099 , n59100 , n59101 , n59102 , n59103 , n59104 , n59105 , n59106 , 
     n59107 , n59108 , n59109 , n59110 , n59111 , n59112 , n59113 , n59114 , n59115 , n59116 , 
     n59117 , n59118 , n59119 , n59120 , n59121 , n59122 , n59123 , n59124 , n59125 , n59126 , 
     n59127 , n59128 , n59129 , n59130 , n59131 , n59132 , n59133 , n59134 , n59135 , n59136 , 
     n59137 , n59138 , n59139 , n59140 , n59141 , n59142 , n59143 , n59144 , n59145 , n59146 , 
     n59147 , n59148 , n59149 , n59150 , n59151 , n59152 , n59153 , n59154 , n59155 , n59156 , 
     n59157 , n59158 , n59159 , n59160 , n59161 , n59162 , n59163 , n59164 , n59165 , n59166 , 
     n59167 , n59168 , n59169 , n59170 , n59171 , n59172 , n59173 , n59174 , n59175 , n59176 , 
     n59177 , n59178 , n59179 , n59180 , n59181 , n59182 , n59183 , n59184 , n59185 , n59186 , 
     n59187 , n59188 , n59189 , n59190 , n59191 , n59192 , n59193 , n59194 , n59195 , n59196 , 
     n59197 , n59198 , n59199 , n59200 , n59201 , n59202 , n59203 , n59204 , n59205 , n59206 , 
     n59207 , n59208 , n59209 , n59210 , n59211 , n59212 , n59213 , n59214 , n59215 , n59216 , 
     n59217 , n59218 , n59219 , n59220 , n59221 , n59222 , n59223 , n59224 , n59225 , n59226 , 
     n59227 , n59228 , n59229 , n59230 , n59231 , n59232 , n59233 , n59234 , n59235 , n59236 , 
     n59237 , n59238 , n59239 , n59240 , n59241 , n59242 , n59243 , n59244 , n59245 , n59246 , 
     n59247 , n59248 , n59249 , n59250 , n59251 , n59252 , n59253 , n59254 , n59255 , n59256 , 
     n59257 , n59258 , n59259 , n59260 , n59261 , n59262 , n59263 , n59264 , n59265 , n59266 , 
     n59267 , n59268 , n59269 , n59270 , n59271 , n59272 , n59273 , n59274 , n59275 , n59276 , 
     n59277 , n59278 , n59279 , n59280 , n59281 , n59282 , n59283 , n59284 , n59285 , n59286 , 
     n59287 , n59288 , n59289 , n59290 , n59291 , n59292 , n59293 , n59294 , n59295 , n59296 , 
     n59297 , n59298 , n59299 , n59300 , n59301 , n59302 , n59303 , n59304 , n59305 , n59306 , 
     n59307 , n59308 , n59309 , n59310 , n59311 , n59312 , n59313 , n59314 , n59315 , n59316 , 
     n59317 , n59318 , n59319 , n59320 , n59321 , n59322 , n59323 , n59324 , n59325 , n59326 , 
     n59327 , n59328 , n59329 , n59330 , n59331 , n59332 , n59333 , n59334 , n59335 , n59336 , 
     n59337 , n59338 , n59339 , n59340 , n59341 , n59342 , n59343 , n59344 , n59345 , n59346 , 
     n59347 , n59348 , n59349 , n59350 , n59351 , n59352 , n59353 , n59354 , n59355 , n59356 , 
     n59357 , n59358 , n59359 , n59360 , n59361 , n59362 , n59363 , n59364 , n59365 , n59366 , 
     n59367 , n59368 , n59369 , n59370 , n59371 , n59372 , n59373 , n59374 , n59375 , n59376 , 
     n59377 , n59378 , n59379 , n59380 , n59381 , n59382 , n59383 , n59384 , n59385 , n59386 , 
     n59387 , n59388 , n59389 , n59390 , n59391 , n59392 , n59393 , n59394 , n59395 , n59396 , 
     n59397 , n59398 , n59399 , n59400 , n59401 , n59402 , n59403 , n59404 , n59405 , n59406 , 
     n59407 , n59408 , n59409 , n59410 , n59411 , n59412 , n59413 , n59414 , n59415 , n59416 , 
     n59417 , n59418 , n59419 , n59420 , n59421 , n59422 , n59423 , n59424 , n59425 , n59426 , 
     n59427 , n59428 , n59429 , n59430 , n59431 , n59432 , n59433 , n59434 , n59435 , n59436 , 
     n59437 , n59438 , n59439 , n59440 , n59441 , n59442 , n59443 , n59444 , n59445 , n59446 , 
     n59447 , n59448 , n59449 , n59450 , n59451 , n59452 , n59453 , n59454 , n59455 , n59456 , 
     n59457 , n59458 , n59459 , n59460 , n59461 , n59462 , n59463 , n59464 , n59465 , n59466 , 
     n59467 , n59468 , n59469 , n59470 , n59471 , n59472 , n59473 , n59474 , n59475 , n59476 , 
     n59477 , n59478 , n59479 , n59480 , n59481 , n59482 , n59483 , n59484 , n59485 , n59486 , 
     n59487 , n59488 , n59489 , n59490 , n59491 , n59492 , n59493 , n59494 , n59495 , n59496 , 
     n59497 , n59498 , n59499 , n59500 , n59501 , n59502 , n59503 , n59504 , n59505 , n59506 , 
     n59507 , n59508 , n59509 , n59510 , n59511 , n59512 , n59513 , n59514 , n59515 , n59516 , 
     n59517 , n59518 , n59519 , n59520 , n59521 , n59522 , n59523 , n59524 , n59525 , n59526 , 
     n59527 , n59528 , n59529 , n59530 , n59531 , n59532 , n59533 , n59534 , n59535 , n59536 , 
     n59537 , n59538 , n59539 , n59540 , n59541 , n59542 , n59543 , n59544 , n59545 , n59546 , 
     n59547 , n59548 , n59549 , n59550 , n59551 , n59552 , n59553 , n59554 , n59555 , n59556 , 
     n59557 , n59558 , n59559 , n59560 , n59561 , n59562 , n59563 , n59564 , n59565 , n59566 , 
     n59567 , n59568 , n59569 , n59570 , n59571 , n59572 , n59573 , n59574 , n59575 , n59576 , 
     n59577 , n59578 , n59579 , n59580 , n59581 , n59582 , n59583 , n59584 , n59585 , n59586 , 
     n59587 , n59588 , n59589 , n59590 , n59591 , n59592 , n59593 , n59594 , n59595 , n59596 , 
     n59597 , n59598 , n59599 , n59600 , n59601 , n59602 , n59603 , n59604 , n59605 , n59606 , 
     n59607 , n59608 , n59609 , n59610 , n59611 , n59612 , n59613 , n59614 , n59615 , n59616 , 
     n59617 , n59618 , n59619 , n59620 , n59621 , n59622 , n59623 , n59624 , n59625 , n59626 , 
     n59627 , n59628 , n59629 , n59630 , n59631 , n59632 , n59633 , n59634 , n59635 , n59636 , 
     n59637 , n59638 , n59639 , n59640 , n59641 , n59642 , n59643 , n59644 , n59645 , n59646 , 
     n59647 , n59648 , n59649 , n59650 , n59651 , n59652 , n59653 , n59654 , n59655 , n59656 , 
     n59657 , n59658 , n59659 , n59660 , n59661 , n59662 , n59663 , n59664 , n59665 , n59666 , 
     n59667 , n59668 , n59669 , n59670 , n59671 , n59672 , n59673 , n59674 , n59675 , n59676 , 
     n59677 , n59678 , n59679 , n59680 , n59681 , n59682 , n59683 , n59684 , n59685 , n59686 , 
     n59687 , n59688 , n59689 , n59690 , n59691 , n59692 , n59693 , n59694 , n59695 , n59696 , 
     n59697 , n59698 , n59699 , n59700 , n59701 , n59702 , n59703 , n59704 , n59705 , n59706 , 
     n59707 , n59708 , n59709 , n59710 , n59711 , n59712 , n59713 , n59714 , n59715 , n59716 , 
     n59717 , n59718 , n59719 , n59720 , n59721 , n59722 , n59723 , n59724 , n59725 , n59726 , 
     n59727 , n59728 , n59729 , n59730 , n59731 , n59732 , n59733 , n59734 , n59735 , n59736 , 
     n59737 , n59738 , n59739 , n59740 , n59741 , n59742 , n59743 , n59744 , n59745 , n59746 , 
     n59747 , n59748 , n59749 , n59750 , n59751 , n59752 , n59753 , n59754 , n59755 , n59756 , 
     n59757 , n59758 , n59759 , n59760 , n59761 , n59762 , n59763 , n59764 , n59765 , n59766 , 
     n59767 , n59768 , n59769 , n59770 , n59771 , n59772 , n59773 , n59774 , n59775 , n59776 , 
     n59777 , n59778 , n59779 , n59780 , n59781 , n59782 , n59783 , n59784 , n59785 , n59786 , 
     n59787 , n59788 , n59789 , n59790 , n59791 , n59792 , n59793 , n59794 , n59795 , n59796 , 
     n59797 , n59798 , n59799 , n59800 , n59801 , n59802 , n59803 , n59804 , n59805 , n59806 , 
     n59807 , n59808 , n59809 , n59810 , n59811 , n59812 , n59813 , n59814 , n59815 , n59816 , 
     n59817 , n59818 , n59819 , n59820 , n59821 , n59822 , n59823 , n59824 , n59825 , n59826 , 
     n59827 , n59828 , n59829 , n59830 , n59831 , n59832 , n59833 , n59834 , n59835 , n59836 , 
     n59837 , n59838 , n59839 , n59840 , n59841 , n59842 , n59843 , n59844 , n59845 , n59846 , 
     n59847 , n59848 , n59849 , n59850 , n59851 , n59852 , n59853 , n59854 , n59855 , n59856 , 
     n59857 , n59858 , n59859 , n59860 , n59861 , n59862 , n59863 , n59864 , n59865 , n59866 , 
     n59867 , n59868 , n59869 , n59870 , n59871 , n59872 , n59873 , n59874 , n59875 , n59876 , 
     n59877 , n59878 , n59879 , n59880 , n59881 , n59882 , n59883 , n59884 , n59885 , n59886 , 
     n59887 , n59888 , n59889 , n59890 , n59891 , n59892 , n59893 , n59894 , n59895 , n59896 , 
     n59897 , n59898 , n59899 , n59900 , n59901 , n59902 , n59903 , n59904 , n59905 , n59906 , 
     n59907 , n59908 , n59909 , n59910 , n59911 , n59912 , n59913 , n59914 , n59915 , n59916 , 
     n59917 , n59918 , n59919 , n59920 , n59921 , n59922 , n59923 , n59924 , n59925 , n59926 , 
     n59927 , n59928 , n59929 , n59930 , n59931 , n59932 , n59933 , n59934 , n59935 , n59936 , 
     n59937 , n59938 , n59939 , n59940 , n59941 , n59942 , n59943 , n59944 , n59945 , n59946 , 
     n59947 , n59948 , n59949 , n59950 , n59951 , n59952 , n59953 , n59954 , n59955 , n59956 , 
     n59957 , n59958 , n59959 , n59960 , n59961 , n59962 , n59963 , n59964 , n59965 , n59966 , 
     n59967 , n59968 , n59969 , n59970 , n59971 , n59972 , n59973 , n59974 , n59975 , n59976 , 
     n59977 , n59978 , n59979 , n59980 , n59981 , n59982 , n59983 , n59984 , n59985 , n59986 , 
     n59987 , n59988 , n59989 , n59990 , n59991 , n59992 , n59993 , n59994 , n59995 , n59996 , 
     n59997 , n59998 , n59999 , n60000 , n60001 , n60002 , n60003 , n60004 , n60005 , n60006 , 
     n60007 , n60008 , n60009 , n60010 , n60011 , n60012 , n60013 , n60014 , n60015 , n60016 , 
     n60017 , n60018 , n60019 , n60020 , n60021 , n60022 , n60023 , n60024 , n60025 , n60026 , 
     n60027 , n60028 , n60029 , n60030 , n60031 , n60032 , n60033 , n60034 , n60035 , n60036 , 
     n60037 , n60038 , n60039 , n60040 , n60041 , n60042 , n60043 , n60044 , n60045 , n60046 , 
     n60047 , n60048 , n60049 , n60050 , n60051 , n60052 , n60053 , n60054 , n60055 , n60056 , 
     n60057 , n60058 , n60059 , n60060 , n60061 , n60062 , n60063 , n60064 , n60065 , n60066 , 
     n60067 , n60068 , n60069 , n60070 , n60071 , n60072 , n60073 , n60074 , n60075 , n60076 , 
     n60077 , n60078 , n60079 , n60080 , n60081 , n60082 , n60083 , n60084 , n60085 , n60086 , 
     n60087 , n60088 , n60089 , n60090 , n60091 , n60092 , n60093 , n60094 , n60095 , n60096 , 
     n60097 , n60098 , n60099 , n60100 , n60101 , n60102 , n60103 , n60104 , n60105 , n60106 , 
     n60107 , n60108 , n60109 , n60110 , n60111 , n60112 , n60113 , n60114 , n60115 , n60116 , 
     n60117 , n60118 , n60119 , n60120 , n60121 , n60122 , n60123 , n60124 , n60125 , n60126 , 
     n60127 , n60128 , n60129 , n60130 , n60131 , n60132 , n60133 , n60134 , n60135 , n60136 , 
     n60137 , n60138 , n60139 , n60140 , n60141 , n60142 , n60143 , n60144 , n60145 , n60146 , 
     n60147 , n60148 , n60149 , n60150 , n60151 , n60152 , n60153 , n60154 , n60155 , n60156 , 
     n60157 , n60158 , n60159 , n60160 , n60161 , n60162 , n60163 , n60164 , n60165 , n60166 , 
     n60167 , n60168 , n60169 , n60170 , n60171 , n60172 , n60173 , n60174 , n60175 , n60176 , 
     n60177 , n60178 , n60179 , n60180 , n60181 , n60182 , n60183 , n60184 , n60185 , n60186 , 
     n60187 , n60188 , n60189 , n60190 , n60191 , n60192 , n60193 , n60194 , n60195 , n60196 , 
     n60197 , n60198 , n60199 , n60200 , n60201 , n60202 , n60203 , n60204 , n60205 , n60206 , 
     n60207 , n60208 , n60209 , n60210 , n60211 , n60212 , n60213 , n60214 , n60215 , n60216 , 
     n60217 , n60218 , n60219 , n60220 , n60221 , n60222 , n60223 , n60224 , n60225 , n60226 , 
     n60227 , n60228 , n60229 , n60230 , n60231 , n60232 , n60233 , n60234 , n60235 , n60236 , 
     n60237 , n60238 , n60239 , n60240 , n60241 , n60242 , n60243 , n60244 , n60245 , n60246 , 
     n60247 , n60248 , n60249 , n60250 , n60251 , n60252 , n60253 , n60254 , n60255 , n60256 , 
     n60257 , n60258 , n60259 , n60260 , n60261 , n60262 , n60263 , n60264 , n60265 , n60266 , 
     n60267 , n60268 , n60269 , n60270 , n60271 , n60272 , n60273 , n60274 , n60275 , n60276 , 
     n60277 , n60278 , n60279 , n60280 , n60281 , n60282 , n60283 , n60284 , n60285 , n60286 , 
     n60287 , n60288 , n60289 , n60290 , n60291 , n60292 , n60293 , n60294 , n60295 , n60296 , 
     n60297 , n60298 , n60299 , n60300 , n60301 , n60302 , n60303 , n60304 , n60305 , n60306 , 
     n60307 , n60308 , n60309 , n60310 , n60311 , n60312 , n60313 , n60314 , n60315 , n60316 , 
     n60317 , n60318 , n60319 , n60320 , n60321 , n60322 , n60323 , n60324 , n60325 , n60326 , 
     n60327 , n60328 , n60329 , n60330 , n60331 , n60332 , n60333 , n60334 , n60335 , n60336 , 
     n60337 , n60338 , n60339 , n60340 , n60341 , n60342 , n60343 , n60344 , n60345 , n60346 , 
     n60347 , n60348 , n60349 , n60350 , n60351 , n60352 , n60353 , n60354 , n60355 , n60356 , 
     n60357 , n60358 , n60359 , n60360 , n60361 , n60362 , n60363 , n60364 , n60365 , n60366 , 
     n60367 , n60368 , n60369 , n60370 , n60371 , n60372 , n60373 , n60374 , n60375 , n60376 , 
     n60377 , n60378 , n60379 , n60380 , n60381 , n60382 , n60383 , n60384 , n60385 , n60386 , 
     n60387 , n60388 , n60389 , n60390 , n60391 , n60392 , n60393 , n60394 , n60395 , n60396 , 
     n60397 , n60398 , n60399 , n60400 , n60401 , n60402 , n60403 , n60404 , n60405 , n60406 , 
     n60407 , n60408 , n60409 , n60410 , n60411 , n60412 , n60413 , n60414 , n60415 , n60416 , 
     n60417 , n60418 , n60419 , n60420 , n60421 , n60422 , n60423 , n60424 , n60425 , n60426 , 
     n60427 , n60428 , n60429 , n60430 , n60431 , n60432 , n60433 , n60434 , n60435 , n60436 , 
     n60437 , n60438 , n60439 , n60440 , n60441 , n60442 , n60443 , n60444 , n60445 , n60446 , 
     n60447 , n60448 , n60449 , n60450 , n60451 , n60452 , n60453 , n60454 , n60455 , n60456 , 
     n60457 , n60458 , n60459 , n60460 , n60461 , n60462 , n60463 , n60464 , n60465 , n60466 , 
     n60467 , n60468 , n60469 , n60470 , n60471 , n60472 , n60473 , n60474 , n60475 , n60476 , 
     n60477 , n60478 , n60479 , n60480 , n60481 , n60482 , n60483 , n60484 , n60485 , n60486 , 
     n60487 , n60488 , n60489 , n60490 , n60491 , n60492 , n60493 , n60494 , n60495 , n60496 , 
     n60497 , n60498 , n60499 , n60500 , n60501 , n60502 , n60503 , n60504 , n60505 , n60506 , 
     n60507 , n60508 , n60509 , n60510 , n60511 , n60512 , n60513 , n60514 , n60515 , n60516 , 
     n60517 , n60518 , n60519 , n60520 , n60521 , n60522 , n60523 , n60524 , n60525 , n60526 , 
     n60527 , n60528 , n60529 , n60530 , n60531 , n60532 , n60533 , n60534 , n60535 , n60536 , 
     n60537 , n60538 , n60539 , n60540 , n60541 , n60542 , n60543 , n60544 , n60545 , n60546 , 
     n60547 , n60548 , n60549 , n60550 , n60551 , n60552 , n60553 , n60554 , n60555 , n60556 , 
     n60557 , n60558 , n60559 , n60560 , n60561 , n60562 , n60563 , n60564 , n60565 , n60566 , 
     n60567 , n60568 , n60569 , n60570 , n60571 , n60572 , n60573 , n60574 , n60575 , n60576 , 
     n60577 , n60578 , n60579 , n60580 , n60581 , n60582 , n60583 , n60584 , n60585 , n60586 , 
     n60587 , n60588 , n60589 , n60590 , n60591 , n60592 , n60593 , n60594 , n60595 , n60596 , 
     n60597 , n60598 , n60599 , n60600 , n60601 , n60602 , n60603 , n60604 , n60605 , n60606 , 
     n60607 , n60608 , n60609 , n60610 , n60611 , n60612 , n60613 , n60614 , n60615 , n60616 , 
     n60617 , n60618 , n60619 , n60620 , n60621 , n60622 , n60623 , n60624 , n60625 , n60626 , 
     n60627 , n60628 , n60629 , n60630 , n60631 , n60632 , n60633 , n60634 , n60635 , n60636 , 
     n60637 , n60638 , n60639 , n60640 , n60641 , n60642 , n60643 , n60644 , n60645 , n60646 , 
     n60647 , n60648 , n60649 , n60650 , n60651 , n60652 , n60653 , n60654 , n60655 , n60656 , 
     n60657 , n60658 , n60659 , n60660 , n60661 , n60662 , n60663 , n60664 , n60665 , n60666 , 
     n60667 , n60668 , n60669 , n60670 , n60671 , n60672 , n60673 , n60674 , n60675 , n60676 , 
     n60677 , n60678 , n60679 , n60680 , n60681 , n60682 , n60683 , n60684 , n60685 , n60686 , 
     n60687 , n60688 , n60689 , n60690 , n60691 , n60692 , n60693 , n60694 , n60695 , n60696 , 
     n60697 , n60698 , n60699 , n60700 , n60701 , n60702 , n60703 , n60704 , n60705 , n60706 , 
     n60707 , n60708 , n60709 , n60710 , n60711 , n60712 , n60713 , n60714 , n60715 , n60716 , 
     n60717 , n60718 , n60719 , n60720 , n60721 , n60722 , n60723 , n60724 , n60725 , n60726 , 
     n60727 , n60728 , n60729 , n60730 , n60731 , n60732 , n60733 , n60734 , n60735 , n60736 , 
     n60737 , n60738 , n60739 , n60740 , n60741 , n60742 , n60743 , n60744 , n60745 , n60746 , 
     n60747 , n60748 , n60749 , n60750 , n60751 , n60752 , n60753 , n60754 , n60755 , n60756 , 
     n60757 , n60758 , n60759 , n60760 , n60761 , n60762 , n60763 , n60764 , n60765 , n60766 , 
     n60767 , n60768 , n60769 , n60770 , n60771 , n60772 , n60773 , n60774 , n60775 , n60776 , 
     n60777 , n60778 , n60779 , n60780 , n60781 , n60782 , n60783 , n60784 , n60785 , n60786 , 
     n60787 , n60788 , n60789 , n60790 , n60791 , n60792 , n60793 , n60794 , n60795 , n60796 , 
     n60797 , n60798 , n60799 , n60800 , n60801 , n60802 , n60803 , n60804 , n60805 , n60806 , 
     n60807 , n60808 , n60809 , n60810 , n60811 , n60812 , n60813 , n60814 , n60815 , n60816 , 
     n60817 , n60818 , n60819 , n60820 , n60821 , n60822 , n60823 , n60824 , n60825 , n60826 , 
     n60827 , n60828 , n60829 , n60830 , n60831 , n60832 , n60833 , n60834 , n60835 , n60836 , 
     n60837 , n60838 , n60839 , n60840 , n60841 , n60842 , n60843 , n60844 , n60845 , n60846 , 
     n60847 , n60848 , n60849 , n60850 , n60851 , n60852 , n60853 , n60854 , n60855 , n60856 , 
     n60857 , n60858 , n60859 , n60860 , n60861 , n60862 , n60863 , n60864 , n60865 , n60866 , 
     n60867 , n60868 , n60869 , n60870 , n60871 , n60872 , n60873 , n60874 , n60875 , n60876 , 
     n60877 , n60878 , n60879 , n60880 , n60881 , n60882 , n60883 , n60884 , n60885 , n60886 , 
     n60887 , n60888 , n60889 , n60890 , n60891 , n60892 , n60893 , n60894 , n60895 , n60896 , 
     n60897 , n60898 , n60899 , n60900 , n60901 , n60902 , n60903 , n60904 , n60905 , n60906 , 
     n60907 , n60908 , n60909 , n60910 , n60911 , n60912 , n60913 , n60914 , n60915 , n60916 , 
     n60917 , n60918 , n60919 , n60920 , n60921 , n60922 , n60923 , n60924 , n60925 , n60926 , 
     n60927 , n60928 , n60929 , n60930 , n60931 , n60932 , n60933 , n60934 , n60935 , n60936 , 
     n60937 , n60938 , n60939 , n60940 , n60941 , n60942 , n60943 , n60944 , n60945 , n60946 , 
     n60947 , n60948 , n60949 , n60950 , n60951 , n60952 , n60953 , n60954 , n60955 , n60956 , 
     n60957 , n60958 , n60959 , n60960 , n60961 , n60962 , n60963 , n60964 , n60965 , n60966 , 
     n60967 , n60968 , n60969 , n60970 , n60971 , n60972 , n60973 , n60974 , n60975 , n60976 , 
     n60977 , n60978 , n60979 , n60980 , n60981 , n60982 , n60983 , n60984 , n60985 , n60986 , 
     n60987 , n60988 , n60989 , n60990 , n60991 , n60992 , n60993 , n60994 , n60995 , n60996 , 
     n60997 , n60998 , n60999 , n61000 , n61001 , n61002 , n61003 , n61004 , n61005 , n61006 , 
     n61007 , n61008 , n61009 , n61010 , n61011 , n61012 , n61013 , n61014 , n61015 , n61016 , 
     n61017 , n61018 , n61019 , n61020 , n61021 , n61022 , n61023 , n61024 , n61025 , n61026 , 
     n61027 , n61028 , n61029 , n61030 , n61031 , n61032 , n61033 , n61034 , n61035 , n61036 , 
     n61037 , n61038 , n61039 , n61040 , n61041 , n61042 , n61043 , n61044 , n61045 , n61046 , 
     n61047 , n61048 , n61049 , n61050 , n61051 , n61052 , n61053 , n61054 , n61055 , n61056 , 
     n61057 , n61058 , n61059 , n61060 , n61061 , n61062 , n61063 , n61064 , n61065 , n61066 , 
     n61067 , n61068 , n61069 , n61070 , n61071 , n61072 , n61073 , n61074 , n61075 , n61076 , 
     n61077 , n61078 , n61079 , n61080 , n61081 , n61082 , n61083 , n61084 , n61085 , n61086 , 
     n61087 , n61088 , n61089 , n61090 , n61091 , n61092 , n61093 , n61094 , n61095 , n61096 , 
     n61097 , n61098 , n61099 , n61100 , n61101 , n61102 , n61103 , n61104 , n61105 , n61106 , 
     n61107 , n61108 , n61109 , n61110 , n61111 , n61112 , n61113 , n61114 , n61115 , n61116 , 
     n61117 , n61118 , n61119 , n61120 , n61121 , n61122 , n61123 , n61124 , n61125 , n61126 , 
     n61127 , n61128 , n61129 , n61130 , n61131 , n61132 , n61133 , n61134 , n61135 , n61136 , 
     n61137 , n61138 , n61139 , n61140 , n61141 , n61142 , n61143 , n61144 , n61145 , n61146 , 
     n61147 , n61148 , n61149 , n61150 , n61151 , n61152 , n61153 , n61154 , n61155 , n61156 , 
     n61157 , n61158 , n61159 , n61160 , n61161 , n61162 , n61163 , n61164 , n61165 , n61166 , 
     n61167 , n61168 , n61169 , n61170 , n61171 , n61172 , n61173 , n61174 , n61175 , n61176 , 
     n61177 , n61178 , n61179 , n61180 , n61181 , n61182 , n61183 , n61184 , n61185 , n61186 , 
     n61187 , n61188 , n61189 , n61190 , n61191 , n61192 , n61193 , n61194 , n61195 , n61196 , 
     n61197 , n61198 , n61199 , n61200 , n61201 , n61202 , n61203 , n61204 , n61205 , n61206 , 
     n61207 , n61208 , n61209 , n61210 , n61211 , n61212 , n61213 , n61214 , n61215 , n61216 , 
     n61217 , n61218 , n61219 , n61220 , n61221 , n61222 , n61223 , n61224 , n61225 , n61226 , 
     n61227 , n61228 , n61229 , n61230 , n61231 , n61232 , n61233 , n61234 , n61235 , n61236 , 
     n61237 , n61238 , n61239 , n61240 , n61241 , n61242 , n61243 , n61244 , n61245 , n61246 , 
     n61247 , n61248 , n61249 , n61250 , n61251 , n61252 , n61253 , n61254 , n61255 , n61256 , 
     n61257 , n61258 , n61259 , n61260 , n61261 , n61262 , n61263 , n61264 , n61265 , n61266 , 
     n61267 , n61268 , n61269 , n61270 , n61271 , n61272 , n61273 , n61274 , n61275 , n61276 , 
     n61277 , n61278 , n61279 , n61280 , n61281 , n61282 , n61283 , n61284 , n61285 , n61286 , 
     n61287 , n61288 , n61289 , n61290 , n61291 , n61292 , n61293 , n61294 , n61295 , n61296 , 
     n61297 , n61298 , n61299 , n61300 , n61301 , n61302 , n61303 , n61304 , n61305 , n61306 , 
     n61307 , n61308 , n61309 , n61310 , n61311 , n61312 , n61313 , n61314 , n61315 , n61316 , 
     n61317 , n61318 , n61319 , n61320 , n61321 , n61322 , n61323 , n61324 , n61325 , n61326 , 
     n61327 , n61328 , n61329 , n61330 , n61331 , n61332 , n61333 , n61334 , n61335 , n61336 , 
     n61337 , n61338 , n61339 , n61340 , n61341 , n61342 , n61343 , n61344 , n61345 , n61346 , 
     n61347 , n61348 , n61349 , n61350 , n61351 , n61352 , n61353 , n61354 , n61355 , n61356 , 
     n61357 , n61358 , n61359 , n61360 , n61361 , n61362 , n61363 , n61364 , n61365 , n61366 , 
     n61367 , n61368 , n61369 , n61370 , n61371 , n61372 , n61373 , n61374 , n61375 , n61376 , 
     n61377 , n61378 , n61379 , n61380 , n61381 , n61382 , n61383 , n61384 , n61385 , n61386 , 
     n61387 , n61388 , n61389 , n61390 , n61391 , n61392 , n61393 , n61394 , n61395 , n61396 , 
     n61397 , n61398 , n61399 , n61400 , n61401 , n61402 , n61403 , n61404 , n61405 , n61406 , 
     n61407 , n61408 , n61409 , n61410 , n61411 , n61412 , n61413 , n61414 , n61415 , n61416 , 
     n61417 , n61418 , n61419 , n61420 , n61421 , n61422 , n61423 , n61424 , n61425 , n61426 , 
     n61427 , n61428 , n61429 , n61430 , n61431 , n61432 , n61433 , n61434 , n61435 , n61436 , 
     n61437 , n61438 , n61439 , n61440 , n61441 , n61442 , n61443 , n61444 , n61445 , n61446 , 
     n61447 , n61448 , n61449 , n61450 , n61451 , n61452 , n61453 , n61454 , n61455 , n61456 , 
     n61457 , n61458 , n61459 , n61460 , n61461 , n61462 , n61463 , n61464 , n61465 , n61466 , 
     n61467 , n61468 , n61469 , n61470 , n61471 , n61472 , n61473 , n61474 , n61475 , n61476 , 
     n61477 , n61478 , n61479 , n61480 , n61481 , n61482 , n61483 , n61484 , n61485 , n61486 , 
     n61487 , n61488 , n61489 , n61490 , n61491 , n61492 , n61493 , n61494 , n61495 , n61496 , 
     n61497 , n61498 , n61499 , n61500 , n61501 , n61502 , n61503 , n61504 , n61505 , n61506 , 
     n61507 , n61508 , n61509 , n61510 , n61511 , n61512 , n61513 , n61514 , n61515 , n61516 , 
     n61517 , n61518 , n61519 , n61520 , n61521 , n61522 , n61523 , n61524 , n61525 , n61526 , 
     n61527 , n61528 , n61529 , n61530 , n61531 , n61532 , n61533 , n61534 , n61535 , n61536 , 
     n61537 , n61538 , n61539 , n61540 , n61541 , n61542 , n61543 , n61544 , n61545 , n61546 , 
     n61547 , n61548 , n61549 , n61550 , n61551 , n61552 , n61553 , n61554 , n61555 , n61556 , 
     n61557 , n61558 , n61559 , n61560 , n61561 , n61562 , n61563 , n61564 , n61565 , n61566 , 
     n61567 , n61568 , n61569 , n61570 , n61571 , n61572 , n61573 , n61574 , n61575 , n61576 , 
     n61577 , n61578 , n61579 , n61580 , n61581 , n61582 , n61583 , n61584 , n61585 , n61586 , 
     n61587 , n61588 , n61589 , n61590 , n61591 , n61592 , n61593 , n61594 , n61595 , n61596 , 
     n61597 , n61598 , n61599 , n61600 , n61601 , n61602 , n61603 , n61604 , n61605 , n61606 , 
     n61607 , n61608 , n61609 , n61610 , n61611 , n61612 , n61613 , n61614 , n61615 , n61616 , 
     n61617 , n61618 , n61619 , n61620 , n61621 , n61622 , n61623 , n61624 , n61625 , n61626 , 
     n61627 , n61628 , n61629 , n61630 , n61631 , n61632 , n61633 , n61634 , n61635 , n61636 , 
     n61637 , n61638 , n61639 , n61640 , n61641 , n61642 , n61643 , n61644 , n61645 , n61646 , 
     n61647 , n61648 , n61649 , n61650 , n61651 , n61652 , n61653 , n61654 , n61655 , n61656 , 
     n61657 , n61658 , n61659 , n61660 , n61661 , n61662 , n61663 , n61664 , n61665 , n61666 , 
     n61667 , n61668 , n61669 , n61670 , n61671 , n61672 , n61673 , n61674 , n61675 , n61676 , 
     n61677 , n61678 , n61679 , n61680 , n61681 , n61682 , n61683 , n61684 , n61685 , n61686 , 
     n61687 , n61688 , n61689 , n61690 , n61691 , n61692 , n61693 , n61694 , n61695 , n61696 , 
     n61697 , n61698 , n61699 , n61700 , n61701 , n61702 , n61703 , n61704 , n61705 , n61706 , 
     n61707 , n61708 , n61709 , n61710 , n61711 , n61712 , n61713 , n61714 , n61715 , n61716 , 
     n61717 , n61718 , n61719 , n61720 , n61721 , n61722 , n61723 , n61724 , n61725 , n61726 , 
     n61727 , n61728 , n61729 , n61730 , n61731 , n61732 , n61733 , n61734 , n61735 , n61736 , 
     n61737 , n61738 , n61739 , n61740 , n61741 , n61742 , n61743 , n61744 , n61745 , n61746 , 
     n61747 , n61748 , n61749 , n61750 , n61751 , n61752 , n61753 , n61754 , n61755 , n61756 , 
     n61757 , n61758 , n61759 , n61760 , n61761 , n61762 , n61763 , n61764 , n61765 , n61766 , 
     n61767 , n61768 , n61769 , n61770 , n61771 , n61772 , n61773 , n61774 , n61775 , n61776 , 
     n61777 , n61778 , n61779 , n61780 , n61781 , n61782 , n61783 , n61784 , n61785 , n61786 , 
     n61787 , n61788 , n61789 , n61790 , n61791 , n61792 , n61793 , n61794 , n61795 , n61796 , 
     n61797 , n61798 , n61799 , n61800 , n61801 , n61802 , n61803 , n61804 , n61805 , n61806 , 
     n61807 , n61808 , n61809 , n61810 , n61811 , n61812 , n61813 , n61814 , n61815 , n61816 , 
     n61817 , n61818 , n61819 , n61820 , n61821 , n61822 , n61823 , n61824 , n61825 , n61826 , 
     n61827 , n61828 , n61829 , n61830 , n61831 , n61832 , n61833 , n61834 , n61835 , n61836 , 
     n61837 , n61838 , n61839 , n61840 , n61841 , n61842 , n61843 , n61844 , n61845 , n61846 , 
     n61847 , n61848 , n61849 , n61850 , n61851 , n61852 , n61853 , n61854 , n61855 , n61856 , 
     n61857 , n61858 , n61859 , n61860 , n61861 , n61862 , n61863 , n61864 , n61865 , n61866 , 
     n61867 , n61868 , n61869 , n61870 , n61871 , n61872 , n61873 , n61874 , n61875 , n61876 , 
     n61877 , n61878 , n61879 , n61880 , n61881 , n61882 , n61883 , n61884 , n61885 , n61886 , 
     n61887 , n61888 , n61889 , n61890 , n61891 , n61892 , n61893 , n61894 , n61895 , n61896 , 
     n61897 , n61898 , n61899 , n61900 , n61901 , n61902 , n61903 , n61904 , n61905 , n61906 , 
     n61907 , n61908 , n61909 , n61910 , n61911 , n61912 , n61913 , n61914 , n61915 , n61916 , 
     n61917 , n61918 , n61919 , n61920 , n61921 , n61922 , n61923 , n61924 , n61925 , n61926 , 
     n61927 , n61928 , n61929 , n61930 , n61931 , n61932 , n61933 , n61934 , n61935 , n61936 , 
     n61937 , n61938 , n61939 , n61940 , n61941 , n61942 , n61943 , n61944 , n61945 , n61946 , 
     n61947 , n61948 , n61949 , n61950 , n61951 , n61952 , n61953 , n61954 , n61955 , n61956 , 
     n61957 , n61958 , n61959 , n61960 , n61961 , n61962 , n61963 , n61964 , n61965 , n61966 , 
     n61967 , n61968 , n61969 , n61970 , n61971 , n61972 , n61973 , n61974 , n61975 , n61976 , 
     n61977 , n61978 , n61979 , n61980 , n61981 , n61982 , n61983 , n61984 , n61985 , n61986 , 
     n61987 , n61988 , n61989 , n61990 , n61991 , n61992 , n61993 , n61994 , n61995 , n61996 , 
     n61997 , n61998 , n61999 , n62000 , n62001 , n62002 , n62003 , n62004 , n62005 , n62006 , 
     n62007 , n62008 , n62009 , n62010 , n62011 , n62012 , n62013 , n62014 , n62015 , n62016 , 
     n62017 , n62018 , n62019 , n62020 , n62021 , n62022 , n62023 , n62024 , n62025 , n62026 , 
     n62027 , n62028 , n62029 , n62030 , n62031 , n62032 , n62033 , n62034 , n62035 , n62036 , 
     n62037 , n62038 , n62039 , n62040 , n62041 , n62042 , n62043 , n62044 , n62045 , n62046 , 
     n62047 , n62048 , n62049 , n62050 , n62051 , n62052 , n62053 , n62054 , n62055 , n62056 , 
     n62057 , n62058 , n62059 , n62060 , n62061 , n62062 , n62063 , n62064 , n62065 , n62066 , 
     n62067 , n62068 , n62069 , n62070 , n62071 , n62072 , n62073 , n62074 , n62075 , n62076 , 
     n62077 , n62078 , n62079 , n62080 , n62081 , n62082 , n62083 , n62084 , n62085 , n62086 , 
     n62087 , n62088 , n62089 , n62090 , n62091 , n62092 , n62093 , n62094 , n62095 , n62096 , 
     n62097 , n62098 , n62099 , n62100 , n62101 , n62102 , n62103 , n62104 , n62105 , n62106 , 
     n62107 , n62108 , n62109 , n62110 , n62111 , n62112 , n62113 , n62114 , n62115 , n62116 , 
     n62117 , n62118 , n62119 , n62120 , n62121 , n62122 , n62123 , n62124 , n62125 , n62126 , 
     n62127 , n62128 , n62129 , n62130 , n62131 , n62132 , n62133 , n62134 , n62135 , n62136 , 
     n62137 , n62138 , n62139 , n62140 , n62141 , n62142 , n62143 , n62144 , n62145 , n62146 , 
     n62147 , n62148 , n62149 , n62150 , n62151 , n62152 , n62153 , n62154 , n62155 , n62156 , 
     n62157 , n62158 , n62159 , n62160 , n62161 , n62162 , n62163 , n62164 , n62165 , n62166 , 
     n62167 , n62168 , n62169 , n62170 , n62171 , n62172 , n62173 , n62174 , n62175 , n62176 , 
     n62177 , n62178 , n62179 , n62180 , n62181 , n62182 , n62183 , n62184 , n62185 , n62186 , 
     n62187 , n62188 , n62189 , n62190 , n62191 , n62192 , n62193 , n62194 , n62195 , n62196 , 
     n62197 , n62198 , n62199 , n62200 , n62201 , n62202 , n62203 , n62204 , n62205 , n62206 , 
     n62207 , n62208 , n62209 , n62210 , n62211 , n62212 , n62213 , n62214 , n62215 , n62216 , 
     n62217 , n62218 , n62219 , n62220 , n62221 , n62222 , n62223 , n62224 , n62225 , n62226 , 
     n62227 , n62228 , n62229 , n62230 , n62231 , n62232 , n62233 , n62234 , n62235 , n62236 , 
     n62237 , n62238 , n62239 , n62240 , n62241 , n62242 , n62243 , n62244 , n62245 , n62246 , 
     n62247 , n62248 , n62249 , n62250 , n62251 , n62252 , n62253 , n62254 , n62255 , n62256 , 
     n62257 , n62258 , n62259 , n62260 , n62261 , n62262 , n62263 , n62264 , n62265 , n62266 , 
     n62267 , n62268 , n62269 , n62270 , n62271 , n62272 , n62273 , n62274 , n62275 , n62276 , 
     n62277 , n62278 , n62279 , n62280 , n62281 , n62282 , n62283 , n62284 , n62285 , n62286 , 
     n62287 , n62288 , n62289 , n62290 , n62291 , n62292 , n62293 , n62294 , n62295 , n62296 , 
     n62297 , n62298 , n62299 , n62300 , n62301 , n62302 , n62303 , n62304 , n62305 , n62306 , 
     n62307 , n62308 , n62309 , n62310 , n62311 , n62312 , n62313 , n62314 , n62315 , n62316 , 
     n62317 , n62318 , n62319 , n62320 , n62321 , n62322 , n62323 , n62324 , n62325 , n62326 , 
     n62327 , n62328 , n62329 , n62330 , n62331 , n62332 , n62333 , n62334 , n62335 , n62336 , 
     n62337 , n62338 , n62339 , n62340 , n62341 , n62342 , n62343 , n62344 , n62345 , n62346 , 
     n62347 , n62348 , n62349 , n62350 , n62351 , n62352 , n62353 , n62354 , n62355 , n62356 , 
     n62357 , n62358 , n62359 , n62360 , n62361 , n62362 , n62363 , n62364 , n62365 , n62366 , 
     n62367 , n62368 , n62369 , n62370 , n62371 , n62372 , n62373 , n62374 , n62375 , n62376 , 
     n62377 , n62378 , n62379 , n62380 , n62381 , n62382 , n62383 , n62384 , n62385 , n62386 , 
     n62387 , n62388 , n62389 , n62390 , n62391 , n62392 , n62393 , n62394 , n62395 , n62396 , 
     n62397 , n62398 , n62399 , n62400 , n62401 , n62402 , n62403 , n62404 , n62405 , n62406 , 
     n62407 , n62408 , n62409 , n62410 , n62411 , n62412 , n62413 , n62414 , n62415 , n62416 , 
     n62417 , n62418 , n62419 , n62420 , n62421 , n62422 , n62423 , n62424 , n62425 , n62426 , 
     n62427 , n62428 , n62429 , n62430 , n62431 , n62432 , n62433 , n62434 , n62435 , n62436 , 
     n62437 , n62438 , n62439 , n62440 , n62441 , n62442 , n62443 , n62444 , n62445 , n62446 , 
     n62447 , n62448 , n62449 , n62450 , n62451 , n62452 , n62453 , n62454 , n62455 , n62456 , 
     n62457 , n62458 , n62459 , n62460 , n62461 , n62462 , n62463 , n62464 , n62465 , n62466 , 
     n62467 , n62468 , n62469 , n62470 , n62471 , n62472 , n62473 , n62474 , n62475 , n62476 , 
     n62477 , n62478 , n62479 , n62480 , n62481 , n62482 , n62483 , n62484 , n62485 , n62486 , 
     n62487 , n62488 , n62489 , n62490 , n62491 , n62492 , n62493 , n62494 , n62495 , n62496 , 
     n62497 , n62498 , n62499 , n62500 , n62501 , n62502 , n62503 , n62504 , n62505 , n62506 , 
     n62507 , n62508 , n62509 , n62510 , n62511 , n62512 , n62513 , n62514 , n62515 , n62516 , 
     n62517 , n62518 , n62519 , n62520 , n62521 , n62522 , n62523 , n62524 , n62525 , n62526 , 
     n62527 , n62528 , n62529 , n62530 , n62531 , n62532 , n62533 , n62534 , n62535 , n62536 , 
     n62537 , n62538 , n62539 , n62540 , n62541 , n62542 , n62543 , n62544 , n62545 , n62546 , 
     n62547 , n62548 , n62549 , n62550 , n62551 , n62552 , n62553 , n62554 , n62555 , n62556 , 
     n62557 , n62558 , n62559 , n62560 , n62561 , n62562 , n62563 , n62564 , n62565 , n62566 , 
     n62567 , n62568 , n62569 , n62570 , n62571 , n62572 , n62573 , n62574 , n62575 , n62576 , 
     n62577 , n62578 , n62579 , n62580 , n62581 , n62582 , n62583 , n62584 , n62585 , n62586 , 
     n62587 , n62588 , n62589 , n62590 , n62591 , n62592 , n62593 , n62594 , n62595 , n62596 , 
     n62597 , n62598 , n62599 , n62600 , n62601 , n62602 , n62603 , n62604 , n62605 , n62606 , 
     n62607 , n62608 , n62609 , n62610 , n62611 , n62612 , n62613 , n62614 , n62615 , n62616 , 
     n62617 , n62618 , n62619 , n62620 , n62621 , n62622 , n62623 , n62624 , n62625 , n62626 , 
     n62627 , n62628 , n62629 , n62630 , n62631 , n62632 , n62633 , n62634 , n62635 , n62636 , 
     n62637 , n62638 , n62639 , n62640 , n62641 , n62642 , n62643 , n62644 , n62645 , n62646 , 
     n62647 , n62648 , n62649 , n62650 , n62651 , n62652 , n62653 , n62654 , n62655 , n62656 , 
     n62657 , n62658 , n62659 , n62660 , n62661 , n62662 , n62663 , n62664 , n62665 , n62666 , 
     n62667 , n62668 , n62669 , n62670 , n62671 , n62672 , n62673 , n62674 , n62675 , n62676 , 
     n62677 , n62678 , n62679 , n62680 , n62681 , n62682 , n62683 , n62684 , n62685 , n62686 , 
     n62687 , n62688 , n62689 , n62690 , n62691 , n62692 , n62693 , n62694 , n62695 , n62696 , 
     n62697 , n62698 , n62699 , n62700 , n62701 , n62702 , n62703 , n62704 , n62705 , n62706 , 
     n62707 , n62708 , n62709 , n62710 , n62711 , n62712 , n62713 , n62714 , n62715 , n62716 , 
     n62717 , n62718 , n62719 , n62720 , n62721 , n62722 , n62723 , n62724 , n62725 , n62726 , 
     n62727 , n62728 , n62729 , n62730 , n62731 , n62732 , n62733 , n62734 , n62735 , n62736 , 
     n62737 , n62738 , n62739 , n62740 , n62741 , n62742 , n62743 , n62744 , n62745 , n62746 , 
     n62747 , n62748 , n62749 , n62750 , n62751 , n62752 , n62753 , n62754 , n62755 , n62756 , 
     n62757 , n62758 , n62759 , n62760 , n62761 , n62762 , n62763 , n62764 , n62765 , n62766 , 
     n62767 , n62768 , n62769 , n62770 , n62771 , n62772 , n62773 , n62774 , n62775 , n62776 , 
     n62777 , n62778 , n62779 , n62780 , n62781 , n62782 , n62783 , n62784 , n62785 , n62786 , 
     n62787 , n62788 , n62789 , n62790 , n62791 , n62792 , n62793 , n62794 , n62795 , n62796 , 
     n62797 , n62798 , n62799 , n62800 , n62801 , n62802 , n62803 , n62804 , n62805 , n62806 , 
     n62807 , n62808 , n62809 , n62810 , n62811 , n62812 , n62813 , n62814 , n62815 , n62816 , 
     n62817 , n62818 , n62819 , n62820 , n62821 , n62822 , n62823 , n62824 , n62825 , n62826 , 
     n62827 , n62828 , n62829 , n62830 , n62831 , n62832 , n62833 , n62834 , n62835 , n62836 , 
     n62837 , n62838 , n62839 , n62840 , n62841 , n62842 , n62843 , n62844 , n62845 , n62846 , 
     n62847 , n62848 , n62849 , n62850 , n62851 , n62852 , n62853 , n62854 , n62855 , n62856 , 
     n62857 , n62858 , n62859 , n62860 , n62861 , n62862 , n62863 , n62864 , n62865 , n62866 , 
     n62867 , n62868 , n62869 , n62870 , n62871 , n62872 , n62873 , n62874 , n62875 , n62876 , 
     n62877 , n62878 , n62879 , n62880 , n62881 , n62882 , n62883 , n62884 , n62885 , n62886 , 
     n62887 , n62888 , n62889 , n62890 , n62891 , n62892 , n62893 , n62894 , n62895 , n62896 , 
     n62897 , n62898 , n62899 , n62900 , n62901 , n62902 , n62903 , n62904 , n62905 , n62906 , 
     n62907 , n62908 , n62909 , n62910 , n62911 , n62912 , n62913 , n62914 , n62915 , n62916 , 
     n62917 , n62918 , n62919 , n62920 , n62921 , n62922 , n62923 , n62924 , n62925 , n62926 , 
     n62927 , n62928 , n62929 , n62930 , n62931 , n62932 , n62933 , n62934 , n62935 , n62936 , 
     n62937 , n62938 , n62939 , n62940 , n62941 , n62942 , n62943 , n62944 , n62945 , n62946 , 
     n62947 , n62948 , n62949 , n62950 , n62951 , n62952 , n62953 , n62954 , n62955 , n62956 , 
     n62957 , n62958 , n62959 , n62960 , n62961 , n62962 , n62963 , n62964 , n62965 , n62966 , 
     n62967 , n62968 , n62969 , n62970 , n62971 , n62972 , n62973 , n62974 , n62975 , n62976 , 
     n62977 , n62978 , n62979 , n62980 , n62981 , n62982 , n62983 , n62984 , n62985 , n62986 , 
     n62987 , n62988 , n62989 , n62990 , n62991 , n62992 , n62993 , n62994 , n62995 , n62996 , 
     n62997 , n62998 , n62999 , n63000 , n63001 , n63002 , n63003 , n63004 , n63005 , n63006 , 
     n63007 , n63008 , n63009 , n63010 , n63011 , n63012 , n63013 , n63014 , n63015 , n63016 , 
     n63017 , n63018 , n63019 , n63020 , n63021 , n63022 , n63023 , n63024 , n63025 , n63026 , 
     n63027 , n63028 , n63029 , n63030 , n63031 , n63032 , n63033 , n63034 , n63035 , n63036 , 
     n63037 , n63038 , n63039 , n63040 , n63041 , n63042 , n63043 , n63044 , n63045 , n63046 , 
     n63047 , n63048 , n63049 , n63050 , n63051 , n63052 , n63053 , n63054 , n63055 , n63056 , 
     n63057 , n63058 , n63059 , n63060 , n63061 , n63062 , n63063 , n63064 , n63065 , n63066 , 
     n63067 , n63068 , n63069 , n63070 , n63071 , n63072 , n63073 , n63074 , n63075 , n63076 , 
     n63077 , n63078 , n63079 , n63080 , n63081 , n63082 , n63083 , n63084 , n63085 , n63086 , 
     n63087 , n63088 , n63089 , n63090 , n63091 , n63092 , n63093 , n63094 , n63095 , n63096 , 
     n63097 , n63098 , n63099 , n63100 , n63101 , n63102 , n63103 , n63104 , n63105 , n63106 , 
     n63107 , n63108 , n63109 , n63110 , n63111 , n63112 , n63113 , n63114 , n63115 , n63116 , 
     n63117 , n63118 , n63119 , n63120 , n63121 , n63122 , n63123 , n63124 , n63125 , n63126 , 
     n63127 , n63128 , n63129 , n63130 , n63131 , n63132 , n63133 , n63134 , n63135 , n63136 , 
     n63137 , n63138 , n63139 , n63140 , n63141 , n63142 , n63143 , n63144 , n63145 , n63146 , 
     n63147 , n63148 , n63149 , n63150 , n63151 , n63152 , n63153 , n63154 , n63155 , n63156 , 
     n63157 , n63158 , n63159 , n63160 , n63161 , n63162 , n63163 , n63164 , n63165 , n63166 , 
     n63167 , n63168 , n63169 , n63170 , n63171 , n63172 , n63173 , n63174 , n63175 , n63176 , 
     n63177 , n63178 , n63179 , n63180 , n63181 , n63182 , n63183 , n63184 , n63185 , n63186 , 
     n63187 , n63188 , n63189 , n63190 , n63191 , n63192 , n63193 , n63194 , n63195 , n63196 , 
     n63197 , n63198 , n63199 , n63200 , n63201 , n63202 , n63203 , n63204 , n63205 , n63206 , 
     n63207 , n63208 , n63209 , n63210 , n63211 , n63212 , n63213 , n63214 , n63215 , n63216 , 
     n63217 , n63218 , n63219 , n63220 , n63221 , n63222 , n63223 , n63224 , n63225 , n63226 , 
     n63227 , n63228 , n63229 , n63230 , n63231 , n63232 , n63233 , n63234 , n63235 , n63236 , 
     n63237 , n63238 , n63239 , n63240 , n63241 , n63242 , n63243 , n63244 , n63245 , n63246 , 
     n63247 , n63248 , n63249 , n63250 , n63251 , n63252 , n63253 , n63254 , n63255 , n63256 , 
     n63257 , n63258 , n63259 , n63260 , n63261 , n63262 , n63263 , n63264 , n63265 , n63266 , 
     n63267 , n63268 , n63269 , n63270 , n63271 , n63272 , n63273 , n63274 , n63275 , n63276 , 
     n63277 , n63278 , n63279 , n63280 , n63281 , n63282 , n63283 , n63284 , n63285 , n63286 , 
     n63287 , n63288 , n63289 , n63290 , n63291 , n63292 , n63293 , n63294 , n63295 , n63296 , 
     n63297 , n63298 , n63299 , n63300 , n63301 , n63302 , n63303 , n63304 , n63305 , n63306 , 
     n63307 , n63308 , n63309 , n63310 , n63311 , n63312 , n63313 , n63314 , n63315 , n63316 , 
     n63317 , n63318 , n63319 , n63320 , n63321 , n63322 , n63323 , n63324 , n63325 , n63326 , 
     n63327 , n63328 , n63329 , n63330 , n63331 , n63332 , n63333 , n63334 , n63335 , n63336 , 
     n63337 , n63338 , n63339 , n63340 , n63341 , n63342 , n63343 , n63344 , n63345 , n63346 , 
     n63347 , n63348 , n63349 , n63350 , n63351 , n63352 , n63353 , n63354 , n63355 , n63356 , 
     n63357 , n63358 , n63359 , n63360 , n63361 , n63362 , n63363 , n63364 , n63365 , n63366 , 
     n63367 , n63368 , n63369 , n63370 , n63371 , n63372 , n63373 , n63374 , n63375 , n63376 , 
     n63377 , n63378 , n63379 , n63380 , n63381 , n63382 , n63383 , n63384 , n63385 , n63386 , 
     n63387 , n63388 , n63389 , n63390 , n63391 , n63392 , n63393 , n63394 , n63395 , n63396 , 
     n63397 , n63398 , n63399 , n63400 , n63401 , n63402 , n63403 , n63404 , n63405 , n63406 , 
     n63407 , n63408 , n63409 , n63410 , n63411 , n63412 , n63413 , n63414 , n63415 , n63416 , 
     n63417 , n63418 , n63419 , n63420 , n63421 , n63422 , n63423 , n63424 , n63425 , n63426 , 
     n63427 , n63428 , n63429 , n63430 , n63431 , n63432 , n63433 , n63434 , n63435 , n63436 , 
     n63437 , n63438 , n63439 , n63440 , n63441 , n63442 , n63443 , n63444 , n63445 , n63446 , 
     n63447 , n63448 , n63449 , n63450 , n63451 , n63452 , n63453 , n63454 , n63455 , n63456 , 
     n63457 , n63458 , n63459 , n63460 , n63461 , n63462 , n63463 , n63464 , n63465 , n63466 , 
     n63467 , n63468 , n63469 , n63470 , n63471 , n63472 , n63473 , n63474 , n63475 , n63476 , 
     n63477 , n63478 , n63479 , n63480 , n63481 , n63482 , n63483 , n63484 , n63485 , n63486 , 
     n63487 , n63488 , n63489 , n63490 , n63491 , n63492 , n63493 , n63494 , n63495 , n63496 , 
     n63497 , n63498 , n63499 , n63500 , n63501 , n63502 , n63503 , n63504 , n63505 , n63506 , 
     n63507 , n63508 , n63509 , n63510 , n63511 , n63512 , n63513 , n63514 , n63515 , n63516 , 
     n63517 , n63518 , n63519 , n63520 , n63521 , n63522 , n63523 , n63524 , n63525 , n63526 , 
     n63527 , n63528 , n63529 , n63530 , n63531 , n63532 , n63533 , n63534 , n63535 , n63536 , 
     n63537 , n63538 , n63539 , n63540 , n63541 , n63542 , n63543 , n63544 , n63545 , n63546 , 
     n63547 , n63548 , n63549 , n63550 , n63551 , n63552 , n63553 , n63554 , n63555 , n63556 , 
     n63557 , n63558 , n63559 , n63560 , n63561 , n63562 , n63563 , n63564 , n63565 , n63566 , 
     n63567 , n63568 , n63569 , n63570 , n63571 , n63572 , n63573 , n63574 , n63575 , n63576 , 
     n63577 , n63578 , n63579 , n63580 , n63581 , n63582 , n63583 , n63584 , n63585 , n63586 , 
     n63587 , n63588 , n63589 , n63590 , n63591 , n63592 , n63593 , n63594 , n63595 , n63596 , 
     n63597 , n63598 , n63599 , n63600 , n63601 , n63602 , n63603 , n63604 , n63605 , n63606 , 
     n63607 , n63608 , n63609 , n63610 , n63611 , n63612 , n63613 , n63614 , n63615 , n63616 , 
     n63617 , n63618 , n63619 , n63620 , n63621 , n63622 , n63623 , n63624 , n63625 , n63626 , 
     n63627 , n63628 , n63629 , n63630 , n63631 , n63632 , n63633 , n63634 , n63635 , n63636 , 
     n63637 , n63638 , n63639 , n63640 , n63641 , n63642 , n63643 , n63644 , n63645 , n63646 , 
     n63647 , n63648 , n63649 , n63650 , n63651 , n63652 , n63653 , n63654 , n63655 , n63656 , 
     n63657 , n63658 , n63659 , n63660 , n63661 , n63662 , n63663 , n63664 , n63665 , n63666 , 
     n63667 , n63668 , n63669 , n63670 , n63671 , n63672 , n63673 , n63674 , n63675 , n63676 , 
     n63677 , n63678 , n63679 , n63680 , n63681 , n63682 , n63683 , n63684 , n63685 , n63686 , 
     n63687 , n63688 , n63689 , n63690 , n63691 , n63692 , n63693 , n63694 , n63695 , n63696 , 
     n63697 , n63698 , n63699 , n63700 , n63701 , n63702 , n63703 , n63704 , n63705 , n63706 , 
     n63707 , n63708 , n63709 , n63710 , n63711 , n63712 , n63713 , n63714 , n63715 , n63716 , 
     n63717 , n63718 , n63719 , n63720 , n63721 , n63722 , n63723 , n63724 , n63725 , n63726 , 
     n63727 , n63728 , n63729 , n63730 , n63731 , n63732 , n63733 , n63734 , n63735 , n63736 , 
     n63737 , n63738 , n63739 , n63740 , n63741 , n63742 , n63743 , n63744 , n63745 , n63746 , 
     n63747 , n63748 , n63749 , n63750 , n63751 , n63752 , n63753 , n63754 , n63755 , n63756 , 
     n63757 , n63758 , n63759 , n63760 , n63761 , n63762 , n63763 , n63764 , n63765 , n63766 , 
     n63767 , n63768 , n63769 , n63770 , n63771 , n63772 , n63773 , n63774 , n63775 , n63776 , 
     n63777 , n63778 , n63779 , n63780 , n63781 , n63782 , n63783 , n63784 , n63785 , n63786 , 
     n63787 , n63788 , n63789 , n63790 , n63791 , n63792 , n63793 , n63794 , n63795 , n63796 , 
     n63797 , n63798 , n63799 , n63800 , n63801 , n63802 , n63803 , n63804 , n63805 , n63806 , 
     n63807 , n63808 , n63809 , n63810 , n63811 , n63812 , n63813 , n63814 , n63815 , n63816 , 
     n63817 , n63818 , n63819 , n63820 , n63821 , n63822 , n63823 , n63824 , n63825 , n63826 , 
     n63827 , n63828 , n63829 , n63830 , n63831 , n63832 , n63833 , n63834 , n63835 , n63836 , 
     n63837 , n63838 , n63839 , n63840 , n63841 , n63842 , n63843 , n63844 , n63845 , n63846 , 
     n63847 , n63848 , n63849 , n63850 , n63851 , n63852 , n63853 , n63854 , n63855 , n63856 , 
     n63857 , n63858 , n63859 , n63860 , n63861 , n63862 , n63863 , n63864 , n63865 , n63866 , 
     n63867 , n63868 , n63869 , n63870 , n63871 , n63872 , n63873 , n63874 , n63875 , n63876 , 
     n63877 , n63878 , n63879 , n63880 , n63881 , n63882 , n63883 , n63884 , n63885 , n63886 , 
     n63887 , n63888 , n63889 , n63890 , n63891 , n63892 , n63893 , n63894 , n63895 , n63896 , 
     n63897 , n63898 , n63899 , n63900 , n63901 , n63902 , n63903 , n63904 , n63905 , n63906 , 
     n63907 , n63908 , n63909 , n63910 , n63911 , n63912 , n63913 , n63914 , n63915 , n63916 , 
     n63917 , n63918 , n63919 , n63920 , n63921 , n63922 , n63923 , n63924 , n63925 , n63926 , 
     n63927 , n63928 , n63929 , n63930 , n63931 , n63932 , n63933 , n63934 , n63935 , n63936 , 
     n63937 , n63938 , n63939 , n63940 , n63941 , n63942 , n63943 , n63944 , n63945 , n63946 , 
     n63947 , n63948 , n63949 , n63950 , n63951 , n63952 , n63953 , n63954 , n63955 , n63956 , 
     n63957 , n63958 , n63959 , n63960 , n63961 , n63962 , n63963 , n63964 , n63965 , n63966 , 
     n63967 , n63968 , n63969 , n63970 , n63971 , n63972 , n63973 , n63974 , n63975 , n63976 , 
     n63977 , n63978 , n63979 , n63980 , n63981 , n63982 , n63983 , n63984 , n63985 , n63986 , 
     n63987 , n63988 , n63989 , n63990 , n63991 , n63992 , n63993 , n63994 , n63995 , n63996 , 
     n63997 , n63998 , n63999 , n64000 , n64001 , n64002 , n64003 , n64004 , n64005 , n64006 , 
     n64007 , n64008 , n64009 , n64010 , n64011 , n64012 , n64013 , n64014 , n64015 , n64016 , 
     n64017 , n64018 , n64019 , n64020 , n64021 , n64022 , n64023 , n64024 , n64025 , n64026 , 
     n64027 , n64028 , n64029 , n64030 , n64031 , n64032 , n64033 , n64034 , n64035 , n64036 , 
     n64037 , n64038 , n64039 , n64040 , n64041 , n64042 , n64043 , n64044 , n64045 , n64046 , 
     n64047 , n64048 , n64049 , n64050 , n64051 , n64052 , n64053 , n64054 , n64055 , n64056 , 
     n64057 , n64058 , n64059 , n64060 , n64061 , n64062 , n64063 , n64064 , n64065 , n64066 , 
     n64067 , n64068 , n64069 , n64070 , n64071 , n64072 , n64073 , n64074 , n64075 , n64076 , 
     n64077 , n64078 , n64079 , n64080 , n64081 , n64082 , n64083 , n64084 , n64085 , n64086 , 
     n64087 , n64088 , n64089 , n64090 , n64091 , n64092 , n64093 , n64094 , n64095 , n64096 , 
     n64097 , n64098 , n64099 , n64100 , n64101 , n64102 , n64103 , n64104 , n64105 , n64106 , 
     n64107 , n64108 , n64109 , n64110 , n64111 , n64112 , n64113 , n64114 , n64115 , n64116 , 
     n64117 , n64118 , n64119 , n64120 , n64121 , n64122 , n64123 , n64124 , n64125 , n64126 , 
     n64127 , n64128 , n64129 , n64130 , n64131 , n64132 , n64133 , n64134 , n64135 , n64136 , 
     n64137 , n64138 , n64139 , n64140 , n64141 , n64142 , n64143 , n64144 , n64145 , n64146 , 
     n64147 , n64148 , n64149 , n64150 , n64151 , n64152 , n64153 , n64154 , n64155 , n64156 , 
     n64157 , n64158 , n64159 , n64160 , n64161 , n64162 , n64163 , n64164 , n64165 , n64166 , 
     n64167 , n64168 , n64169 , n64170 , n64171 , n64172 , n64173 , n64174 , n64175 , n64176 , 
     n64177 , n64178 , n64179 , n64180 , n64181 , n64182 , n64183 , n64184 , n64185 , n64186 , 
     n64187 , n64188 , n64189 , n64190 , n64191 , n64192 , n64193 , n64194 , n64195 , n64196 , 
     n64197 , n64198 , n64199 , n64200 , n64201 , n64202 , n64203 , n64204 , n64205 , n64206 , 
     n64207 , n64208 , n64209 , n64210 , n64211 , n64212 , n64213 , n64214 , n64215 , n64216 , 
     n64217 , n64218 , n64219 , n64220 , n64221 , n64222 , n64223 , n64224 , n64225 , n64226 , 
     n64227 , n64228 , n64229 , n64230 , n64231 , n64232 , n64233 , n64234 , n64235 , n64236 , 
     n64237 , n64238 , n64239 , n64240 , n64241 , n64242 , n64243 , n64244 , n64245 , n64246 , 
     n64247 , n64248 , n64249 , n64250 , n64251 , n64252 , n64253 , n64254 , n64255 , n64256 , 
     n64257 , n64258 , n64259 , n64260 , n64261 , n64262 , n64263 , n64264 , n64265 , n64266 , 
     n64267 , n64268 , n64269 , n64270 , n64271 , n64272 , n64273 , n64274 , n64275 , n64276 , 
     n64277 , n64278 , n64279 , n64280 , n64281 , n64282 , n64283 , n64284 , n64285 , n64286 , 
     n64287 , n64288 , n64289 , n64290 , n64291 , n64292 , n64293 , n64294 , n64295 , n64296 , 
     n64297 , n64298 , n64299 , n64300 , n64301 , n64302 , n64303 , n64304 , n64305 , n64306 , 
     n64307 , n64308 , n64309 , n64310 , n64311 , n64312 , n64313 , n64314 , n64315 , n64316 , 
     n64317 , n64318 , n64319 , n64320 , n64321 , n64322 , n64323 , n64324 , n64325 , n64326 , 
     n64327 , n64328 , n64329 , n64330 , n64331 , n64332 , n64333 , n64334 , n64335 , n64336 , 
     n64337 , n64338 , n64339 , n64340 , n64341 , n64342 , n64343 , n64344 , n64345 , n64346 , 
     n64347 , n64348 , n64349 , n64350 , n64351 , n64352 , n64353 , n64354 , n64355 , n64356 , 
     n64357 , n64358 , n64359 , n64360 , n64361 , n64362 , n64363 , n64364 , n64365 , n64366 , 
     n64367 , n64368 , n64369 , n64370 , n64371 , n64372 , n64373 , n64374 , n64375 , n64376 , 
     n64377 , n64378 , n64379 , n64380 , n64381 , n64382 , n64383 , n64384 , n64385 , n64386 , 
     n64387 , n64388 , n64389 , n64390 , n64391 , n64392 , n64393 , n64394 , n64395 , n64396 , 
     n64397 , n64398 , n64399 , n64400 , n64401 , n64402 , n64403 , n64404 , n64405 , n64406 , 
     n64407 , n64408 , n64409 , n64410 , n64411 , n64412 , n64413 , n64414 , n64415 , n64416 , 
     n64417 , n64418 , n64419 , n64420 , n64421 , n64422 , n64423 , n64424 , n64425 , n64426 , 
     n64427 , n64428 , n64429 , n64430 , n64431 , n64432 , n64433 , n64434 , n64435 , n64436 , 
     n64437 , n64438 , n64439 , n64440 , n64441 , n64442 , n64443 , n64444 , n64445 , n64446 , 
     n64447 , n64448 , n64449 , n64450 , n64451 , n64452 , n64453 , n64454 , n64455 , n64456 , 
     n64457 , n64458 , n64459 , n64460 , n64461 , n64462 , n64463 , n64464 , n64465 , n64466 , 
     n64467 , n64468 , n64469 , n64470 , n64471 , n64472 , n64473 , n64474 , n64475 , n64476 , 
     n64477 , n64478 , n64479 , n64480 , n64481 , n64482 , n64483 , n64484 , n64485 , n64486 , 
     n64487 , n64488 , n64489 , n64490 , n64491 , n64492 , n64493 , n64494 , n64495 , n64496 , 
     n64497 , n64498 , n64499 , n64500 , n64501 , n64502 , n64503 , n64504 , n64505 , n64506 , 
     n64507 , n64508 , n64509 , n64510 , n64511 , n64512 , n64513 , n64514 , n64515 , n64516 , 
     n64517 , n64518 , n64519 , n64520 , n64521 , n64522 , n64523 , n64524 , n64525 , n64526 , 
     n64527 , n64528 , n64529 , n64530 , n64531 , n64532 , n64533 , n64534 , n64535 , n64536 , 
     n64537 , n64538 , n64539 , n64540 , n64541 , n64542 , n64543 , n64544 , n64545 , n64546 , 
     n64547 , n64548 , n64549 , n64550 , n64551 , n64552 , n64553 , n64554 , n64555 , n64556 , 
     n64557 , n64558 , n64559 , n64560 , n64561 , n64562 , n64563 , n64564 , n64565 , n64566 , 
     n64567 , n64568 , n64569 , n64570 , n64571 , n64572 , n64573 , n64574 , n64575 , n64576 , 
     n64577 , n64578 , n64579 , n64580 , n64581 , n64582 , n64583 , n64584 , n64585 , n64586 , 
     n64587 , n64588 , n64589 , n64590 , n64591 , n64592 , n64593 , n64594 , n64595 , n64596 , 
     n64597 , n64598 , n64599 , n64600 , n64601 , n64602 , n64603 , n64604 , n64605 , n64606 , 
     n64607 , n64608 , n64609 , n64610 , n64611 , n64612 , n64613 , n64614 , n64615 , n64616 , 
     n64617 , n64618 , n64619 , n64620 , n64621 , n64622 , n64623 , n64624 , n64625 , n64626 , 
     n64627 , n64628 , n64629 , n64630 , n64631 , n64632 , n64633 , n64634 , n64635 , n64636 , 
     n64637 , n64638 , n64639 , n64640 , n64641 , n64642 , n64643 , n64644 , n64645 , n64646 , 
     n64647 , n64648 , n64649 , n64650 , n64651 , n64652 , n64653 , n64654 , n64655 , n64656 , 
     n64657 , n64658 , n64659 , n64660 , n64661 , n64662 , n64663 , n64664 , n64665 , n64666 , 
     n64667 , n64668 , n64669 , n64670 , n64671 , n64672 , n64673 , n64674 , n64675 , n64676 , 
     n64677 , n64678 , n64679 , n64680 , n64681 , n64682 , n64683 , n64684 , n64685 , n64686 , 
     n64687 , n64688 , n64689 , n64690 , n64691 , n64692 , n64693 , n64694 , n64695 , n64696 , 
     n64697 , n64698 , n64699 , n64700 , n64701 , n64702 , n64703 , n64704 , n64705 , n64706 , 
     n64707 , n64708 , n64709 , n64710 , n64711 , n64712 , n64713 , n64714 , n64715 , n64716 , 
     n64717 , n64718 , n64719 , n64720 , n64721 , n64722 , n64723 , n64724 , n64725 , n64726 , 
     n64727 , n64728 , n64729 , n64730 , n64731 , n64732 , n64733 , n64734 , n64735 , n64736 , 
     n64737 , n64738 , n64739 , n64740 , n64741 , n64742 , n64743 , n64744 , n64745 , n64746 , 
     n64747 , n64748 , n64749 , n64750 , n64751 , n64752 , n64753 , n64754 , n64755 , n64756 , 
     n64757 , n64758 , n64759 , n64760 , n64761 , n64762 , n64763 , n64764 , n64765 , n64766 , 
     n64767 , n64768 , n64769 , n64770 , n64771 , n64772 , n64773 , n64774 , n64775 , n64776 , 
     n64777 , n64778 , n64779 , n64780 , n64781 , n64782 , n64783 , n64784 , n64785 , n64786 , 
     n64787 , n64788 , n64789 , n64790 , n64791 , n64792 , n64793 , n64794 , n64795 , n64796 , 
     n64797 , n64798 , n64799 , n64800 , n64801 , n64802 , n64803 , n64804 , n64805 , n64806 , 
     n64807 , n64808 , n64809 , n64810 , n64811 , n64812 , n64813 , n64814 , n64815 , n64816 , 
     n64817 , n64818 , n64819 , n64820 , n64821 , n64822 , n64823 , n64824 , n64825 , n64826 , 
     n64827 , n64828 , n64829 , n64830 , n64831 , n64832 , n64833 , n64834 , n64835 , n64836 , 
     n64837 , n64838 , n64839 , n64840 , n64841 , n64842 , n64843 , n64844 , n64845 , n64846 , 
     n64847 , n64848 , n64849 , n64850 , n64851 , n64852 , n64853 , n64854 , n64855 , n64856 , 
     n64857 , n64858 , n64859 , n64860 , n64861 , n64862 , n64863 , n64864 , n64865 , n64866 , 
     n64867 , n64868 , n64869 , n64870 , n64871 , n64872 , n64873 , n64874 , n64875 , n64876 , 
     n64877 , n64878 , n64879 , n64880 , n64881 , n64882 , n64883 , n64884 , n64885 , n64886 , 
     n64887 , n64888 , n64889 , n64890 , n64891 , n64892 , n64893 , n64894 , n64895 , n64896 , 
     n64897 , n64898 ;
buf ( RI21a19c60_2 , n0 );
buf ( RI21a5daf0_1 , n1 );
buf ( RI2107e620_463 , n2 );
buf ( RI21a139f0_68 , n3 );
buf ( RI21084368_418 , n4 );
buf ( RI21079850_497 , n5 );
buf ( RI21a12820_78 , n6 );
buf ( RI210beb08_292 , n7 );
buf ( RI21a12898_77 , n8 );
buf ( RI210beb80_291 , n9 );
buf ( RI21a12910_76 , n10 );
buf ( RI210bf3f0_290 , n11 );
buf ( RI21a12988_75 , n12 );
buf ( RI210bf468_289 , n13 );
buf ( RI21a13090_74 , n14 );
buf ( RI210bf4e0_288 , n15 );
buf ( RI21a13108_73 , n16 );
buf ( RI210bf558_287 , n17 );
buf ( RI21a13180_72 , n18 );
buf ( RI210bfdc8_286 , n19 );
buf ( RI21a131f8_71 , n20 );
buf ( RI210bfe40_285 , n21 );
buf ( RI21a13270_70 , n22 );
buf ( RI210bfeb8_284 , n23 );
buf ( RI21a132e8_69 , n24 );
buf ( RI210bff30_283 , n25 );
buf ( RI21a116c8_87 , n26 );
buf ( RI210bd6e0_301 , n27 );
buf ( RI21a11dd0_86 , n28 );
buf ( RI210bd758_300 , n29 );
buf ( RI21a11e48_85 , n30 );
buf ( RI210bd7d0_299 , n31 );
buf ( RI21a11ec0_84 , n32 );
buf ( RI210be040_298 , n33 );
buf ( RI21a11f38_83 , n34 );
buf ( RI210be0b8_297 , n35 );
buf ( RI21a11fb0_82 , n36 );
buf ( RI210be130_296 , n37 );
buf ( RI21a12028_81 , n38 );
buf ( RI210be1a8_295 , n39 );
buf ( RI21a12730_80 , n40 );
buf ( RI210bea18_294 , n41 );
buf ( RI21a127a8_79 , n42 );
buf ( RI210bea90_293 , n43 );
buf ( RI21077f00_507 , n44 );
buf ( RI21077f78_506 , n45 );
buf ( RI21078a40_505 , n46 );
buf ( RI21078ab8_504 , n47 );
buf ( RI21078b30_503 , n48 );
buf ( RI21078ba8_502 , n49 );
buf ( RI21078c20_501 , n50 );
buf ( RI21078c98_500 , n51 );
buf ( RI21079760_499 , n52 );
buf ( RI210797d8_498 , n53 );
buf ( RI21077078_516 , n54 );
buf ( RI210770f0_515 , n55 );
buf ( RI21077168_514 , n56 );
buf ( RI210771e0_513 , n57 );
buf ( RI21077258_512 , n58 );
buf ( RI21077d20_511 , n59 );
buf ( RI21077d98_510 , n60 );
buf ( RI21077e10_509 , n61 );
buf ( RI21077e88_508 , n62 );
buf ( RI2107a660_489 , n63 );
buf ( RI2107a6d8_488 , n64 );
buf ( RI2107b218_486 , n65 );
buf ( RI2107b290_485 , n66 );
buf ( RI2107b308_484 , n67 );
buf ( RI2107b380_483 , n68 );
buf ( RI2107b3f8_482 , n69 );
buf ( RI2107bec0_481 , n70 );
buf ( RI2107bf38_480 , n71 );
buf ( RI2107bfb0_479 , n72 );
buf ( RI2107c028_478 , n73 );
buf ( RI2107c0a0_477 , n74 );
buf ( RI2107cbe0_475 , n75 );
buf ( RI2107cc58_474 , n76 );
buf ( RI2107ccd0_473 , n77 );
buf ( RI2107cd48_472 , n78 );
buf ( RI2107cdc0_471 , n79 );
buf ( RI2107ce38_470 , n80 );
buf ( RI2107d900_469 , n81 );
buf ( RI2107d978_468 , n82 );
buf ( RI2107d9f0_467 , n83 );
buf ( RI2107da68_466 , n84 );
buf ( RI210798c8_496 , n85 );
buf ( RI21079940_495 , n86 );
buf ( RI210799b8_494 , n87 );
buf ( RI2107a480_493 , n88 );
buf ( RI2107a4f8_492 , n89 );
buf ( RI2107a570_491 , n90 );
buf ( RI2107a5e8_490 , n91 );
buf ( RI2107b1a0_487 , n92 );
buf ( RI2107c118_476 , n93 );
buf ( RI2106bde0_608 , n94 );
buf ( GI20478f00_682 , n95 );
buf ( RI2106c0b0_602 , n96 );
buf ( RI2106c128_601 , n97 );
buf ( RI2106c1a0_600 , n98 );
buf ( RI2106c218_599 , n99 );
buf ( RI2106c290_598 , n100 );
buf ( RI2106a238_641 , n101 );
buf ( RI2106a2b0_640 , n102 );
buf ( RI2106a328_639 , n103 );
buf ( RI2106a3a0_638 , n104 );
buf ( RI2106a490_636 , n105 );
buf ( RI2106a508_635 , n106 );
buf ( RI2106a580_634 , n107 );
buf ( RI2106c308_597 , n108 );
buf ( RI2106a5f8_633 , n109 );
buf ( RI2106a670_632 , n110 );
buf ( RI2106a6e8_631 , n111 );
buf ( RI2106a760_630 , n112 );
buf ( RI2106a7d8_629 , n113 );
buf ( RI2106ae68_628 , n114 );
buf ( RI21069a40_645 , n115 );
buf ( RI2106bed0_606 , n116 );
buf ( RI21069ab8_644 , n117 );
buf ( RI2106bf48_605 , n118 );
buf ( RI2106bfc0_604 , n119 );
buf ( RI2106c038_603 , n120 );
buf ( RI2106a148_643 , n121 );
buf ( RI2106a1c0_642 , n122 );
buf ( RI2106a418_637 , n123 );
buf ( RI2106c380_596 , n124 );
buf ( RI2106cbf0_591 , n125 );
buf ( RI2106dd48_567 , n126 );
buf ( RI21073040_543 , n127 );
buf ( RI2106cd58_588 , n128 );
buf ( RI2106deb0_564 , n129 );
buf ( RI21073c70_539 , n130 );
buf ( RI2106cdd0_587 , n131 );
buf ( RI2106df28_563 , n132 );
buf ( RI21073ce8_538 , n133 );
buf ( RI2106ce48_586 , n134 );
buf ( RI2106dfa0_562 , n135 );
buf ( RI21073d60_537 , n136 );
buf ( RI2106cec0_585 , n137 );
buf ( RI2106e018_561 , n138 );
buf ( RI21073dd8_536 , n139 );
buf ( RI2106cf38_584 , n140 );
buf ( RI2106e090_560 , n141 );
buf ( RI210748a0_535 , n142 );
buf ( RI2106cfb0_583 , n143 );
buf ( RI2106e108_559 , n144 );
buf ( RI21074918_534 , n145 );
buf ( RI2106d028_582 , n146 );
buf ( RI21070a48_558 , n147 );
buf ( RI21074990_533 , n148 );
buf ( RI2106d0a0_581 , n149 );
buf ( RI21070ac0_557 , n150 );
buf ( RI21074a08_532 , n151 );
buf ( RI2106d118_580 , n152 );
buf ( RI21071588_556 , n153 );
buf ( RI21074a80_531 , n154 );
buf ( RI2106b138_622 , n155 );
buf ( RI2106b4f8_614 , n156 );
buf ( RI210755c0_529 , n157 );
buf ( RI2106b1b0_621 , n158 );
buf ( RI2106b570_613 , n159 );
buf ( RI21075638_528 , n160 );
buf ( RI2106b228_620 , n161 );
buf ( RI2106bc00_612 , n162 );
buf ( RI210756b0_527 , n163 );
buf ( RI2106d190_579 , n164 );
buf ( RI21071600_555 , n165 );
buf ( RI21075728_526 , n166 );
buf ( RI2106d208_578 , n167 );
buf ( RI21071678_554 , n168 );
buf ( RI210757a0_525 , n169 );
buf ( RI2106d898_577 , n170 );
buf ( RI2106bc78_611 , n171 );
buf ( RI21075818_524 , n172 );
buf ( RI2106d910_576 , n173 );
buf ( RI2106bcf0_610 , n174 );
buf ( RI210762e0_523 , n175 );
buf ( RI2106d988_575 , n176 );
buf ( RI210716f0_553 , n177 );
buf ( RI21076358_522 , n178 );
buf ( RI2106da00_574 , n179 );
buf ( RI210721b8_552 , n180 );
buf ( RI210763d0_521 , n181 );
buf ( RI2106da78_573 , n182 );
buf ( RI2106bd68_609 , n183 );
buf ( RI21076448_520 , n184 );
buf ( RI2106ca10_595 , n185 );
buf ( RI2106db68_571 , n186 );
buf ( RI210722a8_550 , n187 );
buf ( RI2106ca88_594 , n188 );
buf ( RI2106dbe0_570 , n189 );
buf ( RI21072320_549 , n190 );
buf ( RI2106aee0_627 , n191 );
buf ( RI2106dc58_569 , n192 );
buf ( RI21072398_548 , n193 );
buf ( RI2106af58_626 , n194 );
buf ( RI2106dcd0_568 , n195 );
buf ( RI21072e60_547 , n196 );
buf ( RI2106cb00_593 , n197 );
buf ( RI2106b2a0_619 , n198 );
buf ( RI21072ed8_546 , n199 );
buf ( RI2106afd0_625 , n200 );
buf ( RI2106b318_618 , n201 );
buf ( RI21072f50_545 , n202 );
buf ( RI2106cb78_592 , n203 );
buf ( RI2106b390_617 , n204 );
buf ( RI21072fc8_544 , n205 );
buf ( RI2106b048_624 , n206 );
buf ( RI2106b408_616 , n207 );
buf ( RI21073b80_541 , n208 );
buf ( RI2106b0c0_623 , n209 );
buf ( RI2106b480_615 , n210 );
buf ( RI21074af8_530 , n211 );
buf ( RI2106daf0_572 , n212 );
buf ( RI21072230_551 , n213 );
buf ( RI210764c0_519 , n214 );
buf ( RI2107dae0_465 , n215 );
buf ( RI2106cc68_590 , n216 );
buf ( RI2106ddc0_566 , n217 );
buf ( RI210730b8_542 , n218 );
buf ( RI21a0e608_121 , n219 );
buf ( RI210b87a8_334 , n220 );
buf ( RI21a19a08_3 , n221 );
buf ( RI21a0f058_113 , n222 );
buf ( RI210b9b58_326 , n223 );
buf ( RI21a0f0d0_112 , n224 );
buf ( RI210b9bd0_325 , n225 );
buf ( RI21a0f850_110 , n226 );
buf ( RI210b9c48_324 , n227 );
buf ( RI21a0f8c8_109 , n228 );
buf ( RI210b9cc0_323 , n229 );
buf ( RI21a0f940_108 , n230 );
buf ( RI210ba530_322 , n231 );
buf ( RI21a0f9b8_107 , n232 );
buf ( RI210ba5a8_321 , n233 );
buf ( RI21a0fa30_106 , n234 );
buf ( RI210ba620_320 , n235 );
buf ( RI21a0faa8_105 , n236 );
buf ( RI210ba698_319 , n237 );
buf ( RI21a101b0_104 , n238 );
buf ( RI210baf08_318 , n239 );
buf ( RI21a10228_103 , n240 );
buf ( RI210baf80_317 , n241 );
buf ( RI21a102a0_102 , n242 );
buf ( RI210baff8_316 , n243 );
buf ( RI21a10318_101 , n244 );
buf ( RI210bb070_315 , n245 );
buf ( RI21a10390_100 , n246 );
buf ( RI210bb8e0_314 , n247 );
buf ( RI21a10408_99 , n248 );
buf ( RI210bb958_313 , n249 );
buf ( RI21a10b10_98 , n250 );
buf ( RI210bb9d0_312 , n251 );
buf ( RI21a10b88_97 , n252 );
buf ( RI210bba48_311 , n253 );
buf ( RI21a10c00_96 , n254 );
buf ( RI210bc2b8_310 , n255 );
buf ( RI21a10c78_95 , n256 );
buf ( RI210bc330_309 , n257 );
buf ( RI21a10cf0_94 , n258 );
buf ( RI210bc3a8_308 , n259 );
buf ( RI21a10d68_93 , n260 );
buf ( RI210bc420_307 , n261 );
buf ( RI21a11470_92 , n262 );
buf ( RI210bcc90_306 , n263 );
buf ( RI21a114e8_91 , n264 );
buf ( RI210bcd08_305 , n265 );
buf ( RI21a0e680_120 , n266 );
buf ( RI210b8820_333 , n267 );
buf ( RI21a0e6f8_119 , n268 );
buf ( RI210b8898_332 , n269 );
buf ( RI21a0e770_118 , n270 );
buf ( RI210b8910_331 , n271 );
buf ( RI21a0e7e8_117 , n272 );
buf ( RI210b9180_330 , n273 );
buf ( RI21a0eef0_116 , n274 );
buf ( RI210b91f8_329 , n275 );
buf ( RI21a0ef68_115 , n276 );
buf ( RI210b9270_328 , n277 );
buf ( RI21a0efe0_114 , n278 );
buf ( RI210b92e8_327 , n279 );
buf ( RI21a0f148_111 , n280 );
buf ( RI21084278_420 , n281 );
buf ( RI210cfcc8_237 , n282 );
buf ( RI210842f0_419 , n283 );
buf ( RI21a11560_90 , n284 );
buf ( RI210bcd80_304 , n285 );
buf ( RI21a19990_4 , n286 );
buf ( RI2106cce0_589 , n287 );
buf ( RI2106de38_565 , n288 );
buf ( RI21073bf8_540 , n289 );
buf ( RI21a19918_5 , n290 );
buf ( RI21a198a0_6 , n291 );
buf ( RI21a19828_7 , n292 );
buf ( RI21a197b0_8 , n293 );
buf ( RI21a190a8_9 , n294 );
buf ( RI21a19030_10 , n295 );
buf ( RI21a18fb8_11 , n296 );
buf ( RI21a18f40_12 , n297 );
buf ( RI21a18ec8_13 , n298 );
buf ( RI21a18e50_14 , n299 );
buf ( RI21a18748_15 , n300 );
buf ( RI21a186d0_16 , n301 );
buf ( RI21a18658_17 , n302 );
buf ( RI21a185e0_18 , n303 );
buf ( RI21a18568_19 , n304 );
buf ( RI21a184f0_20 , n305 );
buf ( RI21a17de8_21 , n306 );
buf ( RI21a17d70_22 , n307 );
buf ( RI21a17cf8_23 , n308 );
buf ( RI21a17c80_24 , n309 );
buf ( RI21a17c08_25 , n310 );
buf ( RI21a17b90_26 , n311 );
buf ( RI21a17488_27 , n312 );
buf ( RI21a17410_28 , n313 );
buf ( RI21a17398_29 , n314 );
buf ( RI21a17320_30 , n315 );
buf ( RI21a172a8_31 , n316 );
buf ( RI21a17230_32 , n317 );
buf ( RI21a16b28_33 , n318 );
buf ( RI21a16ab0_34 , n319 );
buf ( RI2106be58_607 , n320 );
buf ( RI21a14440_60 , n321 );
buf ( RI21a144b8_59 , n322 );
buf ( RI21a145a8_57 , n323 );
buf ( RI21a14cb0_56 , n324 );
buf ( RI21a14d28_55 , n325 );
buf ( RI21a14da0_54 , n326 );
buf ( RI21a14e18_53 , n327 );
buf ( RI21a14e90_52 , n328 );
buf ( RI21a14f08_51 , n329 );
buf ( RI21a15610_50 , n330 );
buf ( RI21a15688_49 , n331 );
buf ( RI21a15700_48 , n332 );
buf ( RI21a157f0_46 , n333 );
buf ( RI21a15868_45 , n334 );
buf ( RI21a15f70_44 , n335 );
buf ( RI21a15fe8_43 , n336 );
buf ( RI21a16060_42 , n337 );
buf ( RI21a160d8_41 , n338 );
buf ( RI21a16150_40 , n339 );
buf ( RI21a161c8_39 , n340 );
buf ( RI21a168d0_38 , n341 );
buf ( RI21a16948_37 , n342 );
buf ( RI21a13a68_67 , n343 );
buf ( RI21a13ae0_66 , n344 );
buf ( RI21a13b58_65 , n345 );
buf ( RI21a13bd0_64 , n346 );
buf ( RI21a13c48_63 , n347 );
buf ( RI21a14350_62 , n348 );
buf ( RI21a143c8_61 , n349 );
buf ( RI21a14530_58 , n350 );
buf ( RI21a15778_47 , n351 );
buf ( RI21a169c0_36 , n352 );
buf ( RI210d6910_193 , n353 );
buf ( RI210cdfb8_248 , n354 );
buf ( GI2046a680_186 , n355 );
buf ( RI210d2d88_218 , n356 );
buf ( RI210d10f0_228 , n357 );
buf ( RI210d1078_229 , n358 );
buf ( RI210d1000_230 , n359 );
buf ( RI210d0790_231 , n360 );
buf ( RI210d0718_232 , n361 );
buf ( RI210d06a0_233 , n362 );
buf ( RI210d0628_234 , n363 );
buf ( RI210cfdb8_235 , n364 );
buf ( RI210d4228_208 , n365 );
buf ( RI210d41b0_209 , n366 );
buf ( RI210d4138_210 , n367 );
buf ( RI210d38c8_211 , n368 );
buf ( RI210d3850_212 , n369 );
buf ( RI210d37d8_213 , n370 );
buf ( RI210d3760_214 , n371 );
buf ( RI210d2ef0_215 , n372 );
buf ( RI210d2e78_216 , n373 );
buf ( RI210d2e00_217 , n374 );
buf ( RI210d2518_219 , n375 );
buf ( RI210d24a0_220 , n376 );
buf ( RI210d2428_221 , n377 );
buf ( RI210d23b0_222 , n378 );
buf ( RI210d1b40_223 , n379 );
buf ( RI210d1ac8_224 , n380 );
buf ( RI210d1a50_225 , n381 );
buf ( RI210d19d8_226 , n382 );
buf ( RI210d1168_227 , n383 );
buf ( RI210d8ff8_178 , n384 );
buf ( RI21a0b7a0_150 , n385 );
buf ( RI21a0e590_122 , n386 );
buf ( RI210d55d8_200 , n387 );
buf ( RI210da3a8_170 , n388 );
buf ( RI21a0c178_143 , n389 );
buf ( RI210d73d8_187 , n390 );
buf ( RI21a0a6c0_158 , n391 );
buf ( RI21a0d438_131 , n392 );
buf ( RI210d5ec0_198 , n393 );
buf ( RI210da498_168 , n394 );
buf ( RI21a0c268_141 , n395 );
buf ( RI210d5560_201 , n396 );
buf ( RI210d9b38_171 , n397 );
buf ( RI21a0c100_144 , n398 );
buf ( RI210d54e8_202 , n399 );
buf ( RI210d9ac0_172 , n400 );
buf ( RI210cf2f0_241 , n401 );
buf ( RI210d4c78_203 , n402 );
buf ( RI210d9a48_173 , n403 );
buf ( RI21a0c088_145 , n404 );
buf ( RI210d4c00_204 , n405 );
buf ( RI210d99d0_174 , n406 );
buf ( RI21a0c010_146 , n407 );
buf ( RI210d4b88_205 , n408 );
buf ( RI210d9160_175 , n409 );
buf ( RI21a0b908_147 , n410 );
buf ( RI210d4b10_206 , n411 );
buf ( RI210d90e8_176 , n412 );
buf ( RI21a0b890_148 , n413 );
buf ( RI210d42a0_207 , n414 );
buf ( RI210d9070_177 , n415 );
buf ( RI21a0b818_149 , n416 );
buf ( RI210d8788_179 , n417 );
buf ( RI21a0b728_151 , n418 );
buf ( RI21a0de88_123 , n419 );
buf ( RI210d8710_180 , n420 );
buf ( RI21a0b6b0_152 , n421 );
buf ( RI21a0de10_124 , n422 );
buf ( RI210d8698_181 , n423 );
buf ( RI21a0afa8_153 , n424 );
buf ( RI21a0dd98_125 , n425 );
buf ( RI210d8620_182 , n426 );
buf ( RI21a0af30_154 , n427 );
buf ( RI21a0dd20_126 , n428 );
buf ( RI210d7db0_183 , n429 );
buf ( RI21a0aeb8_155 , n430 );
buf ( RI21a0dca8_127 , n431 );
buf ( RI210d7d38_184 , n432 );
buf ( RI21a0ae40_156 , n433 );
buf ( RI21a0dc30_128 , n434 );
buf ( RI210ce8a0_246 , n435 );
buf ( RI210cf278_242 , n436 );
buf ( RI21a0d528_129 , n437 );
buf ( RI210d7cc0_185 , n438 );
buf ( RI210cea08_243 , n439 );
buf ( RI210cfc50_238 , n440 );
buf ( RI210ce030_247 , n441 );
buf ( RI21a0adc8_157 , n442 );
buf ( RI21a0d4b0_130 , n443 );
buf ( RI210d7c48_186 , n444 );
buf ( RI210ce990_244 , n445 );
buf ( RI210cf3e0_239 , n446 );
buf ( RI210d7360_188 , n447 );
buf ( RI210ce918_245 , n448 );
buf ( RI210cf368_240 , n449 );
buf ( RI210d72e8_189 , n450 );
buf ( RI21a0a648_159 , n451 );
buf ( RI21a0d3c0_132 , n452 );
buf ( RI210d7270_190 , n453 );
buf ( RI21a0a5d0_160 , n454 );
buf ( RI21a0d348_133 , n455 );
buf ( RI210d6a00_191 , n456 );
buf ( RI21a0a558_161 , n457 );
buf ( RI21a0d2d0_134 , n458 );
buf ( RI210d6988_192 , n459 );
buf ( RI21a09e50_162 , n460 );
buf ( RI21a0cbc8_135 , n461 );
buf ( RI21a09dd8_163 , n462 );
buf ( RI21a0cb50_136 , n463 );
buf ( RI210d6898_194 , n464 );
buf ( RI21a09478_164 , n465 );
buf ( RI21a0cad8_137 , n466 );
buf ( RI210d6028_195 , n467 );
buf ( RI210dadf8_165 , n468 );
buf ( RI21a0ca60_138 , n469 );
buf ( RI210d5fb0_196 , n470 );
buf ( RI210dad80_166 , n471 );
buf ( RI21a0c9e8_139 , n472 );
buf ( RI21a16a38_35 , n473 );
buf ( RI210d5650_199 , n474 );
buf ( RI210da420_169 , n475 );
buf ( RI21a0c1f0_142 , n476 );
buf ( RI210d5f38_197 , n477 );
buf ( RI210da510_167 , n478 );
buf ( RI21a0c970_140 , n479 );
buf ( RI21a11650_88 , n480 );
buf ( RI21a115d8_89 , n481 );
buf ( RI210cfd40_236 , n482 );
buf ( RI210c9b48_275 , n483 );
buf ( RI210ca3b8_274 , n484 );
buf ( RI210ca4a8_272 , n485 );
buf ( RI210ca520_271 , n486 );
buf ( RI210cad90_270 , n487 );
buf ( RI210cae08_269 , n488 );
buf ( RI210cae80_268 , n489 );
buf ( RI210caef8_267 , n490 );
buf ( RI210cb768_266 , n491 );
buf ( RI210cb7e0_265 , n492 );
buf ( RI210cb858_264 , n493 );
buf ( RI210cb8d0_263 , n494 );
buf ( RI210cc1b8_261 , n495 );
buf ( RI210cc230_260 , n496 );
buf ( RI210cc2a8_259 , n497 );
buf ( RI210ccb18_258 , n498 );
buf ( RI210ccb90_257 , n499 );
buf ( RI210ccc08_256 , n500 );
buf ( RI210ccc80_255 , n501 );
buf ( RI210cd4f0_254 , n502 );
buf ( RI210cd568_253 , n503 );
buf ( RI210cd5e0_252 , n504 );
buf ( RI210c07a0_282 , n505 );
buf ( RI210c0818_281 , n506 );
buf ( RI210c2078_280 , n507 );
buf ( RI210c9170_279 , n508 );
buf ( RI210c91e8_278 , n509 );
buf ( RI210c9a58_277 , n510 );
buf ( RI210c9ad0_276 , n511 );
buf ( RI210ca430_273 , n512 );
buf ( RI210cc140_262 , n513 );
buf ( RI210cd658_251 , n514 );
buf ( RI2107f4a8_454 , n515 );
buf ( RI210aeb90_395 , n516 );
buf ( GI20471ac0_434 , n517 );
buf ( RI2107f340_457 , n518 );
buf ( RI2107e878_458 , n519 );
buf ( RI21084f20_415 , n520 );
buf ( RI21084458_416 , n521 );
buf ( RI2107e800_459 , n522 );
buf ( RI2107e788_460 , n523 );
buf ( RI2107e710_461 , n524 );
buf ( RI2107e698_462 , n525 );
buf ( RI210843e0_417 , n526 );
buf ( RI210a63a0_396 , n527 );
buf ( RI21086e10_397 , n528 );
buf ( RI21086bb8_398 , n529 );
buf ( RI21086b40_399 , n530 );
buf ( RI21086ac8_400 , n531 );
buf ( RI21086a50_401 , n532 );
buf ( RI210869d8_402 , n533 );
buf ( RI21086960_403 , n534 );
buf ( RI21085e98_404 , n535 );
buf ( RI21085e20_405 , n536 );
buf ( RI21085da8_406 , n537 );
buf ( RI21085d30_407 , n538 );
buf ( RI21085cb8_408 , n539 );
buf ( RI21085c40_409 , n540 );
buf ( RI21085178_410 , n541 );
buf ( RI21085100_411 , n542 );
buf ( RI21085088_412 , n543 );
buf ( RI21085010_413 , n544 );
buf ( RI21084f98_414 , n545 );
buf ( RI210b2538_374 , n546 );
buf ( RI210b43b0_360 , n547 );
buf ( RI210b7f38_335 , n548 );
buf ( RI210afec8_388 , n549 );
buf ( RI210b2628_372 , n550 );
buf ( RI210b4d88_356 , n551 );
buf ( RI21081b18_438 , n552 );
buf ( RI210b6b88_343 , n553 );
buf ( RI210b07b0_386 , n554 );
buf ( RI21081aa0_439 , n555 );
buf ( RI210b5670_354 , n556 );
buf ( RI210afe50_389 , n557 );
buf ( RI21080fd8_440 , n558 );
buf ( RI21083648_424 , n559 );
buf ( RI2107f3b8_456 , n560 );
buf ( RI21080f60_441 , n561 );
buf ( RI210835d0_425 , n562 );
buf ( RI210afdd8_390 , n563 );
buf ( RI21080ee8_442 , n564 );
buf ( RI210b4d10_357 , n565 );
buf ( RI210af568_391 , n566 );
buf ( RI21080e70_443 , n567 );
buf ( RI210b4c98_358 , n568 );
buf ( RI210af4f0_392 , n569 );
buf ( RI21080df8_444 , n570 );
buf ( RI21083558_426 , n571 );
buf ( RI210af478_393 , n572 );
buf ( RI21080d80_445 , n573 );
buf ( RI210834e0_427 , n574 );
buf ( RI210aec08_394 , n575 );
buf ( RI210b25b0_373 , n576 );
buf ( RI210b4428_359 , n577 );
buf ( RI210b1cc8_375 , n578 );
buf ( RI21082a18_428 , n579 );
buf ( RI210b7ec0_336 , n580 );
buf ( RI210802b8_446 , n581 );
buf ( RI210829a0_429 , n582 );
buf ( RI210b7e48_337 , n583 );
buf ( RI21080240_447 , n584 );
buf ( RI21082928_430 , n585 );
buf ( RI210b7dd0_338 , n586 );
buf ( RI210801c8_448 , n587 );
buf ( RI210828b0_431 , n588 );
buf ( RI210b7560_339 , n589 );
buf ( RI21080150_449 , n590 );
buf ( RI21082838_432 , n591 );
buf ( RI210b74e8_340 , n592 );
buf ( RI210800d8_450 , n593 );
buf ( RI210827c0_433 , n594 );
buf ( RI210b7470_341 , n595 );
buf ( RI21080060_451 , n596 );
buf ( RI21081cf8_434 , n597 );
buf ( RI21084200_421 , n598 );
buf ( RI2107f598_452 , n599 );
buf ( RI21081c80_435 , n600 );
buf ( RI21083738_422 , n601 );
buf ( RI210b1c50_376 , n602 );
buf ( RI21081c08_436 , n603 );
buf ( RI210836c0_423 , n604 );
buf ( RI2107f520_453 , n605 );
buf ( RI21081b90_437 , n606 );
buf ( RI210b73f8_342 , n607 );
buf ( RI2107f430_455 , n608 );
buf ( RI210b4338_361 , n609 );
buf ( RI210b6b10_344 , n610 );
buf ( RI210b1bd8_377 , n611 );
buf ( RI210b42c0_362 , n612 );
buf ( RI210b6a98_345 , n613 );
buf ( RI210b1b60_378 , n614 );
buf ( RI210b3a50_363 , n615 );
buf ( RI210b6a20_346 , n616 );
buf ( RI210b12f0_379 , n617 );
buf ( RI210b39d8_364 , n618 );
buf ( RI210b61b0_347 , n619 );
buf ( RI210b1278_380 , n620 );
buf ( RI210b3960_365 , n621 );
buf ( RI210b6138_348 , n622 );
buf ( RI210b1200_381 , n623 );
buf ( RI210b38e8_366 , n624 );
buf ( RI210b60c0_349 , n625 );
buf ( RI210b1188_382 , n626 );
buf ( RI210b3078_367 , n627 );
buf ( RI210b6048_350 , n628 );
buf ( RI210b0918_383 , n629 );
buf ( RI210b3000_368 , n630 );
buf ( RI210b57d8_351 , n631 );
buf ( RI210b08a0_384 , n632 );
buf ( RI210b2f88_369 , n633 );
buf ( RI210b5760_352 , n634 );
buf ( RI210cdec8_250 , n635 );
buf ( RI210aff40_387 , n636 );
buf ( RI210b26a0_371 , n637 );
buf ( RI210b4e00_355 , n638 );
buf ( RI210b0828_385 , n639 );
buf ( RI210b2f10_370 , n640 );
buf ( RI210b56e8_353 , n641 );
buf ( RI210bd668_302 , n642 );
buf ( RI210bcdf8_303 , n643 );
buf ( RI21077000_517 , n644 );
buf ( RI21076538_518 , n645 );
buf ( RI210cdf40_249 , n646 );
buf ( RI2107db58_464 , n647 );
buf ( RI21069950_647 , n648 );
buf ( RI210699c8_646 , n649 );
buf ( n650 , R_61e_1dfaf3c8 );
buf ( n651 , R_8f7_1e09b6c8 );
buf ( n652 , R_714_1dfb8888 );
buf ( n653 , R_951_1e17ef68 );
buf ( n654 , R_28c_1d9fb268 );
buf ( n655 , R_9be_1e183888 );
buf ( n656 , R_9ab_1e1827a8 );
buf ( n657 , R_30f_1d9d04a8 );
buf ( n658 , R_959_1e17f468 );
buf ( n659 , R_b13_1e6b0908 );
buf ( n660 , R_519_1dda4b48 );
buf ( n661 , R_92d_1e09d888 );
buf ( n662 , R_c06_1e6bafe8 );
buf ( n663 , R_8c6_1e099d28 );
buf ( n664 , R_845_1e094788 );
buf ( n665 , R_414_1d9da7c8 );
buf ( n666 , R_313_1d9d0728 );
buf ( n667 , R_518_1dda4aa8 );
buf ( n668 , R_9d9_1e184468 );
buf ( n669 , R_4dd_1dda25c8 );
buf ( n670 , R_59f_1dda9f08 );
buf ( n671 , R_517_1dda4a08 );
buf ( n672 , R_509_1dda4148 );
buf ( n673 , R_508_1dda40a8 );
buf ( n674 , R_401_1d9d9be8 );
buf ( n675 , R_5f9_1ddad748 );
buf ( n676 , R_6ef_1dfb7168 );
buf ( n677 , R_a30_1e187ac8 );
buf ( n678 , R_2b0_1d9fc8e8 );
buf ( n679 , R_77c_1dfbc988 );
buf ( n680 , R_8f1_1e09b308 );
buf ( n681 , R_36a_1d9d4288 );
buf ( n682 , R_507_1dda4008 );
buf ( n683 , R_516_1dda4e68 );
buf ( n684 , R_98e_1e181a88 );
buf ( n685 , R_8d5_1e09a188 );
buf ( n686 , R_498_1dd9faa8 );
buf ( n687 , R_68b_1dfb32e8 );
buf ( n688 , R_773_1dfbc3e8 );
buf ( n689 , R_45b_1d9dd428 );
buf ( n690 , R_48d_1dd9f3c8 );
buf ( n691 , R_5ff_1ddadb08 );
buf ( n692 , R_705_1dfb7f28 );
buf ( n693 , R_644_1dfb0688 );
buf ( n694 , R_63a_1dfb0548 );
buf ( n695 , R_ac7_1e18d928 );
buf ( n696 , R_320_1d9d0f48 );
buf ( n697 , R_737_1dfb9e68 );
buf ( n698 , R_506_1dda4468 );
buf ( n699 , R_647_1dfb0868 );
buf ( n700 , R_b86_1e6bb4e8 );
buf ( n701 , R_883_1e096e48 );
buf ( n702 , R_6a8_1dfb4508 );
buf ( n703 , R_aa5_1e18c3e8 );
buf ( n704 , R_440_1d9dc348 );
buf ( n705 , R_2f9_1d9cf6e8 );
buf ( n706 , R_69c_1dfb3d88 );
buf ( n707 , R_65d_1dfb1628 );
buf ( n708 , R_b0c_1e6b04a8 );
buf ( n709 , R_b20_1e6b1128 );
buf ( n710 , R_a2e_1e189788 );
buf ( n711 , R_905_1e09bf88 );
buf ( n712 , R_a57_1e189328 );
buf ( n713 , R_5f8_1ddad6a8 );
buf ( n714 , R_54c_1dda6b28 );
buf ( n715 , R_bd2_1e6b32e8 );
buf ( n716 , R_aca_1e6ae068 );
buf ( n717 , R_58b_1dda9288 );
buf ( n718 , R_2e3_1d9ce928 );
buf ( n719 , R_3e2_1d9d8d88 );
buf ( n720 , R_8f6_1e09bb28 );
buf ( n721 , R_331_1d9d19e8 );
buf ( n722 , R_97d_1e180ae8 );
buf ( n723 , R_5cd_1ddabbc8 );
buf ( n724 , R_45c_1d9dd4c8 );
buf ( n725 , R_999_1e181c68 );
buf ( n726 , R_b99_1e6b5cc8 );
buf ( n727 , R_948_1e17e9c8 );
buf ( n728 , R_97e_1e181308 );
buf ( n729 , R_ab0_1e18cac8 );
buf ( n730 , R_bb8_1e6b7028 );
buf ( n731 , R_489_1dd9f148 );
buf ( n732 , R_4b6_1dda1268 );
buf ( n733 , R_63f_1dfb0368 );
buf ( n734 , R_3e7_1d9d8ba8 );
buf ( n735 , R_2bd_1d9fd108 );
buf ( n736 , R_81b_1e092d48 );
buf ( n737 , R_b54_1e6b31a8 );
buf ( n738 , R_4df_1dda2708 );
buf ( n739 , R_bab_1e6b6808 );
buf ( n740 , R_431_1d9db9e8 );
buf ( n741 , R_2f2_1d9cf788 );
buf ( n742 , R_601_1ddadc48 );
buf ( n743 , R_6e7_1dfb6c68 );
buf ( n744 , R_bdf_1e6b8888 );
buf ( n745 , R_656_1dfb1bc8 );
buf ( n746 , R_4e0_1dda27a8 );
buf ( n747 , R_4de_1dda2b68 );
buf ( n748 , R_a4e_1e189288 );
buf ( n749 , R_8e1_1e09a908 );
buf ( n750 , R_8f0_1e09b268 );
buf ( n751 , R_299_1d9fba88 );
buf ( n752 , R_292_1d9fb628 );
buf ( n753 , R_4e1_1dda2848 );
buf ( n754 , R_a7f_1e18ac28 );
buf ( n755 , R_c04_1e6b9fa8 );
buf ( n756 , R_3ef_1d9d90a8 );
buf ( n757 , R_5de_1dd9f1e8 );
buf ( n758 , R_878_1e096768 );
buf ( n759 , R_720_1dfb9008 );
buf ( n760 , R_ad6_1e6ae7e8 );
buf ( n761 , R_9a2_1e182708 );
buf ( n762 , R_630_1dfafa08 );
buf ( n763 , R_52f_1dda5908 );
buf ( n764 , R_7a9_1e08e608 );
buf ( n765 , R_976_1e180b88 );
buf ( n766 , R_439_1d9dbee8 );
buf ( n767 , R_604_1ddade28 );
buf ( n768 , R_530_1dda59a8 );
buf ( n769 , R_52e_1dda5d68 );
buf ( n770 , R_7ed_1e091088 );
buf ( n771 , R_3f2_1d9d4c88 );
buf ( n772 , R_3d4_1d9d7fc8 );
buf ( n773 , R_84a_1e094fa8 );
buf ( n774 , R_2de_1d9ceb08 );
buf ( n775 , R_690_1dfb3608 );
buf ( n776 , R_4cd_1dda1bc8 );
buf ( n777 , R_531_1dda5a48 );
buf ( n778 , R_b34_1e6b1da8 );
buf ( n779 , R_5f7_1ddad608 );
buf ( n780 , R_806_1e092528 );
buf ( n781 , R_a5b_1e1895a8 );
buf ( n782 , R_718_1dfb8b08 );
buf ( n783 , R_695_1dfb3928 );
buf ( n784 , R_7af_1e08e9c8 );
buf ( n785 , R_62b_1dfaf6e8 );
buf ( n786 , R_904_1e09bee8 );
buf ( n787 , R_501_1dda3c48 );
buf ( n788 , R_585_1dda8ec8 );
buf ( n789 , R_9cd_1e183ce8 );
buf ( n790 , R_78c_1dfbd388 );
buf ( n791 , R_392_1d9d5b88 );
buf ( n792 , R_4b4_1dda0c28 );
buf ( n793 , R_b44_1e6b27a8 );
buf ( n794 , R_969_1e17fe68 );
buf ( n795 , R_40d_1d9da368 );
buf ( n796 , R_627_1dfaf468 );
buf ( n797 , R_67a_1dfadfc8 );
buf ( n798 , R_45d_1d9dd568 );
buf ( n799 , R_7c1_1e08f508 );
buf ( n800 , R_552_1dda73e8 );
buf ( n801 , R_2bf_1d9fd248 );
buf ( n802 , R_5d4_1ddac028 );
buf ( n803 , R_b77_1e6b4788 );
buf ( n804 , R_3fa_1d9db088 );
buf ( n805 , R_6aa_1dfb4b48 );
buf ( n806 , R_82a_1e093ba8 );
buf ( n807 , R_3aa_1d9d6a88 );
buf ( n808 , R_300_1d9cfb48 );
buf ( n809 , R_405_1d9d9e68 );
buf ( n810 , R_953_1e17f0a8 );
buf ( n811 , R_3cf_1d9d7ca8 );
buf ( n812 , R_ac1_1e18d568 );
buf ( n813 , R_61c_1dfaed88 );
buf ( n814 , R_a99_1e18bc68 );
buf ( n815 , R_4ae_1dda0fe8 );
buf ( n816 , R_aec_1e6af0a8 );
buf ( n817 , R_af8_1e6af828 );
buf ( n818 , R_762_1dfbbe48 );
buf ( n819 , R_3a8_1d9d6448 );
buf ( n820 , R_4ca_1dda1ee8 );
buf ( n821 , R_6b7_1dfb4e68 );
buf ( n822 , R_57c_1dda8928 );
buf ( n823 , R_52b_1dda5688 );
buf ( n824 , R_8ef_1e09b1c8 );
buf ( n825 , R_8c5_1e099788 );
buf ( n826 , R_8ab_1e098748 );
buf ( n827 , R_71c_1dfb8d88 );
buf ( n828 , R_388_1d9d5048 );
buf ( n829 , R_b6e_1e6b46e8 );
buf ( n830 , R_9cc_1e183c48 );
buf ( n831 , R_65b_1dfb14e8 );
buf ( n832 , R_bbd_1e6b7348 );
buf ( n833 , R_3b2_1d9d6f88 );
buf ( n834 , R_862_1e095ea8 );
buf ( n835 , R_4a5_1dda02c8 );
buf ( n836 , R_90f_1e09c5c8 );
buf ( n837 , R_702_1dfb8248 );
buf ( n838 , R_29f_1d9fbe48 );
buf ( n839 , R_72b_1dfb96e8 );
buf ( n840 , R_6f4_1dfb7488 );
buf ( n841 , R_5f2_1dda8a68 );
buf ( n842 , R_a64_1e189b48 );
buf ( n843 , R_2e9_1d9cece8 );
buf ( n844 , R_683_1dfb2de8 );
buf ( n845 , R_2fd_1d9cf968 );
buf ( n846 , R_8b2_1e0990a8 );
buf ( n847 , R_5f0_1ddad1a8 );
buf ( n848 , R_bac_1e6b68a8 );
buf ( n849 , R_642_1dfb0a48 );
buf ( n850 , R_5f6_1d9fbda8 );
buf ( n851 , R_568_1dda7ca8 );
buf ( n852 , R_409_1d9da0e8 );
buf ( n853 , R_5a8_1ddaa4a8 );
buf ( n854 , R_5e3_1ddac988 );
buf ( n855 , R_96b_1e17ffa8 );
buf ( n856 , R_bca_1e6b14e8 );
buf ( n857 , R_3b8_1d9d6e48 );
buf ( n858 , R_789_1dfbd1a8 );
buf ( n859 , R_86a_1e0963a8 );
buf ( n860 , R_416_1ddabc68 );
buf ( n861 , R_903_1e09be48 );
buf ( n862 , R_a2d_1e1878e8 );
buf ( n863 , R_9cb_1e183ba8 );
buf ( n864 , R_59b_1dda9c88 );
buf ( n865 , R_a4c_1e188c48 );
buf ( n866 , R_79c_1dfbdd88 );
buf ( n867 , R_888_1e097168 );
buf ( n868 , R_2a7_1d9fc348 );
buf ( n869 , R_7f3_1e091448 );
buf ( n870 , R_73c_1dfba188 );
buf ( n871 , R_bd1_1e6b7fc8 );
buf ( n872 , R_4a6_1dda0868 );
buf ( n873 , R_3dd_1d9d8568 );
buf ( n874 , R_346_1d9d2c08 );
buf ( n875 , R_4c4_1dda1628 );
buf ( n876 , R_b15_1e6b0a48 );
buf ( n877 , R_5ec_1ddacf28 );
buf ( n878 , R_bb4_1e6b6da8 );
buf ( n879 , R_bed_1e6b9148 );
buf ( n880 , R_7bf_1e08f3c8 );
buf ( n881 , R_344_1d9d25c8 );
buf ( n882 , R_c0b_1e6ba408 );
buf ( n883 , R_6a5_1dfb4328 );
buf ( n884 , R_b8c_1e6b54a8 );
buf ( n885 , R_3a1_1d9d5fe8 );
buf ( n886 , R_7ea_1e09d928 );
buf ( n887 , R_46e_1dd9e568 );
buf ( n888 , R_8ee_1e09b628 );
buf ( n889 , R_697_1dfb3a68 );
buf ( n890 , R_77f_1dfbcb68 );
buf ( n891 , R_391_1d9d55e8 );
buf ( n892 , R_746_1dfb6448 );
buf ( n893 , R_b3b_1e6b2208 );
buf ( n894 , R_7f1_1e091308 );
buf ( n895 , R_410_1d9da548 );
buf ( n896 , R_700_1dfb7c08 );
buf ( n897 , R_58f_1dda9508 );
buf ( n898 , R_582_1dda91e8 );
buf ( n899 , R_793_1dfbd7e8 );
buf ( n900 , R_847_1e0948c8 );
buf ( n901 , R_95e_1e17fc88 );
buf ( n902 , R_560_1dda77a8 );
buf ( n903 , R_9ca_1e184008 );
buf ( n904 , R_397_1d9d59a8 );
buf ( n905 , R_46b_1d9dde28 );
buf ( n906 , R_44e_1d9fc028 );
buf ( n907 , R_6cc_1dfb5b88 );
buf ( n908 , R_62e_1dfafdc8 );
buf ( n909 , R_2b1_1d9fc988 );
buf ( n910 , R_6f9_1dfb77a8 );
buf ( n911 , R_af5_1e6af648 );
buf ( n912 , R_b81_1e6b4dc8 );
buf ( n913 , R_427_1d9db3a8 );
buf ( n914 , R_547_1dda6808 );
buf ( n915 , R_c1d_1e6baf48 );
buf ( n916 , R_a2c_1e187848 );
buf ( n917 , R_355_1d9d3068 );
buf ( n918 , R_857_1e0952c8 );
buf ( n919 , R_413_1d9da728 );
buf ( n920 , R_afa_1e6afe68 );
buf ( n921 , R_adc_1e6ae6a8 );
buf ( n922 , R_5fc_1ddad928 );
buf ( n923 , R_c24_1e6bb3a8 );
buf ( n924 , R_421_1d9dafe8 );
buf ( n925 , R_892_1e17e608 );
buf ( n926 , R_70b_1dfb82e8 );
buf ( n927 , R_aad_1e18c8e8 );
buf ( n928 , R_3ca_1d9d8108 );
buf ( n929 , R_7ac_1e08e7e8 );
buf ( n930 , R_8da_1e09a9a8 );
buf ( n931 , R_400_1d9d9b48 );
buf ( n932 , R_bb0_1e6b6b28 );
buf ( n933 , R_893_1e097848 );
buf ( n934 , R_902_1e09c2a8 );
buf ( n935 , R_a93_1e18b8a8 );
buf ( n936 , R_8cd_1e099c88 );
buf ( n937 , R_861_1e095908 );
buf ( n938 , R_3ea_1d9d9288 );
buf ( n939 , R_915_1e09c988 );
buf ( n940 , R_844_1e0946e8 );
buf ( n941 , R_677_1dfb2668 );
buf ( n942 , R_602_1dfae248 );
buf ( n943 , R_39c_1d9d5cc8 );
buf ( n944 , R_be3_1e6b8b08 );
buf ( n945 , R_bea_1e6b9468 );
buf ( n946 , R_993_1e1818a8 );
buf ( n947 , R_bad_1e6b6948 );
buf ( n948 , R_88d_1e097488 );
buf ( n949 , R_5a2_1ddaa5e8 );
buf ( n950 , R_655_1dfb1128 );
buf ( n951 , R_4ad_1dda07c8 );
buf ( n952 , R_493_1dd9f788 );
buf ( n953 , R_894_1e0978e8 );
buf ( n954 , R_668_1dfb1d08 );
buf ( n955 , R_730_1dfb9a08 );
buf ( n956 , R_7dc_1e0905e8 );
buf ( n957 , R_abd_1e18d2e8 );
buf ( n958 , R_662_1dfb1e48 );
buf ( n959 , R_a7c_1e18aa48 );
buf ( n960 , R_5cf_1ddabd08 );
buf ( n961 , R_328_1d9d1448 );
buf ( n962 , R_741_1dfba4a8 );
buf ( n963 , R_9a6_1e182988 );
buf ( n964 , R_36d_1d9d3f68 );
buf ( n965 , R_308_1d9d0048 );
buf ( n966 , R_95b_1e17f5a8 );
buf ( n967 , R_b63_1e6b3b08 );
buf ( n968 , R_2da_1d9ce888 );
buf ( n969 , R_5dc_1ddac528 );
buf ( n970 , R_49f_1dd9ff08 );
buf ( n971 , R_895_1e097988 );
buf ( n972 , R_761_1dfbb8a8 );
buf ( n973 , R_2e4_1d9ce9c8 );
buf ( n974 , R_ab5_1e18cde8 );
buf ( n975 , R_c28_1e6bb628 );
buf ( n976 , R_8d4_1e09a0e8 );
buf ( n977 , R_a8c_1e18b448 );
buf ( n978 , R_597_1dda9a08 );
buf ( n979 , R_5c4_1ddab628 );
buf ( n980 , R_384_1d9d4dc8 );
buf ( n981 , R_31c_1d9d0cc8 );
buf ( n982 , R_987_1e181128 );
buf ( n983 , R_b2e_1e6b1ee8 );
buf ( n984 , R_2f3_1d9cf328 );
buf ( n985 , R_6cf_1dfb5d68 );
buf ( n986 , R_6e4_1dfb6a88 );
buf ( n987 , R_357_1d9d31a8 );
buf ( n988 , R_3c1_1d9d73e8 );
buf ( n989 , R_5e7_1ddacc08 );
buf ( n990 , R_974_1e180548 );
buf ( n991 , R_61a_1dfaf148 );
buf ( n992 , R_3f8_1d9d9648 );
buf ( n993 , R_802_1e0922a8 );
buf ( n994 , R_593_1dda9788 );
buf ( n995 , R_a69_1e189e68 );
buf ( n996 , R_a87_1e18b128 );
buf ( n997 , R_a5d_1e1896e8 );
buf ( n998 , R_a2b_1e1877a8 );
buf ( n999 , R_671_1dfb22a8 );
buf ( n1000 , R_4cf_1dda1d08 );
buf ( n1001 , R_420_1d9daf48 );
buf ( n1002 , R_6bc_1dfb5188 );
buf ( n1003 , R_43f_1d9dc2a8 );
buf ( n1004 , R_692_1dfb3c48 );
buf ( n1005 , R_80b_1e092348 );
buf ( n1006 , R_882_1e0972a8 );
buf ( n1007 , R_871_1e096308 );
buf ( n1008 , R_2c2_1d9fd928 );
buf ( n1009 , R_2ce_1d9cfa08 );
buf ( n1010 , R_a9c_1e18be48 );
buf ( n1011 , R_768_1dfbbd08 );
buf ( n1012 , R_56d_1dda7fc8 );
buf ( n1013 , R_34c_1d9d2ac8 );
buf ( n1014 , R_b8f_1e6b5688 );
buf ( n1015 , R_b07_1e6b0188 );
buf ( n1016 , R_6b5_1dfb4d28 );
buf ( n1017 , R_5ae_1ddaad68 );
buf ( n1018 , R_2df_1d9ce6a8 );
buf ( n1019 , R_674_1dfb2488 );
buf ( n1020 , R_608_1dfae108 );
buf ( n1021 , R_ad3_1e6ae108 );
buf ( n1022 , R_505_1dda3ec8 );
buf ( n1023 , R_8bf_1e0993c8 );
buf ( n1024 , R_542_1dda69e8 );
buf ( n1025 , R_7f6_1e091b28 );
buf ( n1026 , R_504_1dda3e28 );
buf ( n1027 , R_8a7_1e0984c8 );
buf ( n1028 , R_76a_1dfbc5c8 );
buf ( n1029 , R_937_1e09dec8 );
buf ( n1030 , R_6fb_1dfb78e8 );
buf ( n1031 , R_3b0_1d9d6948 );
buf ( n1032 , R_2c0_1d9fd2e8 );
buf ( n1033 , R_37c_1d9d48c8 );
buf ( n1034 , R_782_1dfbd248 );
buf ( n1035 , R_503_1dda3d88 );
buf ( n1036 , R_82e_1e093e28 );
buf ( n1037 , R_8bb_1e099148 );
buf ( n1038 , R_430_1d9db948 );
buf ( n1039 , R_5cb_1ddaba88 );
buf ( n1040 , R_ae6_1e6af1e8 );
buf ( n1041 , R_7a3_1e08e248 );
buf ( n1042 , R_b78_1e6b4828 );
buf ( n1043 , R_bc9_1e6b7ac8 );
buf ( n1044 , R_380_1d9d4b48 );
buf ( n1045 , R_33d_1d9d2168 );
buf ( n1046 , R_8e0_1e09a868 );
buf ( n1047 , R_3c7_1d9d77a8 );
buf ( n1048 , R_2b2_1d9fcf28 );
buf ( n1049 , R_618_1dfaeb08 );
buf ( n1050 , R_823_1e093248 );
buf ( n1051 , R_89e_1e098428 );
buf ( n1052 , R_502_1dda41e8 );
buf ( n1053 , R_b6f_1e6b4288 );
buf ( n1054 , R_c00_1e6b9d28 );
buf ( n1055 , R_98d_1e1814e8 );
buf ( n1056 , R_28b_1d9fb1c8 );
buf ( n1057 , R_a55_1e1891e8 );
buf ( n1058 , R_3c4_1d9d75c8 );
buf ( n1059 , R_40c_1d9da2c8 );
buf ( n1060 , R_2d2_1d9ce388 );
buf ( n1061 , R_c21_1e6bb1c8 );
buf ( n1062 , R_b3d_1e6b2348 );
buf ( n1063 , R_877_1e0966c8 );
buf ( n1064 , R_855_1e095188 );
buf ( n1065 , R_41d_1d9dad68 );
buf ( n1066 , R_438_1d9dbe48 );
buf ( n1067 , R_2d6_1d9ce608 );
buf ( n1068 , R_7da_1e0909a8 );
buf ( n1069 , R_6f6_1dfb7ac8 );
buf ( n1070 , R_9aa_1e182e88 );
buf ( n1071 , R_b47_1e6b2988 );
buf ( n1072 , R_a2a_1e6b3ce8 );
buf ( n1073 , R_41f_1d9daea8 );
buf ( n1074 , R_ae4_1e6aeba8 );
buf ( n1075 , R_a79_1e18a868 );
buf ( n1076 , R_3a3_1d9d6128 );
buf ( n1077 , R_5bd_1ddab1c8 );
buf ( n1078 , R_301_1d9cfbe8 );
buf ( n1079 , R_298_1d9fb9e8 );
buf ( n1080 , R_bb9_1e6b70c8 );
buf ( n1081 , R_82d_1e093888 );
buf ( n1082 , R_404_1d9d9dc8 );
buf ( n1083 , R_a62_1e189f08 );
buf ( n1084 , R_93c_1e17e248 );
buf ( n1085 , R_62d_1dfaf828 );
buf ( n1086 , R_579_1dda8748 );
buf ( n1087 , R_452_1ddac3e8 );
buf ( n1088 , R_54d_1dda6bc8 );
buf ( n1089 , R_4d9_1dda2348 );
buf ( n1090 , R_4d4_1dda2028 );
buf ( n1091 , R_6c1_1dfb54a8 );
buf ( n1092 , R_379_1d9d46e8 );
buf ( n1093 , R_34e_1d9d3108 );
buf ( n1094 , R_94a_1e097ca8 );
buf ( n1095 , R_74b_1dfbaae8 );
buf ( n1096 , R_ade_1e6aece8 );
buf ( n1097 , R_79f_1e08dfc8 );
buf ( n1098 , R_797_1dfbda68 );
buf ( n1099 , R_943_1e17e6a8 );
buf ( n1100 , R_653_1dfb0fe8 );
buf ( n1101 , R_3d8_1d9d8248 );
buf ( n1102 , R_b61_1e6b39c8 );
buf ( n1103 , R_bc4_1e6b77a8 );
buf ( n1104 , R_a02_1e186308 );
buf ( n1105 , R_368_1d9d3c48 );
buf ( n1106 , R_35e_1d9d3b08 );
buf ( n1107 , R_7fe_1e092028 );
buf ( n1108 , R_499_1dd9fb48 );
buf ( n1109 , R_680_1dfb2c08 );
buf ( n1110 , R_2a8_1d9fc3e8 );
buf ( n1111 , R_6ec_1dfb6f88 );
buf ( n1112 , R_776_1dfbcac8 );
buf ( n1113 , R_b5e_1e6b0368 );
buf ( n1114 , R_635_1dfafd28 );
buf ( n1115 , R_7fa_1e091da8 );
buf ( n1116 , R_af7_1e6af788 );
buf ( n1117 , R_8c4_1e0996e8 );
buf ( n1118 , R_408_1d9da048 );
buf ( n1119 , R_ab9_1e18d068 );
buf ( n1120 , R_6a2_1dfb61c8 );
buf ( n1121 , R_291_1d9fb588 );
buf ( n1122 , R_7b8_1e08ef68 );
buf ( n1123 , R_8b6_1e08e6a8 );
buf ( n1124 , R_48a_1dda0d68 );
buf ( n1125 , R_6c7_1dfb5868 );
buf ( n1126 , R_c10_1e6ba728 );
buf ( n1127 , R_bf1_1e6b93c8 );
buf ( n1128 , R_4d6_1dd9e2e8 );
buf ( n1129 , R_5b3_1ddaab88 );
buf ( n1130 , R_771_1dfbc2a8 );
buf ( n1131 , R_af1_1e6af3c8 );
buf ( n1132 , R_6e1_1dfb68a8 );
buf ( n1133 , R_a9f_1e18c028 );
buf ( n1134 , R_b17_1e6b0b88 );
buf ( n1135 , R_b30_1e6b1b28 );
buf ( n1136 , R_bde_1e6b37e8 );
buf ( n1137 , R_998_1e181bc8 );
buf ( n1138 , R_a4a_1e189008 );
buf ( n1139 , R_48e_1dd9f968 );
buf ( n1140 , R_688_1dfb3108 );
buf ( n1141 , R_810_1e092668 );
buf ( n1142 , R_75c_1dfbb588 );
buf ( n1143 , R_3bb_1d9d7028 );
buf ( n1144 , R_c2e_1e17f008 );
buf ( n1145 , R_5d2_1d9db308 );
buf ( n1146 , R_32e_1d9d1d08 );
buf ( n1147 , R_580_1dda8ba8 );
buf ( n1148 , R_453_1d9dcf28 );
buf ( n1149 , R_83a_1e0913a8 );
buf ( n1150 , R_41e_1d9dc988 );
buf ( n1151 , R_97c_1e180a48 );
buf ( n1152 , R_5b8_1ddaaea8 );
buf ( n1153 , R_363_1d9d3928 );
buf ( n1154 , R_94e_1ddadce8 );
buf ( n1155 , R_7c4_1e08f6e8 );
buf ( n1156 , R_52c_1dda5728 );
buf ( n1157 , R_aa2_1e18c708 );
buf ( n1158 , R_625_1dfaf328 );
buf ( n1159 , R_4b7_1dda0e08 );
buf ( n1160 , R_55d_1dda75c8 );
buf ( n1161 , R_b0e_1e6b0ae8 );
buf ( n1162 , R_425_1d9db268 );
buf ( n1163 , R_30c_1d9d02c8 );
buf ( n1164 , R_3db_1d9d8428 );
buf ( n1165 , R_a48_1e1889c8 );
buf ( n1166 , R_aaf_1e18ca28 );
buf ( n1167 , R_5ad_1ddaa7c8 );
buf ( n1168 , R_589_1dda9148 );
buf ( n1169 , R_338_1d9d1e48 );
buf ( n1170 , R_832_1e0940a8 );
buf ( n1171 , R_790_1dfbd608 );
buf ( n1172 , R_318_1d9d0a48 );
buf ( n1173 , R_869_1e095e08 );
buf ( n1174 , R_6d3_1dfb5fe8 );
buf ( n1175 , R_60c_1dfae388 );
buf ( n1176 , R_56a_1dda82e8 );
buf ( n1177 , R_887_1e0970c8 );
buf ( n1178 , R_815_1e092988 );
buf ( n1179 , R_66b_1dfb1ee8 );
buf ( n1180 , R_a34_1e187d48 );
buf ( n1181 , R_40f_1d9da4a8 );
buf ( n1182 , R_ac3_1e18d6a8 );
buf ( n1183 , R_324_1d9d11c8 );
buf ( n1184 , R_614_1dfae888 );
buf ( n1185 , R_752_1dfbb448 );
buf ( n1186 , R_4c0_1dda13a8 );
buf ( n1187 , R_7d9_1e090408 );
buf ( n1188 , R_ad0_1e18dec8 );
buf ( n1189 , R_bee_1e6b96e8 );
buf ( n1190 , R_736_1dfba2c8 );
buf ( n1191 , R_727_1dfb9468 );
buf ( n1192 , R_a8a_1e18b808 );
buf ( n1193 , R_933_1e09dc48 );
buf ( n1194 , R_8b1_1e098b08 );
buf ( n1195 , R_606_1dfae4c8 );
buf ( n1196 , R_927_1e09d4c8 );
buf ( n1197 , R_a7a_1e18ae08 );
buf ( n1198 , R_333_1d9d1b28 );
buf ( n1199 , R_968_1e17fdc8 );
buf ( n1200 , R_574_1dda8428 );
buf ( n1201 , R_836_1e094328 );
buf ( n1202 , R_757_1dfbb268 );
buf ( n1203 , R_2db_1d9ce428 );
buf ( n1204 , R_af4_1e6af5a8 );
buf ( n1205 , R_454_1d9dcfc8 );
buf ( n1206 , R_412_1d9dab88 );
buf ( n1207 , R_709_1dfb81a8 );
buf ( n1208 , R_8a4_1e0982e8 );
buf ( n1209 , R_c1b_1e6bae08 );
buf ( n1210 , R_846_1e094d28 );
buf ( n1211 , R_3ff_1d9d9aa8 );
buf ( n1212 , R_76e_1dfbdec8 );
buf ( n1213 , R_33f_1d9d22a8 );
buf ( n1214 , R_4af_1dda0908 );
buf ( n1215 , R_a67_1e189d28 );
buf ( n1216 , R_616_1dfaeec8 );
buf ( n1217 , R_b49_1e6b2ac8 );
buf ( n1218 , R_2f4_1d9cf3c8 );
buf ( n1219 , R_426_1d9db808 );
buf ( n1220 , R_2e5_1d9cea68 );
buf ( n1221 , R_bb5_1e6b6e48 );
buf ( n1222 , R_7b6_1e08f328 );
buf ( n1223 , R_751_1dfbaea8 );
buf ( n1224 , R_bd0_1e6b7f28 );
buf ( n1225 , R_610_1dfae608 );
buf ( n1226 , R_918_1e09cb68 );
buf ( n1227 , R_35c_1d9d34c8 );
buf ( n1228 , R_924_1e09d2e8 );
buf ( n1229 , R_912_1e09cca8 );
buf ( n1230 , R_77d_1dfbca28 );
buf ( n1231 , R_774_1dfbc488 );
buf ( n1232 , R_a71_1e18a368 );
buf ( n1233 , R_32d_1d9d1768 );
buf ( n1234 , R_99d_1e181ee8 );
buf ( n1235 , R_87d_1e096a88 );
buf ( n1236 , R_472_1dd9e7e8 );
buf ( n1237 , R_b2a_1e6b1c68 );
buf ( n1238 , R_56f_1dda8108 );
buf ( n1239 , R_b87_1e6b5188 );
buf ( n1240 , R_921_1e09d108 );
buf ( n1241 , R_375_1d9d4468 );
buf ( n1242 , R_576_1dda8ce8 );
buf ( n1243 , R_b82_1e6b5368 );
buf ( n1244 , R_39e_1d9d6308 );
buf ( n1245 , R_856_1e095728 );
buf ( n1246 , R_6c2_1dfb5a48 );
buf ( n1247 , R_2c3_1d9fd4c8 );
buf ( n1248 , R_90b_1e09c348 );
buf ( n1249 , R_92f_1e09d9c8 );
buf ( n1250 , R_38e_1d9d5908 );
buf ( n1251 , R_b9e_1e18d388 );
buf ( n1252 , R_8cc_1e099be8 );
buf ( n1253 , R_860_1e095868 );
buf ( n1254 , R_c09_1e6ba2c8 );
buf ( n1255 , R_b09_1e6b02c8 );
buf ( n1256 , R_521_1dda5048 );
buf ( n1257 , R_b4a_1e6b3068 );
buf ( n1258 , R_88c_1e0973e8 );
buf ( n1259 , R_520_1dda4fa8 );
buf ( n1260 , R_8b5_1e098d88 );
buf ( n1261 , R_b5d_1e6b3748 );
buf ( n1262 , R_843_1e094648 );
buf ( n1263 , R_633_1dfafbe8 );
buf ( n1264 , R_7c2_1e08faa8 );
buf ( n1265 , R_6d8_1dfb6308 );
buf ( n1266 , R_38d_1d9d5368 );
buf ( n1267 , R_7e7_1e090cc8 );
buf ( n1268 , R_bfc_1e6b9aa8 );
buf ( n1269 , R_841_1e094508 );
buf ( n1270 , R_a96_1e18bf88 );
buf ( n1271 , R_7e5_1e090b88 );
buf ( n1272 , R_51f_1dda4f08 );
buf ( n1273 , R_949_1e17ea68 );
buf ( n1274 , R_b5a_1e6b3a68 );
buf ( n1275 , R_2e0_1d9ce748 );
buf ( n1276 , R_acd_1e18dce8 );
buf ( n1277 , R_70f_1dfb8568 );
buf ( n1278 , R_c15_1e6baa48 );
buf ( n1279 , R_310_1d9d0548 );
buf ( n1280 , R_bf5_1e6b9648 );
buf ( n1281 , R_314_1d9d07c8 );
buf ( n1282 , R_6af_1dfb4968 );
buf ( n1283 , R_445_1d9dc668 );
buf ( n1284 , R_658_1dfb1308 );
buf ( n1285 , R_a6c_1e18a048 );
buf ( n1286 , R_2c1_1d9fd388 );
buf ( n1287 , R_2b3_1d9fcac8 );
buf ( n1288 , R_6de_1dfb6bc8 );
buf ( n1289 , R_9b9_1e183068 );
buf ( n1290 , R_6ad_1dfb4828 );
buf ( n1291 , R_548_1dda68a8 );
buf ( n1292 , R_4c9_1dda1948 );
buf ( n1293 , R_51e_1dda5368 );
buf ( n1294 , R_96a_1e180408 );
buf ( n1295 , R_455_1d9dd068 );
buf ( n1296 , R_8d3_1e09a048 );
buf ( n1297 , R_bb1_1e6b6bc8 );
buf ( n1298 , R_7d7_1e0902c8 );
buf ( n1299 , R_6a0_1dfb4008 );
buf ( n1300 , R_b79_1e6b48c8 );
buf ( n1301 , R_565_1dda7ac8 );
buf ( n1302 , R_586_1dda9468 );
buf ( n1303 , R_4a7_1dda0408 );
buf ( n1304 , R_b70_1e6b4328 );
buf ( n1305 , R_661_1dfb18a8 );
buf ( n1306 , R_2d3_1d9fdec8 );
buf ( n1307 , R_ad9_1e6ae4c8 );
buf ( n1308 , R_a85_1e18afe8 );
buf ( n1309 , R_a77_1e18a728 );
buf ( n1310 , R_2d7_1d9ce1a8 );
buf ( n1311 , R_7b3_1e08ec48 );
buf ( n1312 , R_870_1e096268 );
buf ( n1313 , R_43e_1d9dc708 );
buf ( n1314 , R_6db_1dfb64e8 );
buf ( n1315 , R_807_1e0920c8 );
buf ( n1316 , R_a74_1e18a548 );
buf ( n1317 , R_bf9_1e6b98c8 );
buf ( n1318 , R_321_1d9d0fe8 );
buf ( n1319 , R_a53_1e1890a8 );
buf ( n1320 , R_4e3_1dda2988 );
buf ( n1321 , R_831_1e093b08 );
buf ( n1322 , R_66e_1dfb25c8 );
buf ( n1323 , R_ac6_1e18dd88 );
buf ( n1324 , R_55a_1dda78e8 );
buf ( n1325 , R_4c6_1dda1c68 );
buf ( n1326 , R_4e4_1dda2a28 );
buf ( n1327 , R_4e2_1dda2de8 );
buf ( n1328 , R_c22_1e6b55e8 );
buf ( n1329 , R_92c_1e09d7e8 );
buf ( n1330 , R_7c9_1e08fa08 );
buf ( n1331 , R_623_1dfaf1e8 );
buf ( n1332 , R_b58_1e6b3428 );
buf ( n1333 , R_370_1d9d4148 );
buf ( n1334 , R_3be_1d9d7708 );
buf ( n1335 , R_4e5_1dda2ac8 );
buf ( n1336 , R_a03_1e185ea8 );
buf ( n1337 , R_c12_1e6bad68 );
buf ( n1338 , R_456_1d9dd608 );
buf ( n1339 , R_bf2_1e6b9968 );
buf ( n1340 , R_6a7_1dfb4468 );
buf ( n1341 , R_c30_1e6bbb28 );
buf ( n1342 , R_40b_1d9da228 );
buf ( n1343 , R_42f_1d9db8a8 );
buf ( n1344 , R_68d_1dfb3428 );
buf ( n1345 , R_735_1dfb9d28 );
buf ( n1346 , R_78d_1dfbd428 );
buf ( n1347 , R_8df_1e09a7c8 );
buf ( n1348 , R_41c_1d9dacc8 );
buf ( n1349 , R_46f_1dd9e108 );
buf ( n1350 , R_2a9_1d9fc488 );
buf ( n1351 , R_81e_1e093428 );
buf ( n1352 , R_5e0_1ddac7a8 );
buf ( n1353 , R_462_1d9ddd88 );
buf ( n1354 , R_60a_1dfae748 );
buf ( n1355 , R_5a7_1ddaa408 );
buf ( n1356 , R_403_1d9d9d28 );
buf ( n1357 , R_2c6_1d9fdba8 );
buf ( n1358 , R_7e3_1e090a48 );
buf ( n1359 , R_7ee_1e09c528 );
buf ( n1360 , R_706_1dfb84c8 );
buf ( n1361 , R_c17_1e6bab88 );
buf ( n1362 , R_c1f_1e6bb088 );
buf ( n1363 , R_b93_1e6b5908 );
buf ( n1364 , R_854_1e0950e8 );
buf ( n1365 , R_b9f_1e6b6088 );
buf ( n1366 , R_8e5_1e09ab88 );
buf ( n1367 , R_437_1d9dbda8 );
buf ( n1368 , R_612_1dfaec48 );
buf ( n1369 , R_816_1e0931a8 );
buf ( n1370 , R_b19_1e6b0cc8 );
buf ( n1371 , R_73b_1dfba0e8 );
buf ( n1372 , R_a44_1e188748 );
buf ( n1373 , R_93e_1e17e888 );
buf ( n1374 , R_67c_1dfb2988 );
buf ( n1375 , R_992_1e181d08 );
buf ( n1376 , R_494_1dd9f828 );
buf ( n1377 , R_3e0_1d9d8748 );
buf ( n1378 , R_7a7_1e08e4c8 );
buf ( n1379 , R_876_1e096b28 );
buf ( n1380 , R_543_1dda6588 );
buf ( n1381 , R_8ae_1dfbc0c8 );
buf ( n1382 , R_351_1d9d2de8 );
buf ( n1383 , R_457_1d9dd1a8 );
buf ( n1384 , R_bf6_1e6b3f68 );
buf ( n1385 , R_a38_1e187fc8 );
buf ( n1386 , R_6f1_1dfb72a8 );
buf ( n1387 , R_b3e_1e6b28e8 );
buf ( n1388 , R_53e_1dda6768 );
buf ( n1389 , R_ac0_1e18d4c8 );
buf ( n1390 , R_763_1dfbb9e8 );
buf ( n1391 , R_c26_1e6b8ce8 );
buf ( n1392 , R_650_1dfb0e08 );
buf ( n1393 , R_361_1d9d37e8 );
buf ( n1394 , R_aaa_1e187e88 );
buf ( n1395 , R_b10_1e6b0728 );
buf ( n1396 , R_b2c_1e6b18a8 );
buf ( n1397 , R_5a1_1ddaa048 );
buf ( n1398 , R_be7_1e6b8d88 );
buf ( n1399 , R_b26_1e6b19e8 );
buf ( n1400 , R_4a0_1dd9ffa8 );
buf ( n1401 , R_95a_1e17fa08 );
buf ( n1402 , R_909_1e09c208 );
buf ( n1403 , R_463_1d9dd928 );
buf ( n1404 , R_407_1d9d9fa8 );
buf ( n1405 , R_5c5_1ddab6c8 );
buf ( n1406 , R_986_1e181588 );
buf ( n1407 , R_515_1dda48c8 );
buf ( n1408 , R_5c1_1ddab448 );
buf ( n1409 , R_297_1d9fb948 );
buf ( n1410 , R_514_1dda4828 );
buf ( n1411 , R_b4c_1e6b2ca8 );
buf ( n1412 , R_973_1e1804a8 );
buf ( n1413 , R_60e_1dfae9c8 );
buf ( n1414 , R_7d4_1e0900e8 );
buf ( n1415 , R_7c7_1e08f8c8 );
buf ( n1416 , R_513_1dda4788 );
buf ( n1417 , R_65f_1dfb1768 );
buf ( n1418 , R_9b5_1e182de8 );
buf ( n1419 , R_2ee_1d9cf508 );
buf ( n1420 , R_91b_1e09cd48 );
buf ( n1421 , R_af6_1e6afbe8 );
buf ( n1422 , R_83d_1e094288 );
buf ( n1423 , R_8c3_1e099648 );
buf ( n1424 , R_458_1d9dd248 );
buf ( n1425 , R_512_1dda4be8 );
buf ( n1426 , R_ba6_1e6b69e8 );
buf ( n1427 , R_5e5_1ddacac8 );
buf ( n1428 , R_57b_1dda8888 );
buf ( n1429 , R_aeb_1e6af008 );
buf ( n1430 , R_7f4_1e0914e8 );
buf ( n1431 , R_a46_1e188d88 );
buf ( n1432 , R_b8d_1e6b5548 );
buf ( n1433 , R_562_1dda7de8 );
buf ( n1434 , R_745_1dfba728 );
buf ( n1435 , R_557_1dda7208 );
buf ( n1436 , R_464_1d9dd9c8 );
buf ( n1437 , R_835_1e093d88 );
buf ( n1438 , R_49a_1dda00e8 );
buf ( n1439 , R_7d1_1e08ff08 );
buf ( n1440 , R_911_1e09c708 );
buf ( n1441 , R_6e9_1dfb6da8 );
buf ( n1442 , R_723_1dfb91e8 );
buf ( n1443 , R_a95_1e18b9e8 );
buf ( n1444 , R_58d_1dda93c8 );
buf ( n1445 , R_a89_1e18b268 );
buf ( n1446 , R_780_1dfbcc08 );
buf ( n1447 , R_740_1dfba408 );
buf ( n1448 , R_72f_1dfb9968 );
buf ( n1449 , R_828_1e093568 );
buf ( n1450 , R_89c_1e097de8 );
buf ( n1451 , R_a32_1e188108 );
buf ( n1452 , R_840_1e094468 );
buf ( n1453 , R_b37_1e6b1f88 );
buf ( n1454 , R_9db_1e1845a8 );
buf ( n1455 , R_b22_1e6b1768 );
buf ( n1456 , R_9dc_1e184648 );
buf ( n1457 , R_9da_1e184a08 );
buf ( n1458 , R_794_1dfbd888 );
buf ( n1459 , R_33a_1d9d2488 );
buf ( n1460 , R_424_1d9db1c8 );
buf ( n1461 , R_2dc_1d9ce4c8 );
buf ( n1462 , R_a6f_1e18a228 );
buf ( n1463 , R_98c_1e181448 );
buf ( n1464 , R_6b6_1dfb52c8 );
buf ( n1465 , R_908_1e09c168 );
buf ( n1466 , R_9dd_1e1846e8 );
buf ( n1467 , R_965_1e17fbe8 );
buf ( n1468 , R_28a_1d9fb128 );
buf ( n1469 , R_529_1dda5548 );
buf ( n1470 , R_40e_1d9da908 );
buf ( n1471 , R_bcd_1e6b7d48 );
buf ( n1472 , R_476_1dd9ea68 );
buf ( n1473 , R_393_1d9d5728 );
buf ( n1474 , R_a40_1e1884c8 );
buf ( n1475 , R_528_1dda54a8 );
buf ( n1476 , R_2fa_1d9d0188 );
buf ( n1477 , R_a3c_1e188248 );
buf ( n1478 , R_868_1e095d68 );
buf ( n1479 , R_2cf_1d9fdc48 );
buf ( n1480 , R_2c4_1d9fd568 );
buf ( n1481 , R_7cc_1e08fbe8 );
buf ( n1482 , R_8fd_1e09ba88 );
buf ( n1483 , R_3d5_1d9d8068 );
buf ( n1484 , R_b64_1e6b3ba8 );
buf ( n1485 , R_527_1dda5408 );
buf ( n1486 , R_9d1_1e183f68 );
buf ( n1487 , R_46c_1d9ddec8 );
buf ( n1488 , R_2f5_1d9cf468 );
buf ( n1489 , R_839_1e094008 );
buf ( n1490 , R_554_1dda7028 );
buf ( n1491 , R_3ab_1d9d6628 );
buf ( n1492 , R_459_1d9dd2e8 );
buf ( n1493 , R_b4f_1e6b2e88 );
buf ( n1494 , R_886_1e097528 );
buf ( n1495 , R_3e5_1d9d8a68 );
buf ( n1496 , R_52d_1dda57c8 );
buf ( n1497 , R_290_1d9fb4e8 );
buf ( n1498 , R_b7a_1e18cc08 );
buf ( n1499 , R_526_1dda5ae8 );
buf ( n1500 , R_79a_1e098e28 );
buf ( n1501 , R_ba0_1e6b6128 );
buf ( n1502 , R_6d1_1dfb5ea8 );
buf ( n1503 , R_713_1dfb87e8 );
buf ( n1504 , R_685_1dfb2f28 );
buf ( n1505 , R_3fe_1d9d9f08 );
buf ( n1506 , R_638_1dfaff08 );
buf ( n1507 , R_465_1d9dda68 );
buf ( n1508 , R_b91_1e6b57c8 );
buf ( n1509 , R_b53_1e6b3108 );
buf ( n1510 , R_8ad_1e098888 );
buf ( n1511 , R_59e_1dd9e068 );
buf ( n1512 , R_9c5_1e1837e8 );
buf ( n1513 , R_3a9_1d9d64e8 );
buf ( n1514 , R_3b3_1d9d6b28 );
buf ( n1515 , R_2b4_1d9fcb68 );
buf ( n1516 , R_af3_1e6af508 );
buf ( n1517 , R_4f9_1dda3748 );
buf ( n1518 , R_a90_1e18b6c8 );
buf ( n1519 , R_389_1d9d50e8 );
buf ( n1520 , R_a6a_1e18a408 );
buf ( n1521 , R_b1b_1e6b0e08 );
buf ( n1522 , R_4f8_1dda36a8 );
buf ( n1523 , R_b66_1e6b9be8 );
buf ( n1524 , R_9d0_1e183ec8 );
buf ( n1525 , R_2e1_1d9ce7e8 );
buf ( n1526 , R_7d2_1e0904a8 );
buf ( n1527 , R_803_1e091e48 );
buf ( n1528 , R_91e_1e09d428 );
buf ( n1529 , R_4f7_1dda3608 );
buf ( n1530 , R_ab4_1e18cd48 );
buf ( n1531 , R_6ee_1dfb75c8 );
buf ( n1532 , R_c05_1e6ba048 );
buf ( n1533 , R_704_1dfb7e88 );
buf ( n1534 , R_353_1d9d2f28 );
buf ( n1535 , R_ba7_1e6b6588 );
buf ( n1536 , R_87c_1e0969e8 );
buf ( n1537 , R_3f5_1d9d9468 );
buf ( n1538 , R_abc_1e18d248 );
buf ( n1539 , R_a83_1e18aea8 );
buf ( n1540 , R_b40_1e6b2528 );
buf ( n1541 , R_a06_1e186588 );
buf ( n1542 , R_907_1e09c0c8 );
buf ( n1543 , R_664_1dfb1a88 );
buf ( n1544 , R_b71_1e6b43c8 );
buf ( n1545 , R_4f6_1ddad2e8 );
buf ( n1546 , R_8b9_1e099008 );
buf ( n1547 , R_971_1e180368 );
buf ( n1548 , R_64e_1dfb11c8 );
buf ( n1549 , R_679_1dfb27a8 );
buf ( n1550 , R_80c_1e0923e8 );
buf ( n1551 , R_347_1d9d27a8 );
buf ( n1552 , R_b28_1e6b1628 );
buf ( n1553 , R_7cf_1e08fdc8 );
buf ( n1554 , R_8fc_1e09b9e8 );
buf ( n1555 , R_72d_1dfb9828 );
buf ( n1556 , R_9c4_1e183748 );
buf ( n1557 , R_997_1e181b28 );
buf ( n1558 , R_85f_1e0957c8 );
buf ( n1559 , R_2d4_1d9cdfc8 );
buf ( n1560 , R_48f_1dd9f508 );
buf ( n1561 , R_adb_1e6ae608 );
buf ( n1562 , R_3b9_1d9d6ee8 );
buf ( n1563 , R_a51_1e188f68 );
buf ( n1564 , R_8cb_1e099b48 );
buf ( n1565 , R_2d8_1d9ce248 );
buf ( n1566 , R_a72_1e18a908 );
buf ( n1567 , R_7f7_1e0916c8 );
buf ( n1568 , R_4b5_1dda0cc8 );
buf ( n1569 , R_88b_1e097348 );
buf ( n1570 , R_aa7_1e18c528 );
buf ( n1571 , R_699_1dfb3ba8 );
buf ( n1572 , R_68a_1dfb3748 );
buf ( n1573 , R_9cf_1e183e28 );
buf ( n1574 , R_345_1d9d2668 );
buf ( n1575 , R_76b_1dfbbee8 );
buf ( n1576 , R_7aa_1e099328 );
buf ( n1577 , R_5e9_1ddacd48 );
buf ( n1578 , R_a04_1e185f48 );
buf ( n1579 , R_36b_1d9d3e28 );
buf ( n1580 , R_444_1d9dc5c8 );
buf ( n1581 , R_842_1e094aa8 );
buf ( n1582 , R_58a_1dda96e8 );
buf ( n1583 , R_97b_1e1809a8 );
buf ( n1584 , R_5bc_1ddab128 );
buf ( n1585 , R_ae9_1e6aeec8 );
buf ( n1586 , R_74e_1dfbc348 );
buf ( n1587 , R_69b_1dfb3ce8 );
buf ( n1588 , R_783_1dfbcde8 );
buf ( n1589 , R_64d_1dfb0c28 );
buf ( n1590 , R_938_1e17dfc8 );
buf ( n1591 , R_7bd_1e08f288 );
buf ( n1592 , R_7ca_1e08ffa8 );
buf ( n1593 , R_482_1ddac668 );
buf ( n1594 , R_2c7_1d9fd748 );
buf ( n1595 , R_621_1dfaf0a8 );
buf ( n1596 , R_9c3_1e1836a8 );
buf ( n1597 , R_309_1d9d00e8 );
buf ( n1598 , R_5f1_1ddad248 );
buf ( n1599 , R_4b8_1dda0ea8 );
buf ( n1600 , R_bcf_1e6b7e88 );
buf ( n1601 , R_824_1e0932e8 );
buf ( n1602 , R_6e6_1dfb70c8 );
buf ( n1603 , R_7a4_1e08e2e8 );
buf ( n1604 , R_59d_1dda9dc8 );
buf ( n1605 , R_769_1dfbbda8 );
buf ( n1606 , R_38a_1d9d5688 );
buf ( n1607 , R_4cb_1dda1a88 );
buf ( n1608 , R_8d9_1e09a408 );
buf ( n1609 , R_8d2_1e09a4a8 );
buf ( n1610 , R_b24_1e6b13a8 );
buf ( n1611 , R_4ba_1d9d9a08 );
buf ( n1612 , R_bdd_1e6b8748 );
buf ( n1613 , R_398_1d9d5a48 );
buf ( n1614 , R_31d_1d9d0d68 );
buf ( n1615 , R_47a_1dd9ece8 );
buf ( n1616 , R_2ca_1d9ce108 );
buf ( n1617 , R_b03_1e6aff08 );
buf ( n1618 , R_2a0_1d9fbee8 );
buf ( n1619 , R_71f_1dfb8f68 );
buf ( n1620 , R_950_1e17eec8 );
buf ( n1621 , R_9ce_1e184288 );
buf ( n1622 , R_aae_1e6b6c68 );
buf ( n1623 , R_b39_1e6b20c8 );
buf ( n1624 , R_906_1e090ea8 );
buf ( n1625 , R_786_1dfbd4c8 );
buf ( n1626 , R_81c_1e092de8 );
buf ( n1627 , R_94b_1e17eba8 );
buf ( n1628 , R_8fb_1e09b948 );
buf ( n1629 , R_3cb_1d9d7a28 );
buf ( n1630 , R_86f_1e0961c8 );
buf ( n1631 , R_584_1dda8e28 );
buf ( n1632 , R_40a_1d9da688 );
buf ( n1633 , R_954_1e17f148 );
buf ( n1634 , R_944_1e17e748 );
buf ( n1635 , R_bc8_1e6b7a28 );
buf ( n1636 , R_9a1_1e182168 );
buf ( n1637 , R_c02_1e6ba5e8 );
buf ( n1638 , R_967_1e17fd28 );
buf ( n1639 , R_7ff_1e091bc8 );
buf ( n1640 , R_329_1d9d14e8 );
buf ( n1641 , R_ba1_1e6b61c8 );
buf ( n1642 , R_717_1dfb8a68 );
buf ( n1643 , R_aa1_1e18c168 );
buf ( n1644 , R_591_1dda9648 );
buf ( n1645 , R_99c_1e181e48 );
buf ( n1646 , R_a42_1e188b08 );
buf ( n1647 , R_ba8_1e6b6628 );
buf ( n1648 , R_ae1_1e6ae9c8 );
buf ( n1649 , R_9c2_1e183b08 );
buf ( n1650 , R_6bb_1dfb50e8 );
buf ( n1651 , R_41b_1d9dac28 );
buf ( n1652 , R_93d_1e17e2e8 );
buf ( n1653 , R_5b2_1ddaafe8 );
buf ( n1654 , R_5d6_1d9dd388 );
buf ( n1655 , R_402_1d9da188 );
buf ( n1656 , R_4b0_1dda09a8 );
buf ( n1657 , R_549_1dda6948 );
buf ( n1658 , R_53a_1dda64e8 );
buf ( n1659 , R_70d_1dfb8428 );
buf ( n1660 , R_aa4_1e18c348 );
buf ( n1661 , R_798_1dfbdb08 );
buf ( n1662 , R_7fb_1e091948 );
buf ( n1663 , R_32a_1d9d1a88 );
buf ( n1664 , R_a36_1e188388 );
buf ( n1665 , R_5ed_1ddacfc8 );
buf ( n1666 , R_b9a_1e6b6268 );
buf ( n1667 , R_c07_1e6ba188 );
buf ( n1668 , R_47e_1dd9ef68 );
buf ( n1669 , R_ad2_1e6ae568 );
buf ( n1670 , R_39d_1d9d5d68 );
buf ( n1671 , R_83f_1e0943c8 );
buf ( n1672 , R_7eb_1e090f48 );
buf ( n1673 , R_42e_1d9dbd08 );
buf ( n1674 , R_b51_1e6b2fc8 );
buf ( n1675 , R_6b4_1dfb4c88 );
buf ( n1676 , R_694_1dfb3888 );
buf ( n1677 , R_68f_1dfb3568 );
buf ( n1678 , R_777_1dfbc668 );
buf ( n1679 , R_7b0_1e08ea68 );
buf ( n1680 , R_7a0_1e08e068 );
buf ( n1681 , R_75e_1dfbbbc8 );
buf ( n1682 , R_5b7_1ddaae08 );
buf ( n1683 , R_63d_1dfb0228 );
buf ( n1684 , R_636_1dfb02c8 );
buf ( n1685 , R_8de_1e09ac28 );
buf ( n1686 , R_2ef_1d9cf0a8 );
buf ( n1687 , R_302_1d9d4508 );
buf ( n1688 , R_9b8_1e182fc8 );
buf ( n1689 , R_4b2_1dda14e8 );
buf ( n1690 , R_8e4_1e09aae8 );
buf ( n1691 , R_3de_1d9d8b08 );
buf ( n1692 , R_ab8_1e18cfc8 );
buf ( n1693 , R_71b_1dfb8ce8 );
buf ( n1694 , R_c0c_1e6ba4a8 );
buf ( n1695 , R_c2b_1e6bb808 );
buf ( n1696 , R_5ac_1ddaa728 );
buf ( n1697 , R_853_1e095048 );
buf ( n1698 , R_2aa_1d9fca28 );
buf ( n1699 , R_385_1d9d4e68 );
buf ( n1700 , R_436_1d9dc208 );
buf ( n1701 , R_a60_1e1898c8 );
buf ( n1702 , R_7bb_1e08f148 );
buf ( n1703 , R_811_1e092708 );
buf ( n1704 , R_4c5_1dda16c8 );
buf ( n1705 , R_406_1d9da408 );
buf ( n1706 , R_473_1dd9e388 );
buf ( n1707 , R_8aa_1e098ba8 );
buf ( n1708 , R_b7e_1e6b50e8 );
buf ( n1709 , R_7b5_1e08ed88 );
buf ( n1710 , R_5fb_1ddad888 );
buf ( n1711 , R_34d_1d9d2b68 );
buf ( n1712 , R_ae3_1e6aeb08 );
buf ( n1713 , R_6f3_1dfb73e8 );
buf ( n1714 , R_82b_1e093748 );
buf ( n1715 , R_72a_1dfbacc8 );
buf ( n1716 , R_bc3_1e6b7708 );
buf ( n1717 , R_8fa_1e09bda8 );
buf ( n1718 , R_567_1dda7c08 );
buf ( n1719 , R_89f_1e097fc8 );
buf ( n1720 , R_3ed_1d9d8f68 );
buf ( n1721 , R_599_1dda9b48 );
buf ( n1722 , R_851_1e094f08 );
buf ( n1723 , R_2dd_1d9ce568 );
buf ( n1724 , R_4a8_1dda04a8 );
buf ( n1725 , R_8a9_1e098608 );
buf ( n1726 , R_366_1d9d4008 );
buf ( n1727 , R_376_1ddad568 );
buf ( n1728 , R_75d_1dfbb628 );
buf ( n1729 , R_59a_1ddaa0e8 );
buf ( n1730 , R_4c2_1dda19e8 );
buf ( n1731 , R_8be_1e08eba8 );
buf ( n1732 , R_2c5_1d9fd608 );
buf ( n1733 , R_595_1dda98c8 );
buf ( n1734 , R_446_1d9dd108 );
buf ( n1735 , R_6c5_1dfb5728 );
buf ( n1736 , R_5d8_1ddac2a8 );
buf ( n1737 , R_682_1dfb3248 );
buf ( n1738 , R_64b_1dfb0ae8 );
buf ( n1739 , R_791_1dfbd6a8 );
buf ( n1740 , R_b7b_1e6b4a08 );
buf ( n1741 , R_3b1_1d9d69e8 );
buf ( n1742 , R_7e9_1e090e08 );
buf ( n1743 , R_beb_1e6b9008 );
buf ( n1744 , R_6c0_1dfb5408 );
buf ( n1745 , R_8ba_1e0995a8 );
buf ( n1746 , R_a8e_1e17f508 );
buf ( n1747 , R_3c8_1d9d7848 );
buf ( n1748 , R_be4_1e6b8ba8 );
buf ( n1749 , R_544_1dda6628 );
buf ( n1750 , R_53f_1dda6308 );
buf ( n1751 , R_90e_1e09ca28 );
buf ( n1752 , R_381_1d9d4be8 );
buf ( n1753 , R_a3e_1e188888 );
buf ( n1754 , R_6fd_1dfb7a28 );
buf ( n1755 , R_a3a_1e188608 );
buf ( n1756 , R_8c2_1e099aa8 );
buf ( n1757 , R_af0_1e6af328 );
buf ( n1758 , R_296_1d9fb8a8 );
buf ( n1759 , R_b12_1e6b0d68 );
buf ( n1760 , R_ba9_1e6b66c8 );
buf ( n1761 , R_b1d_1e6b0f48 );
buf ( n1762 , R_2b5_1d9fcc08 );
buf ( n1763 , R_6ff_1dfb7b68 );
buf ( n1764 , R_a98_1e18bbc8 );
buf ( n1765 , R_58e_1dda9968 );
buf ( n1766 , R_753_1dfbafe8 );
buf ( n1767 , R_3c5_1d9d7668 );
buf ( n1768 , R_447_1d9dc7a8 );
buf ( n1769 , R_61f_1dfaef68 );
buf ( n1770 , R_54e_1dda28e8 );
buf ( n1771 , R_6f8_1dfb7708 );
buf ( n1772 , R_3a4_1d9d61c8 );
buf ( n1773 , R_423_1d9db128 );
buf ( n1774 , R_6a4_1dfb4288 );
buf ( n1775 , R_b9b_1e6b5e08 );
buf ( n1776 , R_a07_1e186128 );
buf ( n1777 , R_55f_1dda7708 );
buf ( n1778 , R_79d_1dfbde28 );
buf ( n1779 , R_66d_1dfb2028 );
buf ( n1780 , R_5e2_1ddacde8 );
buf ( n1781 , R_48b_1dd9f288 );
buf ( n1782 , R_5ee_1dda3a68 );
buf ( n1783 , R_6c6_1dfb2d48 );
buf ( n1784 , R_3e3_1d9d8928 );
buf ( n1785 , R_b83_1e6b4f08 );
buf ( n1786 , R_533_1dda5b88 );
buf ( n1787 , R_42d_1d9db768 );
buf ( n1788 , R_7e0_1e090868 );
buf ( n1789 , R_696_1dfb3ec8 );
buf ( n1790 , R_3f9_1d9d96e8 );
buf ( n1791 , R_b88_1e6b5228 );
buf ( n1792 , R_758_1dfbb308 );
buf ( n1793 , R_3d2_1d9d8388 );
buf ( n1794 , R_534_1dda5c28 );
buf ( n1795 , R_532_1d9d1308 );
buf ( n1796 , R_867_1e095cc8 );
buf ( n1797 , R_2b6_1d9fd1a8 );
buf ( n1798 , R_775_1dfbc528 );
buf ( n1799 , R_3e8_1d9d8c48 );
buf ( n1800 , R_4d0_1dda1da8 );
buf ( n1801 , R_30d_1d9d0368 );
buf ( n1802 , R_4e7_1dda2c08 );
buf ( n1803 , R_70a_1dfb8748 );
buf ( n1804 , R_a58_1e1893c8 );
buf ( n1805 , R_4e8_1dda2ca8 );
buf ( n1806 , R_4e6_1dda3068 );
buf ( n1807 , R_535_1dda5cc8 );
buf ( n1808 , R_5ea_1dda37e8 );
buf ( n1809 , R_929_1e09d608 );
buf ( n1810 , R_448_1d9dc848 );
buf ( n1811 , R_b0b_1e6b0408 );
buf ( n1812 , R_319_1d9d0ae8 );
buf ( n1813 , R_985_1e180fe8 );
buf ( n1814 , R_32f_1d9d18a8 );
buf ( n1815 , R_4e9_1dda2d48 );
buf ( n1816 , R_b1f_1e6b1088 );
buf ( n1817 , R_495_1dd9f8c8 );
buf ( n1818 , R_63b_1dfb00e8 );
buf ( n1819 , R_536_1dda6268 );
buf ( n1820 , R_3d9_1d9d82e8 );
buf ( n1821 , R_a4f_1e188e28 );
buf ( n1822 , R_470_1dd9e1a8 );
buf ( n1823 , R_2d5_1d9ce068 );
buf ( n1824 , R_3f0_1d9d9148 );
buf ( n1825 , R_acf_1e18de28 );
buf ( n1826 , R_ac2_1e18db08 );
buf ( n1827 , R_9b4_1e182d48 );
buf ( n1828 , R_a05_1e185fe8 );
buf ( n1829 , R_2d9_1d9ce2e8 );
buf ( n1830 , R_8ed_1e09b088 );
buf ( n1831 , R_3f3_1d9d9328 );
buf ( n1832 , R_af2_1e6af968 );
buf ( n1833 , R_44d_1d9dcb68 );
buf ( n1834 , R_645_1dfb0728 );
buf ( n1835 , R_648_1dfb0908 );
buf ( n1836 , R_4a1_1dda0048 );
buf ( n1837 , R_749_1dfba9a8 );
buf ( n1838 , R_2c8_1d9fd7e8 );
buf ( n1839 , R_3bc_1d9d70c8 );
buf ( n1840 , R_3f6_1ddad7e8 );
buf ( n1841 , R_596_1dda9e68 );
buf ( n1842 , R_c01_1e6b9dc8 );
buf ( n1843 , R_734_1dfb9c88 );
buf ( n1844 , R_5a5_1ddaa2c8 );
buf ( n1845 , R_6e3_1dfb69e8 );
buf ( n1846 , R_914_1e09c8e8 );
buf ( n1847 , R_43d_1d9dc168 );
buf ( n1848 , R_2cb_1d9fd9c8 );
buf ( n1849 , R_3d0_1d9d7d48 );
buf ( n1850 , R_b67_1e6b3d88 );
buf ( n1851 , R_b01_1e6afdc8 );
buf ( n1852 , R_37d_1d9d4968 );
buf ( n1853 , R_a80_1e18acc8 );
buf ( n1854 , R_9bd_1e1832e8 );
buf ( n1855 , R_339_1d9d1ee8 );
buf ( n1856 , R_7ad_1e08e888 );
buf ( n1857 , R_972_1e180908 );
buf ( n1858 , R_a22_1e184788 );
buf ( n1859 , R_486_1ddacb68 );
buf ( n1860 , R_5d5_1ddac0c8 );
buf ( n1861 , R_592_1dda9be8 );
buf ( n1862 , R_449_1d9dc8e8 );
buf ( n1863 , R_87b_1e096948 );
buf ( n1864 , R_8f5_1e09b588 );
buf ( n1865 , R_35a_1d9d3888 );
buf ( n1866 , R_37a_1ddab9e8 );
buf ( n1867 , R_991_1e181768 );
buf ( n1868 , R_62a_1dfb1448 );
buf ( n1869 , R_808_1e092168 );
buf ( n1870 , R_3a6_1d9d6808 );
buf ( n1871 , R_b95_1e6b5a48 );
buf ( n1872 , R_83e_1e17e108 );
buf ( n1873 , R_386_1d9d5408 );
buf ( n1874 , R_90d_1e09c488 );
buf ( n1875 , R_931_1e09db08 );
buf ( n1876 , R_ac9_1e18da68 );
buf ( n1877 , R_a31_1e187b68 );
buf ( n1878 , R_640_1dfb0408 );
buf ( n1879 , R_667_1dfb1c68 );
buf ( n1880 , R_6cb_1dfb5ae8 );
buf ( n1881 , R_74a_1e17f288 );
buf ( n1882 , R_676_1dfb2ac8 );
buf ( n1883 , R_372_1d9d4788 );
buf ( n1884 , R_56c_1dda7f28 );
buf ( n1885 , R_334_1d9d1bc8 );
buf ( n1886 , R_31e_1d9fc528 );
buf ( n1887 , R_981_1e180d68 );
buf ( n1888 , R_8ca_1e099fa8 );
buf ( n1889 , R_85e_1e095c28 );
buf ( n1890 , R_bbe_1e6af6e8 );
buf ( n1891 , R_49b_1dd9fc88 );
buf ( n1892 , R_73a_1dfba548 );
buf ( n1893 , R_5fe_1dfaf8c8 );
buf ( n1894 , R_98b_1e1813a8 );
buf ( n1895 , R_88e_1e097a28 );
buf ( n1896 , R_28f_1d9fb448 );
buf ( n1897 , R_9bc_1e183248 );
buf ( n1898 , R_5db_1ddac488 );
buf ( n1899 , R_88a_1e08ee28 );
buf ( n1900 , R_5a6_1ddaa868 );
buf ( n1901 , R_443_1d9dc528 );
buf ( n1902 , R_a0a_1e186808 );
buf ( n1903 , R_358_1d9d3248 );
buf ( n1904 , R_88f_1e0975c8 );
buf ( n1905 , R_acc_1e18dc48 );
buf ( n1906 , R_aac_1e18c848 );
buf ( n1907 , R_2a2_1d9fde28 );
buf ( n1908 , R_8a5_1e098388 );
buf ( n1909 , R_8ec_1e09afe8 );
buf ( n1910 , R_289_1d9fb088 );
buf ( n1911 , R_340_1d9d2348 );
buf ( n1912 , R_c2d_1e6bb948 );
buf ( n1913 , R_964_1e17fb48 );
buf ( n1914 , R_85d_1e095688 );
buf ( n1915 , R_6fa_1dfb7d48 );
buf ( n1916 , R_4d5_1dda20c8 );
buf ( n1917 , R_a5a_1e18b308 );
buf ( n1918 , R_7de_1e090c28 );
buf ( n1919 , R_605_1ddadec8 );
buf ( n1920 , R_311_1d9d05e8 );
buf ( n1921 , R_8a6_1e098928 );
buf ( n1922 , R_a2f_1e187a28 );
buf ( n1923 , R_81f_1e092fc8 );
buf ( n1924 , R_3b6_1d9d7208 );
buf ( n1925 , R_315_1d9d0868 );
buf ( n1926 , R_93f_1e17e428 );
buf ( n1927 , R_5b1_1ddaaa48 );
buf ( n1928 , R_631_1dfafaa8 );
buf ( n1929 , R_890_1e097668 );
buf ( n1930 , R_670_1dfb2208 );
buf ( n1931 , R_b9c_1e6b5ea8 );
buf ( n1932 , R_8e9_1e09ae08 );
buf ( n1933 , R_932_1e093928 );
buf ( n1934 , R_817_1e092ac8 );
buf ( n1935 , R_b60_1e6b3928 );
buf ( n1936 , R_979_1e180868 );
buf ( n1937 , R_8d8_1e09a368 );
buf ( n1938 , R_628_1dfaf508 );
buf ( n1939 , R_729_1dfb95a8 );
buf ( n1940 , R_a92_1e18bd08 );
buf ( n1941 , R_b33_1e6b1d08 );
buf ( n1942 , R_2ab_1d9fc5c8 );
buf ( n1943 , R_5e6_1dd9f6e8 );
buf ( n1944 , R_5c0_1ddab3a8 );
buf ( n1945 , R_600_1ddadba8 );
buf ( n1946 , R_8f4_1e09b4e8 );
buf ( n1947 , R_29d_1d9fbd08 );
buf ( n1948 , R_c11_1e6ba7c8 );
buf ( n1949 , R_4d7_1dda2208 );
buf ( n1950 , R_b43_1e6b2708 );
buf ( n1951 , R_881_1e096d08 );
buf ( n1952 , R_891_1e097708 );
buf ( n1953 , R_8b4_1e098ce8 );
buf ( n1954 , R_6ac_1dfb4788 );
buf ( n1955 , R_2f0_1d9cf148 );
buf ( n1956 , R_ad8_1e6ae428 );
buf ( n1957 , R_9bb_1e1831a8 );
buf ( n1958 , R_bd9_1e6b84c8 );
buf ( n1959 , R_39f_1d9d5ea8 );
buf ( n1960 , R_a5e_1e189c88 );
buf ( n1961 , R_303_1d9cfd28 );
buf ( n1962 , R_6ae_1dfb4dc8 );
buf ( n1963 , R_477_1dd9e608 );
buf ( n1964 , R_6d2_1e0981a8 );
buf ( n1965 , R_38f_1d9d54a8 );
buf ( n1966 , R_4d2_1dda23e8 );
buf ( n1967 , R_82f_1e0939c8 );
buf ( n1968 , R_61d_1dfaee28 );
buf ( n1969 , R_673_1dfb23e8 );
buf ( n1970 , R_578_1dda86a8 );
buf ( n1971 , R_a65_1e189be8 );
buf ( n1972 , R_9a5_1e1823e8 );
buf ( n1973 , R_744_1dfba688 );
buf ( n1974 , R_bfe_1e6ba0e8 );
buf ( n1975 , R_86e_1e096628 );
buf ( n1976 , R_6ce_1e0945a8 );
buf ( n1977 , R_9df_1e184828 );
buf ( n1978 , R_571_1dda8248 );
buf ( n1979 , R_9e0_1e1848c8 );
buf ( n1980 , R_9de_1e184c88 );
buf ( n1981 , R_41a_1ddabee8 );
buf ( n1982 , R_36e_1d9d1588 );
buf ( n1983 , R_6b9_1dfb4fa8 );
buf ( n1984 , R_b72_1e6b4968 );
buf ( n1985 , R_73f_1dfba368 );
buf ( n1986 , R_a4d_1e188ce8 );
buf ( n1987 , R_9e1_1e184968 );
buf ( n1988 , R_2d0_1d9fdce8 );
buf ( n1989 , R_72e_1dfb9dc8 );
buf ( n1990 , R_c25_1e6bb448 );
buf ( n1991 , R_8eb_1e09af48 );
buf ( n1992 , R_6eb_1dfb6ee8 );
buf ( n1993 , R_764_1dfbba88 );
buf ( n1994 , R_9b1_1e182b68 );
buf ( n1995 , R_970_1e1802c8 );
buf ( n1996 , R_bce_1e6b82e8 );
buf ( n1997 , R_325_1d9d1268 );
buf ( n1998 , R_65c_1dfb1588 );
buf ( n1999 , R_643_1dfb05e8 );
buf ( n2000 , R_abf_1e18d428 );
buf ( n2001 , R_a9b_1e18bda8 );
buf ( n2002 , R_b7c_1e6b4aa8 );
buf ( n2003 , R_9ba_1e183608 );
buf ( n2004 , R_bef_1e6b9288 );
buf ( n2005 , R_b14_1e6b09a8 );
buf ( n2006 , R_996_1e181f88 );
buf ( n2007 , R_812_1e092ca8 );
buf ( n2008 , R_4a2_1dda05e8 );
buf ( n2009 , R_6e0_1dfb6808 );
buf ( n2010 , R_490_1dd9f5a8 );
buf ( n2011 , R_711_1dfb86a8 );
buf ( n2012 , R_a86_1e18ba88 );
buf ( n2013 , R_342_1d9d2988 );
buf ( n2014 , R_c0e_1e6baae8 );
buf ( n2015 , R_8e3_1e09aa48 );
buf ( n2016 , R_646_1dfb0cc8 );
buf ( n2017 , R_74d_1dfbac28 );
buf ( n2018 , R_67f_1dfb2b68 );
buf ( n2019 , R_34f_1d9d2ca8 );
buf ( n2020 , R_8f3_1e09b448 );
buf ( n2021 , R_bdc_1e6b86a8 );
buf ( n2022 , R_57f_1dda8b08 );
buf ( n2023 , R_77a_1dfbcd48 );
buf ( n2024 , R_4c1_1dda1448 );
buf ( n2025 , R_b8e_1e6b5ae8 );
buf ( n2026 , R_c29_1e6bb6c8 );
buf ( n2027 , R_875_1e096588 );
buf ( n2028 , R_852_1e0954a8 );
buf ( n2029 , R_6a6_1dfb48c8 );
buf ( n2030 , R_76f_1dfbc168 );
buf ( n2031 , R_984_1e180f48 );
buf ( n2032 , R_39a_1d9d6088 );
buf ( n2033 , R_35f_1d9d36a8 );
buf ( n2034 , R_5d0_1ddabda8 );
buf ( n2035 , R_b65_1e6b3c48 );
buf ( n2036 , R_92b_1e09d748 );
buf ( n2037 , R_3eb_1d9d8e28 );
buf ( n2038 , R_53b_1dda6088 );
buf ( n2039 , R_97a_1e180e08 );
buf ( n2040 , R_369_1d9d3ce8 );
buf ( n2041 , R_7f5_1e091588 );
buf ( n2042 , R_588_1dda90a8 );
buf ( n2043 , R_b6a_1e6b4468 );
buf ( n2044 , R_435_1d9dbc68 );
buf ( n2045 , R_a08_1e1861c8 );
buf ( n2046 , R_7ef_1e0911c8 );
buf ( n2047 , R_781_1dfbcca8 );
buf ( n2048 , R_55c_1dda7528 );
buf ( n2049 , R_3bf_1d9d72a8 );
buf ( n2050 , R_850_1e094e68 );
buf ( n2051 , R_2ea_1d9cf288 );
buf ( n2052 , R_687_1dfb3068 );
buf ( n2053 , R_795_1dfbd928 );
buf ( n2054 , R_382_1d9d5188 );
buf ( n2055 , R_63e_1dfb07c8 );
buf ( n2056 , R_2b7_1d9fcd48 );
buf ( n2057 , R_9b0_1e182ac8 );
buf ( n2058 , R_6dd_1dfb6628 );
buf ( n2059 , R_4be_1dda1768 );
buf ( n2060 , R_bfd_1e6b9b48 );
buf ( n2061 , R_b0d_1e6b0548 );
buf ( n2062 , R_b9d_1e6b5f48 );
buf ( n2063 , R_b3a_1e6b2668 );
buf ( n2064 , R_4b9_1dda0f48 );
buf ( n2065 , R_4bb_1dda1088 );
buf ( n2066 , R_9a0_1e1820c8 );
buf ( n2067 , R_83b_1e094148 );
buf ( n2068 , R_8ea_1e09b3a8 );
buf ( n2069 , R_b21_1e6b11c8 );
buf ( n2070 , R_62f_1dfaf968 );
buf ( n2071 , R_91d_1e09ce88 );
buf ( n2072 , R_483_1dd9ed88 );
buf ( n2073 , R_7c0_1e08f468 );
buf ( n2074 , R_bd5_1e6b8248 );
buf ( n2075 , R_364_1d9d39c8 );
buf ( n2076 , R_322_1d9d2e88 );
buf ( n2077 , R_326_1d9d1808 );
buf ( n2078 , R_99b_1e181da8 );
buf ( n2079 , R_961_1e17f968 );
buf ( n2080 , R_726_1dfb98c8 );
buf ( n2081 , R_a7d_1e18aae8 );
buf ( n2082 , R_826_1e09de28 );
buf ( n2083 , R_89a_1dfb4648 );
buf ( n2084 , R_511_1dda4648 );
buf ( n2085 , R_2fb_1d9cf828 );
buf ( n2086 , R_b5c_1e6b36a8 );
buf ( n2087 , R_8b0_1e098a68 );
buf ( n2088 , R_708_1dfb8108 );
buf ( n2089 , R_603_1ddadd88 );
buf ( n2090 , R_804_1e091ee8 );
buf ( n2091 , R_573_1dda8388 );
buf ( n2092 , R_a56_1e189a08 );
buf ( n2093 , R_510_1dda45a8 );
buf ( n2094 , R_833_1e093c48 );
buf ( n2095 , R_8c1_1e099508 );
buf ( n2096 , R_966_1e180188 );
buf ( n2097 , R_46d_1dd9dfc8 );
buf ( n2098 , R_bcc_1e6b7ca8 );
buf ( n2099 , R_47b_1dd9e888 );
buf ( n2100 , R_aea_1e6af468 );
buf ( n2101 , R_8d1_1e099f08 );
buf ( n2102 , R_57a_1ddaa368 );
buf ( n2103 , R_8f2_1e09b8a8 );
buf ( n2104 , R_b35_1e6b1e48 );
buf ( n2105 , R_b05_1e6b0048 );
buf ( n2106 , R_aa9_1e18c668 );
buf ( n2107 , R_9b7_1e182f28 );
buf ( n2108 , R_3ae_1d9d6d08 );
buf ( n2109 , R_50f_1dda4508 );
buf ( n2110 , R_a23_1e1872a8 );
buf ( n2111 , R_2c9_1d9fd888 );
buf ( n2112 , R_5c6_1d9d7e88 );
buf ( n2113 , R_8bd_1e099288 );
buf ( n2114 , R_4b1_1dda0a48 );
buf ( n2115 , R_b45_1e6b2848 );
buf ( n2116 , R_422_1d9db588 );
buf ( n2117 , R_2cc_1d9fda68 );
buf ( n2118 , R_9d5_1e1841e8 );
buf ( n2119 , R_37e_1d9d4f08 );
buf ( n2120 , R_42c_1d9db6c8 );
buf ( n2121 , R_a7e_1e18b088 );
buf ( n2122 , R_a8d_1e18b4e8 );
buf ( n2123 , R_50e_1dda4968 );
buf ( n2124 , R_626_1dfafb48 );
buf ( n2125 , R_5cc_1ddabb28 );
buf ( n2126 , R_295_1d9fb808 );
buf ( n2127 , R_a9e_1e18c488 );
buf ( n2128 , R_80d_1e092488 );
buf ( n2129 , R_9af_1e182a28 );
buf ( n2130 , R_946_1e17ed88 );
buf ( n2131 , R_a5c_1e189648 );
buf ( n2132 , R_5bb_1ddab088 );
buf ( n2133 , R_3e6_1d9d9008 );
buf ( n2134 , R_ab3_1e18cca8 );
buf ( n2135 , R_a1e_1e187488 );
buf ( n2136 , R_66a_1dfb2348 );
buf ( n2137 , R_7f8_1e091768 );
buf ( n2138 , R_56e_1dda8568 );
buf ( n2139 , R_3c2_1d9d7988 );
buf ( n2140 , R_837_1e093ec8 );
buf ( n2141 , R_866_1e096128 );
buf ( n2142 , R_65a_1dfb1948 );
buf ( n2143 , R_4aa_1dda0ae8 );
buf ( n2144 , R_540_1dda63a8 );
buf ( n2145 , R_61b_1dfaece8 );
buf ( n2146 , R_78a_1dfbd748 );
buf ( n2147 , R_76c_1dfbbf88 );
buf ( n2148 , R_4c7_1dda1808 );
buf ( n2149 , R_47f_1dd9eb08 );
buf ( n2150 , R_34a_1d9d4a08 );
buf ( n2151 , R_b57_1e6b3388 );
buf ( n2152 , R_545_1dda66c8 );
buf ( n2153 , R_c13_1e6ba908 );
buf ( n2154 , R_44c_1d9dcac8 );
buf ( n2155 , R_a0b_1e1863a8 );
buf ( n2156 , R_6d5_1dfb6128 );
buf ( n2157 , R_bf3_1e6b9508 );
buf ( n2158 , R_3ee_1d9d9508 );
buf ( n2159 , R_6d7_1dfb6268 );
buf ( n2160 , R_3d6_1d9d9788 );
buf ( n2161 , R_b06_1e6b05e8 );
buf ( n2162 , R_9d4_1e184148 );
buf ( n2163 , R_33b_1d9d2028 );
buf ( n2164 , R_739_1dfb9fa8 );
buf ( n2165 , R_a0e_1e186a88 );
buf ( n2166 , R_7dd_1e090688 );
buf ( n2167 , R_54f_1dda6d08 );
buf ( n2168 , R_926_1e09dba8 );
buf ( n2169 , R_abb_1e18d1a8 );
buf ( n2170 , R_70e_1dfb89c8 );
buf ( n2171 , R_ba2_1e6b6768 );
buf ( n2172 , R_917_1e09cac8 );
buf ( n2173 , R_923_1e09d248 );
buf ( n2174 , R_784_1dfbce88 );
buf ( n2175 , R_920_1e09d068 );
buf ( n2176 , R_564_1dda7a28 );
buf ( n2177 , R_9a9_1e182668 );
buf ( n2178 , R_bfa_1e6b9e68 );
buf ( n2179 , R_62c_1dfaf788 );
buf ( n2180 , R_8c9_1e099a08 );
buf ( n2181 , R_43c_1d9dc0c8 );
buf ( n2182 , R_b00_1e6afd28 );
buf ( n2183 , R_35d_1d9d3568 );
buf ( n2184 , R_c18_1e6bac28 );
buf ( n2185 , R_306_1d9d0408 );
buf ( n2186 , R_939_1e17e068 );
buf ( n2187 , R_474_1dd9e428 );
buf ( n2188 , R_4a9_1dda0548 );
buf ( n2189 , R_2ac_1d9fc668 );
buf ( n2190 , R_609_1dfae1a8 );
buf ( n2191 , R_94c_1e17ec48 );
buf ( n2192 , R_90a_1e09c7a8 );
buf ( n2193 , R_92e_1e0918a8 );
buf ( n2194 , R_7be_1e08f828 );
buf ( n2195 , R_825_1e093388 );
buf ( n2196 , R_559_1dda7348 );
buf ( n2197 , R_bf7_1e6b9788 );
buf ( n2198 , R_87a_1e096da8 );
buf ( n2199 , R_9d3_1e1840a8 );
buf ( n2200 , R_394_1d9d57c8 );
buf ( n2201 , R_31a_1d9d1088 );
buf ( n2202 , R_69f_1dfb3f68 );
buf ( n2203 , R_787_1dfbd068 );
buf ( n2204 , R_a63_1e189aa8 );
buf ( n2205 , R_9ae_1e183388 );
buf ( n2206 , R_945_1e17e7e8 );
buf ( n2207 , R_537_1dda5e08 );
buf ( n2208 , R_725_1dfb9328 );
buf ( n2209 , R_b68_1e6b3e28 );
buf ( n2210 , R_7a5_1e08e388 );
buf ( n2211 , R_4eb_1dda2e88 );
buf ( n2212 , R_619_1dfaeba8 );
buf ( n2213 , R_800_1e091c68 );
buf ( n2214 , R_be8_1e6b8e28 );
buf ( n2215 , R_4ec_1dda2f28 );
buf ( n2216 , R_4ea_1dda32e8 );
buf ( n2217 , R_2f1_1d9cf1e8 );
buf ( n2218 , R_5d3_1ddabf88 );
buf ( n2219 , R_6da_1dfb6948 );
buf ( n2220 , R_5b6_1ddab268 );
buf ( n2221 , R_3ac_1d9d66c8 );
buf ( n2222 , R_983_1e180ea8 );
buf ( n2223 , R_b73_1e6b4508 );
buf ( n2224 , R_4ed_1dda2fc8 );
buf ( n2225 , R_ada_1e6aea68 );
buf ( n2226 , R_7fc_1e0919e8 );
buf ( n2227 , R_b3c_1e6b22a8 );
buf ( n2228 , R_304_1d9cfdc8 );
buf ( n2229 , R_5ab_1ddaa688 );
buf ( n2230 , R_85c_1e0955e8 );
buf ( n2231 , R_442_1d9dcc08 );
buf ( n2232 , R_3ce_1d9d8608 );
buf ( n2233 , R_ad5_1e6ae248 );
buf ( n2234 , R_ae8_1e6aee28 );
buf ( n2235 , R_3b4_1d9d6bc8 );
buf ( n2236 , R_8b8_1e098f68 );
buf ( n2237 , R_b46_1e6b2de8 );
buf ( n2238 , R_8e8_1e09ad68 );
buf ( n2239 , R_bbf_1e6b7488 );
buf ( n2240 , R_799_1dfbdba8 );
buf ( n2241 , R_778_1dfbc708 );
buf ( n2242 , R_a4b_1e188ba8 );
buf ( n2243 , R_51d_1dda4dc8 );
buf ( n2244 , R_657_1dfb1268 );
buf ( n2245 , R_9d2_1e17f788 );
buf ( n2246 , R_348_1d9d2848 );
buf ( n2247 , R_51c_1dda4d28 );
buf ( n2248 , R_8d7_1e09a2c8 );
buf ( n2249 , R_9b3_1e182ca8 );
buf ( n2250 , R_7db_1e090548 );
buf ( n2251 , R_715_1dfb8928 );
buf ( n2252 , R_68c_1dfb3388 );
buf ( n2253 , R_880_1e096c68 );
buf ( n2254 , R_29c_1d9fbc68 );
buf ( n2255 , R_b7d_1e6b4b48 );
buf ( n2256 , R_51b_1dda4c88 );
buf ( n2257 , R_bba_1e6b7668 );
buf ( n2258 , R_3dc_1d9d84c8 );
buf ( n2259 , R_5a0_1dda9fa8 );
buf ( n2260 , R_75f_1dfbb768 );
buf ( n2261 , R_b7f_1e6b4c88 );
buf ( n2262 , R_b16_1e6b0fe8 );
buf ( n2263 , R_ba3_1e6b6308 );
buf ( n2264 , R_654_1dfb1088 );
buf ( n2265 , R_bc7_1e6b7988 );
buf ( n2266 , R_2a3_1d9fc0c8 );
buf ( n2267 , R_6f0_1dfb7208 );
buf ( n2268 , R_7a1_1e08e108 );
buf ( n2269 , R_371_1d9d41e8 );
buf ( n2270 , R_51a_1dda50e8 );
buf ( n2271 , R_ab7_1e18cf28 );
buf ( n2272 , R_7e6_1e099828 );
buf ( n2273 , R_b6b_1e6b4008 );
buf ( n2274 , R_9ad_1e1828e8 );
buf ( n2275 , R_935_1e09dd88 );
buf ( n2276 , R_b8a_1e6bb768 );
buf ( n2277 , R_69d_1dfb3e28 );
buf ( n2278 , R_45e_1d9ddb08 );
buf ( n2279 , R_a1a_1e187208 );
buf ( n2280 , R_a49_1e188a68 );
buf ( n2281 , R_a09_1e186268 );
buf ( n2282 , R_496_1dd9fe68 );
buf ( n2283 , R_336_1d9d2208 );
buf ( n2284 , R_5df_1ddac708 );
buf ( n2285 , R_5c7_1ddab808 );
buf ( n2286 , R_990_1e1816c8 );
buf ( n2287 , R_6c9_1dfb59a8 );
buf ( n2288 , R_2eb_1d9cee28 );
buf ( n2289 , R_2b8_1d9fcde8 );
buf ( n2290 , R_ae0_1e6ae928 );
buf ( n2291 , R_b2f_1e6b1a88 );
buf ( n2292 , R_84d_1e094c88 );
buf ( n2293 , R_a12_1e186d08 );
buf ( n2294 , R_74f_1dfbad68 );
buf ( n2295 , R_a35_1e187de8 );
buf ( n2296 , R_28e_1d9fb3a8 );
buf ( n2297 , R_81a_1e0936a8 );
buf ( n2298 , R_487_1dd9f008 );
buf ( n2299 , R_c1c_1e6baea8 );
buf ( n2300 , R_7a8_1e08e568 );
buf ( n2301 , R_471_1dd9e248 );
buf ( n2302 , R_766_1e0986a8 );
buf ( n2303 , R_38b_1d9d5228 );
buf ( n2304 , R_a7b_1e18a9a8 );
buf ( n2305 , R_b52_1e6b8568 );
buf ( n2306 , R_9ff_1e185c28 );
buf ( n2307 , R_7b9_1e08f008 );
buf ( n2308 , R_67b_1dfb28e8 );
buf ( n2309 , R_a00_1e185cc8 );
buf ( n2310 , R_9fe_1e6bb9e8 );
buf ( n2311 , R_980_1e180cc8 );
buf ( n2312 , R_874_1e0964e8 );
buf ( n2313 , R_49c_1dd9fd28 );
buf ( n2314 , R_58c_1dda9328 );
buf ( n2315 , R_45f_1d9dd6a8 );
buf ( n2316 , R_98a_1e181808 );
buf ( n2317 , R_8e2_1e09aea8 );
buf ( n2318 , R_6ba_1dfb5548 );
buf ( n2319 , R_bd8_1e6b8428 );
buf ( n2320 , R_a8b_1e18b3a8 );
buf ( n2321 , R_a01_1e185d68 );
buf ( n2322 , R_6b3_1dfb4be8 );
buf ( n2323 , R_60d_1dfae428 );
buf ( n2324 , R_6e8_1dfb6d08 );
buf ( n2325 , R_399_1d9d5ae8 );
buf ( n2326 , R_a16_1e186f88 );
buf ( n2327 , R_bc2_1e6b7b68 );
buf ( n2328 , R_32b_1d9d1628 );
buf ( n2329 , R_434_1d9dbbc8 );
buf ( n2330 , R_a24_1e187348 );
buf ( n2331 , R_377_1d9d45a8 );
buf ( n2332 , R_3cc_1d9d7ac8 );
buf ( n2333 , R_a68_1e189dc8 );
buf ( n2334 , R_963_1e17faa8 );
buf ( n2335 , R_7c5_1e08f788 );
buf ( n2336 , R_615_1dfae928 );
buf ( n2337 , R_8a2_1dfb9b48 );
buf ( n2338 , R_722_1dfb9648 );
buf ( n2339 , R_288_1d9f96e8 );
buf ( n2340 , R_556_1dda7668 );
buf ( n2341 , R_748_1dfba908 );
buf ( n2342 , R_865_1e095b88 );
buf ( n2343 , R_607_1dfae068 );
buf ( n2344 , R_691_1dfb36a8 );
buf ( n2345 , R_978_1e1807c8 );
buf ( n2346 , R_84f_1e094dc8 );
buf ( n2347 , R_2cd_1d9fdb08 );
buf ( n2348 , R_ae2_1e6aef68 );
buf ( n2349 , R_a1f_1e187028 );
buf ( n2350 , R_721_1dfb90a8 );
buf ( n2351 , R_733_1dfb9be8 );
buf ( n2352 , R_9e3_1e184aa8 );
buf ( n2353 , R_9e4_1e184b48 );
buf ( n2354 , R_c23_1e6bb308 );
buf ( n2355 , R_9e2_1e184f08 );
buf ( n2356 , R_7ae_1dfbb1c8 );
buf ( n2357 , R_91a_1e09d1a8 );
buf ( n2358 , R_b84_1e6b4fa8 );
buf ( n2359 , R_b92_1e181088 );
buf ( n2360 , R_ba4_1e6b63a8 );
buf ( n2361 , R_754_1dfbb088 );
buf ( n2362 , R_5a4_1ddaa228 );
buf ( n2363 , R_9a4_1e182348 );
buf ( n2364 , R_b08_1e6b0228 );
buf ( n2365 , R_9e5_1e184be8 );
buf ( n2366 , R_617_1dfaea68 );
buf ( n2367 , R_5ce_1ddac168 );
buf ( n2368 , R_b89_1e6b52c8 );
buf ( n2369 , R_7b2_1e09b128 );
buf ( n2370 , R_460_1d9dd748 );
buf ( n2371 , R_5e4_1ddaca28 );
buf ( n2372 , R_30a_1d9d0688 );
buf ( n2373 , R_a0c_1e186448 );
buf ( n2374 , R_910_1e09c668 );
buf ( n2375 , R_553_1dda6f88 );
buf ( n2376 , R_86d_1e096088 );
buf ( n2377 , R_a0f_1e186628 );
buf ( n2378 , R_719_1dfb8ba8 );
buf ( n2379 , R_b48_1e6b2a28 );
buf ( n2380 , R_316_1d9d0e08 );
buf ( n2381 , R_901_1e09bd08 );
buf ( n2382 , R_611_1dfae6a8 );
buf ( n2383 , R_ac5_1e18d7e8 );
buf ( n2384 , R_6c4_1dfb5688 );
buf ( n2385 , R_53c_1dda6128 );
buf ( n2386 , R_712_1dfb8c48 );
buf ( n2387 , R_2f6_1d9cfc88 );
buf ( n2388 , R_829_1e093608 );
buf ( n2389 , R_89d_1e097e88 );
buf ( n2390 , R_8d0_1e099e68 );
buf ( n2391 , R_8ac_1e0987e8 );
buf ( n2392 , R_8a0_1e098068 );
buf ( n2393 , R_aef_1e6af288 );
buf ( n2394 , R_759_1dfbb3a8 );
buf ( n2395 , R_a6d_1e18a0e8 );
buf ( n2396 , R_6bf_1dfb5368 );
buf ( n2397 , R_982_1e182c08 );
buf ( n2398 , R_bdb_1e6b8608 );
buf ( n2399 , R_684_1dfb2e88 );
buf ( n2400 , R_7b7_1e08eec8 );
buf ( n2401 , R_478_1dd9e6a8 );
buf ( n2402 , R_be1_1e6b89c8 );
buf ( n2403 , R_b55_1e6b3248 );
buf ( n2404 , R_79b_1dfbdce8 );
buf ( n2405 , R_c27_1e6bb588 );
buf ( n2406 , R_96f_1e180228 );
buf ( n2407 , R_42b_1d9db628 );
buf ( n2408 , R_6cd_1dfb5c28 );
buf ( n2409 , R_652_1dfb16c8 );
buf ( n2410 , R_71d_1dfb8e28 );
buf ( n2411 , R_703_1dfb7de8 );
buf ( n2412 , R_a54_1e189148 );
buf ( n2413 , R_4a3_1dda0188 );
buf ( n2414 , R_634_1dfafc88 );
buf ( n2415 , R_2ad_1d9fc708 );
buf ( n2416 , R_4cc_1dda1b28 );
buf ( n2417 , R_2a1_1d9fbf88 );
buf ( n2418 , R_93a_1e0977a8 );
buf ( n2419 , R_a78_1e18a7c8 );
buf ( n2420 , R_c03_1e6b9f08 );
buf ( n2421 , R_72c_1dfb9788 );
buf ( n2422 , R_809_1e092208 );
buf ( n2423 , R_5b0_1ddaa9a8 );
buf ( n2424 , R_44b_1d9dca28 );
buf ( n2425 , R_952_1ddab768 );
buf ( n2426 , R_899_1e097c08 );
buf ( n2427 , R_bd4_1e6b81a8 );
buf ( n2428 , R_a94_1e18b948 );
buf ( n2429 , R_6b1_1dfb4aa8 );
buf ( n2430 , R_491_1dd9f648 );
buf ( n2431 , R_5ca_1d9dae08 );
buf ( n2432 , R_6f5_1dfb7528 );
buf ( n2433 , R_9c9_1e183a68 );
buf ( n2434 , R_75a_1dfbb948 );
buf ( n2435 , R_461_1d9dd7e8 );
buf ( n2436 , R_7c3_1e08f648 );
buf ( n2437 , R_569_1dda7d48 );
buf ( n2438 , R_a75_1e18a5e8 );
buf ( n2439 , R_7ec_1e090fe8 );
buf ( n2440 , R_c20_1e6bb128 );
buf ( n2441 , R_96d_1e1800e8 );
buf ( n2442 , R_54a_1dda6ee8 );
buf ( n2443 , R_b31_1e6b1bc8 );
buf ( n2444 , R_5bf_1ddab308 );
buf ( n2445 , R_900_1e09bc68 );
buf ( n2446 , R_b74_1e6b45a8 );
buf ( n2447 , R_940_1e17e4c8 );
buf ( n2448 , R_8dd_1e09a688 );
buf ( n2449 , R_a88_1e18b1c8 );
buf ( n2450 , R_743_1dfba5e8 );
buf ( n2451 , R_2d1_1d9fdd88 );
buf ( n2452 , R_4b3_1dda0b88 );
buf ( n2453 , R_48c_1dd9f328 );
buf ( n2454 , R_419_1d9daae8 );
buf ( n2455 , R_2ba_1d9fd428 );
buf ( n2456 , R_898_1e097b68 );
buf ( n2457 , R_354_1d9d2fc8 );
buf ( n2458 , R_3c9_1d9d78e8 );
buf ( n2459 , R_afd_1e6afb48 );
buf ( n2460 , R_698_1dfb3b08 );
buf ( n2461 , R_8c8_1e099968 );
buf ( n2462 , R_aff_1e6afc88 );
buf ( n2463 , R_59c_1dda9d28 );
buf ( n2464 , R_43b_1d9dc028 );
buf ( n2465 , R_3e1_1d9d87e8 );
buf ( n2466 , R_7d8_1e090368 );
buf ( n2467 , R_624_1dfaf288 );
buf ( n2468 , R_ace_1e6ae2e8 );
buf ( n2469 , R_294_1d9fb768 );
buf ( n2470 , R_818_1e092b68 );
buf ( n2471 , R_9c8_1e1839c8 );
buf ( n2472 , R_5c8_1ddab8a8 );
buf ( n2473 , R_c2f_1e6bba88 );
buf ( n2474 , R_ba5_1e6b6448 );
buf ( n2475 , R_6d0_1dfb5e08 );
buf ( n2476 , R_820_1e093068 );
buf ( n2477 , R_30e_1d9d0908 );
buf ( n2478 , R_99f_1e182028 );
buf ( n2479 , R_73e_1dfba7c8 );
buf ( n2480 , R_4ef_1dda3108 );
buf ( n2481 , R_451_1d9dcde8 );
buf ( n2482 , R_678_1dfb2708 );
buf ( n2483 , R_663_1dfb19e8 );
buf ( n2484 , R_5fa_1e091128 );
buf ( n2485 , R_312_1d9d0b88 );
buf ( n2486 , R_a45_1e1887e8 );
buf ( n2487 , R_b18_1e6b0c28 );
buf ( n2488 , R_4f0_1dda31a8 );
buf ( n2489 , R_4ee_1dda3568 );
buf ( n2490 , R_7ab_1e08e748 );
buf ( n2491 , R_305_1d9cfe68 );
buf ( n2492 , R_955_1e17f1e8 );
buf ( n2493 , R_373_1d9d4328 );
buf ( n2494 , R_a39_1e188068 );
buf ( n2495 , R_669_1dfb1da8 );
buf ( n2496 , R_3a5_1d9d6268 );
buf ( n2497 , R_c0d_1e6ba548 );
buf ( n2498 , R_4f1_1dda3248 );
buf ( n2499 , R_541_1dda6448 );
buf ( n2500 , R_69a_1dfb4148 );
buf ( n2501 , R_b90_1e6b5728 );
buf ( n2502 , R_99a_1e182208 );
buf ( n2503 , R_960_1e17f8c8 );
buf ( n2504 , R_6a9_1dfb45a8 );
buf ( n2505 , R_4bc_1dda1128 );
buf ( n2506 , R_897_1e097ac8 );
buf ( n2507 , R_701_1dfb7ca8 );
buf ( n2508 , R_36c_1d9d3ec8 );
buf ( n2509 , R_60b_1dfae2e8 );
buf ( n2510 , R_583_1dda8d88 );
buf ( n2511 , R_330_1d9d1948 );
buf ( n2512 , R_bb6_1e6b73e8 );
buf ( n2513 , R_71e_1dfb93c8 );
buf ( n2514 , R_590_1dda95a8 );
buf ( n2515 , R_29e_1dda2668 );
buf ( n2516 , R_b0f_1e6b0688 );
buf ( n2517 , R_a1b_1e186da8 );
buf ( n2518 , R_550_1dda6da8 );
buf ( n2519 , R_ac8_1e18d9c8 );
buf ( n2520 , R_a9d_1e18bee8 );
buf ( n2521 , R_561_1dda7848 );
buf ( n2522 , R_80e_1e092a28 );
buf ( n2523 , R_9b6_1e187708 );
buf ( n2524 , R_5e8_1ddacca8 );
buf ( n2525 , R_613_1dfae7e8 );
buf ( n2526 , R_b6c_1e6b40a8 );
buf ( n2527 , R_3d3_1d9d7f28 );
buf ( n2528 , R_31f_1d9d0ea8 );
buf ( n2529 , R_9c7_1e183928 );
buf ( n2530 , R_5dd_1ddac5c8 );
buf ( n2531 , R_78e_1dfbd9c8 );
buf ( n2532 , R_a13_1e1868a8 );
buf ( n2533 , R_70c_1dfb8388 );
buf ( n2534 , R_885_1e096f88 );
buf ( n2535 , R_85b_1e095548 );
buf ( n2536 , R_8ff_1e09bbc8 );
buf ( n2537 , R_716_1dfb8ec8 );
buf ( n2538 , R_2b9_1d9fce88 );
buf ( n2539 , R_b69_1e6b3ec8 );
buf ( n2540 , R_356_1d9d3608 );
buf ( n2541 , R_2e6_1d9cf008 );
buf ( n2542 , R_484_1dd9ee28 );
buf ( n2543 , R_2ec_1d9ceec8 );
buf ( n2544 , R_acb_1e18dba8 );
buf ( n2545 , R_813_1e092848 );
buf ( n2546 , R_4c3_1dda1588 );
buf ( n2547 , R_a47_1e188928 );
buf ( n2548 , R_81d_1e092e88 );
buf ( n2549 , R_8e7_1e09acc8 );
buf ( n2550 , R_5ef_1ddad108 );
buf ( n2551 , R_896_1e094828 );
buf ( n2552 , R_bec_1e6b90a8 );
buf ( n2553 , R_b2b_1e6b1808 );
buf ( n2554 , R_4ab_1dda0688 );
buf ( n2555 , R_7e4_1e090ae8 );
buf ( n2556 , R_a33_1e187ca8 );
buf ( n2557 , R_47c_1dd9e928 );
buf ( n2558 , R_8d6_1e09a728 );
buf ( n2559 , R_87f_1e096bc8 );
buf ( n2560 , R_5b5_1ddaacc8 );
buf ( n2561 , R_651_1dfb0ea8 );
buf ( n2562 , R_3da_1d9d8888 );
buf ( n2563 , R_538_1dda5ea8 );
buf ( n2564 , R_675_1dfb2528 );
buf ( n2565 , R_60f_1dfae568 );
buf ( n2566 , R_29b_1d9fbbc8 );
buf ( n2567 , R_aa6_1e18c988 );
buf ( n2568 , R_3bd_1d9d7168 );
buf ( n2569 , R_be5_1e6b8c48 );
buf ( n2570 , R_c0a_1e6ba868 );
buf ( n2571 , R_5f5_1ddad4c8 );
buf ( n2572 , R_b4b_1e6b2c08 );
buf ( n2573 , R_7b1_1e08eb08 );
buf ( n2574 , R_95d_1e17f6e8 );
buf ( n2575 , R_a17_1e186b28 );
buf ( n2576 , R_a29_1e187668 );
buf ( n2577 , R_71a_1dfb9148 );
buf ( n2578 , R_693_1dfb37e8 );
buf ( n2579 , R_77b_1dfbc8e8 );
buf ( n2580 , R_9c6_1e183d88 );
buf ( n2581 , R_3a7_1d9d63a8 );
buf ( n2582 , R_bc0_1e6b7528 );
buf ( n2583 , R_68e_1dfb39c8 );
buf ( n2584 , R_335_1d9d1c68 );
buf ( n2585 , R_5eb_1ddace88 );
buf ( n2586 , R_ad7_1e6ae388 );
buf ( n2587 , R_765_1dfbbb28 );
buf ( n2588 , R_387_1d9d4fa8 );
buf ( n2589 , R_9a8_1e1825c8 );
buf ( n2590 , R_632_1dfb0048 );
buf ( n2591 , R_6e5_1dfb6b28 );
buf ( n2592 , R_772_1dfbc848 );
buf ( n2593 , R_995_1e1819e8 );
buf ( n2594 , R_7d6_1e090728 );
buf ( n2595 , R_598_1dda9aa8 );
buf ( n2596 , R_a70_1e18a2c8 );
buf ( n2597 , R_a25_1e1873e8 );
buf ( n2598 , R_bbb_1e6b7208 );
buf ( n2599 , R_6f2_1dfb7848 );
buf ( n2600 , R_a41_1e188568 );
buf ( n2601 , R_a66_1e18a188 );
buf ( n2602 , R_a3d_1e1882e8 );
buf ( n2603 , R_341_1d9d23e8 );
buf ( n2604 , R_594_1dda9828 );
buf ( n2605 , R_4fe_1dda5868 );
buf ( n2606 , R_480_1dd9eba8 );
buf ( n2607 , R_6ab_1dfb46e8 );
buf ( n2608 , R_84c_1e094be8 );
buf ( n2609 , R_660_1dfb1808 );
buf ( n2610 , R_a20_1e1870c8 );
buf ( n2611 , R_abe_1e6b64e8 );
buf ( n2612 , R_566_1dda8068 );
buf ( n2613 , R_7c8_1e08f968 );
buf ( n2614 , R_5c2_1d9fc2a8 );
buf ( n2615 , R_989_1e181268 );
buf ( n2616 , R_8a8_1e098568 );
buf ( n2617 , R_2a4_1d9fc168 );
buf ( n2618 , R_7d5_1e090188 );
buf ( n2619 , R_8fe_1e09c028 );
buf ( n2620 , R_3b7_1d9d6da8 );
buf ( n2621 , R_6b8_1dfb4f08 );
buf ( n2622 , R_8b3_1e098c48 );
buf ( n2623 , R_94f_1e17ee28 );
buf ( n2624 , R_9fb_1e1859a8 );
buf ( n2625 , R_a10_1e1866c8 );
buf ( n2626 , R_b36_1e6b23e8 );
buf ( n2627 , R_aa0_1e18c0c8 );
buf ( n2628 , R_c1a_1e6bb268 );
buf ( n2629 , R_82c_1e0937e8 );
buf ( n2630 , R_4d1_1dda1e48 );
buf ( n2631 , R_6fc_1dfb7988 );
buf ( n2632 , R_9fa_1e185e08 );
buf ( n2633 , R_9fc_1e185a48 );
buf ( n2634 , R_a0d_1e1864e8 );
buf ( n2635 , R_be2_1e6b8f68 );
buf ( n2636 , R_b02_1e6b8068 );
buf ( n2637 , R_a28_1e1875c8 );
buf ( n2638 , R_4fd_1dda39c8 );
buf ( n2639 , R_5fd_1ddad9c8 );
buf ( n2640 , R_873_1e096448 );
buf ( n2641 , R_9fd_1e185ae8 );
buf ( n2642 , R_a6b_1e189fa8 );
buf ( n2643 , R_aa3_1e18c2a8 );
buf ( n2644 , R_738_1dfb9f08 );
buf ( n2645 , R_805_1e091f88 );
buf ( n2646 , R_2f7_1d9cf5a8 );
buf ( n2647 , R_5ba_1ddab4e8 );
buf ( n2648 , R_57d_1dda89c8 );
buf ( n2649 , R_475_1dd9e4c8 );
buf ( n2650 , R_433_1d9dbb28 );
buf ( n2651 , R_aed_1e6af148 );
buf ( n2652 , R_4fc_1dda3928 );
buf ( n2653 , R_3a0_1d9d5f48 );
buf ( n2654 , R_3f7_1d9d95a8 );
buf ( n2655 , R_367_1d9d3ba8 );
buf ( n2656 , R_947_1e17e928 );
buf ( n2657 , R_b1a_1e6b1268 );
buf ( n2658 , R_525_1dda52c8 );
buf ( n2659 , R_50d_1dda43c8 );
buf ( n2660 , R_390_1d9d5548 );
buf ( n2661 , R_6fe_1dfb7fc8 );
buf ( n2662 , R_6f7_1dfb7668 );
buf ( n2663 , R_2ae_1d9fcca8 );
buf ( n2664 , R_864_1e095ae8 );
buf ( n2665 , R_9e7_1e184d28 );
buf ( n2666 , R_524_1dda5228 );
buf ( n2667 , R_50c_1dda4328 );
buf ( n2668 , R_9e6_1e185188 );
buf ( n2669 , R_9e8_1e184dc8 );
buf ( n2670 , R_9b2_1e183108 );
buf ( n2671 , R_7e2_1dfbaf48 );
buf ( n2672 , R_622_1dfaf648 );
buf ( n2673 , R_b4e_1e184508 );
buf ( n2674 , R_a91_1e18b768 );
buf ( n2675 , R_a84_1e18af48 );
buf ( n2676 , R_4ce_1dda2168 );
buf ( n2677 , R_bb2_1e6b7168 );
buf ( n2678 , R_523_1dda5188 );
buf ( n2679 , R_50b_1dda4288 );
buf ( n2680 , R_9e9_1e184e68 );
buf ( n2681 , R_4f3_1dda3388 );
buf ( n2682 , R_4fb_1dda3888 );
buf ( n2683 , R_4f2_1ddad068 );
buf ( n2684 , R_4f4_1dda3428 );
buf ( n2685 , R_55e_1dda7b68 );
buf ( n2686 , R_84e_1e095228 );
buf ( n2687 , R_a76_1e18ab88 );
buf ( n2688 , R_5c9_1ddab948 );
buf ( n2689 , R_343_1d9d2528 );
buf ( n2690 , R_a73_1e18a4a8 );
buf ( n2691 , R_7cd_1e08fc88 );
buf ( n2692 , R_522_1dda55e8 );
buf ( n2693 , R_50a_1dda46e8 );
buf ( n2694 , R_4f5_1dda34c8 );
buf ( n2695 , R_396_1d9d5e08 );
buf ( n2696 , R_7f9_1e091808 );
buf ( n2697 , R_681_1dfb2ca8 );
buf ( n2698 , R_37b_1d9d4828 );
buf ( n2699 , R_639_1dfaffa8 );
buf ( n2700 , R_76d_1dfbc028 );
buf ( n2701 , R_78b_1dfbd2e8 );
buf ( n2702 , R_6a3_1dfb41e8 );
buf ( n2703 , R_9ac_1e182848 );
buf ( n2704 , R_86c_1e095fe8 );
buf ( n2705 , R_c08_1e6ba228 );
buf ( n2706 , R_2fc_1d9cf8c8 );
buf ( n2707 , R_7f0_1e091268 );
buf ( n2708 , R_c31_1e6bbbc8 );
buf ( n2709 , R_a52_1e189508 );
buf ( n2710 , R_ab2_1e18d108 );
buf ( n2711 , R_28d_1d9fb308 );
buf ( n2712 , R_bcb_1e6b7c08 );
buf ( n2713 , R_4fa_1dda3f68 );
buf ( n2714 , R_2bb_1d9fcfc8 );
buf ( n2715 , R_b3f_1e6b2488 );
buf ( n2716 , R_a27_1e187528 );
buf ( n2717 , R_362_1d9d3d88 );
buf ( n2718 , R_497_1dd9fa08 );
buf ( n2719 , R_64f_1dfb0d68 );
buf ( n2720 , R_bd7_1e6b8388 );
buf ( n2721 , R_b75_1e6b4648 );
buf ( n2722 , R_98f_1e181628 );
buf ( n2723 , R_6ed_1dfb7028 );
buf ( n2724 , R_7d3_1e090048 );
buf ( n2725 , R_b27_1e6b1588 );
buf ( n2726 , R_39b_1d9d5c28 );
buf ( n2727 , R_8cf_1e099dc8 );
buf ( n2728 , R_689_1dfb31a8 );
buf ( n2729 , R_7c6_1e08fd28 );
buf ( n2730 , R_b2d_1e6b1948 );
buf ( n2731 , R_92a_1e092f28 );
buf ( n2732 , R_66c_1dfb1f88 );
buf ( n2733 , R_956_1e6b00e8 );
buf ( n2734 , R_b96_1e18ce88 );
buf ( n2735 , R_bae_1e6b6ee8 );
buf ( n2736 , R_94d_1e17ece8 );
buf ( n2737 , R_785_1dfbcf28 );
buf ( n2738 , R_6e2_1dfb6e48 );
buf ( n2739 , R_65e_1dfb5cc8 );
buf ( n2740 , R_42a_1d9dba88 );
buf ( n2741 , R_7e8_1e090d68 );
buf ( n2742 , R_b4d_1e6b2d48 );
buf ( n2743 , R_bff_1e6b9c88 );
buf ( n2744 , R_3c0_1d9d7348 );
buf ( n2745 , R_44a_1d9dce88 );
buf ( n2746 , R_2fe_1d9cff08 );
buf ( n2747 , R_383_1d9d4d28 );
buf ( n2748 , R_928_1e09d568 );
buf ( n2749 , R_488_1dd9f0a8 );
buf ( n2750 , R_5aa_1ddaaae8 );
buf ( n2751 , R_3fd_1d9d9968 );
buf ( n2752 , R_7d0_1e08fe68 );
buf ( n2753 , R_7b4_1e08ece8 );
buf ( n2754 , R_4d8_1dda22a8 );
buf ( n2755 , R_418_1d9daa48 );
buf ( n2756 , R_a43_1e1886a8 );
buf ( n2757 , R_327_1d9d13a8 );
buf ( n2758 , R_849_1e094a08 );
buf ( n2759 , R_b5f_1e6b3888 );
buf ( n2760 , R_4d3_1dda1f88 );
buf ( n2761 , R_a97_1e18bb28 );
buf ( n2762 , R_aba_1e18d608 );
buf ( n2763 , R_ab1_1e18cb68 );
buf ( n2764 , R_97f_1e180c28 );
buf ( n2765 , R_788_1dfbd108 );
buf ( n2766 , R_a1c_1e186e48 );
buf ( n2767 , R_b11_1e6b07c8 );
buf ( n2768 , R_a37_1e187f28 );
buf ( n2769 , R_801_1e091d08 );
buf ( n2770 , R_581_1dda8c48 );
buf ( n2771 , R_49d_1dd9fdc8 );
buf ( n2772 , R_56b_1dda7e88 );
buf ( n2773 , R_4da_1dda3ce8 );
buf ( n2774 , R_7f2_1e09d6a8 );
buf ( n2775 , R_53d_1dda61c8 );
buf ( n2776 , R_3df_1d9d86a8 );
buf ( n2777 , R_429_1d9db4e8 );
buf ( n2778 , R_8dc_1e09a5e8 );
buf ( n2779 , R_a14_1e186948 );
buf ( n2780 , R_9d6_1e186088 );
buf ( n2781 , R_add_1e6ae748 );
buf ( n2782 , R_b6d_1e6b4148 );
buf ( n2783 , R_c1e_1e6b4e68 );
buf ( n2784 , R_7fd_1e091a88 );
buf ( n2785 , R_859_1e095408 );
buf ( n2786 , R_b23_1e6b1308 );
buf ( n2787 , R_afc_1e6afaa8 );
buf ( n2788 , R_913_1e09c848 );
buf ( n2789 , R_450_1d9dcd48 );
buf ( n2790 , R_7cb_1e08fb48 );
buf ( n2791 , R_b38_1e6b2028 );
buf ( n2792 , R_a26_1e187988 );
buf ( n2793 , R_74c_1dfbab88 );
buf ( n2794 , R_35b_1d9d3428 );
buf ( n2795 , R_962_1e17ff08 );
buf ( n2796 , R_2e7_1d9ceba8 );
buf ( n2797 , R_8c0_1e099468 );
buf ( n2798 , R_8c7_1e0998c8 );
buf ( n2799 , R_afe_1e6b5d68 );
buf ( n2800 , R_977_1e180728 );
buf ( n2801 , R_925_1e09d388 );
buf ( n2802 , R_919_1e09cc08 );
buf ( n2803 , R_728_1dfb9508 );
buf ( n2804 , R_43a_1d9dc488 );
buf ( n2805 , R_bf0_1e6b9328 );
buf ( n2806 , R_9a3_1e1822a8 );
buf ( n2807 , R_3af_1d9d68a8 );
buf ( n2808 , R_930_1e09da68 );
buf ( n2809 , R_90c_1e09c3e8 );
buf ( n2810 , R_5a9_1ddaa548 );
buf ( n2811 , R_659_1dfb13a8 );
buf ( n2812 , R_c0f_1e6ba688 );
buf ( n2813 , R_307_1d9cffa8 );
buf ( n2814 , R_8bc_1e0991e8 );
buf ( n2815 , R_2ed_1d9cef68 );
buf ( n2816 , R_770_1dfbc208 );
buf ( n2817 , R_34b_1d9d2a28 );
buf ( n2818 , R_37f_1d9d4aa8 );
buf ( n2819 , R_5f4_1ddad428 );
buf ( n2820 , R_779_1dfbc7a8 );
buf ( n2821 , R_46a_1dd9f468 );
buf ( n2822 , R_be0_1e6b8928 );
buf ( n2823 , R_bd3_1e6b8108 );
buf ( n2824 , R_466_1d9d9c88 );
buf ( n2825 , R_77e_1dfbcfc8 );
buf ( n2826 , R_575_1dda84c8 );
buf ( n2827 , R_4ff_1dda3b08 );
buf ( n2828 , R_a18_1e186bc8 );
buf ( n2829 , R_bda_1e6b8a68 );
buf ( n2830 , R_31b_1d9d0c28 );
buf ( n2831 , R_3c6_1d9d7c08 );
buf ( n2832 , R_792_1dfbdc48 );
buf ( n2833 , R_54b_1dda6a88 );
buf ( n2834 , R_6bd_1dfb5228 );
buf ( n2835 , R_b50_1e6b2f28 );
buf ( n2836 , R_a61_1e189968 );
buf ( n2837 , R_b8b_1e6b5408 );
buf ( n2838 , R_b80_1e6b4d28 );
buf ( n2839 , R_33c_1d9d20c8 );
buf ( n2840 , R_3c3_1d9d7528 );
buf ( n2841 , R_666_1dfb20c8 );
buf ( n2842 , R_c2a_1e6bbc68 );
buf ( n2843 , R_359_1d9d32e8 );
buf ( n2844 , R_415_1d9da868 );
buf ( n2845 , R_5da_1ddac8e8 );
buf ( n2846 , R_577_1dda8608 );
buf ( n2847 , R_637_1dfafe68 );
buf ( n2848 , R_9f7_1e185728 );
buf ( n2849 , R_570_1dda81a8 );
buf ( n2850 , R_9f6_1e185b88 );
buf ( n2851 , R_9f8_1e1857c8 );
buf ( n2852 , R_a6e_1e18a688 );
buf ( n2853 , R_73d_1dfba228 );
buf ( n2854 , R_293_1d9fb6c8 );
buf ( n2855 , R_884_1e096ee8 );
buf ( n2856 , R_3a2_1d9d6588 );
buf ( n2857 , R_9f9_1e185868 );
buf ( n2858 , R_957_1e17f328 );
buf ( n2859 , R_ab6_1e6b5fe8 );
buf ( n2860 , R_760_1dfbb808 );
buf ( n2861 , R_a21_1e187168 );
buf ( n2862 , R_bb7_1e6b6f88 );
buf ( n2863 , R_9eb_1e184fa8 );
buf ( n2864 , R_a3f_1e188428 );
buf ( n2865 , R_747_1dfba868 );
buf ( n2866 , R_4bf_1dda1308 );
buf ( n2867 , R_3d7_1d9d81a8 );
buf ( n2868 , R_4a4_1dda0228 );
buf ( n2869 , R_441_1d9dc3e8 );
buf ( n2870 , R_7ce_1e090228 );
buf ( n2871 , R_85a_1e0959a8 );
buf ( n2872 , R_66f_1dfb2168 );
buf ( n2873 , R_9ea_1e185408 );
buf ( n2874 , R_9ec_1e185048 );
buf ( n2875 , R_a3b_1e1881a8 );
buf ( n2876 , R_ad4_1e6ae1a8 );
buf ( n2877 , R_b94_1e6b59a8 );
buf ( n2878 , R_467_1d9ddba8 );
buf ( n2879 , R_96e_1e180688 );
buf ( n2880 , R_323_1d9d1128 );
buf ( n2881 , R_6ea_1dfb7348 );
buf ( n2882 , R_6ca_1dfb5f48 );
buf ( n2883 , R_9ed_1e1850e8 );
buf ( n2884 , R_ae7_1e6aed88 );
buf ( n2885 , R_830_1e093a68 );
buf ( n2886 , R_6d9_1dfb63a8 );
buf ( n2887 , R_8e6_1e08f0a8 );
buf ( n2888 , R_6a1_1dfb40a8 );
buf ( n2889 , R_710_1dfb8608 );
buf ( n2890 , R_b41_1e6b25c8 );
buf ( n2891 , R_732_1dfba048 );
buf ( n2892 , R_6df_1dfb6768 );
buf ( n2893 , R_a11_1e186768 );
buf ( n2894 , R_a8f_1e18b628 );
buf ( n2895 , R_b97_1e6b5b88 );
buf ( n2896 , R_bc6_1e6b7de8 );
buf ( n2897 , R_4db_1dda2488 );
buf ( n2898 , R_9d7_1e184328 );
buf ( n2899 , R_b29_1e6b16c8 );
buf ( n2900 , R_57e_1dda8f68 );
buf ( n2901 , R_29a_1d9fbb28 );
buf ( n2902 , R_36f_1d9d40a8 );
buf ( n2903 , R_3e4_1d9d89c8 );
buf ( n2904 , R_7bc_1e08f1e8 );
buf ( n2905 , R_87e_1e097028 );
buf ( n2906 , R_b1c_1e6b0ea8 );
buf ( n2907 , R_aab_1e18c7a8 );
buf ( n2908 , R_96c_1e180048 );
buf ( n2909 , R_551_1dda6e48 );
buf ( n2910 , R_6d4_1dfb6088 );
buf ( n2911 , R_2af_1d9fc848 );
buf ( n2912 , R_479_1dd9e748 );
buf ( n2913 , R_5a3_1ddaa188 );
buf ( n2914 , R_672_1dfb2848 );
buf ( n2915 , R_587_1dda9008 );
buf ( n2916 , R_767_1dfbbc68 );
buf ( n2917 , R_395_1d9d5868 );
buf ( n2918 , R_3e9_1d9d8ce8 );
buf ( n2919 , R_2f8_1d9cf648 );
buf ( n2920 , R_64c_1dfb0b88 );
buf ( n2921 , R_5e1_1ddac848 );
buf ( n2922 , R_3fc_1d9d98c8 );
buf ( n2923 , R_468_1d9ddc48 );
buf ( n2924 , R_3ba_1d9d7488 );
buf ( n2925 , R_55b_1dda7488 );
buf ( n2926 , R_67e_1dfb2fc8 );
buf ( n2927 , R_8b7_1e098ec8 );
buf ( n2928 , R_879_1e096808 );
buf ( n2929 , R_b5b_1e6b3608 );
buf ( n2930 , R_a82_1e18b588 );
buf ( n2931 , R_ae5_1e6aec48 );
buf ( n2932 , R_84b_1e094b48 );
buf ( n2933 , R_99e_1e182488 );
buf ( n2934 , R_6dc_1dfb6588 );
buf ( n2935 , R_3ad_1d9d6768 );
buf ( n2936 , R_a59_1e189468 );
buf ( n2937 , R_b62_1e6ba368 );
buf ( n2938 , R_731_1dfb9aa8 );
buf ( n2939 , R_3f1_1d9d91e8 );
buf ( n2940 , R_620_1dfaf008 );
buf ( n2941 , R_67d_1dfb2a28 );
buf ( n2942 , R_adf_1e6ae888 );
buf ( n2943 , R_349_1d9d28e8 );
buf ( n2944 , R_3d1_1d9d7de8 );
buf ( n2945 , R_3f4_1d9d93c8 );
buf ( n2946 , R_80a_1e0927a8 );
buf ( n2947 , R_350_1d9d2d48 );
buf ( n2948 , R_a50_1e188ec8 );
buf ( n2949 , R_bc1_1e6b75c8 );
buf ( n2950 , R_b85_1e6b5048 );
buf ( n2951 , R_5d7_1ddac208 );
buf ( n2952 , R_7a2_1ddada68 );
buf ( n2953 , R_539_1dda5f48 );
buf ( n2954 , R_bbc_1e6b72a8 );
buf ( n2955 , R_c14_1e6ba9a8 );
buf ( n2956 , R_6c8_1dfb5908 );
buf ( n2957 , R_4c8_1dda18a8 );
buf ( n2958 , R_360_1d9d3748 );
buf ( n2959 , R_2e2_1d9ced88 );
buf ( n2960 , R_936_1e17e388 );
buf ( n2961 , R_9f3_1e1854a8 );
buf ( n2962 , R_b25_1e6b1448 );
buf ( n2963 , R_b0a_1e6b0868 );
buf ( n2964 , R_b56_1e6b87e8 );
buf ( n2965 , R_bf4_1e6b95a8 );
buf ( n2966 , R_95f_1e17f828 );
buf ( n2967 , R_3b5_1d9d6c68 );
buf ( n2968 , R_52a_1dda5fe8 );
buf ( n2969 , R_9f2_1e185908 );
buf ( n2970 , R_9f4_1e185548 );
buf ( n2971 , R_686_1dfb34c8 );
buf ( n2972 , R_2bc_1d9fd068 );
buf ( n2973 , R_7a6_1e08e928 );
buf ( n2974 , R_9ef_1e185228 );
buf ( n2975 , R_b1e_1e6b78e8 );
buf ( n2976 , R_bfb_1e6b9a08 );
buf ( n2977 , R_378_1d9d4648 );
buf ( n2978 , R_9ee_1e185688 );
buf ( n2979 , R_9f0_1e1852c8 );
buf ( n2980 , R_9f5_1e1855e8 );
buf ( n2981 , R_4bd_1dda11c8 );
buf ( n2982 , R_5af_1ddaa908 );
buf ( n2983 , R_822_1e097f28 );
buf ( n2984 , R_872_1e0968a8 );
buf ( n2985 , R_9f1_1e185368 );
buf ( n2986 , R_337_1d9d1da8 );
buf ( n2987 , R_707_1dfb8068 );
buf ( n2988 , R_755_1dfbb128 );
buf ( n2989 , R_8f9_1e09b808 );
buf ( n2990 , R_432_1d9dbf88 );
buf ( n2991 , R_8af_1e0989c8 );
buf ( n2992 , R_bc5_1e6b7848 );
buf ( n2993 , R_934_1e09dce8 );
buf ( n2994 , R_469_1d9ddce8 );
buf ( n2995 , R_572_1dda87e8 );
buf ( n2996 , R_863_1e095a48 );
buf ( n2997 , R_958_1e17f3c8 );
buf ( n2998 , R_742_1dfbaa48 );
buf ( n2999 , R_2a5_1d9fc208 );
buf ( n3000 , R_a9a_1e18c208 );
buf ( n3001 , R_af9_1e6af8c8 );
buf ( n3002 , R_9c1_1e183568 );
buf ( n3003 , R_83c_1e0941e8 );
buf ( n3004 , R_a81_1e18ad68 );
buf ( n3005 , R_c19_1e6bacc8 );
buf ( n3006 , R_91c_1e09cde8 );
buf ( n3007 , R_4ac_1dda0728 );
buf ( n3008 , R_bf8_1e6b9828 );
buf ( n3009 , R_5be_1dda7168 );
buf ( n3010 , R_93b_1e17e1a8 );
buf ( n3011 , R_63c_1dfb0188 );
buf ( n3012 , R_7e1_1e090908 );
buf ( n3013 , R_7ba_1e08f5a8 );
buf ( n3014 , R_6b2_1dfb5048 );
buf ( n3015 , R_4dc_1dda2528 );
buf ( n3016 , R_79e_1e08e428 );
buf ( n3017 , R_492_1dd9fbe8 );
buf ( n3018 , R_750_1dfbae08 );
buf ( n3019 , R_9d8_1e1843c8 );
buf ( n3020 , R_365_1d9d3a68 );
buf ( n3021 , R_994_1e181948 );
buf ( n3022 , R_95c_1e17f648 );
buf ( n3023 , R_2ff_1d9cfaa8 );
buf ( n3024 , R_89b_1e097d48 );
buf ( n3025 , R_827_1e0934c8 );
buf ( n3026 , R_332_1d9d1f88 );
buf ( n3027 , R_9a7_1e182528 );
buf ( n3028 , R_834_1e093ce8 );
buf ( n3029 , R_30b_1d9d0228 );
buf ( n3030 , R_86b_1e095f48 );
buf ( n3031 , R_649_1dfb09a8 );
buf ( n3032 , R_a1d_1e186ee8 );
buf ( n3033 , R_b59_1e6b34c8 );
buf ( n3034 , R_bb3_1e6b6d08 );
buf ( n3035 , R_796_1e08e1a8 );
buf ( n3036 , R_941_1e17e568 );
buf ( n3037 , R_be9_1e6b8ec8 );
buf ( n3038 , R_485_1dd9eec8 );
buf ( n3039 , R_317_1d9d09a8 );
buf ( n3040 , R_8a3_1e098248 );
buf ( n3041 , R_49e_1dda0368 );
buf ( n3042 , R_9c0_1e1834c8 );
buf ( n3043 , R_32c_1d9d16c8 );
buf ( n3044 , R_6d6_1dfb66c8 );
buf ( n3045 , R_a15_1e1869e8 );
buf ( n3046 , R_33e_1d9d2708 );
buf ( n3047 , R_38c_1d9d52c8 );
buf ( n3048 , R_75b_1dfbb4e8 );
buf ( n3049 , R_ac4_1e18d748 );
buf ( n3050 , R_5d9_1ddac348 );
buf ( n3051 , R_546_1dda6c68 );
buf ( n3052 , R_2be_1d9fd6a8 );
buf ( n3053 , R_b76_1e6b4be8 );
buf ( n3054 , R_975_1e1805e8 );
buf ( n3055 , R_5c3_1ddab588 );
buf ( n3056 , R_500_1dda3ba8 );
buf ( n3057 , R_889_1e097208 );
buf ( n3058 , R_988_1e1811c8 );
buf ( n3059 , R_c2c_1e6bb8a8 );
buf ( n3060 , R_b98_1e6b5c28 );
buf ( n3061 , R_47d_1dd9e9c8 );
buf ( n3062 , R_417_1d9da9a8 );
buf ( n3063 , R_819_1e092c08 );
buf ( n3064 , R_8f8_1e09b768 );
buf ( n3065 , R_942_1e17eb08 );
buf ( n3066 , R_ad1_1e6adfc8 );
buf ( n3067 , R_8ce_1e09a228 );
buf ( n3068 , R_563_1dda7988 );
buf ( n3069 , R_2e8_1d9cec48 );
buf ( n3070 , R_838_1e093f68 );
buf ( n3071 , R_aee_1e187c08 );
buf ( n3072 , R_641_1dfb04a8 );
buf ( n3073 , R_c16_1e6b41e8 );
buf ( n3074 , R_6c3_1dfb55e8 );
buf ( n3075 , R_5f3_1ddad388 );
buf ( n3076 , R_558_1dda72a8 );
buf ( n3077 , R_821_1e093108 );
buf ( n3078 , R_a5f_1e189828 );
buf ( n3079 , R_3cd_1d9d7b68 );
buf ( n3080 , R_80f_1e0925c8 );
buf ( n3081 , R_724_1dfb9288 );
buf ( n3082 , R_848_1e094968 );
buf ( n3083 , R_9bf_1e183428 );
buf ( n3084 , R_a19_1e186c68 );
buf ( n3085 , R_baf_1e6b6a88 );
buf ( n3086 , R_64a_1dfb0f48 );
buf ( n3087 , R_aa8_1e18c5c8 );
buf ( n3088 , R_6be_1dfb57c8 );
buf ( n3089 , R_481_1dd9ec48 );
buf ( n3090 , R_428_1d9db448 );
buf ( n3091 , R_be6_1e6b91e8 );
buf ( n3092 , R_44f_1d9dcca8 );
buf ( n3093 , R_5b4_1ddaac28 );
buf ( n3094 , R_629_1dfaf5a8 );
buf ( n3095 , R_78f_1dfbd568 );
buf ( n3096 , R_91f_1e09cfc8 );
buf ( n3097 , R_858_1e095368 );
buf ( n3098 , R_afb_1e6afa08 );
buf ( n3099 , R_3fb_1d9d9828 );
buf ( n3100 , R_922_1e091628 );
buf ( n3101 , R_916_1e09cf28 );
buf ( n3102 , R_8a1_1e098108 );
buf ( n3103 , R_8db_1e09a548 );
buf ( n3104 , R_b32_1e6b2168 );
buf ( n3105 , R_411_1d9da5e8 );
buf ( n3106 , R_6b0_1dfb4a08 );
buf ( n3107 , R_5d1_1ddabe48 );
buf ( n3108 , R_7df_1e0907c8 );
buf ( n3109 , R_b04_1e6affa8 );
buf ( n3110 , R_45a_1d9dd888 );
buf ( n3111 , R_814_1e0928e8 );
buf ( n3112 , R_665_1dfb1b28 );
buf ( n3113 , R_69e_1dfb43c8 );
buf ( n3114 , R_b42_1e6b2b68 );
buf ( n3115 , R_555_1dda70c8 );
buf ( n3116 , R_374_1d9d43c8 );
buf ( n3117 , R_352_1d9d3388 );
buf ( n3118 , R_2a6_1d9fc7a8 );
buf ( n3119 , R_756_1dfbb6c8 );
buf ( n3120 , R_bd6_1e6b3568 );
buf ( n3121 , R_baa_1e18d888 );
buf ( n3122 , R_5b9_1ddaaf48 );
buf ( n3123 , R_3ec_1d9d8ec8 );
buf ( R_61e_1dfaf3c8 , C0 );
buf ( R_8f7_1e09b6c8 , n10614 );
buf ( R_714_1dfb8888 , n10616 );
buf ( R_951_1e17ef68 , n10620 );
buf ( R_28c_1d9fb268 , n11371 );
buf ( R_9be_1e183888 , C0 );
buf ( R_9ab_1e1827a8 , n11372 );
buf ( R_30f_1d9d04a8 , n11373 );
buf ( R_959_1e17f468 , n16580 );
buf ( R_b13_1e6b0908 , n16581 );
buf ( R_519_1dda4b48 , n23930 );
buf ( R_92d_1e09d888 , n31013 );
buf ( R_c06_1e6bafe8 , C0 );
buf ( R_8c6_1e099d28 , C0 );
buf ( R_845_1e094788 , n31181 );
buf ( R_414_1d9da7c8 , n31182 );
buf ( R_313_1d9d0728 , n31183 );
buf ( R_518_1dda4aa8 , n31184 );
buf ( R_9d9_1e184468 , n34338 );
buf ( R_4dd_1dda25c8 , n34396 );
buf ( R_59f_1dda9f08 , n34397 );
buf ( R_517_1dda4a08 , n34398 );
buf ( R_509_1dda4148 , n34465 );
buf ( R_508_1dda40a8 , n34466 );
buf ( R_401_1d9d9be8 , n34536 );
buf ( R_5f9_1ddad748 , n34543 );
buf ( R_6ef_1dfb7168 , n34544 );
buf ( R_a30_1e187ac8 , n34545 );
buf ( R_2b0_1d9fc8e8 , n34546 );
buf ( R_77c_1dfbc988 , n34547 );
buf ( R_8f1_1e09b308 , n34617 );
buf ( R_36a_1d9d4288 , C0 );
buf ( R_507_1dda4008 , n34618 );
buf ( R_516_1dda4e68 , C0 );
buf ( R_98e_1e181a88 , C0 );
buf ( R_8d5_1e09a188 , n34728 );
buf ( R_498_1dd9faa8 , n34729 );
buf ( R_68b_1dfb32e8 , n34730 );
buf ( R_773_1dfbc3e8 , n34731 );
buf ( R_45b_1d9dd428 , n34732 );
buf ( R_48d_1dd9f3c8 , n34801 );
buf ( R_5ff_1ddadb08 , n34802 );
buf ( R_705_1dfb7f28 , n34813 );
buf ( R_644_1dfb0688 , n34814 );
buf ( R_63a_1dfb0548 , C0 );
buf ( R_ac7_1e18d928 , n34815 );
buf ( R_320_1d9d0f48 , n34816 );
buf ( R_737_1dfb9e68 , n34817 );
buf ( R_506_1dda4468 , C0 );
buf ( R_647_1dfb0868 , n34818 );
buf ( R_b86_1e6bb4e8 , C0 );
buf ( R_883_1e096e48 , n34819 );
buf ( R_6a8_1dfb4508 , n34820 );
buf ( R_aa5_1e18c3e8 , n37859 );
buf ( R_440_1d9dc348 , n37860 );
buf ( R_2f9_1d9cf6e8 , n37865 );
buf ( R_69c_1dfb3d88 , n37866 );
buf ( R_65d_1dfb1628 , n37871 );
buf ( R_b0c_1e6b04a8 , n37872 );
buf ( R_b20_1e6b1128 , n37873 );
buf ( R_a2e_1e189788 , C0 );
buf ( R_905_1e09bf88 , n37939 );
buf ( R_a57_1e189328 , n37940 );
buf ( R_5f8_1ddad6a8 , n37941 );
buf ( R_54c_1dda6b28 , n37942 );
buf ( R_bd2_1e6b32e8 , C0 );
buf ( R_aca_1e6ae068 , C0 );
buf ( R_58b_1dda9288 , n37943 );
buf ( R_2e3_1d9ce928 , n37944 );
buf ( R_3e2_1d9d8d88 , C0 );
buf ( R_8f6_1e09bb28 , C0 );
buf ( R_331_1d9d19e8 , n39299 );
buf ( R_97d_1e180ae8 , n39304 );
buf ( R_5cd_1ddabbc8 , n39370 );
buf ( R_45c_1d9dd4c8 , n39371 );
buf ( R_999_1e181c68 , n39376 );
buf ( R_b99_1e6b5cc8 , n39474 );
buf ( R_948_1e17e9c8 , n39475 );
buf ( R_97e_1e181308 , C0 );
buf ( R_ab0_1e18cac8 , n39476 );
buf ( R_bb8_1e6b7028 , n39477 );
buf ( R_489_1dd9f148 , n39543 );
buf ( R_4b6_1dda1268 , C0 );
buf ( R_63f_1dfb0368 , n39544 );
buf ( R_3e7_1d9d8ba8 , n39545 );
buf ( R_2bd_1d9fd108 , n39550 );
buf ( R_81b_1e092d48 , n39551 );
buf ( R_b54_1e6b31a8 , n39552 );
buf ( R_4df_1dda2708 , n39553 );
buf ( R_bab_1e6b6808 , n39554 );
buf ( R_431_1d9db9e8 , n39620 );
buf ( R_2f2_1d9cf788 , C0 );
buf ( R_601_1ddadc48 , n39625 );
buf ( R_6e7_1dfb6c68 , n39626 );
buf ( R_bdf_1e6b8888 , n39627 );
buf ( R_656_1dfb1bc8 , C0 );
buf ( R_4e0_1dda27a8 , n39628 );
buf ( R_4de_1dda2b68 , C0 );
buf ( R_a4e_1e189288 , C0 );
buf ( R_8e1_1e09a908 , n39727 );
buf ( R_8f0_1e09b268 , n39728 );
buf ( R_299_1d9fba88 , n39735 );
buf ( R_292_1d9fb628 , n39742 );
buf ( R_4e1_1dda2848 , n39774 );
buf ( R_a7f_1e18ac28 , n39775 );
buf ( R_c04_1e6b9fa8 , n39776 );
buf ( R_3ef_1d9d90a8 , n39777 );
buf ( R_5de_1dd9f1e8 , C0 );
buf ( R_878_1e096768 , n39778 );
buf ( R_720_1dfb9008 , n39779 );
buf ( R_ad6_1e6ae7e8 , C0 );
buf ( R_9a2_1e182708 , C0 );
buf ( R_630_1dfafa08 , n39780 );
buf ( R_52f_1dda5908 , n39781 );
buf ( R_7a9_1e08e608 , n39850 );
buf ( R_976_1e180b88 , C0 );
buf ( R_439_1d9dbee8 , n39927 );
buf ( R_604_1ddade28 , n39928 );
buf ( R_530_1dda59a8 , n39929 );
buf ( R_52e_1dda5d68 , C0 );
buf ( R_7ed_1e091088 , n39987 );
buf ( R_3f2_1d9d4c88 , C0 );
buf ( R_3d4_1d9d7fc8 , n39988 );
buf ( R_84a_1e094fa8 , C0 );
buf ( R_2de_1d9ceb08 , C0 );
buf ( R_690_1dfb3608 , n39989 );
buf ( R_4cd_1dda1bc8 , n40055 );
buf ( R_531_1dda5a48 , n40147 );
buf ( R_b34_1e6b1da8 , n40148 );
buf ( R_5f7_1ddad608 , n40149 );
buf ( R_806_1e092528 , C0 );
buf ( R_a5b_1e1895a8 , n40150 );
buf ( R_718_1dfb8b08 , n40151 );
buf ( R_695_1dfb3928 , n42642 );
buf ( R_7af_1e08e9c8 , n42643 );
buf ( R_62b_1dfaf6e8 , n42644 );
buf ( R_904_1e09bee8 , n42645 );
buf ( R_501_1dda3c48 , n42677 );
buf ( R_585_1dda8ec8 , n42711 );
buf ( R_9cd_1e183ce8 , n42716 );
buf ( R_78c_1dfbd388 , n42717 );
buf ( R_392_1d9d5b88 , C0 );
buf ( R_4b4_1dda0c28 , n42718 );
buf ( R_b44_1e6b27a8 , n42719 );
buf ( R_969_1e17fe68 , n42724 );
buf ( R_40d_1d9da368 , n42790 );
buf ( R_627_1dfaf468 , n42791 );
buf ( R_67a_1dfadfc8 , C0 );
buf ( R_45d_1d9dd568 , n42822 );
buf ( R_7c1_1e08f508 , n42943 );
buf ( R_552_1dda73e8 , C0 );
buf ( R_2bf_1d9fd248 , n42944 );
buf ( R_5d4_1ddac028 , n42945 );
buf ( R_b77_1e6b4788 , n42946 );
buf ( R_3fa_1d9db088 , C0 );
buf ( R_6aa_1dfb4b48 , C0 );
buf ( R_82a_1e093ba8 , C0 );
buf ( R_3aa_1d9d6a88 , C0 );
buf ( R_300_1d9cfb48 , n42947 );
buf ( R_405_1d9d9e68 , n43013 );
buf ( R_953_1e17f0a8 , n43014 );
buf ( R_3cf_1d9d7ca8 , n43015 );
buf ( R_ac1_1e18d568 , n43119 );
buf ( R_61c_1dfaed88 , n43120 );
buf ( R_a99_1e18bc68 , n43188 );
buf ( R_4ae_1dda0fe8 , C0 );
buf ( R_aec_1e6af0a8 , n43189 );
buf ( R_af8_1e6af828 , n43190 );
buf ( R_762_1dfbbe48 , C0 );
buf ( R_3a8_1d9d6448 , n43191 );
buf ( R_4ca_1dda1ee8 , C0 );
buf ( R_6b7_1dfb4e68 , n43192 );
buf ( R_57c_1dda8928 , n43193 );
buf ( R_52b_1dda5688 , n43194 );
buf ( R_8ef_1e09b1c8 , n43195 );
buf ( R_8c5_1e099788 , n43226 );
buf ( R_8ab_1e098748 , n43227 );
buf ( R_71c_1dfb8d88 , n43228 );
buf ( R_388_1d9d5048 , n43229 );
buf ( R_b6e_1e6b46e8 , C0 );
buf ( R_9cc_1e183c48 , n43230 );
buf ( R_65b_1dfb14e8 , n43231 );
buf ( R_bbd_1e6b7348 , n43266 );
buf ( R_3b2_1d9d6f88 , C0 );
buf ( R_862_1e095ea8 , C0 );
buf ( R_4a5_1dda02c8 , n43297 );
buf ( R_90f_1e09c5c8 , n43298 );
buf ( R_702_1dfb8248 , C0 );
buf ( R_29f_1d9fbe48 , n43299 );
buf ( R_72b_1dfb96e8 , n43300 );
buf ( R_6f4_1dfb7488 , n43301 );
buf ( R_5f2_1dda8a68 , C0 );
buf ( R_a64_1e189b48 , n43302 );
buf ( R_2e9_1d9cece8 , n43307 );
buf ( R_683_1dfb2de8 , n43308 );
buf ( R_2fd_1d9cf968 , n43313 );
buf ( R_8b2_1e0990a8 , C0 );
buf ( R_5f0_1ddad1a8 , n43314 );
buf ( R_bac_1e6b68a8 , n43315 );
buf ( R_642_1dfb0a48 , C0 );
buf ( R_5f6_1d9fbda8 , C0 );
buf ( R_568_1dda7ca8 , n43316 );
buf ( R_409_1d9da0e8 , n43382 );
buf ( R_5a8_1ddaa4a8 , n43383 );
buf ( R_5e3_1ddac988 , n43384 );
buf ( R_96b_1e17ffa8 , n43385 );
buf ( R_bca_1e6b14e8 , C0 );
buf ( R_3b8_1d9d6e48 , n43386 );
buf ( R_789_1dfbd1a8 , n43485 );
buf ( R_86a_1e0963a8 , C0 );
buf ( R_416_1ddabc68 , C0 );
buf ( R_903_1e09be48 , n43486 );
buf ( R_a2d_1e1878e8 , n43495 );
buf ( R_9cb_1e183ba8 , n43496 );
buf ( R_59b_1dda9c88 , n43497 );
buf ( R_a4c_1e188c48 , n43498 );
buf ( R_79c_1dfbdd88 , n43499 );
buf ( R_888_1e097168 , n43500 );
buf ( R_2a7_1d9fc348 , n43501 );
buf ( R_7f3_1e091448 , n43502 );
buf ( R_73c_1dfba188 , n43503 );
buf ( R_bd1_1e6b7fc8 , n43584 );
buf ( R_4a6_1dda0868 , C0 );
buf ( R_3dd_1d9d8568 , n43593 );
buf ( R_346_1d9d2c08 , C0 );
buf ( R_4c4_1dda1628 , n43594 );
buf ( R_b15_1e6b0a48 , n43663 );
buf ( R_5ec_1ddacf28 , n43664 );
buf ( R_bb4_1e6b6da8 , n43665 );
buf ( R_bed_1e6b9148 , n43742 );
buf ( R_7bf_1e08f3c8 , n43743 );
buf ( R_344_1d9d25c8 , n43744 );
buf ( R_c0b_1e6ba408 , n43745 );
buf ( R_6a5_1dfb4328 , n43969 );
buf ( R_b8c_1e6b54a8 , n43970 );
buf ( R_3a1_1d9d5fe8 , n43979 );
buf ( R_7ea_1e09d928 , C0 );
buf ( R_46e_1dd9e568 , C0 );
buf ( R_8ee_1e09b628 , C0 );
buf ( R_697_1dfb3a68 , n43980 );
buf ( R_77f_1dfbcb68 , n43981 );
buf ( R_391_1d9d55e8 , n43990 );
buf ( R_746_1dfb6448 , C0 );
buf ( R_b3b_1e6b2208 , n43991 );
buf ( R_7f1_1e091308 , n44023 );
buf ( R_410_1d9da548 , n44024 );
buf ( R_700_1dfb7c08 , n44025 );
buf ( R_58f_1dda9508 , n44026 );
buf ( R_582_1dda91e8 , C0 );
buf ( R_793_1dfbd7e8 , n44027 );
buf ( R_847_1e0948c8 , n44028 );
buf ( R_95e_1e17fc88 , C0 );
buf ( R_560_1dda77a8 , n44029 );
buf ( R_9ca_1e184008 , C0 );
buf ( R_397_1d9d59a8 , n44030 );
buf ( R_46b_1d9dde28 , n44031 );
buf ( R_44e_1d9fc028 , C0 );
buf ( R_6cc_1dfb5b88 , n44032 );
buf ( R_62e_1dfafdc8 , C0 );
buf ( R_2b1_1d9fc988 , n44037 );
buf ( R_6f9_1dfb77a8 , n44046 );
buf ( R_af5_1e6af648 , n44114 );
buf ( R_b81_1e6b4dc8 , n44150 );
buf ( R_427_1d9db3a8 , n44151 );
buf ( R_547_1dda6808 , n44152 );
buf ( R_c1d_1e6baf48 , n44221 );
buf ( R_a2c_1e187848 , n44222 );
buf ( R_355_1d9d3068 , n44857 );
buf ( R_857_1e0952c8 , n44858 );
buf ( R_413_1d9da728 , n44859 );
buf ( R_afa_1e6afe68 , C0 );
buf ( R_adc_1e6ae6a8 , n44860 );
buf ( R_5fc_1ddad928 , n44861 );
buf ( R_c24_1e6bb3a8 , n44862 );
buf ( R_421_1d9dafe8 , n44893 );
buf ( R_892_1e17e608 , C0 );
buf ( R_70b_1dfb82e8 , n44894 );
buf ( R_aad_1e18c8e8 , n44962 );
buf ( R_3ca_1d9d8108 , C0 );
buf ( R_7ac_1e08e7e8 , n44963 );
buf ( R_8da_1e09a9a8 , C0 );
buf ( R_400_1d9d9b48 , n44964 );
buf ( R_bb0_1e6b6b28 , n44965 );
buf ( R_893_1e097848 , n44966 );
buf ( R_902_1e09c2a8 , C0 );
buf ( R_a93_1e18b8a8 , n44967 );
buf ( R_8cd_1e099c88 , n45033 );
buf ( R_861_1e095908 , n45065 );
buf ( R_3ea_1d9d9288 , C0 );
buf ( R_915_1e09c988 , n45132 );
buf ( R_844_1e0946e8 , n45133 );
buf ( R_677_1dfb2668 , n45134 );
buf ( R_602_1dfae248 , C0 );
buf ( R_39c_1d9d5cc8 , n45135 );
buf ( R_be3_1e6b8b08 , n45136 );
buf ( R_bea_1e6b9468 , C0 );
buf ( R_993_1e1818a8 , n45137 );
buf ( R_bad_1e6b6948 , n45223 );
buf ( R_88d_1e097488 , n45323 );
buf ( R_5a2_1ddaa5e8 , C0 );
buf ( R_655_1dfb1128 , n45328 );
buf ( R_4ad_1dda07c8 , n45398 );
buf ( R_493_1dd9f788 , n45399 );
buf ( R_894_1e0978e8 , n45400 );
buf ( R_668_1dfb1d08 , n45401 );
buf ( R_730_1dfb9a08 , n45402 );
buf ( R_7dc_1e0905e8 , n45403 );
buf ( R_abd_1e18d2e8 , n45471 );
buf ( R_662_1dfb1e48 , C0 );
buf ( R_a7c_1e18aa48 , n45472 );
buf ( R_5cf_1ddabd08 , n45473 );
buf ( R_328_1d9d1448 , n45474 );
buf ( R_741_1dfba4a8 , n45483 );
buf ( R_9a6_1e182988 , C0 );
buf ( R_36d_1d9d3f68 , n45521 );
buf ( R_308_1d9d0048 , n45522 );
buf ( R_95b_1e17f5a8 , n45523 );
buf ( R_b63_1e6b3b08 , n45524 );
buf ( R_2da_1d9ce888 , C0 );
buf ( R_5dc_1ddac528 , n45525 );
buf ( R_49f_1dd9ff08 , n45526 );
buf ( R_895_1e097988 , n45593 );
buf ( R_761_1dfbb8a8 , n45624 );
buf ( R_2e4_1d9ce9c8 , n45625 );
buf ( R_ab5_1e18cde8 , n45693 );
buf ( R_c28_1e6bb628 , n45694 );
buf ( R_8d4_1e09a0e8 , n45695 );
buf ( R_a8c_1e18b448 , n45696 );
buf ( R_597_1dda9a08 , n45697 );
buf ( R_5c4_1ddab628 , n45698 );
buf ( R_384_1d9d4dc8 , n45699 );
buf ( R_31c_1d9d0cc8 , n45700 );
buf ( R_987_1e181128 , n45701 );
buf ( R_b2e_1e6b1ee8 , C0 );
buf ( R_2f3_1d9cf328 , n45702 );
buf ( R_6cf_1dfb5d68 , n45703 );
buf ( R_6e4_1dfb6a88 , n45704 );
buf ( R_357_1d9d31a8 , n45705 );
buf ( R_3c1_1d9d73e8 , n45714 );
buf ( R_5e7_1ddacc08 , n45715 );
buf ( R_974_1e180548 , n45716 );
buf ( R_61a_1dfaf148 , C0 );
buf ( R_3f8_1d9d9648 , n45717 );
buf ( R_802_1e0922a8 , C0 );
buf ( R_593_1dda9788 , n45718 );
buf ( R_a69_1e189e68 , n45804 );
buf ( R_a87_1e18b128 , n45805 );
buf ( R_a5d_1e1896e8 , n45840 );
buf ( R_a2b_1e1877a8 , n45841 );
buf ( R_671_1dfb22a8 , n45846 );
buf ( R_4cf_1dda1d08 , n45847 );
buf ( R_420_1d9daf48 , n45848 );
buf ( R_6bc_1dfb5188 , n45849 );
buf ( R_43f_1d9dc2a8 , n45850 );
buf ( R_692_1dfb3c48 , C0 );
buf ( R_80b_1e092348 , n45851 );
buf ( R_882_1e0972a8 , C0 );
buf ( R_871_1e096308 , n45918 );
buf ( R_2c2_1d9fd928 , C0 );
buf ( R_2ce_1d9cfa08 , C0 );
buf ( R_a9c_1e18be48 , n45919 );
buf ( R_768_1dfbbd08 , n45920 );
buf ( R_56d_1dda7fc8 , n45987 );
buf ( R_34c_1d9d2ac8 , n45988 );
buf ( R_b8f_1e6b5688 , n45989 );
buf ( R_b07_1e6b0188 , n45990 );
buf ( R_6b5_1dfb4d28 , n46050 );
buf ( R_5ae_1ddaad68 , C0 );
buf ( R_2df_1d9ce6a8 , n46051 );
buf ( R_674_1dfb2488 , n46052 );
buf ( R_608_1dfae108 , n46053 );
buf ( R_ad3_1e6ae108 , n46054 );
buf ( R_505_1dda3ec8 , n46121 );
buf ( R_8bf_1e0993c8 , n46122 );
buf ( R_542_1dda69e8 , C0 );
buf ( R_7f6_1e091b28 , C0 );
buf ( R_504_1dda3e28 , n46123 );
buf ( R_8a7_1e0984c8 , n46124 );
buf ( R_76a_1dfbc5c8 , C0 );
buf ( R_937_1e09dec8 , n46125 );
buf ( R_6fb_1dfb78e8 , n46126 );
buf ( R_3b0_1d9d6948 , n46127 );
buf ( R_2c0_1d9fd2e8 , n46128 );
buf ( R_37c_1d9d48c8 , n46129 );
buf ( R_782_1dfbd248 , C0 );
buf ( R_503_1dda3d88 , n46130 );
buf ( R_82e_1e093e28 , C0 );
buf ( R_8bb_1e099148 , n46131 );
buf ( R_430_1d9db948 , n46132 );
buf ( R_5cb_1ddaba88 , n46133 );
buf ( R_ae6_1e6af1e8 , C0 );
buf ( R_7a3_1e08e248 , n46134 );
buf ( R_b78_1e6b4828 , n46135 );
buf ( R_bc9_1e6b7ac8 , n46204 );
buf ( R_380_1d9d4b48 , n46205 );
buf ( R_33d_1d9d2168 , n46261 );
buf ( R_8e0_1e09a868 , n46262 );
buf ( R_3c7_1d9d77a8 , n46263 );
buf ( R_2b2_1d9fcf28 , C0 );
buf ( R_618_1dfaeb08 , n46264 );
buf ( R_823_1e093248 , n46265 );
buf ( R_89e_1e098428 , C0 );
buf ( R_502_1dda41e8 , C0 );
buf ( R_b6f_1e6b4288 , n46266 );
buf ( R_c00_1e6b9d28 , n46267 );
buf ( R_98d_1e1814e8 , n46272 );
buf ( R_28b_1d9fb1c8 , n46281 );
buf ( R_a55_1e1891e8 , n46316 );
buf ( R_3c4_1d9d75c8 , n46317 );
buf ( R_40c_1d9da2c8 , n46318 );
buf ( R_2d2_1d9ce388 , C0 );
buf ( R_c21_1e6bb1c8 , n46387 );
buf ( R_b3d_1e6b2348 , n46480 );
buf ( R_877_1e0966c8 , n46481 );
buf ( R_855_1e095188 , n46513 );
buf ( R_41d_1d9dad68 , n46544 );
buf ( R_438_1d9dbe48 , n46545 );
buf ( R_2d6_1d9ce608 , C0 );
buf ( R_7da_1e0909a8 , C0 );
buf ( R_6f6_1dfb7ac8 , C0 );
buf ( R_9aa_1e182e88 , C0 );
buf ( R_b47_1e6b2988 , n46546 );
buf ( R_a2a_1e6b3ce8 , C0 );
buf ( R_41f_1d9daea8 , n46547 );
buf ( R_ae4_1e6aeba8 , n46548 );
buf ( R_a79_1e18a868 , n46583 );
buf ( R_3a3_1d9d6128 , n46584 );
buf ( R_5bd_1ddab1c8 , n46651 );
buf ( R_301_1d9cfbe8 , n46656 );
buf ( R_298_1d9fb9e8 , n46663 );
buf ( R_bb9_1e6b70c8 , n46698 );
buf ( R_82d_1e093888 , n46730 );
buf ( R_404_1d9d9dc8 , n46731 );
buf ( R_a62_1e189f08 , C0 );
buf ( R_93c_1e17e248 , n46732 );
buf ( R_62d_1dfaf828 , n46737 );
buf ( R_579_1dda8748 , n46804 );
buf ( R_452_1ddac3e8 , C0 );
buf ( R_54d_1dda6bc8 , n46836 );
buf ( R_4d9_1dda2348 , n46902 );
buf ( R_4d4_1dda2028 , n46903 );
buf ( R_6c1_1dfb54a8 , n46963 );
buf ( R_379_1d9d46e8 , n46972 );
buf ( R_34e_1d9d3108 , C0 );
buf ( R_94a_1e097ca8 , C0 );
buf ( R_74b_1dfbaae8 , n46973 );
buf ( R_ade_1e6aece8 , C0 );
buf ( R_79f_1e08dfc8 , n46974 );
buf ( R_797_1dfbda68 , n46975 );
buf ( R_943_1e17e6a8 , n46976 );
buf ( R_653_1dfb0fe8 , n46977 );
buf ( R_3d8_1d9d8248 , n46978 );
buf ( R_b61_1e6b39c8 , n47014 );
buf ( R_bc4_1e6b77a8 , n47015 );
buf ( R_a02_1e186308 , C0 );
buf ( R_368_1d9d3c48 , n47016 );
buf ( R_35e_1d9d3b08 , C0 );
buf ( R_7fe_1e092028 , C0 );
buf ( R_499_1dd9fb48 , n47082 );
buf ( R_680_1dfb2c08 , n47083 );
buf ( R_2a8_1d9fc3e8 , n47084 );
buf ( R_6ec_1dfb6f88 , n47085 );
buf ( R_776_1dfbcac8 , C0 );
buf ( R_b5e_1e6b0368 , C0 );
buf ( R_635_1dfafd28 , n47090 );
buf ( R_7fa_1e091da8 , C0 );
buf ( R_af7_1e6af788 , n47091 );
buf ( R_8c4_1e0996e8 , n47092 );
buf ( R_408_1d9da048 , n47093 );
buf ( R_ab9_1e18d068 , n47128 );
buf ( R_6a2_1dfb61c8 , C0 );
buf ( R_291_1d9fb588 , n47135 );
buf ( R_7b8_1e08ef68 , n47136 );
buf ( R_8b6_1e08e6a8 , C0 );
buf ( R_48a_1dda0d68 , C0 );
buf ( R_6c7_1dfb5868 , n47137 );
buf ( R_c10_1e6ba728 , n47138 );
buf ( R_bf1_1e6b93c8 , n47174 );
buf ( R_4d6_1dd9e2e8 , C0 );
buf ( R_5b3_1ddaab88 , n47175 );
buf ( R_771_1dfbc2a8 , n47206 );
buf ( R_af1_1e6af3c8 , n47243 );
buf ( R_6e1_1dfb68a8 , n47252 );
buf ( R_a9f_1e18c028 , n47253 );
buf ( R_b17_1e6b0b88 , n47254 );
buf ( R_b30_1e6b1b28 , n47255 );
buf ( R_bde_1e6b37e8 , C0 );
buf ( R_998_1e181bc8 , n47256 );
buf ( R_a4a_1e189008 , C0 );
buf ( R_48e_1dd9f968 , C0 );
buf ( R_688_1dfb3108 , n47257 );
buf ( R_810_1e092668 , n47258 );
buf ( R_75c_1dfbb588 , n47259 );
buf ( R_3bb_1d9d7028 , n47260 );
buf ( R_c2e_1e17f008 , C0 );
buf ( R_5d2_1d9db308 , C0 );
buf ( R_32e_1d9d1d08 , C0 );
buf ( R_580_1dda8ba8 , n47261 );
buf ( R_453_1d9dcf28 , n47262 );
buf ( R_83a_1e0913a8 , C0 );
buf ( R_41e_1d9dc988 , C0 );
buf ( R_97c_1e180a48 , n47263 );
buf ( R_5b8_1ddaaea8 , n47264 );
buf ( R_363_1d9d3928 , n47265 );
buf ( R_94e_1ddadce8 , C0 );
buf ( R_7c4_1e08f6e8 , n47266 );
buf ( R_52c_1dda5728 , n47267 );
buf ( R_aa2_1e18c708 , C0 );
buf ( R_625_1dfaf328 , n47272 );
buf ( R_4b7_1dda0e08 , n47273 );
buf ( R_55d_1dda75c8 , n47305 );
buf ( R_b0e_1e6b0ae8 , C0 );
buf ( R_425_1d9db268 , n47336 );
buf ( R_30c_1d9d02c8 , n47337 );
buf ( R_3db_1d9d8428 , n47338 );
buf ( R_a48_1e1889c8 , n47339 );
buf ( R_aaf_1e18ca28 , n47340 );
buf ( R_5ad_1ddaa7c8 , n47407 );
buf ( R_589_1dda9148 , n47474 );
buf ( R_338_1d9d1e48 , n47475 );
buf ( R_832_1e0940a8 , C0 );
buf ( R_790_1dfbd608 , n47476 );
buf ( R_318_1d9d0a48 , n47477 );
buf ( R_869_1e095e08 , n47544 );
buf ( R_6d3_1dfb5fe8 , n47545 );
buf ( R_60c_1dfae388 , n47546 );
buf ( R_56a_1dda82e8 , C0 );
buf ( R_887_1e0970c8 , n47547 );
buf ( R_815_1e092988 , n47579 );
buf ( R_66b_1dfb1ee8 , n47580 );
buf ( R_a34_1e187d48 , n47581 );
buf ( R_40f_1d9da4a8 , n47582 );
buf ( R_ac3_1e18d6a8 , n47583 );
buf ( R_324_1d9d11c8 , n47584 );
buf ( R_614_1dfae888 , n47585 );
buf ( R_752_1dfbb448 , C0 );
buf ( R_4c0_1dda13a8 , n47586 );
buf ( R_7d9_1e090408 , n47617 );
buf ( R_ad0_1e18dec8 , n47618 );
buf ( R_bee_1e6b96e8 , C0 );
buf ( R_736_1dfba2c8 , C0 );
buf ( R_727_1dfb9468 , n47619 );
buf ( R_a8a_1e18b808 , C0 );
buf ( R_933_1e09dc48 , n47620 );
buf ( R_8b1_1e098b08 , n47686 );
buf ( R_606_1dfae4c8 , C0 );
buf ( R_927_1e09d4c8 , n47687 );
buf ( R_a7a_1e18ae08 , C0 );
buf ( R_333_1d9d1b28 , n47688 );
buf ( R_968_1e17fdc8 , n47689 );
buf ( R_574_1dda8428 , n47690 );
buf ( R_836_1e094328 , C0 );
buf ( R_757_1dfbb268 , n47691 );
buf ( R_2db_1d9ce428 , n47692 );
buf ( R_af4_1e6af5a8 , n47693 );
buf ( R_454_1d9dcfc8 , n47694 );
buf ( R_412_1d9dab88 , C0 );
buf ( R_709_1dfb81a8 , n47703 );
buf ( R_8a4_1e0982e8 , n47704 );
buf ( R_c1b_1e6bae08 , n47705 );
buf ( R_846_1e094d28 , C0 );
buf ( R_3ff_1d9d9aa8 , n47706 );
buf ( R_76e_1dfbdec8 , C0 );
buf ( R_33f_1d9d22a8 , n47707 );
buf ( R_4af_1dda0908 , n47708 );
buf ( R_a67_1e189d28 , n47709 );
buf ( R_616_1dfaeec8 , C0 );
buf ( R_b49_1e6b2ac8 , n47801 );
buf ( R_2f4_1d9cf3c8 , n47802 );
buf ( R_426_1d9db808 , C0 );
buf ( R_2e5_1d9cea68 , n47807 );
buf ( R_bb5_1e6b6e48 , n47842 );
buf ( R_7b6_1e08f328 , C0 );
buf ( R_751_1dfbaea8 , n47873 );
buf ( R_bd0_1e6b7f28 , n47874 );
buf ( R_610_1dfae608 , n47875 );
buf ( R_918_1e09cb68 , n47876 );
buf ( R_35c_1d9d34c8 , n47877 );
buf ( R_924_1e09d2e8 , n47878 );
buf ( R_912_1e09cca8 , C0 );
buf ( R_77d_1dfbca28 , n47909 );
buf ( R_774_1dfbc488 , n47910 );
buf ( R_a71_1e18a368 , n47978 );
buf ( R_32d_1d9d1768 , n48016 );
buf ( R_99d_1e181ee8 , n48021 );
buf ( R_87d_1e096a88 , n48088 );
buf ( R_472_1dd9e7e8 , C0 );
buf ( R_b2a_1e6b1c68 , C0 );
buf ( R_56f_1dda8108 , n48089 );
buf ( R_b87_1e6b5188 , n48090 );
buf ( R_921_1e09d108 , n48157 );
buf ( R_375_1d9d4468 , n48166 );
buf ( R_576_1dda8ce8 , C0 );
buf ( R_b82_1e6b5368 , C0 );
buf ( R_39e_1d9d6308 , C0 );
buf ( R_856_1e095728 , C0 );
buf ( R_6c2_1dfb5a48 , C0 );
buf ( R_2c3_1d9fd4c8 , n48167 );
buf ( R_90b_1e09c348 , n48168 );
buf ( R_92f_1e09d9c8 , n48169 );
buf ( R_38e_1d9d5908 , C0 );
buf ( R_b9e_1e18d388 , C0 );
buf ( R_8cc_1e099be8 , n48170 );
buf ( R_860_1e095868 , n48171 );
buf ( R_c09_1e6ba2c8 , n48207 );
buf ( R_b09_1e6b02c8 , n48243 );
buf ( R_521_1dda5048 , n48310 );
buf ( R_b4a_1e6b3068 , C0 );
buf ( R_88c_1e0973e8 , n48311 );
buf ( R_520_1dda4fa8 , n48312 );
buf ( R_8b5_1e098d88 , n48378 );
buf ( R_b5d_1e6b3748 , n48447 );
buf ( R_843_1e094648 , n48448 );
buf ( R_633_1dfafbe8 , n48449 );
buf ( R_7c2_1e08faa8 , C0 );
buf ( R_6d8_1dfb6308 , n48450 );
buf ( R_38d_1d9d5368 , n48459 );
buf ( R_7e7_1e090cc8 , n48460 );
buf ( R_bfc_1e6b9aa8 , n48461 );
buf ( R_841_1e094508 , n48493 );
buf ( R_a96_1e18bf88 , C0 );
buf ( R_7e5_1e090b88 , n48539 );
buf ( R_51f_1dda4f08 , n48540 );
buf ( R_949_1e17ea68 , n48572 );
buf ( R_b5a_1e6b3a68 , C0 );
buf ( R_2e0_1d9ce748 , n48573 );
buf ( R_acd_1e18dce8 , n48608 );
buf ( R_70f_1dfb8568 , n48609 );
buf ( R_c15_1e6baa48 , n48645 );
buf ( R_310_1d9d0548 , n48646 );
buf ( R_bf5_1e6b9648 , n48715 );
buf ( R_314_1d9d07c8 , n48716 );
buf ( R_6af_1dfb4968 , n48717 );
buf ( R_445_1d9dc668 , n48790 );
buf ( R_658_1dfb1308 , n48791 );
buf ( R_a6c_1e18a048 , n48792 );
buf ( R_2c1_1d9fd388 , n48797 );
buf ( R_2b3_1d9fcac8 , n48798 );
buf ( R_6de_1dfb6bc8 , C0 );
buf ( R_9b9_1e183068 , n48803 );
buf ( R_6ad_1dfb4828 , n48863 );
buf ( R_548_1dda68a8 , n48864 );
buf ( R_4c9_1dda1948 , n48930 );
buf ( R_51e_1dda5368 , C0 );
buf ( R_96a_1e180408 , C0 );
buf ( R_455_1d9dd068 , n48996 );
buf ( R_8d3_1e09a048 , n48997 );
buf ( R_bb1_1e6b6bc8 , n49032 );
buf ( R_7d7_1e0902c8 , n49033 );
buf ( R_6a0_1dfb4008 , n49034 );
buf ( R_b79_1e6b48c8 , n49103 );
buf ( R_565_1dda7ac8 , n49170 );
buf ( R_586_1dda9468 , C0 );
buf ( R_4a7_1dda0408 , n49171 );
buf ( R_b70_1e6b4328 , n49172 );
buf ( R_661_1dfb18a8 , n49177 );
buf ( R_2d3_1d9fdec8 , n49178 );
buf ( R_ad9_1e6ae4c8 , n49246 );
buf ( R_a85_1e18afe8 , n49281 );
buf ( R_a77_1e18a728 , n49282 );
buf ( R_2d7_1d9ce1a8 , n49283 );
buf ( R_7b3_1e08ec48 , n49284 );
buf ( R_870_1e096268 , n49285 );
buf ( R_43e_1d9dc708 , C0 );
buf ( R_6db_1dfb64e8 , n49286 );
buf ( R_807_1e0920c8 , n49287 );
buf ( R_a74_1e18a548 , n49288 );
buf ( R_bf9_1e6b98c8 , n49324 );
buf ( R_321_1d9d0fe8 , n49329 );
buf ( R_a53_1e1890a8 , n49330 );
buf ( R_4e3_1dda2988 , n49331 );
buf ( R_831_1e093b08 , n49398 );
buf ( R_66e_1dfb25c8 , C0 );
buf ( R_ac6_1e18dd88 , C0 );
buf ( R_55a_1dda78e8 , C0 );
buf ( R_4c6_1dda1c68 , C0 );
buf ( R_4e4_1dda2a28 , n49399 );
buf ( R_4e2_1dda2de8 , C0 );
buf ( R_c22_1e6b55e8 , C0 );
buf ( R_92c_1e09d7e8 , n49400 );
buf ( R_7c9_1e08fa08 , n49431 );
buf ( R_623_1dfaf1e8 , n49432 );
buf ( R_b58_1e6b3428 , n49433 );
buf ( R_370_1d9d4148 , n49434 );
buf ( R_3be_1d9d7708 , C0 );
buf ( R_4e5_1dda2ac8 , n49466 );
buf ( R_a03_1e185ea8 , n49467 );
buf ( R_c12_1e6bad68 , C0 );
buf ( R_456_1d9dd608 , C0 );
buf ( R_bf2_1e6b9968 , C0 );
buf ( R_6a7_1dfb4468 , n49468 );
buf ( R_c30_1e6bbb28 , n49469 );
buf ( R_40b_1d9da228 , n49470 );
buf ( R_42f_1d9db8a8 , n49471 );
buf ( R_68d_1dfb3428 , n49531 );
buf ( R_735_1dfb9d28 , n49540 );
buf ( R_78d_1dfbd428 , n49606 );
buf ( R_8df_1e09a7c8 , n49607 );
buf ( R_41c_1d9dacc8 , n49608 );
buf ( R_46f_1dd9e108 , n49609 );
buf ( R_2a9_1d9fc488 , n49614 );
buf ( R_81e_1e093428 , C0 );
buf ( R_5e0_1ddac7a8 , n49615 );
buf ( R_462_1d9ddd88 , C0 );
buf ( R_60a_1dfae748 , C0 );
buf ( R_5a7_1ddaa408 , n49616 );
buf ( R_403_1d9d9d28 , n49617 );
buf ( R_2c6_1d9fdba8 , C0 );
buf ( R_7e3_1e090a48 , n49618 );
buf ( R_7ee_1e09c528 , C0 );
buf ( R_706_1dfb84c8 , C0 );
buf ( R_c17_1e6bab88 , n49619 );
buf ( R_c1f_1e6bb088 , n49620 );
buf ( R_b93_1e6b5908 , n49621 );
buf ( R_854_1e0950e8 , n49622 );
buf ( R_b9f_1e6b6088 , n49623 );
buf ( R_8e5_1e09ab88 , n49654 );
buf ( R_437_1d9dbda8 , n49655 );
buf ( R_612_1dfaec48 , C0 );
buf ( R_816_1e0931a8 , C0 );
buf ( R_b19_1e6b0cc8 , n49691 );
buf ( R_73b_1dfba0e8 , n49692 );
buf ( R_a44_1e188748 , n49693 );
buf ( R_93e_1e17e888 , C0 );
buf ( R_67c_1dfb2988 , n49694 );
buf ( R_992_1e181d08 , C0 );
buf ( R_494_1dd9f828 , n49695 );
buf ( R_3e0_1d9d8748 , n49696 );
buf ( R_7a7_1e08e4c8 , n49697 );
buf ( R_876_1e096b28 , C0 );
buf ( R_543_1dda6588 , n49698 );
buf ( R_8ae_1dfbc0c8 , C0 );
buf ( R_351_1d9d2de8 , n49736 );
buf ( R_457_1d9dd1a8 , n49737 );
buf ( R_bf6_1e6b3f68 , C0 );
buf ( R_a38_1e187fc8 , n49738 );
buf ( R_6f1_1dfb72a8 , n49747 );
buf ( R_b3e_1e6b28e8 , C0 );
buf ( R_53e_1dda6768 , C0 );
buf ( R_ac0_1e18d4c8 , n49748 );
buf ( R_763_1dfbb9e8 , n49749 );
buf ( R_c26_1e6b8ce8 , C0 );
buf ( R_650_1dfb0e08 , n49750 );
buf ( R_361_1d9d37e8 , n49788 );
buf ( R_aaa_1e187e88 , C0 );
buf ( R_b10_1e6b0728 , n49789 );
buf ( R_b2c_1e6b18a8 , n49790 );
buf ( R_5a1_1ddaa048 , n49822 );
buf ( R_be7_1e6b8d88 , n49823 );
buf ( R_b26_1e6b19e8 , C0 );
buf ( R_4a0_1dd9ffa8 , n49824 );
buf ( R_95a_1e17fa08 , C0 );
buf ( R_909_1e09c208 , n49890 );
buf ( R_463_1d9dd928 , n49891 );
buf ( R_407_1d9d9fa8 , n49892 );
buf ( R_5c5_1ddab6c8 , n49894 );
buf ( R_986_1e181588 , C0 );
buf ( R_515_1dda48c8 , n49926 );
buf ( R_5c1_1ddab448 , n49958 );
buf ( R_297_1d9fb948 , n49965 );
buf ( R_514_1dda4828 , n49966 );
buf ( R_b4c_1e6b2ca8 , n49967 );
buf ( R_973_1e1804a8 , n49968 );
buf ( R_60e_1dfae9c8 , C0 );
buf ( R_7d4_1e0900e8 , n49969 );
buf ( R_7c7_1e08f8c8 , n49970 );
buf ( R_513_1dda4788 , n49971 );
buf ( R_65f_1dfb1768 , n49972 );
buf ( R_9b5_1e182de8 , n49977 );
buf ( R_2ee_1d9cf508 , C0 );
buf ( R_91b_1e09cd48 , n49978 );
buf ( R_af6_1e6afbe8 , C0 );
buf ( R_83d_1e094288 , n50045 );
buf ( R_8c3_1e099648 , n50046 );
buf ( R_458_1d9dd248 , n50047 );
buf ( R_512_1dda4be8 , C0 );
buf ( R_ba6_1e6b69e8 , C0 );
buf ( R_5e5_1ddacac8 , n50078 );
buf ( R_57b_1dda8888 , n50079 );
buf ( R_aeb_1e6af008 , n50080 );
buf ( R_7f4_1e0914e8 , n50081 );
buf ( R_a46_1e188d88 , C0 );
buf ( R_b8d_1e6b5548 , n50117 );
buf ( R_562_1dda7de8 , C0 );
buf ( R_745_1dfba728 , n50126 );
buf ( R_557_1dda7208 , n50127 );
buf ( R_464_1d9dd9c8 , n50128 );
buf ( R_835_1e093d88 , n50160 );
buf ( R_49a_1dda00e8 , C0 );
buf ( R_7d1_1e08ff08 , n50191 );
buf ( R_911_1e09c708 , n50223 );
buf ( R_6e9_1dfb6da8 , n50232 );
buf ( R_723_1dfb91e8 , n50233 );
buf ( R_a95_1e18b9e8 , n50268 );
buf ( R_58d_1dda93c8 , n50300 );
buf ( R_a89_1e18b268 , n50335 );
buf ( R_780_1dfbcc08 , n50336 );
buf ( R_740_1dfba408 , n50337 );
buf ( R_72f_1dfb9968 , n50338 );
buf ( R_828_1e093568 , n50339 );
buf ( R_89c_1e097de8 , n50340 );
buf ( R_a32_1e188108 , C0 );
buf ( R_840_1e094468 , n50341 );
buf ( R_b37_1e6b1f88 , n50342 );
buf ( R_9db_1e1845a8 , n50343 );
buf ( R_b22_1e6b1768 , C0 );
buf ( R_9dc_1e184648 , n50344 );
buf ( R_9da_1e184a08 , C0 );
buf ( R_794_1dfbd888 , n50345 );
buf ( R_33a_1d9d2488 , C0 );
buf ( R_424_1d9db1c8 , n50346 );
buf ( R_2dc_1d9ce4c8 , n50347 );
buf ( R_a6f_1e18a228 , n50348 );
buf ( R_98c_1e181448 , n50349 );
buf ( R_6b6_1dfb52c8 , C0 );
buf ( R_908_1e09c168 , n50350 );
buf ( R_9dd_1e1846e8 , n50475 );
buf ( R_965_1e17fbe8 , n50480 );
buf ( R_28a_1d9fb128 , n50489 );
buf ( R_529_1dda5548 , n50521 );
buf ( R_40e_1d9da908 , C0 );
buf ( R_bcd_1e6b7d48 , n50557 );
buf ( R_476_1dd9ea68 , C0 );
buf ( R_393_1d9d5728 , n50558 );
buf ( R_a40_1e1884c8 , n50559 );
buf ( R_528_1dda54a8 , n50560 );
buf ( R_2fa_1d9d0188 , C0 );
buf ( R_a3c_1e188248 , n50561 );
buf ( R_868_1e095d68 , n50562 );
buf ( R_2cf_1d9fdc48 , n50563 );
buf ( R_2c4_1d9fd568 , n50564 );
buf ( R_7cc_1e08fbe8 , n50565 );
buf ( R_8fd_1e09ba88 , n50596 );
buf ( R_3d5_1d9d8068 , n50605 );
buf ( R_b64_1e6b3ba8 , n50606 );
buf ( R_527_1dda5408 , n50607 );
buf ( R_9d1_1e183f68 , n50612 );
buf ( R_46c_1d9ddec8 , n50613 );
buf ( R_2f5_1d9cf468 , n50618 );
buf ( R_839_1e094008 , n50650 );
buf ( R_554_1dda7028 , n50651 );
buf ( R_3ab_1d9d6628 , n50652 );
buf ( R_459_1d9dd2e8 , n50683 );
buf ( R_b4f_1e6b2e88 , n50684 );
buf ( R_886_1e097528 , C0 );
buf ( R_3e5_1d9d8a68 , n50693 );
buf ( R_52d_1dda57c8 , n50760 );
buf ( R_290_1d9fb4e8 , n50767 );
buf ( R_b7a_1e18cc08 , C0 );
buf ( R_526_1dda5ae8 , C0 );
buf ( R_79a_1e098e28 , C0 );
buf ( R_ba0_1e6b6128 , n50768 );
buf ( R_6d1_1dfb5ea8 , n50777 );
buf ( R_713_1dfb87e8 , n50778 );
buf ( R_685_1dfb2f28 , n50838 );
buf ( R_3fe_1d9d9f08 , C0 );
buf ( R_638_1dfaff08 , n50839 );
buf ( R_465_1d9dda68 , n50870 );
buf ( R_b91_1e6b57c8 , n50872 );
buf ( R_b53_1e6b3108 , n50873 );
buf ( R_8ad_1e098888 , n50904 );
buf ( R_59e_1dd9e068 , C0 );
buf ( R_9c5_1e1837e8 , n50909 );
buf ( R_3a9_1d9d64e8 , n50918 );
buf ( R_3b3_1d9d6b28 , n50919 );
buf ( R_2b4_1d9fcb68 , n50920 );
buf ( R_af3_1e6af508 , n50921 );
buf ( R_4f9_1dda3748 , n50953 );
buf ( R_a90_1e18b6c8 , n50954 );
buf ( R_389_1d9d50e8 , n50963 );
buf ( R_a6a_1e18a408 , C0 );
buf ( R_b1b_1e6b0e08 , n50964 );
buf ( R_4f8_1dda36a8 , n50965 );
buf ( R_b66_1e6b9be8 , C0 );
buf ( R_9d0_1e183ec8 , n50966 );
buf ( R_2e1_1d9ce7e8 , n50971 );
buf ( R_7d2_1e0904a8 , C0 );
buf ( R_803_1e091e48 , n50972 );
buf ( R_91e_1e09d428 , C0 );
buf ( R_4f7_1dda3608 , n50973 );
buf ( R_ab4_1e18cd48 , n50974 );
buf ( R_6ee_1dfb75c8 , C0 );
buf ( R_c05_1e6ba048 , n51010 );
buf ( R_704_1dfb7e88 , n51011 );
buf ( R_353_1d9d2f28 , n51012 );
buf ( R_ba7_1e6b6588 , n51013 );
buf ( R_87c_1e0969e8 , n51014 );
buf ( R_3f5_1d9d9468 , n51023 );
buf ( R_abc_1e18d248 , n51024 );
buf ( R_a83_1e18aea8 , n51025 );
buf ( R_b40_1e6b2528 , n51026 );
buf ( R_a06_1e186588 , C0 );
buf ( R_907_1e09c0c8 , n51027 );
buf ( R_664_1dfb1a88 , n51028 );
buf ( R_b71_1e6b43c8 , n51064 );
buf ( R_4f6_1ddad2e8 , C0 );
buf ( R_8b9_1e099008 , n51095 );
buf ( R_971_1e180368 , n51100 );
buf ( R_64e_1dfb11c8 , C0 );
buf ( R_679_1dfb27a8 , n51105 );
buf ( R_80c_1e0923e8 , n51106 );
buf ( R_347_1d9d27a8 , n51107 );
buf ( R_b28_1e6b1628 , n51108 );
buf ( R_7cf_1e08fdc8 , n51109 );
buf ( R_8fc_1e09b9e8 , n51110 );
buf ( R_72d_1dfb9828 , n51119 );
buf ( R_9c4_1e183748 , n51120 );
buf ( R_997_1e181b28 , n51121 );
buf ( R_85f_1e0957c8 , n51122 );
buf ( R_2d4_1d9cdfc8 , n51123 );
buf ( R_48f_1dd9f508 , n51124 );
buf ( R_adb_1e6ae608 , n51125 );
buf ( R_3b9_1d9d6ee8 , n51134 );
buf ( R_a51_1e188f68 , n51202 );
buf ( R_8cb_1e099b48 , n51203 );
buf ( R_2d8_1d9ce248 , n51204 );
buf ( R_a72_1e18a908 , C0 );
buf ( R_7f7_1e0916c8 , n51205 );
buf ( R_4b5_1dda0cc8 , n51236 );
buf ( R_88b_1e097348 , n51237 );
buf ( R_aa7_1e18c528 , n51238 );
buf ( R_699_1dfb3ba8 , n51298 );
buf ( R_68a_1dfb3748 , C0 );
buf ( R_9cf_1e183e28 , n51299 );
buf ( R_345_1d9d2668 , n51349 );
buf ( R_76b_1dfbbee8 , n51350 );
buf ( R_7aa_1e099328 , C0 );
buf ( R_5e9_1ddacd48 , n51381 );
buf ( R_a04_1e185f48 , n51382 );
buf ( R_36b_1d9d3e28 , n51383 );
buf ( R_444_1d9dc5c8 , n51384 );
buf ( R_842_1e094aa8 , C0 );
buf ( R_58a_1dda96e8 , C0 );
buf ( R_97b_1e1809a8 , n51385 );
buf ( R_5bc_1ddab128 , n51386 );
buf ( R_ae9_1e6aeec8 , n51421 );
buf ( R_74e_1dfbc348 , C0 );
buf ( R_69b_1dfb3ce8 , n51422 );
buf ( R_783_1dfbcde8 , n51423 );
buf ( R_64d_1dfb0c28 , n51428 );
buf ( R_938_1e17dfc8 , n51429 );
buf ( R_7bd_1e08f288 , n51460 );
buf ( R_7ca_1e08ffa8 , C0 );
buf ( R_482_1ddac668 , C0 );
buf ( R_2c7_1d9fd748 , n51461 );
buf ( R_621_1dfaf0a8 , n51466 );
buf ( R_9c3_1e1836a8 , n51467 );
buf ( R_309_1d9d00e8 , n51472 );
buf ( R_5f1_1ddad248 , n51504 );
buf ( R_4b8_1dda0ea8 , n51505 );
buf ( R_bcf_1e6b7e88 , n51506 );
buf ( R_824_1e0932e8 , n51507 );
buf ( R_6e6_1dfb70c8 , C0 );
buf ( R_7a4_1e08e2e8 , n51508 );
buf ( R_59d_1dda9dc8 , n51540 );
buf ( R_769_1dfbbda8 , n51606 );
buf ( R_38a_1d9d5688 , C0 );
buf ( R_4cb_1dda1a88 , n51607 );
buf ( R_8d9_1e09a408 , n51638 );
buf ( R_8d2_1e09a4a8 , C0 );
buf ( R_b24_1e6b13a8 , n51639 );
buf ( R_4ba_1d9d9a08 , C0 );
buf ( R_bdd_1e6b8748 , n51675 );
buf ( R_398_1d9d5a48 , n51676 );
buf ( R_31d_1d9d0d68 , n51681 );
buf ( R_47a_1dd9ece8 , C0 );
buf ( R_2ca_1d9ce108 , C0 );
buf ( R_b03_1e6aff08 , n51682 );
buf ( R_2a0_1d9fbee8 , n51683 );
buf ( R_71f_1dfb8f68 , n51684 );
buf ( R_950_1e17eec8 , n51685 );
buf ( R_9ce_1e184288 , C0 );
buf ( R_aae_1e6b6c68 , C0 );
buf ( R_b39_1e6b20c8 , n51721 );
buf ( R_906_1e090ea8 , C0 );
buf ( R_786_1dfbd4c8 , C0 );
buf ( R_81c_1e092de8 , n51722 );
buf ( R_94b_1e17eba8 , n51723 );
buf ( R_8fb_1e09b948 , n51724 );
buf ( R_3cb_1d9d7a28 , n51725 );
buf ( R_86f_1e0961c8 , n51726 );
buf ( R_584_1dda8e28 , n51727 );
buf ( R_40a_1d9da688 , C0 );
buf ( R_954_1e17f148 , n51728 );
buf ( R_944_1e17e748 , n51729 );
buf ( R_bc8_1e6b7a28 , n51730 );
buf ( R_9a1_1e182168 , n51735 );
buf ( R_c02_1e6ba5e8 , C0 );
buf ( R_967_1e17fd28 , n51736 );
buf ( R_7ff_1e091bc8 , n51737 );
buf ( R_329_1d9d14e8 , n51775 );
buf ( R_ba1_1e6b61c8 , n51810 );
buf ( R_717_1dfb8a68 , n51811 );
buf ( R_aa1_1e18c168 , n51846 );
buf ( R_591_1dda9648 , n51878 );
buf ( R_99c_1e181e48 , n51879 );
buf ( R_a42_1e188b08 , C0 );
buf ( R_ba8_1e6b6628 , n51880 );
buf ( R_ae1_1e6ae9c8 , n51915 );
buf ( R_9c2_1e183b08 , C0 );
buf ( R_6bb_1dfb50e8 , n51916 );
buf ( R_41b_1d9dac28 , n51917 );
buf ( R_93d_1e17e2e8 , n51949 );
buf ( R_5b2_1ddaafe8 , C0 );
buf ( R_5d6_1d9dd388 , C0 );
buf ( R_402_1d9da188 , C0 );
buf ( R_4b0_1dda09a8 , n51950 );
buf ( R_549_1dda6948 , n52017 );
buf ( R_53a_1dda64e8 , C0 );
buf ( R_70d_1dfb8428 , n52026 );
buf ( R_aa4_1e18c348 , n52027 );
buf ( R_798_1dfbdb08 , n52028 );
buf ( R_7fb_1e091948 , n52029 );
buf ( R_32a_1d9d1a88 , C0 );
buf ( R_a36_1e188388 , C0 );
buf ( R_5ed_1ddacfc8 , n52061 );
buf ( R_b9a_1e6b6268 , C0 );
buf ( R_c07_1e6ba188 , n52062 );
buf ( R_47e_1dd9ef68 , C0 );
buf ( R_ad2_1e6ae568 , C0 );
buf ( R_39d_1d9d5d68 , n52071 );
buf ( R_83f_1e0943c8 , n52072 );
buf ( R_7eb_1e090f48 , n52073 );
buf ( R_42e_1d9dbd08 , C0 );
buf ( R_b51_1e6b2fc8 , n52105 );
buf ( R_6b4_1dfb4c88 , n52106 );
buf ( R_694_1dfb3888 , n52107 );
buf ( R_68f_1dfb3568 , n52108 );
buf ( R_777_1dfbc668 , n52109 );
buf ( R_7b0_1e08ea68 , n52110 );
buf ( R_7a0_1e08e068 , n52111 );
buf ( R_75e_1dfbbbc8 , C0 );
buf ( R_5b7_1ddaae08 , n52112 );
buf ( R_63d_1dfb0228 , n52117 );
buf ( R_636_1dfb02c8 , C0 );
buf ( R_8de_1e09ac28 , C0 );
buf ( R_2ef_1d9cf0a8 , n52118 );
buf ( R_302_1d9d4508 , C0 );
buf ( R_9b8_1e182fc8 , n52119 );
buf ( R_4b2_1dda14e8 , C0 );
buf ( R_8e4_1e09aae8 , n52120 );
buf ( R_3de_1d9d8b08 , C0 );
buf ( R_ab8_1e18cfc8 , n52121 );
buf ( R_71b_1dfb8ce8 , n52122 );
buf ( R_c0c_1e6ba4a8 , n52123 );
buf ( R_c2b_1e6bb808 , n52124 );
buf ( R_5ac_1ddaa728 , n52125 );
buf ( R_853_1e095048 , n52126 );
buf ( R_2aa_1d9fca28 , C0 );
buf ( R_385_1d9d4e68 , n52135 );
buf ( R_436_1d9dc208 , C0 );
buf ( R_a60_1e1898c8 , n52136 );
buf ( R_7bb_1e08f148 , n52137 );
buf ( R_811_1e092708 , n52204 );
buf ( R_4c5_1dda16c8 , n52235 );
buf ( R_406_1d9da408 , C0 );
buf ( R_473_1dd9e388 , n52236 );
buf ( R_8aa_1e098ba8 , C0 );
buf ( R_b7e_1e6b50e8 , C0 );
buf ( R_7b5_1e08ed88 , n52267 );
buf ( R_5fb_1ddad888 , n52268 );
buf ( R_34d_1d9d2b68 , n52318 );
buf ( R_ae3_1e6aeb08 , n52319 );
buf ( R_6f3_1dfb73e8 , n52320 );
buf ( R_82b_1e093748 , n52321 );
buf ( R_72a_1dfbacc8 , C0 );
buf ( R_bc3_1e6b7708 , n52322 );
buf ( R_8fa_1e09bda8 , C0 );
buf ( R_567_1dda7c08 , n52323 );
buf ( R_89f_1e097fc8 , n52324 );
buf ( R_3ed_1d9d8f68 , n52333 );
buf ( R_599_1dda9b48 , n52365 );
buf ( R_851_1e094f08 , n52397 );
buf ( R_2dd_1d9ce568 , n52402 );
buf ( R_4a8_1dda04a8 , n52403 );
buf ( R_8a9_1e098608 , n52434 );
buf ( R_366_1d9d4008 , C0 );
buf ( R_376_1ddad568 , C0 );
buf ( R_75d_1dfbb628 , n52465 );
buf ( R_59a_1ddaa0e8 , C0 );
buf ( R_4c2_1dda19e8 , C0 );
buf ( R_8be_1e08eba8 , C0 );
buf ( R_2c5_1d9fd608 , n52470 );
buf ( R_595_1dda98c8 , n52502 );
buf ( R_446_1d9dd108 , C0 );
buf ( R_6c5_1dfb5728 , n52562 );
buf ( R_5d8_1ddac2a8 , n52563 );
buf ( R_682_1dfb3248 , C0 );
buf ( R_64b_1dfb0ae8 , n52564 );
buf ( R_791_1dfbd6a8 , n52595 );
buf ( R_b7b_1e6b4a08 , n52596 );
buf ( R_3b1_1d9d69e8 , n52605 );
buf ( R_7e9_1e090e08 , n52636 );
buf ( R_beb_1e6b9008 , n52637 );
buf ( R_6c0_1dfb5408 , n52638 );
buf ( R_8ba_1e0995a8 , C0 );
buf ( R_a8e_1e17f508 , C0 );
buf ( R_3c8_1d9d7848 , n52639 );
buf ( R_be4_1e6b8ba8 , n52640 );
buf ( R_544_1dda6628 , n52641 );
buf ( R_53f_1dda6308 , n52642 );
buf ( R_90e_1e09ca28 , C0 );
buf ( R_381_1d9d4be8 , n52651 );
buf ( R_a3e_1e188888 , C0 );
buf ( R_6fd_1dfb7a28 , n52660 );
buf ( R_a3a_1e188608 , C0 );
buf ( R_8c2_1e099aa8 , C0 );
buf ( R_af0_1e6af328 , n52661 );
buf ( R_296_1d9fb8a8 , n52668 );
buf ( R_b12_1e6b0d68 , C0 );
buf ( R_ba9_1e6b66c8 , n52703 );
buf ( R_b1d_1e6b0f48 , n52739 );
buf ( R_2b5_1d9fcc08 , n52744 );
buf ( R_6ff_1dfb7b68 , n52745 );
buf ( R_a98_1e18bbc8 , n52746 );
buf ( R_58e_1dda9968 , C0 );
buf ( R_753_1dfbafe8 , n52747 );
buf ( R_3c5_1d9d7668 , n52756 );
buf ( R_447_1d9dc7a8 , n52757 );
buf ( R_61f_1dfaef68 , n52758 );
buf ( R_54e_1dda28e8 , C0 );
buf ( R_6f8_1dfb7708 , n52759 );
buf ( R_3a4_1d9d61c8 , n52760 );
buf ( R_423_1d9db128 , n52761 );
buf ( R_6a4_1dfb4288 , n52762 );
buf ( R_b9b_1e6b5e08 , n52763 );
buf ( R_a07_1e186128 , n52764 );
buf ( R_55f_1dda7708 , n52765 );
buf ( R_79d_1dfbde28 , n52796 );
buf ( R_66d_1dfb2028 , n52801 );
buf ( R_5e2_1ddacde8 , C0 );
buf ( R_48b_1dd9f288 , n52802 );
buf ( R_5ee_1dda3a68 , C0 );
buf ( R_6c6_1dfb2d48 , C0 );
buf ( R_3e3_1d9d8928 , n52803 );
buf ( R_b83_1e6b4f08 , n52804 );
buf ( R_533_1dda5b88 , n52805 );
buf ( R_42d_1d9db768 , n52836 );
buf ( R_7e0_1e090868 , n52837 );
buf ( R_696_1dfb3ec8 , C0 );
buf ( R_3f9_1d9d96e8 , n52852 );
buf ( R_b88_1e6b5228 , n52853 );
buf ( R_758_1dfbb308 , n52854 );
buf ( R_3d2_1d9d8388 , C0 );
buf ( R_534_1dda5c28 , n52855 );
buf ( R_532_1d9d1308 , C0 );
buf ( R_867_1e095cc8 , n52856 );
buf ( R_2b6_1d9fd1a8 , C0 );
buf ( R_775_1dfbc528 , n52922 );
buf ( R_3e8_1d9d8c48 , n52923 );
buf ( R_4d0_1dda1da8 , n52924 );
buf ( R_30d_1d9d0368 , n52929 );
buf ( R_4e7_1dda2c08 , n52930 );
buf ( R_70a_1dfb8748 , C0 );
buf ( R_a58_1e1893c8 , n52931 );
buf ( R_4e8_1dda2ca8 , n52932 );
buf ( R_4e6_1dda3068 , C0 );
buf ( R_535_1dda5cc8 , n52972 );
buf ( R_5ea_1dda37e8 , C0 );
buf ( R_929_1e09d608 , n53004 );
buf ( R_448_1d9dc848 , n53005 );
buf ( R_b0b_1e6b0408 , n53006 );
buf ( R_319_1d9d0ae8 , n53011 );
buf ( R_985_1e180fe8 , n53016 );
buf ( R_32f_1d9d18a8 , n53017 );
buf ( R_4e9_1dda2d48 , n53049 );
buf ( R_b1f_1e6b1088 , n53050 );
buf ( R_495_1dd9f8c8 , n53081 );
buf ( R_63b_1dfb00e8 , n53082 );
buf ( R_536_1dda6268 , C0 );
buf ( R_3d9_1d9d82e8 , n53091 );
buf ( R_a4f_1e188e28 , n53092 );
buf ( R_470_1dd9e1a8 , n53093 );
buf ( R_2d5_1d9ce068 , n53098 );
buf ( R_3f0_1d9d9148 , n53099 );
buf ( R_acf_1e18de28 , n53100 );
buf ( R_ac2_1e18db08 , C0 );
buf ( R_9b4_1e182d48 , n53101 );
buf ( R_a05_1e185fe8 , n53146 );
buf ( R_2d9_1d9ce2e8 , n53151 );
buf ( R_8ed_1e09b088 , n53182 );
buf ( R_3f3_1d9d9328 , n53183 );
buf ( R_af2_1e6af968 , C0 );
buf ( R_44d_1d9dcb68 , n53214 );
buf ( R_645_1dfb0728 , n53219 );
buf ( R_648_1dfb0908 , n53220 );
buf ( R_4a1_1dda0048 , n53251 );
buf ( R_749_1dfba9a8 , n53260 );
buf ( R_2c8_1d9fd7e8 , n53261 );
buf ( R_3bc_1d9d70c8 , n53262 );
buf ( R_3f6_1ddad7e8 , C0 );
buf ( R_596_1dda9e68 , C0 );
buf ( R_c01_1e6b9dc8 , n53298 );
buf ( R_734_1dfb9c88 , n53299 );
buf ( R_5a5_1ddaa2c8 , n53331 );
buf ( R_6e3_1dfb69e8 , n53332 );
buf ( R_914_1e09c8e8 , n53333 );
buf ( R_43d_1d9dc168 , n53364 );
buf ( R_2cb_1d9fd9c8 , n53365 );
buf ( R_3d0_1d9d7d48 , n53366 );
buf ( R_b67_1e6b3d88 , n53367 );
buf ( R_b01_1e6afdc8 , n53402 );
buf ( R_37d_1d9d4968 , n53411 );
buf ( R_a80_1e18acc8 , n53412 );
buf ( R_9bd_1e1832e8 , n53417 );
buf ( R_339_1d9d1ee8 , n53455 );
buf ( R_7ad_1e08e888 , n53486 );
buf ( R_972_1e180908 , C0 );
buf ( R_a22_1e184788 , C0 );
buf ( R_486_1ddacb68 , C0 );
buf ( R_5d5_1ddac0c8 , n53517 );
buf ( R_592_1dda9be8 , C0 );
buf ( R_449_1d9dc8e8 , n53548 );
buf ( R_87b_1e096948 , n53549 );
buf ( R_8f5_1e09b588 , n53580 );
buf ( R_35a_1d9d3888 , C0 );
buf ( R_37a_1ddab9e8 , C0 );
buf ( R_991_1e181768 , n53585 );
buf ( R_62a_1dfb1448 , C0 );
buf ( R_808_1e092168 , n53586 );
buf ( R_3a6_1d9d6808 , C0 );
buf ( R_b95_1e6b5a48 , n53591 );
buf ( R_83e_1e17e108 , C0 );
buf ( R_386_1d9d5408 , C0 );
buf ( R_90d_1e09c488 , n53658 );
buf ( R_931_1e09db08 , n53690 );
buf ( R_ac9_1e18da68 , n53758 );
buf ( R_a31_1e187b68 , n53818 );
buf ( R_640_1dfb0408 , n53819 );
buf ( R_667_1dfb1c68 , n53820 );
buf ( R_6cb_1dfb5ae8 , n53821 );
buf ( R_74a_1e17f288 , C0 );
buf ( R_676_1dfb2ac8 , C0 );
buf ( R_372_1d9d4788 , C0 );
buf ( R_56c_1dda7f28 , n53822 );
buf ( R_334_1d9d1bc8 , n53823 );
buf ( R_31e_1d9fc528 , C0 );
buf ( R_981_1e180d68 , n53828 );
buf ( R_8ca_1e099fa8 , C0 );
buf ( R_85e_1e095c28 , C0 );
buf ( R_bbe_1e6af6e8 , C0 );
buf ( R_49b_1dd9fc88 , n53829 );
buf ( R_73a_1dfba548 , C0 );
buf ( R_5fe_1dfaf8c8 , C0 );
buf ( R_98b_1e1813a8 , n53830 );
buf ( R_88e_1e097a28 , C0 );
buf ( R_28f_1d9fb448 , n53837 );
buf ( R_9bc_1e183248 , n53838 );
buf ( R_5db_1ddac488 , n53839 );
buf ( R_88a_1e08ee28 , C0 );
buf ( R_5a6_1ddaa868 , C0 );
buf ( R_443_1d9dc528 , n53840 );
buf ( R_a0a_1e186808 , C0 );
buf ( R_358_1d9d3248 , n53841 );
buf ( R_88f_1e0975c8 , n53842 );
buf ( R_acc_1e18dc48 , n53843 );
buf ( R_aac_1e18c848 , n53844 );
buf ( R_2a2_1d9fde28 , C0 );
buf ( R_8a5_1e098388 , n53853 );
buf ( R_8ec_1e09afe8 , n53854 );
buf ( R_289_1d9fb088 , n53863 );
buf ( R_340_1d9d2348 , n53864 );
buf ( R_c2d_1e6bb948 , n53879 );
buf ( R_964_1e17fb48 , n53880 );
buf ( R_85d_1e095688 , n53912 );
buf ( R_6fa_1dfb7d48 , C0 );
buf ( R_4d5_1dda20c8 , n53943 );
buf ( R_a5a_1e18b308 , C0 );
buf ( R_7de_1e090c28 , C0 );
buf ( R_605_1ddadec8 , n53948 );
buf ( R_311_1d9d05e8 , n53953 );
buf ( R_8a6_1e098928 , C0 );
buf ( R_a2f_1e187a28 , n53954 );
buf ( R_81f_1e092fc8 , n53955 );
buf ( R_3b6_1d9d7208 , C0 );
buf ( R_315_1d9d0868 , n53960 );
buf ( R_93f_1e17e428 , n53961 );
buf ( R_5b1_1ddaaa48 , n53993 );
buf ( R_631_1dfafaa8 , n53998 );
buf ( R_890_1e097668 , n53999 );
buf ( R_670_1dfb2208 , n54000 );
buf ( R_b9c_1e6b5ea8 , n54001 );
buf ( R_8e9_1e09ae08 , n54032 );
buf ( R_932_1e093928 , C0 );
buf ( R_817_1e092ac8 , n54033 );
buf ( R_b60_1e6b3928 , n54034 );
buf ( R_979_1e180868 , n54039 );
buf ( R_8d8_1e09a368 , n54040 );
buf ( R_628_1dfaf508 , n54041 );
buf ( R_729_1dfb95a8 , n54050 );
buf ( R_a92_1e18bd08 , C0 );
buf ( R_b33_1e6b1d08 , n54051 );
buf ( R_2ab_1d9fc5c8 , n54052 );
buf ( R_5e6_1dd9f6e8 , C0 );
buf ( R_5c0_1ddab3a8 , n54053 );
buf ( R_600_1ddadba8 , n54054 );
buf ( R_8f4_1e09b4e8 , n54055 );
buf ( R_29d_1d9fbd08 , n54063 );
buf ( R_c11_1e6ba7c8 , n54099 );
buf ( R_4d7_1dda2208 , n54100 );
buf ( R_b43_1e6b2708 , n54101 );
buf ( R_881_1e096d08 , n54133 );
buf ( R_891_1e097708 , n54165 );
buf ( R_8b4_1e098ce8 , n54166 );
buf ( R_6ac_1dfb4788 , n54167 );
buf ( R_2f0_1d9cf148 , n54168 );
buf ( R_ad8_1e6ae428 , n54169 );
buf ( R_9bb_1e1831a8 , n54170 );
buf ( R_bd9_1e6b84c8 , n54206 );
buf ( R_39f_1d9d5ea8 , n54207 );
buf ( R_a5e_1e189c88 , C0 );
buf ( R_303_1d9cfd28 , n54208 );
buf ( R_6ae_1dfb4dc8 , C0 );
buf ( R_477_1dd9e608 , n54209 );
buf ( R_6d2_1e0981a8 , C0 );
buf ( R_38f_1d9d54a8 , n54210 );
buf ( R_4d2_1dda23e8 , C0 );
buf ( R_82f_1e0939c8 , n54211 );
buf ( R_61d_1dfaee28 , n54216 );
buf ( R_673_1dfb23e8 , n54217 );
buf ( R_578_1dda86a8 , n54218 );
buf ( R_a65_1e189be8 , n54253 );
buf ( R_9a5_1e1823e8 , n54258 );
buf ( R_744_1dfba688 , n54259 );
buf ( R_bfe_1e6ba0e8 , C0 );
buf ( R_86e_1e096628 , C0 );
buf ( R_6ce_1e0945a8 , C0 );
buf ( R_9df_1e184828 , n54260 );
buf ( R_571_1dda8248 , n54292 );
buf ( R_9e0_1e1848c8 , n54293 );
buf ( R_9de_1e184c88 , C0 );
buf ( R_41a_1ddabee8 , C0 );
buf ( R_36e_1d9d1588 , C0 );
buf ( R_6b9_1dfb4fa8 , n54353 );
buf ( R_b72_1e6b4968 , C0 );
buf ( R_73f_1dfba368 , n54354 );
buf ( R_a4d_1e188ce8 , n54389 );
buf ( R_9e1_1e184968 , n54442 );
buf ( R_2d0_1d9fdce8 , n54443 );
buf ( R_72e_1dfb9dc8 , C0 );
buf ( R_c25_1e6bb448 , n54479 );
buf ( R_8eb_1e09af48 , n54480 );
buf ( R_6eb_1dfb6ee8 , n54481 );
buf ( R_764_1dfbba88 , n54482 );
buf ( R_9b1_1e182b68 , n54487 );
buf ( R_970_1e1802c8 , n54488 );
buf ( R_bce_1e6b82e8 , C0 );
buf ( R_325_1d9d1268 , n54526 );
buf ( R_65c_1dfb1588 , n54527 );
buf ( R_643_1dfb05e8 , n54528 );
buf ( R_abf_1e18d428 , n54529 );
buf ( R_a9b_1e18bda8 , n54530 );
buf ( R_b7c_1e6b4aa8 , n54531 );
buf ( R_9ba_1e183608 , C0 );
buf ( R_bef_1e6b9288 , n54532 );
buf ( R_b14_1e6b09a8 , n54533 );
buf ( R_996_1e181f88 , C0 );
buf ( R_812_1e092ca8 , C0 );
buf ( R_4a2_1dda05e8 , C0 );
buf ( R_6e0_1dfb6808 , n54534 );
buf ( R_490_1dd9f5a8 , n54535 );
buf ( R_711_1dfb86a8 , n54544 );
buf ( R_a86_1e18ba88 , C0 );
buf ( R_342_1d9d2988 , C0 );
buf ( R_c0e_1e6baae8 , C0 );
buf ( R_8e3_1e09aa48 , n54545 );
buf ( R_646_1dfb0cc8 , C0 );
buf ( R_74d_1dfbac28 , n54560 );
buf ( R_67f_1dfb2b68 , n54561 );
buf ( R_34f_1d9d2ca8 , n54562 );
buf ( R_8f3_1e09b448 , n54563 );
buf ( R_bdc_1e6b86a8 , n54564 );
buf ( R_57f_1dda8b08 , n54565 );
buf ( R_77a_1dfbcd48 , C0 );
buf ( R_4c1_1dda1448 , n54596 );
buf ( R_b8e_1e6b5ae8 , C0 );
buf ( R_c29_1e6bb6c8 , n54632 );
buf ( R_875_1e096588 , n54664 );
buf ( R_852_1e0954a8 , C0 );
buf ( R_6a6_1dfb48c8 , C0 );
buf ( R_76f_1dfbc168 , n54665 );
buf ( R_984_1e180f48 , n54666 );
buf ( R_39a_1d9d6088 , C0 );
buf ( R_35f_1d9d36a8 , n54667 );
buf ( R_5d0_1ddabda8 , n54668 );
buf ( R_b65_1e6b3c48 , n54704 );
buf ( R_92b_1e09d748 , n54705 );
buf ( R_3eb_1d9d8e28 , n54706 );
buf ( R_53b_1dda6088 , n54707 );
buf ( R_97a_1e180e08 , C0 );
buf ( R_369_1d9d3ce8 , n54745 );
buf ( R_7f5_1e091588 , n54777 );
buf ( R_588_1dda90a8 , n54778 );
buf ( R_b6a_1e6b4468 , C0 );
buf ( R_435_1d9dbc68 , n54809 );
buf ( R_a08_1e1861c8 , n54810 );
buf ( R_7ef_1e0911c8 , n54811 );
buf ( R_781_1dfbcca8 , n54877 );
buf ( R_55c_1dda7528 , n54878 );
buf ( R_3bf_1d9d72a8 , n54879 );
buf ( R_850_1e094e68 , n54880 );
buf ( R_2ea_1d9cf288 , C0 );
buf ( R_687_1dfb3068 , n54881 );
buf ( R_795_1dfbd928 , n54912 );
buf ( R_382_1d9d5188 , C0 );
buf ( R_63e_1dfb07c8 , C0 );
buf ( R_2b7_1d9fcd48 , n54913 );
buf ( R_9b0_1e182ac8 , n54914 );
buf ( R_6dd_1dfb6628 , n54923 );
buf ( R_4be_1dda1768 , C0 );
buf ( R_bfd_1e6b9b48 , n54959 );
buf ( R_b0d_1e6b0548 , n54995 );
buf ( R_b9d_1e6b5f48 , n55030 );
buf ( R_b3a_1e6b2668 , C0 );
buf ( R_4b9_1dda0f48 , n55061 );
buf ( R_4bb_1dda1088 , n55062 );
buf ( R_9a0_1e1820c8 , n55063 );
buf ( R_83b_1e094148 , n55064 );
buf ( R_8ea_1e09b3a8 , C0 );
buf ( R_b21_1e6b11c8 , n55100 );
buf ( R_62f_1dfaf968 , n55101 );
buf ( R_91d_1e09ce88 , n55133 );
buf ( R_483_1dd9ed88 , n55134 );
buf ( R_7c0_1e08f468 , n55135 );
buf ( R_bd5_1e6b8248 , n55171 );
buf ( R_364_1d9d39c8 , n55172 );
buf ( R_322_1d9d2e88 , C0 );
buf ( R_326_1d9d1808 , C0 );
buf ( R_99b_1e181da8 , n55173 );
buf ( R_961_1e17f968 , n55178 );
buf ( R_726_1dfb98c8 , C0 );
buf ( R_a7d_1e18aae8 , n55213 );
buf ( R_826_1e09de28 , C0 );
buf ( R_89a_1dfb4648 , C0 );
buf ( R_511_1dda4648 , n55245 );
buf ( R_2fb_1d9cf828 , n55246 );
buf ( R_b5c_1e6b36a8 , n55247 );
buf ( R_8b0_1e098a68 , n55248 );
buf ( R_708_1dfb8108 , n55249 );
buf ( R_603_1ddadd88 , n55250 );
buf ( R_804_1e091ee8 , n55251 );
buf ( R_573_1dda8388 , n55252 );
buf ( R_a56_1e189a08 , C0 );
buf ( R_510_1dda45a8 , n55253 );
buf ( R_833_1e093c48 , n55254 );
buf ( R_8c1_1e099508 , n55285 );
buf ( R_966_1e180188 , C0 );
buf ( R_46d_1dd9dfc8 , n55316 );
buf ( R_bcc_1e6b7ca8 , n55317 );
buf ( R_47b_1dd9e888 , n55318 );
buf ( R_aea_1e6af468 , C0 );
buf ( R_8d1_1e099f08 , n55349 );
buf ( R_57a_1ddaa368 , C0 );
buf ( R_8f2_1e09b8a8 , C0 );
buf ( R_b35_1e6b1e48 , n55385 );
buf ( R_b05_1e6b0048 , n55421 );
buf ( R_aa9_1e18c668 , n55456 );
buf ( R_9b7_1e182f28 , n55457 );
buf ( R_3ae_1d9d6d08 , C0 );
buf ( R_50f_1dda4508 , n55458 );
buf ( R_a23_1e1872a8 , n55459 );
buf ( R_2c9_1d9fd888 , n55464 );
buf ( R_5c6_1d9d7e88 , C0 );
buf ( R_8bd_1e099288 , n55495 );
buf ( R_4b1_1dda0a48 , n55526 );
buf ( R_b45_1e6b2848 , n55595 );
buf ( R_422_1d9db588 , C0 );
buf ( R_2cc_1d9fda68 , n55596 );
buf ( R_9d5_1e1841e8 , n55601 );
buf ( R_37e_1d9d4f08 , C0 );
buf ( R_42c_1d9db6c8 , n55602 );
buf ( R_a7e_1e18b088 , C0 );
buf ( R_a8d_1e18b4e8 , n55660 );
buf ( R_50e_1dda4968 , C0 );
buf ( R_626_1dfafb48 , C0 );
buf ( R_5cc_1ddabb28 , n55661 );
buf ( R_295_1d9fb808 , n55668 );
buf ( R_a9e_1e18c488 , C0 );
buf ( R_80d_1e092488 , n55700 );
buf ( R_9af_1e182a28 , n55701 );
buf ( R_946_1e17ed88 , C0 );
buf ( R_a5c_1e189648 , n55702 );
buf ( R_5bb_1ddab088 , n55703 );
buf ( R_3e6_1d9d9008 , C0 );
buf ( R_ab3_1e18cca8 , n55704 );
buf ( R_a1e_1e187488 , C0 );
buf ( R_66a_1dfb2348 , C0 );
buf ( R_7f8_1e091768 , n55705 );
buf ( R_56e_1dda8568 , C0 );
buf ( R_3c2_1d9d7988 , C0 );
buf ( R_837_1e093ec8 , n55706 );
buf ( R_866_1e096128 , C0 );
buf ( R_65a_1dfb1948 , C0 );
buf ( R_4aa_1dda0ae8 , C0 );
buf ( R_540_1dda63a8 , n55707 );
buf ( R_61b_1dfaece8 , n55708 );
buf ( R_78a_1dfbd748 , C0 );
buf ( R_76c_1dfbbf88 , n55709 );
buf ( R_4c7_1dda1808 , n55710 );
buf ( R_47f_1dd9eb08 , n55711 );
buf ( R_34a_1d9d4a08 , C0 );
buf ( R_b57_1e6b3388 , n55712 );
buf ( R_545_1dda66c8 , n55744 );
buf ( R_c13_1e6ba908 , n55745 );
buf ( R_44c_1d9dcac8 , n55746 );
buf ( R_a0b_1e1863a8 , n55747 );
buf ( R_6d5_1dfb6128 , n55756 );
buf ( R_bf3_1e6b9508 , n55757 );
buf ( R_3ee_1d9d9508 , C0 );
buf ( R_6d7_1dfb6268 , n55758 );
buf ( R_3d6_1d9d9788 , C0 );
buf ( R_b06_1e6b05e8 , C0 );
buf ( R_9d4_1e184148 , n55759 );
buf ( R_33b_1d9d2028 , n55760 );
buf ( R_739_1dfb9fa8 , n55769 );
buf ( R_a0e_1e186a88 , C0 );
buf ( R_7dd_1e090688 , n55848 );
buf ( R_54f_1dda6d08 , n55849 );
buf ( R_926_1e09dba8 , C0 );
buf ( R_abb_1e18d1a8 , n55850 );
buf ( R_70e_1dfb89c8 , C0 );
buf ( R_ba2_1e6b6768 , C0 );
buf ( R_917_1e09cac8 , n55851 );
buf ( R_923_1e09d248 , n55852 );
buf ( R_784_1dfbce88 , n55853 );
buf ( R_920_1e09d068 , n55854 );
buf ( R_564_1dda7a28 , n55855 );
buf ( R_9a9_1e182668 , n55860 );
buf ( R_bfa_1e6b9e68 , C0 );
buf ( R_62c_1dfaf788 , n55861 );
buf ( R_8c9_1e099a08 , n55892 );
buf ( R_43c_1d9dc0c8 , n55893 );
buf ( R_b00_1e6afd28 , n55894 );
buf ( R_35d_1d9d3568 , n55935 );
buf ( R_c18_1e6bac28 , n55936 );
buf ( R_306_1d9d0408 , C0 );
buf ( R_939_1e17e068 , n55968 );
buf ( R_474_1dd9e428 , n55969 );
buf ( R_4a9_1dda0548 , n56000 );
buf ( R_2ac_1d9fc668 , n56001 );
buf ( R_609_1dfae1a8 , n56006 );
buf ( R_94c_1e17ec48 , n56007 );
buf ( R_90a_1e09c7a8 , C0 );
buf ( R_92e_1e0918a8 , C0 );
buf ( R_7be_1e08f828 , C0 );
buf ( R_825_1e093388 , n56036 );
buf ( R_559_1dda7348 , n56068 );
buf ( R_bf7_1e6b9788 , n56069 );
buf ( R_87a_1e096da8 , C0 );
buf ( R_9d3_1e1840a8 , n56070 );
buf ( R_394_1d9d57c8 , n56071 );
buf ( R_31a_1d9d1088 , C0 );
buf ( R_69f_1dfb3f68 , n56072 );
buf ( R_787_1dfbd068 , n56073 );
buf ( R_a63_1e189aa8 , n56074 );
buf ( R_9ae_1e183388 , C0 );
buf ( R_945_1e17e7e8 , n56106 );
buf ( R_537_1dda5e08 , n56107 );
buf ( R_725_1dfb9328 , n56116 );
buf ( R_b68_1e6b3e28 , n56117 );
buf ( R_7a5_1e08e388 , n56146 );
buf ( R_4eb_1dda2e88 , n56147 );
buf ( R_619_1dfaeba8 , n56152 );
buf ( R_800_1e091c68 , n56153 );
buf ( R_be8_1e6b8e28 , n56154 );
buf ( R_4ec_1dda2f28 , n56155 );
buf ( R_4ea_1dda32e8 , C0 );
buf ( R_2f1_1d9cf1e8 , n56160 );
buf ( R_5d3_1ddabf88 , n56161 );
buf ( R_6da_1dfb6948 , C0 );
buf ( R_5b6_1ddab268 , C0 );
buf ( R_3ac_1d9d66c8 , n56162 );
buf ( R_983_1e180ea8 , n56163 );
buf ( R_b73_1e6b4508 , n56164 );
buf ( R_4ed_1dda2fc8 , n56196 );
buf ( R_ada_1e6aea68 , C0 );
buf ( R_7fc_1e0919e8 , n56197 );
buf ( R_b3c_1e6b22a8 , n56198 );
buf ( R_304_1d9cfdc8 , n56199 );
buf ( R_5ab_1ddaa688 , n56200 );
buf ( R_85c_1e0955e8 , n56201 );
buf ( R_442_1d9dcc08 , C0 );
buf ( R_3ce_1d9d8608 , C0 );
buf ( R_ad5_1e6ae248 , n56236 );
buf ( R_ae8_1e6aee28 , n56237 );
buf ( R_3b4_1d9d6bc8 , n56238 );
buf ( R_8b8_1e098f68 , n56239 );
buf ( R_b46_1e6b2de8 , C0 );
buf ( R_8e8_1e09ad68 , n56240 );
buf ( R_bbf_1e6b7488 , n56241 );
buf ( R_799_1dfbdba8 , n56272 );
buf ( R_778_1dfbc708 , n56273 );
buf ( R_a4b_1e188ba8 , n56274 );
buf ( R_51d_1dda4dc8 , n56306 );
buf ( R_657_1dfb1268 , n56307 );
buf ( R_9d2_1e17f788 , C0 );
buf ( R_348_1d9d2848 , n56308 );
buf ( R_51c_1dda4d28 , n56309 );
buf ( R_8d7_1e09a2c8 , n56310 );
buf ( R_9b3_1e182ca8 , n56311 );
buf ( R_7db_1e090548 , n56312 );
buf ( R_715_1dfb8928 , n56321 );
buf ( R_68c_1dfb3388 , n56322 );
buf ( R_880_1e096c68 , n56323 );
buf ( R_29c_1d9fbc68 , n56328 );
buf ( R_b7d_1e6b4b48 , n56364 );
buf ( R_51b_1dda4c88 , n56365 );
buf ( R_bba_1e6b7668 , C0 );
buf ( R_3dc_1d9d84c8 , n56366 );
buf ( R_5a0_1dda9fa8 , n56367 );
buf ( R_75f_1dfbb768 , n56368 );
buf ( R_b7f_1e6b4c88 , n56369 );
buf ( R_b16_1e6b0fe8 , C0 );
buf ( R_ba3_1e6b6308 , n56370 );
buf ( R_654_1dfb1088 , n56371 );
buf ( R_bc7_1e6b7988 , n56372 );
buf ( R_2a3_1d9fc0c8 , n56373 );
buf ( R_6f0_1dfb7208 , n56374 );
buf ( R_7a1_1e08e108 , n56435 );
buf ( R_371_1d9d41e8 , n56473 );
buf ( R_51a_1dda50e8 , C0 );
buf ( R_ab7_1e18cf28 , n56474 );
buf ( R_7e6_1e099828 , C0 );
buf ( R_b6b_1e6b4008 , n56475 );
buf ( R_9ad_1e1828e8 , n56480 );
buf ( R_935_1e09dd88 , n56512 );
buf ( R_b8a_1e6bb768 , C0 );
buf ( R_69d_1dfb3e28 , n56572 );
buf ( R_45e_1d9ddb08 , C0 );
buf ( R_a1a_1e187208 , C0 );
buf ( R_a49_1e188a68 , n56607 );
buf ( R_a09_1e186268 , n56652 );
buf ( R_496_1dd9fe68 , C0 );
buf ( R_336_1d9d2208 , C0 );
buf ( R_5df_1ddac708 , n56653 );
buf ( R_5c7_1ddab808 , n56654 );
buf ( R_990_1e1816c8 , n56655 );
buf ( R_6c9_1dfb59a8 , n56715 );
buf ( R_2eb_1d9cee28 , n56716 );
buf ( R_2b8_1d9fcde8 , n56717 );
buf ( R_ae0_1e6ae928 , n56718 );
buf ( R_b2f_1e6b1a88 , n56719 );
buf ( R_84d_1e094c88 , n56751 );
buf ( R_a12_1e186d08 , C0 );
buf ( R_74f_1dfbad68 , n56752 );
buf ( R_a35_1e187de8 , n56787 );
buf ( R_28e_1d9fb3a8 , n56794 );
buf ( R_81a_1e0936a8 , C0 );
buf ( R_487_1dd9f008 , n56795 );
buf ( R_c1c_1e6baea8 , n56796 );
buf ( R_7a8_1e08e568 , n56797 );
buf ( R_471_1dd9e248 , n56828 );
buf ( R_766_1e0986a8 , C0 );
buf ( R_38b_1d9d5228 , n56829 );
buf ( R_a7b_1e18a9a8 , n56830 );
buf ( R_b52_1e6b8568 , C0 );
buf ( R_9ff_1e185c28 , n56831 );
buf ( R_7b9_1e08f008 , n56862 );
buf ( R_67b_1dfb28e8 , n56863 );
buf ( R_a00_1e185cc8 , n56864 );
buf ( R_9fe_1e6bb9e8 , C0 );
buf ( R_980_1e180cc8 , n56865 );
buf ( R_874_1e0964e8 , n56866 );
buf ( R_49c_1dd9fd28 , n56867 );
buf ( R_58c_1dda9328 , n56868 );
buf ( R_45f_1d9dd6a8 , n56869 );
buf ( R_98a_1e181808 , C0 );
buf ( R_8e2_1e09aea8 , C0 );
buf ( R_6ba_1dfb5548 , C0 );
buf ( R_bd8_1e6b8428 , n56870 );
buf ( R_a8b_1e18b3a8 , n56871 );
buf ( R_a01_1e185d68 , n56980 );
buf ( R_6b3_1dfb4be8 , n56981 );
buf ( R_60d_1dfae428 , n56986 );
buf ( R_6e8_1dfb6d08 , n56987 );
buf ( R_399_1d9d5ae8 , n56996 );
buf ( R_a16_1e186f88 , C0 );
buf ( R_bc2_1e6b7b68 , C0 );
buf ( R_32b_1d9d1628 , n56997 );
buf ( R_434_1d9dbbc8 , n56998 );
buf ( R_a24_1e187348 , n56999 );
buf ( R_377_1d9d45a8 , n57000 );
buf ( R_3cc_1d9d7ac8 , n57001 );
buf ( R_a68_1e189dc8 , n57002 );
buf ( R_963_1e17faa8 , n57003 );
buf ( R_7c5_1e08f788 , n57034 );
buf ( R_615_1dfae928 , n57039 );
buf ( R_8a2_1dfb9b48 , C0 );
buf ( R_722_1dfb9648 , C0 );
buf ( R_288_1d9f96e8 , n57048 );
buf ( R_556_1dda7668 , C0 );
buf ( R_748_1dfba908 , n57049 );
buf ( R_865_1e095b88 , n57081 );
buf ( R_607_1dfae068 , n57082 );
buf ( R_691_1dfb36a8 , n57142 );
buf ( R_978_1e1807c8 , n57143 );
buf ( R_84f_1e094dc8 , n57144 );
buf ( R_2cd_1d9fdb08 , n57149 );
buf ( R_ae2_1e6aef68 , C0 );
buf ( R_a1f_1e187028 , n57150 );
buf ( R_721_1dfb90a8 , n57159 );
buf ( R_733_1dfb9be8 , n57160 );
buf ( R_9e3_1e184aa8 , n57161 );
buf ( R_9e4_1e184b48 , n57162 );
buf ( R_c23_1e6bb308 , n57163 );
buf ( R_9e2_1e184f08 , C0 );
buf ( R_7ae_1dfbb1c8 , C0 );
buf ( R_91a_1e09d1a8 , C0 );
buf ( R_b84_1e6b4fa8 , n57164 );
buf ( R_b92_1e181088 , C0 );
buf ( R_ba4_1e6b63a8 , n57165 );
buf ( R_754_1dfbb088 , n57166 );
buf ( R_5a4_1ddaa228 , n57167 );
buf ( R_9a4_1e182348 , n57168 );
buf ( R_b08_1e6b0228 , n57169 );
buf ( R_9e5_1e184be8 , n57214 );
buf ( R_617_1dfaea68 , n57215 );
buf ( R_5ce_1ddac168 , C0 );
buf ( R_b89_1e6b52c8 , n57251 );
buf ( R_7b2_1e09b128 , C0 );
buf ( R_460_1d9dd748 , n57252 );
buf ( R_5e4_1ddaca28 , n57253 );
buf ( R_30a_1d9d0688 , C0 );
buf ( R_a0c_1e186448 , n57254 );
buf ( R_910_1e09c668 , n57255 );
buf ( R_553_1dda6f88 , n57256 );
buf ( R_86d_1e096088 , n57288 );
buf ( R_a0f_1e186628 , n57289 );
buf ( R_719_1dfb8ba8 , n57298 );
buf ( R_b48_1e6b2a28 , n57299 );
buf ( R_316_1d9d0e08 , C0 );
buf ( R_901_1e09bd08 , n57330 );
buf ( R_611_1dfae6a8 , n57335 );
buf ( R_ac5_1e18d7e8 , n57403 );
buf ( R_6c4_1dfb5688 , n57404 );
buf ( R_53c_1dda6128 , n57405 );
buf ( R_712_1dfb8c48 , C0 );
buf ( R_2f6_1d9cfc88 , C0 );
buf ( R_829_1e093608 , n57437 );
buf ( R_89d_1e097e88 , n57493 );
buf ( R_8d0_1e099e68 , n57494 );
buf ( R_8ac_1e0987e8 , n57495 );
buf ( R_8a0_1e098068 , n57496 );
buf ( R_aef_1e6af288 , n57497 );
buf ( R_759_1dfbb3a8 , n57528 );
buf ( R_a6d_1e18a0e8 , n57596 );
buf ( R_6bf_1dfb5368 , n57597 );
buf ( R_982_1e182c08 , C0 );
buf ( R_bdb_1e6b8608 , n57598 );
buf ( R_684_1dfb2e88 , n57599 );
buf ( R_7b7_1e08eec8 , n57600 );
buf ( R_478_1dd9e6a8 , n57601 );
buf ( R_be1_1e6b89c8 , n57637 );
buf ( R_b55_1e6b3248 , n57673 );
buf ( R_79b_1dfbdce8 , n57674 );
buf ( R_c27_1e6bb588 , n57675 );
buf ( R_96f_1e180228 , n57676 );
buf ( R_42b_1d9db628 , n57677 );
buf ( R_6cd_1dfb5c28 , n57686 );
buf ( R_652_1dfb16c8 , C0 );
buf ( R_71d_1dfb8e28 , n57695 );
buf ( R_703_1dfb7de8 , n57696 );
buf ( R_a54_1e189148 , n57697 );
buf ( R_4a3_1dda0188 , n57698 );
buf ( R_634_1dfafc88 , n57699 );
buf ( R_2ad_1d9fc708 , n57704 );
buf ( R_4cc_1dda1b28 , n57705 );
buf ( R_2a1_1d9fbf88 , n58610 );
buf ( R_93a_1e0977a8 , C0 );
buf ( R_a78_1e18a7c8 , n58611 );
buf ( R_c03_1e6b9f08 , n58612 );
buf ( R_72c_1dfb9788 , n58613 );
buf ( R_809_1e092208 , n58645 );
buf ( R_5b0_1ddaa9a8 , n58646 );
buf ( R_44b_1d9dca28 , n58647 );
buf ( R_952_1ddab768 , C0 );
buf ( R_899_1e097c08 , n58679 );
buf ( R_bd4_1e6b81a8 , n58680 );
buf ( R_a94_1e18b948 , n58681 );
buf ( R_6b1_1dfb4aa8 , n58741 );
buf ( R_491_1dd9f648 , n58772 );
buf ( R_5ca_1d9dae08 , C0 );
buf ( R_6f5_1dfb7528 , n58781 );
buf ( R_9c9_1e183a68 , n58786 );
buf ( R_75a_1dfbb948 , C0 );
buf ( R_461_1d9dd7e8 , n58817 );
buf ( R_7c3_1e08f648 , n58818 );
buf ( R_569_1dda7d48 , n58885 );
buf ( R_a75_1e18a5e8 , n58920 );
buf ( R_7ec_1e090fe8 , n58921 );
buf ( R_c20_1e6bb128 , n58922 );
buf ( R_96d_1e1800e8 , n58927 );
buf ( R_54a_1dda6ee8 , C0 );
buf ( R_b31_1e6b1bc8 , n58963 );
buf ( R_5bf_1ddab308 , n58964 );
buf ( R_900_1e09bc68 , n58965 );
buf ( R_b74_1e6b45a8 , n58966 );
buf ( R_940_1e17e4c8 , n58967 );
buf ( R_8dd_1e09a688 , n58998 );
buf ( R_a88_1e18b1c8 , n58999 );
buf ( R_743_1dfba5e8 , n59000 );
buf ( R_2d1_1d9fdd88 , n59005 );
buf ( R_4b3_1dda0b88 , n59006 );
buf ( R_48c_1dd9f328 , n59007 );
buf ( R_419_1d9daae8 , n59038 );
buf ( R_2ba_1d9fd428 , C0 );
buf ( R_898_1e097b68 , n59039 );
buf ( R_354_1d9d2fc8 , n59040 );
buf ( R_3c9_1d9d78e8 , n59049 );
buf ( R_afd_1e6afb48 , n59084 );
buf ( R_698_1dfb3b08 , n59085 );
buf ( R_8c8_1e099968 , n59086 );
buf ( R_aff_1e6afc88 , n59087 );
buf ( R_59c_1dda9d28 , n59088 );
buf ( R_43b_1d9dc028 , n59089 );
buf ( R_3e1_1d9d87e8 , n59098 );
buf ( R_7d8_1e090368 , n59099 );
buf ( R_624_1dfaf288 , n59100 );
buf ( R_ace_1e6ae2e8 , C0 );
buf ( R_294_1d9fb768 , n59107 );
buf ( R_818_1e092b68 , n59108 );
buf ( R_9c8_1e1839c8 , n59109 );
buf ( R_5c8_1ddab8a8 , n59110 );
buf ( R_c2f_1e6bba88 , n59111 );
buf ( R_ba5_1e6b6448 , n59146 );
buf ( R_6d0_1dfb5e08 , n59147 );
buf ( R_820_1e093068 , n59148 );
buf ( R_30e_1d9d0908 , C0 );
buf ( R_99f_1e182028 , n59149 );
buf ( R_73e_1dfba7c8 , C0 );
buf ( R_4ef_1dda3108 , n59150 );
buf ( R_451_1d9dcde8 , n59179 );
buf ( R_678_1dfb2708 , n59180 );
buf ( R_663_1dfb19e8 , n59181 );
buf ( R_5fa_1e091128 , C0 );
buf ( R_312_1d9d0b88 , C0 );
buf ( R_a45_1e1887e8 , n59216 );
buf ( R_b18_1e6b0c28 , n59217 );
buf ( R_4f0_1dda31a8 , n59218 );
buf ( R_4ee_1dda3568 , C0 );
buf ( R_7ab_1e08e748 , n59219 );
buf ( R_305_1d9cfe68 , n59224 );
buf ( R_955_1e17f1e8 , n59229 );
buf ( R_373_1d9d4328 , n59230 );
buf ( R_a39_1e188068 , n59265 );
buf ( R_669_1dfb1da8 , n59270 );
buf ( R_3a5_1d9d6268 , n59279 );
buf ( R_c0d_1e6ba548 , n59315 );
buf ( R_4f1_1dda3248 , n59347 );
buf ( R_541_1dda6448 , n59379 );
buf ( R_69a_1dfb4148 , C0 );
buf ( R_b90_1e6b5728 , n59380 );
buf ( R_99a_1e182208 , C0 );
buf ( R_960_1e17f8c8 , n59381 );
buf ( R_6a9_1dfb45a8 , n59441 );
buf ( R_4bc_1dda1128 , n59442 );
buf ( R_897_1e097ac8 , n59443 );
buf ( R_701_1dfb7ca8 , n59452 );
buf ( R_36c_1d9d3ec8 , n59453 );
buf ( R_60b_1dfae2e8 , n59454 );
buf ( R_583_1dda8d88 , n59455 );
buf ( R_330_1d9d1948 , n59456 );
buf ( R_bb6_1e6b73e8 , C0 );
buf ( R_71e_1dfb93c8 , C0 );
buf ( R_590_1dda95a8 , n59457 );
buf ( R_29e_1dda2668 , C0 );
buf ( R_b0f_1e6b0688 , n59458 );
buf ( R_a1b_1e186da8 , n59459 );
buf ( R_550_1dda6da8 , n59460 );
buf ( R_ac8_1e18d9c8 , n59461 );
buf ( R_a9d_1e18bee8 , n59529 );
buf ( R_561_1dda7848 , n59561 );
buf ( R_80e_1e092a28 , C0 );
buf ( R_9b6_1e187708 , C0 );
buf ( R_5e8_1ddacca8 , n59562 );
buf ( R_613_1dfae7e8 , n59563 );
buf ( R_b6c_1e6b40a8 , n59564 );
buf ( R_3d3_1d9d7f28 , n59565 );
buf ( R_31f_1d9d0ea8 , n59566 );
buf ( R_9c7_1e183928 , n59567 );
buf ( R_5dd_1ddac5c8 , n59598 );
buf ( R_78e_1dfbd9c8 , C0 );
buf ( R_a13_1e1868a8 , n59599 );
buf ( R_70c_1dfb8388 , n59600 );
buf ( R_885_1e096f88 , n59632 );
buf ( R_85b_1e095548 , n59633 );
buf ( R_8ff_1e09bbc8 , n59634 );
buf ( R_716_1dfb8ec8 , C0 );
buf ( R_2b9_1d9fce88 , n59639 );
buf ( R_b69_1e6b3ec8 , n59675 );
buf ( R_356_1d9d3608 , C0 );
buf ( R_2e6_1d9cf008 , C0 );
buf ( R_484_1dd9ee28 , n59676 );
buf ( R_2ec_1d9ceec8 , n59677 );
buf ( R_acb_1e18dba8 , n59678 );
buf ( R_813_1e092848 , n59679 );
buf ( R_4c3_1dda1588 , n59680 );
buf ( R_a47_1e188928 , n59681 );
buf ( R_81d_1e092e88 , n59713 );
buf ( R_8e7_1e09acc8 , n59714 );
buf ( R_5ef_1ddad108 , n59715 );
buf ( R_896_1e094828 , C0 );
buf ( R_bec_1e6b90a8 , n59716 );
buf ( R_b2b_1e6b1808 , n59717 );
buf ( R_4ab_1dda0688 , n59718 );
buf ( R_7e4_1e090ae8 , n59719 );
buf ( R_a33_1e187ca8 , n59720 );
buf ( R_47c_1dd9e928 , n59721 );
buf ( R_8d6_1e09a728 , C0 );
buf ( R_87f_1e096bc8 , n59722 );
buf ( R_5b5_1ddaacc8 , n59754 );
buf ( R_651_1dfb0ea8 , n59759 );
buf ( R_3da_1d9d8888 , C0 );
buf ( R_538_1dda5ea8 , n59760 );
buf ( R_675_1dfb2528 , n59765 );
buf ( R_60f_1dfae568 , n59766 );
buf ( R_29b_1d9fbbc8 , n59773 );
buf ( R_aa6_1e18c988 , C0 );
buf ( R_3bd_1d9d7168 , n59782 );
buf ( R_be5_1e6b8c48 , n59818 );
buf ( R_c0a_1e6ba868 , C0 );
buf ( R_5f5_1ddad4c8 , n59850 );
buf ( R_b4b_1e6b2c08 , n59851 );
buf ( R_7b1_1e08eb08 , n59882 );
buf ( R_95d_1e17f6e8 , n59887 );
buf ( R_a17_1e186b28 , n59888 );
buf ( R_a29_1e187668 , n59897 );
buf ( R_71a_1dfb9148 , C0 );
buf ( R_693_1dfb37e8 , n59898 );
buf ( R_77b_1dfbc8e8 , n59899 );
buf ( R_9c6_1e183d88 , C0 );
buf ( R_3a7_1d9d63a8 , n59900 );
buf ( R_bc0_1e6b7528 , n59901 );
buf ( R_68e_1dfb39c8 , C0 );
buf ( R_335_1d9d1c68 , n59939 );
buf ( R_5eb_1ddace88 , n59940 );
buf ( R_ad7_1e6ae388 , n59941 );
buf ( R_765_1dfbbb28 , n59972 );
buf ( R_387_1d9d4fa8 , n59973 );
buf ( R_9a8_1e1825c8 , n59974 );
buf ( R_632_1dfb0048 , C0 );
buf ( R_6e5_1dfb6b28 , n59983 );
buf ( R_772_1dfbc848 , C0 );
buf ( R_995_1e1819e8 , n59988 );
buf ( R_7d6_1e090728 , C0 );
buf ( R_598_1dda9aa8 , n59989 );
buf ( R_a70_1e18a2c8 , n59990 );
buf ( R_a25_1e1873e8 , n60035 );
buf ( R_bbb_1e6b7208 , n60036 );
buf ( R_6f2_1dfb7848 , C0 );
buf ( R_a41_1e188568 , n60071 );
buf ( R_a66_1e18a188 , C0 );
buf ( R_a3d_1e1882e8 , n60106 );
buf ( R_341_1d9d23e8 , n60144 );
buf ( R_594_1dda9828 , n60145 );
buf ( R_4fe_1dda5868 , C0 );
buf ( R_480_1dd9eba8 , n60146 );
buf ( R_6ab_1dfb46e8 , n60147 );
buf ( R_84c_1e094be8 , n60148 );
buf ( R_660_1dfb1808 , n60149 );
buf ( R_a20_1e1870c8 , n60150 );
buf ( R_abe_1e6b64e8 , C0 );
buf ( R_566_1dda8068 , C0 );
buf ( R_7c8_1e08f968 , n60151 );
buf ( R_5c2_1d9fc2a8 , C0 );
buf ( R_989_1e181268 , n60156 );
buf ( R_8a8_1e098568 , n60157 );
buf ( R_2a4_1d9fc168 , n60158 );
buf ( R_7d5_1e090188 , n60189 );
buf ( R_8fe_1e09c028 , C0 );
buf ( R_3b7_1d9d6da8 , n60190 );
buf ( R_6b8_1dfb4f08 , n60191 );
buf ( R_8b3_1e098c48 , n60192 );
buf ( R_94f_1e17ee28 , n60193 );
buf ( R_9fb_1e1859a8 , n60194 );
buf ( R_a10_1e1866c8 , n60195 );
buf ( R_b36_1e6b23e8 , C0 );
buf ( R_aa0_1e18c0c8 , n60196 );
buf ( R_c1a_1e6bb268 , C0 );
buf ( R_82c_1e0937e8 , n60197 );
buf ( R_4d1_1dda1e48 , n60228 );
buf ( R_6fc_1dfb7988 , n60229 );
buf ( R_9fa_1e185e08 , C0 );
buf ( R_9fc_1e185a48 , n60230 );
buf ( R_a0d_1e1864e8 , n60275 );
buf ( R_be2_1e6b8f68 , C0 );
buf ( R_b02_1e6b8068 , C0 );
buf ( R_a28_1e1875c8 , n60276 );
buf ( R_4fd_1dda39c8 , n60308 );
buf ( R_5fd_1ddad9c8 , n61213 );
buf ( R_873_1e096448 , n61214 );
buf ( R_9fd_1e185ae8 , n61259 );
buf ( R_a6b_1e189fa8 , n61260 );
buf ( R_aa3_1e18c2a8 , n61261 );
buf ( R_738_1dfb9f08 , n61262 );
buf ( R_805_1e091f88 , n61294 );
buf ( R_2f7_1d9cf5a8 , n61295 );
buf ( R_5ba_1ddab4e8 , C0 );
buf ( R_57d_1dda89c8 , n61327 );
buf ( R_475_1dd9e4c8 , n61358 );
buf ( R_433_1d9dbb28 , n61359 );
buf ( R_aed_1e6af148 , n61394 );
buf ( R_4fc_1dda3928 , n61395 );
buf ( R_3a0_1d9d5f48 , n61396 );
buf ( R_3f7_1d9d95a8 , n61397 );
buf ( R_367_1d9d3ba8 , n61398 );
buf ( R_947_1e17e928 , n61399 );
buf ( R_b1a_1e6b1268 , C0 );
buf ( R_525_1dda52c8 , n61431 );
buf ( R_50d_1dda43c8 , n61463 );
buf ( R_390_1d9d5548 , n61464 );
buf ( R_6fe_1dfb7fc8 , C0 );
buf ( R_6f7_1dfb7668 , n61465 );
buf ( R_2ae_1d9fcca8 , C0 );
buf ( R_864_1e095ae8 , n61466 );
buf ( R_9e7_1e184d28 , n61467 );
buf ( R_524_1dda5228 , n61468 );
buf ( R_50c_1dda4328 , n61469 );
buf ( R_9e6_1e185188 , C0 );
buf ( R_9e8_1e184dc8 , n61470 );
buf ( R_9b2_1e183108 , C0 );
buf ( R_7e2_1dfbaf48 , C0 );
buf ( R_622_1dfaf648 , C0 );
buf ( R_b4e_1e184508 , C0 );
buf ( R_a91_1e18b768 , n61501 );
buf ( R_a84_1e18af48 , n61502 );
buf ( R_4ce_1dda2168 , C0 );
buf ( R_bb2_1e6b7168 , C0 );
buf ( R_523_1dda5188 , n61503 );
buf ( R_50b_1dda4288 , n61504 );
buf ( R_9e9_1e184e68 , n61549 );
buf ( R_4f3_1dda3388 , n61550 );
buf ( R_4fb_1dda3888 , n61551 );
buf ( R_4f2_1ddad068 , C0 );
buf ( R_4f4_1dda3428 , n61552 );
buf ( R_55e_1dda7b68 , C0 );
buf ( R_84e_1e095228 , C0 );
buf ( R_a76_1e18ab88 , C0 );
buf ( R_5c9_1ddab948 , n61561 );
buf ( R_343_1d9d2528 , n61562 );
buf ( R_a73_1e18a4a8 , n61563 );
buf ( R_7cd_1e08fc88 , n61594 );
buf ( R_522_1dda55e8 , C0 );
buf ( R_50a_1dda46e8 , C0 );
buf ( R_4f5_1dda34c8 , n61626 );
buf ( R_396_1d9d5e08 , C0 );
buf ( R_7f9_1e091808 , n61658 );
buf ( R_681_1dfb2ca8 , n61718 );
buf ( R_37b_1d9d4828 , n61719 );
buf ( R_639_1dfaffa8 , n61724 );
buf ( R_76d_1dfbc028 , n61755 );
buf ( R_78b_1dfbd2e8 , n61756 );
buf ( R_6a3_1dfb41e8 , n61757 );
buf ( R_9ac_1e182848 , n61758 );
buf ( R_86c_1e095fe8 , n61759 );
buf ( R_c08_1e6ba228 , n61760 );
buf ( R_2fc_1d9cf8c8 , n61761 );
buf ( R_7f0_1e091268 , n61762 );
buf ( R_c31_1e6bbbc8 , n61769 );
buf ( R_a52_1e189508 , C0 );
buf ( R_ab2_1e18d108 , C0 );
buf ( R_28d_1d9fb308 , n61776 );
buf ( R_bcb_1e6b7c08 , n61777 );
buf ( R_4fa_1dda3f68 , C0 );
buf ( R_2bb_1d9fcfc8 , n61778 );
buf ( R_b3f_1e6b2488 , n61779 );
buf ( R_a27_1e187528 , n61780 );
buf ( R_362_1d9d3d88 , C0 );
buf ( R_497_1dd9fa08 , n61781 );
buf ( R_64f_1dfb0d68 , n61782 );
buf ( R_bd7_1e6b8388 , n61783 );
buf ( R_b75_1e6b4648 , n61819 );
buf ( R_98f_1e181628 , n61820 );
buf ( R_6ed_1dfb7028 , n61829 );
buf ( R_7d3_1e090048 , n61830 );
buf ( R_b27_1e6b1588 , n61831 );
buf ( R_39b_1d9d5c28 , n61832 );
buf ( R_8cf_1e099dc8 , n61833 );
buf ( R_689_1dfb31a8 , n61893 );
buf ( R_7c6_1e08fd28 , C0 );
buf ( R_b2d_1e6b1948 , n61929 );
buf ( R_92a_1e092f28 , C0 );
buf ( R_66c_1dfb1f88 , n61930 );
buf ( R_956_1e6b00e8 , C0 );
buf ( R_b96_1e18ce88 , C0 );
buf ( R_bae_1e6b6ee8 , C0 );
buf ( R_94d_1e17ece8 , n61962 );
buf ( R_785_1dfbcf28 , n61993 );
buf ( R_6e2_1dfb6e48 , C0 );
buf ( R_65e_1dfb5cc8 , C0 );
buf ( R_42a_1d9dba88 , C0 );
buf ( R_7e8_1e090d68 , n61994 );
buf ( R_b4d_1e6b2d48 , n62030 );
buf ( R_bff_1e6b9c88 , n62031 );
buf ( R_3c0_1d9d7348 , n62032 );
buf ( R_44a_1d9dce88 , C0 );
buf ( R_2fe_1d9cff08 , C0 );
buf ( R_383_1d9d4d28 , n62033 );
buf ( R_928_1e09d568 , n62034 );
buf ( R_488_1dd9f0a8 , n62035 );
buf ( R_5aa_1ddaaae8 , C0 );
buf ( R_3fd_1d9d9968 , n62066 );
buf ( R_7d0_1e08fe68 , n62067 );
buf ( R_7b4_1e08ece8 , n62068 );
buf ( R_4d8_1dda22a8 , n62069 );
buf ( R_418_1d9daa48 , n62070 );
buf ( R_a43_1e1886a8 , n62071 );
buf ( R_327_1d9d13a8 , n62072 );
buf ( R_849_1e094a08 , n62104 );
buf ( R_b5f_1e6b3888 , n62105 );
buf ( R_4d3_1dda1f88 , n62106 );
buf ( R_a97_1e18bb28 , n62107 );
buf ( R_aba_1e18d608 , C0 );
buf ( R_ab1_1e18cb68 , n62142 );
buf ( R_97f_1e180c28 , n62143 );
buf ( R_788_1dfbd108 , n62144 );
buf ( R_a1c_1e186e48 , n62145 );
buf ( R_b11_1e6b07c8 , n62181 );
buf ( R_a37_1e187f28 , n62182 );
buf ( R_801_1e091d08 , n62214 );
buf ( R_581_1dda8c48 , n62246 );
buf ( R_49d_1dd9fdc8 , n62277 );
buf ( R_56b_1dda7e88 , n62278 );
buf ( R_4da_1dda3ce8 , C0 );
buf ( R_7f2_1e09d6a8 , C0 );
buf ( R_53d_1dda61c8 , n62310 );
buf ( R_3df_1d9d86a8 , n62311 );
buf ( R_429_1d9db4e8 , n62342 );
buf ( R_8dc_1e09a5e8 , n62343 );
buf ( R_a14_1e186948 , n62344 );
buf ( R_9d6_1e186088 , C0 );
buf ( R_add_1e6ae748 , n62379 );
buf ( R_b6d_1e6b4148 , n62415 );
buf ( R_c1e_1e6b4e68 , C0 );
buf ( R_7fd_1e091a88 , n62447 );
buf ( R_859_1e095408 , n62479 );
buf ( R_b23_1e6b1308 , n62480 );
buf ( R_afc_1e6afaa8 , n62481 );
buf ( R_913_1e09c848 , n62482 );
buf ( R_450_1d9dcd48 , n62483 );
buf ( R_7cb_1e08fb48 , n62484 );
buf ( R_b38_1e6b2028 , n62485 );
buf ( R_a26_1e187988 , C0 );
buf ( R_74c_1dfbab88 , n62486 );
buf ( R_35b_1d9d3428 , n62487 );
buf ( R_962_1e17ff08 , C0 );
buf ( R_2e7_1d9ceba8 , n62488 );
buf ( R_8c0_1e099468 , n62489 );
buf ( R_8c7_1e0998c8 , n62490 );
buf ( R_afe_1e6b5d68 , C0 );
buf ( R_977_1e180728 , n62491 );
buf ( R_925_1e09d388 , n62523 );
buf ( R_919_1e09cc08 , n62555 );
buf ( R_728_1dfb9508 , n62556 );
buf ( R_43a_1d9dc488 , C0 );
buf ( R_bf0_1e6b9328 , n62557 );
buf ( R_9a3_1e1822a8 , n62558 );
buf ( R_3af_1d9d68a8 , n62559 );
buf ( R_930_1e09da68 , n62560 );
buf ( R_90c_1e09c3e8 , n62561 );
buf ( R_5a9_1ddaa548 , n62593 );
buf ( R_659_1dfb13a8 , n62598 );
buf ( R_c0f_1e6ba688 , n62599 );
buf ( R_307_1d9cffa8 , n62600 );
buf ( R_8bc_1e0991e8 , n62601 );
buf ( R_2ed_1d9cef68 , n62606 );
buf ( R_770_1dfbc208 , n62607 );
buf ( R_34b_1d9d2a28 , n62608 );
buf ( R_37f_1d9d4aa8 , n62609 );
buf ( R_5f4_1ddad428 , n62610 );
buf ( R_779_1dfbc7a8 , n62641 );
buf ( R_46a_1dd9f468 , C0 );
buf ( R_be0_1e6b8928 , n62642 );
buf ( R_bd3_1e6b8108 , n62643 );
buf ( R_466_1d9d9c88 , C0 );
buf ( R_77e_1dfbcfc8 , C0 );
buf ( R_575_1dda84c8 , n62675 );
buf ( R_4ff_1dda3b08 , n62676 );
buf ( R_a18_1e186bc8 , n62677 );
buf ( R_bda_1e6b8a68 , C0 );
buf ( R_31b_1d9d0c28 , n62678 );
buf ( R_3c6_1d9d7c08 , C0 );
buf ( R_792_1dfbdc48 , C0 );
buf ( R_54b_1dda6a88 , n62679 );
buf ( R_6bd_1dfb5228 , n62739 );
buf ( R_b50_1e6b2f28 , n62740 );
buf ( R_a61_1e189968 , n62775 );
buf ( R_b8b_1e6b5408 , n62776 );
buf ( R_b80_1e6b4d28 , n62777 );
buf ( R_33c_1d9d20c8 , n62778 );
buf ( R_3c3_1d9d7528 , n62779 );
buf ( R_666_1dfb20c8 , C0 );
buf ( R_c2a_1e6bbc68 , C0 );
buf ( R_359_1d9d32e8 , n62817 );
buf ( R_415_1d9da868 , n62848 );
buf ( R_5da_1ddac8e8 , C0 );
buf ( R_577_1dda8608 , n62849 );
buf ( R_637_1dfafe68 , n62850 );
buf ( R_9f7_1e185728 , n62851 );
buf ( R_570_1dda81a8 , n62852 );
buf ( R_9f6_1e185b88 , C0 );
buf ( R_9f8_1e1857c8 , n62853 );
buf ( R_a6e_1e18a688 , C0 );
buf ( R_73d_1dfba228 , n62862 );
buf ( R_293_1d9fb6c8 , n62869 );
buf ( R_884_1e096ee8 , n62870 );
buf ( R_3a2_1d9d6588 , C0 );
buf ( R_9f9_1e185868 , n62915 );
buf ( R_957_1e17f328 , n62916 );
buf ( R_ab6_1e6b5fe8 , C0 );
buf ( R_760_1dfbb808 , n62917 );
buf ( R_a21_1e187168 , n62962 );
buf ( R_bb7_1e6b6f88 , n62963 );
buf ( R_9eb_1e184fa8 , n62964 );
buf ( R_a3f_1e188428 , n62965 );
buf ( R_747_1dfba868 , n62966 );
buf ( R_4bf_1dda1308 , n62967 );
buf ( R_3d7_1d9d81a8 , n62968 );
buf ( R_4a4_1dda0228 , n62969 );
buf ( R_441_1d9dc3e8 , n63000 );
buf ( R_7ce_1e090228 , C0 );
buf ( R_85a_1e0959a8 , C0 );
buf ( R_66f_1dfb2168 , n63001 );
buf ( R_9ea_1e185408 , C0 );
buf ( R_9ec_1e185048 , n63002 );
buf ( R_a3b_1e1881a8 , n63003 );
buf ( R_ad4_1e6ae1a8 , n63004 );
buf ( R_b94_1e6b59a8 , n63005 );
buf ( R_467_1d9ddba8 , n63006 );
buf ( R_96e_1e180688 , C0 );
buf ( R_323_1d9d1128 , n63007 );
buf ( R_6ea_1dfb7348 , C0 );
buf ( R_6ca_1dfb5f48 , C0 );
buf ( R_9ed_1e1850e8 , n63052 );
buf ( R_ae7_1e6aed88 , n63053 );
buf ( R_830_1e093a68 , n63054 );
buf ( R_6d9_1dfb63a8 , n63063 );
buf ( R_8e6_1e08f0a8 , C0 );
buf ( R_6a1_1dfb40a8 , n63123 );
buf ( R_710_1dfb8608 , n63124 );
buf ( R_b41_1e6b25c8 , n63160 );
buf ( R_732_1dfba048 , C0 );
buf ( R_6df_1dfb6768 , n63161 );
buf ( R_a11_1e186768 , n63206 );
buf ( R_a8f_1e18b628 , n63207 );
buf ( R_b97_1e6b5b88 , n63208 );
buf ( R_bc6_1e6b7de8 , C0 );
buf ( R_4db_1dda2488 , n63209 );
buf ( R_9d7_1e184328 , n63210 );
buf ( R_b29_1e6b16c8 , n63246 );
buf ( R_57e_1dda8f68 , C0 );
buf ( R_29a_1d9fbb28 , n63253 );
buf ( R_36f_1d9d40a8 , n63254 );
buf ( R_3e4_1d9d89c8 , n63255 );
buf ( R_7bc_1e08f1e8 , n63256 );
buf ( R_87e_1e097028 , C0 );
buf ( R_b1c_1e6b0ea8 , n63257 );
buf ( R_aab_1e18c7a8 , n63258 );
buf ( R_96c_1e180048 , n63259 );
buf ( R_551_1dda6e48 , n63291 );
buf ( R_6d4_1dfb6088 , n63292 );
buf ( R_2af_1d9fc848 , n63293 );
buf ( R_479_1dd9e748 , n63324 );
buf ( R_5a3_1ddaa188 , n63325 );
buf ( R_672_1dfb2848 , C0 );
buf ( R_587_1dda9008 , n63326 );
buf ( R_767_1dfbbc68 , n63327 );
buf ( R_395_1d9d5868 , n63336 );
buf ( R_3e9_1d9d8ce8 , n63345 );
buf ( R_2f8_1d9cf648 , n63346 );
buf ( R_64c_1dfb0b88 , n63347 );
buf ( R_5e1_1ddac848 , n63378 );
buf ( R_3fc_1d9d98c8 , n63379 );
buf ( R_468_1d9ddc48 , n63380 );
buf ( R_3ba_1d9d7488 , C0 );
buf ( R_55b_1dda7488 , n63381 );
buf ( R_67e_1dfb2fc8 , C0 );
buf ( R_8b7_1e098ec8 , n63382 );
buf ( R_879_1e096808 , n63414 );
buf ( R_b5b_1e6b3608 , n63415 );
buf ( R_a82_1e18b588 , C0 );
buf ( R_ae5_1e6aec48 , n63450 );
buf ( R_84b_1e094b48 , n63451 );
buf ( R_99e_1e182488 , C0 );
buf ( R_6dc_1dfb6588 , n63452 );
buf ( R_3ad_1d9d6768 , n63461 );
buf ( R_a59_1e189468 , n63496 );
buf ( R_b62_1e6ba368 , C0 );
buf ( R_731_1dfb9aa8 , n63505 );
buf ( R_3f1_1d9d91e8 , n63514 );
buf ( R_620_1dfaf008 , n63515 );
buf ( R_67d_1dfb2a28 , n63520 );
buf ( R_adf_1e6ae888 , n63521 );
buf ( R_349_1d9d28e8 , n63559 );
buf ( R_3d1_1d9d7de8 , n63568 );
buf ( R_3f4_1d9d93c8 , n63569 );
buf ( R_80a_1e0927a8 , C0 );
buf ( R_350_1d9d2d48 , n63570 );
buf ( R_a50_1e188ec8 , n63571 );
buf ( R_bc1_1e6b75c8 , n63606 );
buf ( R_b85_1e6b5048 , n63642 );
buf ( R_5d7_1ddac208 , n63643 );
buf ( R_7a2_1ddada68 , C0 );
buf ( R_539_1dda5f48 , n63675 );
buf ( R_bbc_1e6b72a8 , n63676 );
buf ( R_c14_1e6ba9a8 , n63677 );
buf ( R_6c8_1dfb5908 , n63678 );
buf ( R_4c8_1dda18a8 , n63679 );
buf ( R_360_1d9d3748 , n63680 );
buf ( R_2e2_1d9ced88 , C0 );
buf ( R_936_1e17e388 , C0 );
buf ( R_9f3_1e1854a8 , n63681 );
buf ( R_b25_1e6b1448 , n63717 );
buf ( R_b0a_1e6b0868 , C0 );
buf ( R_b56_1e6b87e8 , C0 );
buf ( R_bf4_1e6b95a8 , n63718 );
buf ( R_95f_1e17f828 , n63719 );
buf ( R_3b5_1d9d6c68 , n63728 );
buf ( R_52a_1dda5fe8 , C0 );
buf ( R_9f2_1e185908 , C0 );
buf ( R_9f4_1e185548 , n63729 );
buf ( R_686_1dfb34c8 , C0 );
buf ( R_2bc_1d9fd068 , n63730 );
buf ( R_7a6_1e08e928 , C0 );
buf ( R_9ef_1e185228 , n63731 );
buf ( R_b1e_1e6b78e8 , C0 );
buf ( R_bfb_1e6b9a08 , n63732 );
buf ( R_378_1d9d4648 , n63733 );
buf ( R_9ee_1e185688 , C0 );
buf ( R_9f0_1e1852c8 , n63734 );
buf ( R_9f5_1e1855e8 , n63779 );
buf ( R_4bd_1dda11c8 , n63808 );
buf ( R_5af_1ddaa908 , n63809 );
buf ( R_822_1e097f28 , C0 );
buf ( R_872_1e0968a8 , C0 );
buf ( R_9f1_1e185368 , n63854 );
buf ( R_337_1d9d1da8 , n63855 );
buf ( R_707_1dfb8068 , n63856 );
buf ( R_755_1dfbb128 , n63887 );
buf ( R_8f9_1e09b808 , n63918 );
buf ( R_432_1d9dbf88 , C0 );
buf ( R_8af_1e0989c8 , n63919 );
buf ( R_bc5_1e6b7848 , n63955 );
buf ( R_934_1e09dce8 , n63956 );
buf ( R_469_1d9ddce8 , n63987 );
buf ( R_572_1dda87e8 , C0 );
buf ( R_863_1e095a48 , n63988 );
buf ( R_958_1e17f3c8 , n63989 );
buf ( R_742_1dfbaa48 , C0 );
buf ( R_2a5_1d9fc208 , n63994 );
buf ( R_a9a_1e18c208 , C0 );
buf ( R_af9_1e6af8c8 , n64029 );
buf ( R_9c1_1e183568 , n64034 );
buf ( R_83c_1e0941e8 , n64035 );
buf ( R_a81_1e18ad68 , n64070 );
buf ( R_c19_1e6bacc8 , n64106 );
buf ( R_91c_1e09cde8 , n64107 );
buf ( R_4ac_1dda0728 , n64108 );
buf ( R_bf8_1e6b9828 , n64109 );
buf ( R_5be_1dda7168 , C0 );
buf ( R_93b_1e17e1a8 , n64110 );
buf ( R_63c_1dfb0188 , n64111 );
buf ( R_7e1_1e090908 , n64142 );
buf ( R_7ba_1e08f5a8 , C0 );
buf ( R_6b2_1dfb5048 , C0 );
buf ( R_4dc_1dda2528 , n64143 );
buf ( R_79e_1e08e428 , C0 );
buf ( R_492_1dd9fbe8 , C0 );
buf ( R_750_1dfbae08 , n64144 );
buf ( R_9d8_1e1843c8 , n64145 );
buf ( R_365_1d9d3a68 , n64183 );
buf ( R_994_1e181948 , n64184 );
buf ( R_95c_1e17f648 , n64185 );
buf ( R_2ff_1d9cfaa8 , n64186 );
buf ( R_89b_1e097d48 , n64187 );
buf ( R_827_1e0934c8 , n64188 );
buf ( R_332_1d9d1f88 , C0 );
buf ( R_9a7_1e182528 , n64189 );
buf ( R_834_1e093ce8 , n64190 );
buf ( R_30b_1d9d0228 , n64191 );
buf ( R_86b_1e095f48 , n64192 );
buf ( R_649_1dfb09a8 , n64197 );
buf ( R_a1d_1e186ee8 , n64242 );
buf ( R_b59_1e6b34c8 , n64278 );
buf ( R_bb3_1e6b6d08 , n64279 );
buf ( R_796_1e08e1a8 , C0 );
buf ( R_941_1e17e568 , n64311 );
buf ( R_be9_1e6b8ec8 , n64347 );
buf ( R_485_1dd9eec8 , n64378 );
buf ( R_317_1d9d09a8 , n64379 );
buf ( R_8a3_1e098248 , n64380 );
buf ( R_49e_1dda0368 , C0 );
buf ( R_9c0_1e1834c8 , n64381 );
buf ( R_32c_1d9d16c8 , n64382 );
buf ( R_6d6_1dfb66c8 , C0 );
buf ( R_a15_1e1869e8 , n64427 );
buf ( R_33e_1d9d2708 , C0 );
buf ( R_38c_1d9d52c8 , n64428 );
buf ( R_75b_1dfbb4e8 , n64429 );
buf ( R_ac4_1e18d748 , n64430 );
buf ( R_5d9_1ddac348 , n64461 );
buf ( R_546_1dda6c68 , C0 );
buf ( R_2be_1d9fd6a8 , C0 );
buf ( R_b76_1e6b4be8 , C0 );
buf ( R_975_1e1805e8 , n64466 );
buf ( R_5c3_1ddab588 , n64467 );
buf ( R_500_1dda3ba8 , n64468 );
buf ( R_889_1e097208 , n64500 );
buf ( R_988_1e1811c8 , n64501 );
buf ( R_c2c_1e6bb8a8 , n64502 );
buf ( R_b98_1e6b5c28 , n64503 );
buf ( R_47d_1dd9e9c8 , n64534 );
buf ( R_417_1d9da9a8 , n64535 );
buf ( R_819_1e092c08 , n64567 );
buf ( R_8f8_1e09b768 , n64568 );
buf ( R_942_1e17eb08 , C0 );
buf ( R_ad1_1e6adfc8 , n64603 );
buf ( R_8ce_1e09a228 , C0 );
buf ( R_563_1dda7988 , n64604 );
buf ( R_2e8_1d9cec48 , n64605 );
buf ( R_838_1e093f68 , n64606 );
buf ( R_aee_1e187c08 , C0 );
buf ( R_641_1dfb04a8 , n64611 );
buf ( R_c16_1e6b41e8 , C0 );
buf ( R_6c3_1dfb55e8 , n64612 );
buf ( R_5f3_1ddad388 , n64613 );
buf ( R_558_1dda72a8 , n64614 );
buf ( R_821_1e093108 , n64646 );
buf ( R_a5f_1e189828 , n64647 );
buf ( R_3cd_1d9d7b68 , n64656 );
buf ( R_80f_1e0925c8 , n64657 );
buf ( R_724_1dfb9288 , n64658 );
buf ( R_848_1e094968 , n64659 );
buf ( R_9bf_1e183428 , n64660 );
buf ( R_a19_1e186c68 , n64705 );
buf ( R_baf_1e6b6a88 , n64706 );
buf ( R_64a_1dfb0f48 , C0 );
buf ( R_aa8_1e18c5c8 , n64707 );
buf ( R_6be_1dfb57c8 , C0 );
buf ( R_481_1dd9ec48 , n64738 );
buf ( R_428_1d9db448 , n64739 );
buf ( R_be6_1e6b91e8 , C0 );
buf ( R_44f_1d9dcca8 , n64740 );
buf ( R_5b4_1ddaac28 , n64741 );
buf ( R_629_1dfaf5a8 , n64746 );
buf ( R_78f_1dfbd568 , n64747 );
buf ( R_91f_1e09cfc8 , n64748 );
buf ( R_858_1e095368 , n64749 );
buf ( R_afb_1e6afa08 , n64750 );
buf ( R_3fb_1d9d9828 , n64751 );
buf ( R_922_1e091628 , C0 );
buf ( R_916_1e09cf28 , C0 );
buf ( R_8a1_1e098108 , n64760 );
buf ( R_8db_1e09a548 , n64761 );
buf ( R_b32_1e6b2168 , C0 );
buf ( R_411_1d9da5e8 , n64792 );
buf ( R_6b0_1dfb4a08 , n64793 );
buf ( R_5d1_1ddabe48 , n64824 );
buf ( R_7df_1e0907c8 , n64825 );
buf ( R_b04_1e6affa8 , n64826 );
buf ( R_45a_1d9dd888 , C0 );
buf ( R_814_1e0928e8 , n64827 );
buf ( R_665_1dfb1b28 , n64832 );
buf ( R_69e_1dfb43c8 , C0 );
buf ( R_b42_1e6b2b68 , C0 );
buf ( R_555_1dda70c8 , n64864 );
buf ( R_374_1d9d43c8 , n64865 );
buf ( R_352_1d9d3388 , C0 );
buf ( R_2a6_1d9fc7a8 , C0 );
buf ( R_756_1dfbb6c8 , C0 );
buf ( R_bd6_1e6b3568 , C0 );
buf ( R_baa_1e18d888 , C0 );
buf ( R_5b9_1ddaaf48 , n64897 );
buf ( R_3ec_1d9d8ec8 , n64898 );
buf ( n10613 , RI21a19c60_2);
buf ( n10614 , n10613 );
buf ( n10615 , RI21a5daf0_1);
buf ( n10616 , n10615 );
buf ( n10617 , RI2107e620_463);
not ( n10618 , n10617 );
buf ( n10619 , n10618 );
buf ( n10620 , n10619 );
buf ( n10621 , RI21a139f0_68);
buf ( n10622 , n10621 );
buf ( n10623 , RI21084368_418);
buf ( n10624 , n10623 );
xor ( n10625 , n10622 , n10624 );
buf ( n10626 , n10625 );
buf ( n10627 , n10626 );
buf ( n10628 , RI21079850_497);
buf ( n10629 , n10628 );
xor ( n10630 , n10627 , n10629 );
buf ( n10631 , n10630 );
buf ( n10632 , n10631 );
buf ( n10633 , n10632 );
not ( n10634 , n10633 );
buf ( n10635 , n10634 );
buf ( n10636 , n10635 );
not ( n10637 , n10636 );
buf ( n10638 , RI21a12820_78);
buf ( n10639 , n10638 );
buf ( n10640 , RI210beb08_292);
buf ( n10641 , n10640 );
and ( n10642 , n10639 , n10641 );
buf ( n10643 , RI21a12898_77);
buf ( n10644 , n10643 );
buf ( n10645 , RI210beb80_291);
buf ( n10646 , n10645 );
and ( n10647 , n10644 , n10646 );
buf ( n10648 , RI21a12910_76);
buf ( n10649 , n10648 );
buf ( n10650 , RI210bf3f0_290);
buf ( n10651 , n10650 );
and ( n10652 , n10649 , n10651 );
buf ( n10653 , RI21a12988_75);
buf ( n10654 , n10653 );
buf ( n10655 , RI210bf468_289);
buf ( n10656 , n10655 );
and ( n10657 , n10654 , n10656 );
buf ( n10658 , RI21a13090_74);
buf ( n10659 , n10658 );
buf ( n10660 , RI210bf4e0_288);
buf ( n10661 , n10660 );
and ( n10662 , n10659 , n10661 );
buf ( n10663 , RI21a13108_73);
buf ( n10664 , n10663 );
buf ( n10665 , RI210bf558_287);
buf ( n10666 , n10665 );
and ( n10667 , n10664 , n10666 );
buf ( n10668 , RI21a13180_72);
buf ( n10669 , n10668 );
buf ( n10670 , RI210bfdc8_286);
buf ( n10671 , n10670 );
and ( n10672 , n10669 , n10671 );
buf ( n10673 , RI21a131f8_71);
buf ( n10674 , n10673 );
buf ( n10675 , RI210bfe40_285);
buf ( n10676 , n10675 );
and ( n10677 , n10674 , n10676 );
buf ( n10678 , RI21a13270_70);
buf ( n10679 , n10678 );
buf ( n10680 , RI210bfeb8_284);
buf ( n10681 , n10680 );
and ( n10682 , n10679 , n10681 );
buf ( n10683 , RI21a132e8_69);
buf ( n10684 , n10683 );
buf ( n10685 , RI210bff30_283);
buf ( n10686 , n10685 );
and ( n10687 , n10684 , n10686 );
buf ( n10688 , RI21a116c8_87);
buf ( n10689 , n10688 );
buf ( n10690 , RI210bd6e0_301);
buf ( n10691 , n10690 );
and ( n10692 , n10689 , n10691 );
buf ( n10693 , RI21a11dd0_86);
buf ( n10694 , n10693 );
buf ( n10695 , RI210bd758_300);
buf ( n10696 , n10695 );
and ( n10697 , n10694 , n10696 );
buf ( n10698 , RI21a11e48_85);
buf ( n10699 , n10698 );
buf ( n10700 , RI210bd7d0_299);
buf ( n10701 , n10700 );
and ( n10702 , n10699 , n10701 );
buf ( n10703 , RI21a11ec0_84);
buf ( n10704 , n10703 );
buf ( n10705 , RI210be040_298);
buf ( n10706 , n10705 );
and ( n10707 , n10704 , n10706 );
buf ( n10708 , RI21a11f38_83);
buf ( n10709 , n10708 );
buf ( n10710 , RI210be0b8_297);
buf ( n10711 , n10710 );
and ( n10712 , n10709 , n10711 );
buf ( n10713 , RI21a11fb0_82);
buf ( n10714 , n10713 );
buf ( n10715 , RI210be130_296);
buf ( n10716 , n10715 );
and ( n10717 , n10714 , n10716 );
buf ( n10718 , RI21a12028_81);
buf ( n10719 , n10718 );
buf ( n10720 , RI210be1a8_295);
buf ( n10721 , n10720 );
and ( n10722 , n10719 , n10721 );
buf ( n10723 , RI21a12730_80);
buf ( n10724 , n10723 );
buf ( n10725 , RI210bea18_294);
buf ( n10726 , n10725 );
and ( n10727 , n10724 , n10726 );
buf ( n10728 , RI21a127a8_79);
buf ( n10729 , n10728 );
buf ( n10730 , RI210bea90_293);
buf ( n10731 , n10730 );
and ( n10732 , n10729 , n10731 );
and ( n10733 , n10622 , n10624 );
and ( n10734 , n10731 , n10733 );
and ( n10735 , n10729 , n10733 );
or ( n10736 , n10732 , n10734 , n10735 );
and ( n10737 , n10726 , n10736 );
and ( n10738 , n10724 , n10736 );
or ( n10739 , n10727 , n10737 , n10738 );
and ( n10740 , n10721 , n10739 );
and ( n10741 , n10719 , n10739 );
or ( n10742 , n10722 , n10740 , n10741 );
and ( n10743 , n10716 , n10742 );
and ( n10744 , n10714 , n10742 );
or ( n10745 , n10717 , n10743 , n10744 );
and ( n10746 , n10711 , n10745 );
and ( n10747 , n10709 , n10745 );
or ( n10748 , n10712 , n10746 , n10747 );
and ( n10749 , n10706 , n10748 );
and ( n10750 , n10704 , n10748 );
or ( n10751 , n10707 , n10749 , n10750 );
and ( n10752 , n10701 , n10751 );
and ( n10753 , n10699 , n10751 );
or ( n10754 , n10702 , n10752 , n10753 );
and ( n10755 , n10696 , n10754 );
and ( n10756 , n10694 , n10754 );
or ( n10757 , n10697 , n10755 , n10756 );
and ( n10758 , n10691 , n10757 );
and ( n10759 , n10689 , n10757 );
or ( n10760 , n10692 , n10758 , n10759 );
and ( n10761 , n10686 , n10760 );
and ( n10762 , n10684 , n10760 );
or ( n10763 , n10687 , n10761 , n10762 );
and ( n10764 , n10681 , n10763 );
and ( n10765 , n10679 , n10763 );
or ( n10766 , n10682 , n10764 , n10765 );
and ( n10767 , n10676 , n10766 );
and ( n10768 , n10674 , n10766 );
or ( n10769 , n10677 , n10767 , n10768 );
and ( n10770 , n10671 , n10769 );
and ( n10771 , n10669 , n10769 );
or ( n10772 , n10672 , n10770 , n10771 );
and ( n10773 , n10666 , n10772 );
and ( n10774 , n10664 , n10772 );
or ( n10775 , n10667 , n10773 , n10774 );
and ( n10776 , n10661 , n10775 );
and ( n10777 , n10659 , n10775 );
or ( n10778 , n10662 , n10776 , n10777 );
and ( n10779 , n10656 , n10778 );
and ( n10780 , n10654 , n10778 );
or ( n10781 , n10657 , n10779 , n10780 );
and ( n10782 , n10651 , n10781 );
and ( n10783 , n10649 , n10781 );
or ( n10784 , n10652 , n10782 , n10783 );
and ( n10785 , n10646 , n10784 );
and ( n10786 , n10644 , n10784 );
or ( n10787 , n10647 , n10785 , n10786 );
and ( n10788 , n10641 , n10787 );
and ( n10789 , n10639 , n10787 );
or ( n10790 , n10642 , n10788 , n10789 );
buf ( n10791 , n10790 );
buf ( n10792 , n10791 );
xor ( n10793 , n10639 , n10641 );
xor ( n10794 , n10793 , n10787 );
buf ( n10795 , n10794 );
buf ( n10796 , n10795 );
buf ( n10797 , RI21077f00_507);
buf ( n10798 , n10797 );
not ( n10799 , n10798 );
and ( n10800 , n10796 , n10799 );
xor ( n10801 , n10644 , n10646 );
xor ( n10802 , n10801 , n10784 );
buf ( n10803 , n10802 );
buf ( n10804 , n10803 );
buf ( n10805 , RI21077f78_506);
buf ( n10806 , n10805 );
not ( n10807 , n10806 );
and ( n10808 , n10804 , n10807 );
xor ( n10809 , n10649 , n10651 );
xor ( n10810 , n10809 , n10781 );
buf ( n10811 , n10810 );
buf ( n10812 , n10811 );
buf ( n10813 , RI21078a40_505);
buf ( n10814 , n10813 );
not ( n10815 , n10814 );
and ( n10816 , n10812 , n10815 );
xor ( n10817 , n10654 , n10656 );
xor ( n10818 , n10817 , n10778 );
buf ( n10819 , n10818 );
buf ( n10820 , n10819 );
buf ( n10821 , RI21078ab8_504);
buf ( n10822 , n10821 );
not ( n10823 , n10822 );
and ( n10824 , n10820 , n10823 );
xor ( n10825 , n10659 , n10661 );
xor ( n10826 , n10825 , n10775 );
buf ( n10827 , n10826 );
buf ( n10828 , n10827 );
buf ( n10829 , RI21078b30_503);
buf ( n10830 , n10829 );
not ( n10831 , n10830 );
and ( n10832 , n10828 , n10831 );
xor ( n10833 , n10664 , n10666 );
xor ( n10834 , n10833 , n10772 );
buf ( n10835 , n10834 );
buf ( n10836 , n10835 );
buf ( n10837 , RI21078ba8_502);
buf ( n10838 , n10837 );
not ( n10839 , n10838 );
and ( n10840 , n10836 , n10839 );
xor ( n10841 , n10669 , n10671 );
xor ( n10842 , n10841 , n10769 );
buf ( n10843 , n10842 );
buf ( n10844 , n10843 );
buf ( n10845 , RI21078c20_501);
buf ( n10846 , n10845 );
not ( n10847 , n10846 );
and ( n10848 , n10844 , n10847 );
xor ( n10849 , n10674 , n10676 );
xor ( n10850 , n10849 , n10766 );
buf ( n10851 , n10850 );
buf ( n10852 , n10851 );
buf ( n10853 , RI21078c98_500);
buf ( n10854 , n10853 );
not ( n10855 , n10854 );
and ( n10856 , n10852 , n10855 );
xor ( n10857 , n10679 , n10681 );
xor ( n10858 , n10857 , n10763 );
buf ( n10859 , n10858 );
buf ( n10860 , n10859 );
buf ( n10861 , RI21079760_499);
buf ( n10862 , n10861 );
not ( n10863 , n10862 );
and ( n10864 , n10860 , n10863 );
xor ( n10865 , n10684 , n10686 );
xor ( n10866 , n10865 , n10760 );
buf ( n10867 , n10866 );
buf ( n10868 , n10867 );
buf ( n10869 , RI210797d8_498);
buf ( n10870 , n10869 );
not ( n10871 , n10870 );
and ( n10872 , n10868 , n10871 );
xor ( n10873 , n10689 , n10691 );
xor ( n10874 , n10873 , n10757 );
buf ( n10875 , n10874 );
buf ( n10876 , n10875 );
buf ( n10877 , RI21077078_516);
buf ( n10878 , n10877 );
not ( n10879 , n10878 );
and ( n10880 , n10876 , n10879 );
xor ( n10881 , n10694 , n10696 );
xor ( n10882 , n10881 , n10754 );
buf ( n10883 , n10882 );
buf ( n10884 , n10883 );
buf ( n10885 , RI210770f0_515);
buf ( n10886 , n10885 );
not ( n10887 , n10886 );
and ( n10888 , n10884 , n10887 );
xor ( n10889 , n10699 , n10701 );
xor ( n10890 , n10889 , n10751 );
buf ( n10891 , n10890 );
buf ( n10892 , n10891 );
buf ( n10893 , RI21077168_514);
buf ( n10894 , n10893 );
not ( n10895 , n10894 );
and ( n10896 , n10892 , n10895 );
xor ( n10897 , n10704 , n10706 );
xor ( n10898 , n10897 , n10748 );
buf ( n10899 , n10898 );
buf ( n10900 , n10899 );
buf ( n10901 , RI210771e0_513);
buf ( n10902 , n10901 );
not ( n10903 , n10902 );
and ( n10904 , n10900 , n10903 );
xor ( n10905 , n10709 , n10711 );
xor ( n10906 , n10905 , n10745 );
buf ( n10907 , n10906 );
buf ( n10908 , n10907 );
buf ( n10909 , RI21077258_512);
buf ( n10910 , n10909 );
not ( n10911 , n10910 );
and ( n10912 , n10908 , n10911 );
xor ( n10913 , n10714 , n10716 );
xor ( n10914 , n10913 , n10742 );
buf ( n10915 , n10914 );
buf ( n10916 , n10915 );
buf ( n10917 , RI21077d20_511);
buf ( n10918 , n10917 );
not ( n10919 , n10918 );
and ( n10920 , n10916 , n10919 );
xor ( n10921 , n10719 , n10721 );
xor ( n10922 , n10921 , n10739 );
buf ( n10923 , n10922 );
buf ( n10924 , n10923 );
buf ( n10925 , RI21077d98_510);
buf ( n10926 , n10925 );
not ( n10927 , n10926 );
and ( n10928 , n10924 , n10927 );
xor ( n10929 , n10724 , n10726 );
xor ( n10930 , n10929 , n10736 );
buf ( n10931 , n10930 );
buf ( n10932 , n10931 );
buf ( n10933 , RI21077e10_509);
buf ( n10934 , n10933 );
not ( n10935 , n10934 );
and ( n10936 , n10932 , n10935 );
xor ( n10937 , n10729 , n10731 );
xor ( n10938 , n10937 , n10733 );
buf ( n10939 , n10938 );
buf ( n10940 , n10939 );
buf ( n10941 , RI21077e88_508);
buf ( n10942 , n10941 );
not ( n10943 , n10942 );
and ( n10944 , n10940 , n10943 );
not ( n10945 , n10629 );
or ( n10946 , n10627 , n10945 );
and ( n10947 , n10943 , n10946 );
and ( n10948 , n10940 , n10946 );
or ( n10949 , n10944 , n10947 , n10948 );
and ( n10950 , n10935 , n10949 );
and ( n10951 , n10932 , n10949 );
or ( n10952 , n10936 , n10950 , n10951 );
and ( n10953 , n10927 , n10952 );
and ( n10954 , n10924 , n10952 );
or ( n10955 , n10928 , n10953 , n10954 );
and ( n10956 , n10919 , n10955 );
and ( n10957 , n10916 , n10955 );
or ( n10958 , n10920 , n10956 , n10957 );
and ( n10959 , n10911 , n10958 );
and ( n10960 , n10908 , n10958 );
or ( n10961 , n10912 , n10959 , n10960 );
and ( n10962 , n10903 , n10961 );
and ( n10963 , n10900 , n10961 );
or ( n10964 , n10904 , n10962 , n10963 );
and ( n10965 , n10895 , n10964 );
and ( n10966 , n10892 , n10964 );
or ( n10967 , n10896 , n10965 , n10966 );
and ( n10968 , n10887 , n10967 );
and ( n10969 , n10884 , n10967 );
or ( n10970 , n10888 , n10968 , n10969 );
and ( n10971 , n10879 , n10970 );
and ( n10972 , n10876 , n10970 );
or ( n10973 , n10880 , n10971 , n10972 );
and ( n10974 , n10871 , n10973 );
and ( n10975 , n10868 , n10973 );
or ( n10976 , n10872 , n10974 , n10975 );
and ( n10977 , n10863 , n10976 );
and ( n10978 , n10860 , n10976 );
or ( n10979 , n10864 , n10977 , n10978 );
and ( n10980 , n10855 , n10979 );
and ( n10981 , n10852 , n10979 );
or ( n10982 , n10856 , n10980 , n10981 );
and ( n10983 , n10847 , n10982 );
and ( n10984 , n10844 , n10982 );
or ( n10985 , n10848 , n10983 , n10984 );
and ( n10986 , n10839 , n10985 );
and ( n10987 , n10836 , n10985 );
or ( n10988 , n10840 , n10986 , n10987 );
and ( n10989 , n10831 , n10988 );
and ( n10990 , n10828 , n10988 );
or ( n10991 , n10832 , n10989 , n10990 );
and ( n10992 , n10823 , n10991 );
and ( n10993 , n10820 , n10991 );
or ( n10994 , n10824 , n10992 , n10993 );
and ( n10995 , n10815 , n10994 );
and ( n10996 , n10812 , n10994 );
or ( n10997 , n10816 , n10995 , n10996 );
and ( n10998 , n10807 , n10997 );
and ( n10999 , n10804 , n10997 );
or ( n11000 , n10808 , n10998 , n10999 );
and ( n11001 , n10799 , n11000 );
and ( n11002 , n10796 , n11000 );
or ( n11003 , n10800 , n11001 , n11002 );
or ( n11004 , n10792 , n11003 );
not ( n11005 , n11004 );
buf ( n11006 , n11005 );
buf ( n11007 , n11006 );
not ( n11008 , n11007 );
xor ( n11009 , n10940 , n10943 );
xor ( n11010 , n11009 , n10946 );
buf ( n11011 , n11010 );
buf ( n11012 , n11011 );
and ( n11013 , n11008 , n11012 );
not ( n11014 , n11012 );
not ( n11015 , n10632 );
xor ( n11016 , n11014 , n11015 );
and ( n11017 , n11016 , n11007 );
or ( n11018 , n11013 , n11017 );
buf ( n11019 , n11018 );
not ( n11020 , n11019 );
buf ( n11021 , n11020 );
buf ( n11022 , n11021 );
not ( n11023 , n11022 );
or ( n11024 , n10637 , n11023 );
not ( n11025 , n11007 );
xor ( n11026 , n10932 , n10935 );
xor ( n11027 , n11026 , n10949 );
buf ( n11028 , n11027 );
buf ( n11029 , n11028 );
and ( n11030 , n11025 , n11029 );
not ( n11031 , n11029 );
and ( n11032 , n11014 , n11015 );
xor ( n11033 , n11031 , n11032 );
and ( n11034 , n11033 , n11007 );
or ( n11035 , n11030 , n11034 );
buf ( n11036 , n11035 );
not ( n11037 , n11036 );
buf ( n11038 , n11037 );
buf ( n11039 , n11038 );
not ( n11040 , n11039 );
or ( n11041 , n11024 , n11040 );
not ( n11042 , n11007 );
xor ( n11043 , n10924 , n10927 );
xor ( n11044 , n11043 , n10952 );
buf ( n11045 , n11044 );
buf ( n11046 , n11045 );
and ( n11047 , n11042 , n11046 );
not ( n11048 , n11046 );
and ( n11049 , n11031 , n11032 );
xor ( n11050 , n11048 , n11049 );
and ( n11051 , n11050 , n11007 );
or ( n11052 , n11047 , n11051 );
buf ( n11053 , n11052 );
not ( n11054 , n11053 );
buf ( n11055 , n11054 );
buf ( n11056 , n11055 );
not ( n11057 , n11056 );
or ( n11058 , n11041 , n11057 );
not ( n11059 , n11007 );
xor ( n11060 , n10916 , n10919 );
xor ( n11061 , n11060 , n10955 );
buf ( n11062 , n11061 );
buf ( n11063 , n11062 );
and ( n11064 , n11059 , n11063 );
not ( n11065 , n11063 );
and ( n11066 , n11048 , n11049 );
xor ( n11067 , n11065 , n11066 );
and ( n11068 , n11067 , n11007 );
or ( n11069 , n11064 , n11068 );
buf ( n11070 , n11069 );
not ( n11071 , n11070 );
buf ( n11072 , n11071 );
buf ( n11073 , n11072 );
not ( n11074 , n11073 );
or ( n11075 , n11058 , n11074 );
not ( n11076 , n11007 );
xor ( n11077 , n10908 , n10911 );
xor ( n11078 , n11077 , n10958 );
buf ( n11079 , n11078 );
buf ( n11080 , n11079 );
and ( n11081 , n11076 , n11080 );
not ( n11082 , n11080 );
and ( n11083 , n11065 , n11066 );
xor ( n11084 , n11082 , n11083 );
and ( n11085 , n11084 , n11007 );
or ( n11086 , n11081 , n11085 );
buf ( n11087 , n11086 );
not ( n11088 , n11087 );
buf ( n11089 , n11088 );
buf ( n11090 , n11089 );
not ( n11091 , n11090 );
or ( n11092 , n11075 , n11091 );
not ( n11093 , n11007 );
xor ( n11094 , n10900 , n10903 );
xor ( n11095 , n11094 , n10961 );
buf ( n11096 , n11095 );
buf ( n11097 , n11096 );
and ( n11098 , n11093 , n11097 );
not ( n11099 , n11097 );
and ( n11100 , n11082 , n11083 );
xor ( n11101 , n11099 , n11100 );
and ( n11102 , n11101 , n11007 );
or ( n11103 , n11098 , n11102 );
buf ( n11104 , n11103 );
not ( n11105 , n11104 );
buf ( n11106 , n11105 );
buf ( n11107 , n11106 );
not ( n11108 , n11107 );
or ( n11109 , n11092 , n11108 );
not ( n11110 , n11007 );
xor ( n11111 , n10892 , n10895 );
xor ( n11112 , n11111 , n10964 );
buf ( n11113 , n11112 );
buf ( n11114 , n11113 );
and ( n11115 , n11110 , n11114 );
not ( n11116 , n11114 );
and ( n11117 , n11099 , n11100 );
xor ( n11118 , n11116 , n11117 );
and ( n11119 , n11118 , n11007 );
or ( n11120 , n11115 , n11119 );
buf ( n11121 , n11120 );
not ( n11122 , n11121 );
buf ( n11123 , n11122 );
buf ( n11124 , n11123 );
not ( n11125 , n11124 );
or ( n11126 , n11109 , n11125 );
not ( n11127 , n11007 );
xor ( n11128 , n10884 , n10887 );
xor ( n11129 , n11128 , n10967 );
buf ( n11130 , n11129 );
buf ( n11131 , n11130 );
and ( n11132 , n11127 , n11131 );
not ( n11133 , n11131 );
and ( n11134 , n11116 , n11117 );
xor ( n11135 , n11133 , n11134 );
and ( n11136 , n11135 , n11007 );
or ( n11137 , n11132 , n11136 );
buf ( n11138 , n11137 );
not ( n11139 , n11138 );
buf ( n11140 , n11139 );
buf ( n11141 , n11140 );
not ( n11142 , n11141 );
or ( n11143 , n11126 , n11142 );
not ( n11144 , n11007 );
xor ( n11145 , n10876 , n10879 );
xor ( n11146 , n11145 , n10970 );
buf ( n11147 , n11146 );
buf ( n11148 , n11147 );
and ( n11149 , n11144 , n11148 );
not ( n11150 , n11148 );
and ( n11151 , n11133 , n11134 );
xor ( n11152 , n11150 , n11151 );
and ( n11153 , n11152 , n11007 );
or ( n11154 , n11149 , n11153 );
buf ( n11155 , n11154 );
not ( n11156 , n11155 );
buf ( n11157 , n11156 );
buf ( n11158 , n11157 );
not ( n11159 , n11158 );
or ( n11160 , n11143 , n11159 );
not ( n11161 , n11007 );
xor ( n11162 , n10868 , n10871 );
xor ( n11163 , n11162 , n10973 );
buf ( n11164 , n11163 );
buf ( n11165 , n11164 );
and ( n11166 , n11161 , n11165 );
not ( n11167 , n11165 );
and ( n11168 , n11150 , n11151 );
xor ( n11169 , n11167 , n11168 );
and ( n11170 , n11169 , n11007 );
or ( n11171 , n11166 , n11170 );
buf ( n11172 , n11171 );
not ( n11173 , n11172 );
buf ( n11174 , n11173 );
buf ( n11175 , n11174 );
not ( n11176 , n11175 );
or ( n11177 , n11160 , n11176 );
not ( n11178 , n11007 );
xor ( n11179 , n10860 , n10863 );
xor ( n11180 , n11179 , n10976 );
buf ( n11181 , n11180 );
buf ( n11182 , n11181 );
and ( n11183 , n11178 , n11182 );
not ( n11184 , n11182 );
and ( n11185 , n11167 , n11168 );
xor ( n11186 , n11184 , n11185 );
and ( n11187 , n11186 , n11007 );
or ( n11188 , n11183 , n11187 );
buf ( n11189 , n11188 );
not ( n11190 , n11189 );
buf ( n11191 , n11190 );
buf ( n11192 , n11191 );
not ( n11193 , n11192 );
or ( n11194 , n11177 , n11193 );
not ( n11195 , n11007 );
xor ( n11196 , n10852 , n10855 );
xor ( n11197 , n11196 , n10979 );
buf ( n11198 , n11197 );
buf ( n11199 , n11198 );
and ( n11200 , n11195 , n11199 );
not ( n11201 , n11199 );
and ( n11202 , n11184 , n11185 );
xor ( n11203 , n11201 , n11202 );
and ( n11204 , n11203 , n11007 );
or ( n11205 , n11200 , n11204 );
buf ( n11206 , n11205 );
not ( n11207 , n11206 );
buf ( n11208 , n11207 );
buf ( n11209 , n11208 );
not ( n11210 , n11209 );
or ( n11211 , n11194 , n11210 );
not ( n11212 , n11007 );
xor ( n11213 , n10844 , n10847 );
xor ( n11214 , n11213 , n10982 );
buf ( n11215 , n11214 );
buf ( n11216 , n11215 );
and ( n11217 , n11212 , n11216 );
not ( n11218 , n11216 );
and ( n11219 , n11201 , n11202 );
xor ( n11220 , n11218 , n11219 );
and ( n11221 , n11220 , n11007 );
or ( n11222 , n11217 , n11221 );
buf ( n11223 , n11222 );
not ( n11224 , n11223 );
buf ( n11225 , n11224 );
buf ( n11226 , n11225 );
not ( n11227 , n11226 );
or ( n11228 , n11211 , n11227 );
not ( n11229 , n11007 );
xor ( n11230 , n10836 , n10839 );
xor ( n11231 , n11230 , n10985 );
buf ( n11232 , n11231 );
buf ( n11233 , n11232 );
and ( n11234 , n11229 , n11233 );
not ( n11235 , n11233 );
and ( n11236 , n11218 , n11219 );
xor ( n11237 , n11235 , n11236 );
and ( n11238 , n11237 , n11007 );
or ( n11239 , n11234 , n11238 );
buf ( n11240 , n11239 );
not ( n11241 , n11240 );
buf ( n11242 , n11241 );
buf ( n11243 , n11242 );
not ( n11244 , n11243 );
or ( n11245 , n11228 , n11244 );
not ( n11246 , n11007 );
xor ( n11247 , n10828 , n10831 );
xor ( n11248 , n11247 , n10988 );
buf ( n11249 , n11248 );
buf ( n11250 , n11249 );
and ( n11251 , n11246 , n11250 );
not ( n11252 , n11250 );
and ( n11253 , n11235 , n11236 );
xor ( n11254 , n11252 , n11253 );
and ( n11255 , n11254 , n11007 );
or ( n11256 , n11251 , n11255 );
buf ( n11257 , n11256 );
not ( n11258 , n11257 );
buf ( n11259 , n11258 );
buf ( n11260 , n11259 );
not ( n11261 , n11260 );
or ( n11262 , n11245 , n11261 );
not ( n11263 , n11007 );
xor ( n11264 , n10820 , n10823 );
xor ( n11265 , n11264 , n10991 );
buf ( n11266 , n11265 );
buf ( n11267 , n11266 );
and ( n11268 , n11263 , n11267 );
not ( n11269 , n11267 );
and ( n11270 , n11252 , n11253 );
xor ( n11271 , n11269 , n11270 );
and ( n11272 , n11271 , n11007 );
or ( n11273 , n11268 , n11272 );
buf ( n11274 , n11273 );
not ( n11275 , n11274 );
buf ( n11276 , n11275 );
buf ( n11277 , n11276 );
not ( n11278 , n11277 );
or ( n11279 , n11262 , n11278 );
not ( n11280 , n11007 );
xor ( n11281 , n10812 , n10815 );
xor ( n11282 , n11281 , n10994 );
buf ( n11283 , n11282 );
buf ( n11284 , n11283 );
and ( n11285 , n11280 , n11284 );
not ( n11286 , n11284 );
and ( n11287 , n11269 , n11270 );
xor ( n11288 , n11286 , n11287 );
and ( n11289 , n11288 , n11007 );
or ( n11290 , n11285 , n11289 );
buf ( n11291 , n11290 );
not ( n11292 , n11291 );
buf ( n11293 , n11292 );
buf ( n11294 , n11293 );
not ( n11295 , n11294 );
or ( n11296 , n11279 , n11295 );
not ( n11297 , n11007 );
xor ( n11298 , n10804 , n10807 );
xor ( n11299 , n11298 , n10997 );
buf ( n11300 , n11299 );
buf ( n11301 , n11300 );
and ( n11302 , n11297 , n11301 );
not ( n11303 , n11301 );
and ( n11304 , n11286 , n11287 );
xor ( n11305 , n11303 , n11304 );
and ( n11306 , n11305 , n11007 );
or ( n11307 , n11302 , n11306 );
buf ( n11308 , n11307 );
not ( n11309 , n11308 );
buf ( n11310 , n11309 );
buf ( n11311 , n11310 );
not ( n11312 , n11311 );
or ( n11313 , n11296 , n11312 );
not ( n11314 , n11007 );
xor ( n11315 , n10796 , n10799 );
xor ( n11316 , n11315 , n11000 );
buf ( n11317 , n11316 );
buf ( n11318 , n11317 );
and ( n11319 , n11314 , n11318 );
not ( n11320 , n11318 );
and ( n11321 , n11303 , n11304 );
xor ( n11322 , n11320 , n11321 );
and ( n11323 , n11322 , n11007 );
or ( n11324 , n11319 , n11323 );
buf ( n11325 , n11324 );
not ( n11326 , n11325 );
buf ( n11327 , n11326 );
buf ( n11328 , n11327 );
not ( n11329 , n11328 );
or ( n11330 , n11313 , n11329 );
buf ( n11331 , n11330 );
buf ( n11332 , n11331 );
and ( n11333 , n11332 , n11007 );
not ( n11334 , n11333 );
and ( n11335 , n11334 , n11261 );
xor ( n11336 , n11261 , n11007 );
xor ( n11337 , n11244 , n11007 );
xor ( n11338 , n11227 , n11007 );
xor ( n11339 , n11210 , n11007 );
xor ( n11340 , n11193 , n11007 );
xor ( n11341 , n11176 , n11007 );
xor ( n11342 , n11159 , n11007 );
xor ( n11343 , n11142 , n11007 );
xor ( n11344 , n11125 , n11007 );
xor ( n11345 , n11108 , n11007 );
xor ( n11346 , n11091 , n11007 );
xor ( n11347 , n11074 , n11007 );
xor ( n11348 , n11057 , n11007 );
xor ( n11349 , n11040 , n11007 );
xor ( n11350 , n11023 , n11007 );
xor ( n11351 , n10637 , n11007 );
and ( n11352 , n11351 , n11007 );
and ( n11353 , n11350 , n11352 );
and ( n11354 , n11349 , n11353 );
and ( n11355 , n11348 , n11354 );
and ( n11356 , n11347 , n11355 );
and ( n11357 , n11346 , n11356 );
and ( n11358 , n11345 , n11357 );
and ( n11359 , n11344 , n11358 );
and ( n11360 , n11343 , n11359 );
and ( n11361 , n11342 , n11360 );
and ( n11362 , n11341 , n11361 );
and ( n11363 , n11340 , n11362 );
and ( n11364 , n11339 , n11363 );
and ( n11365 , n11338 , n11364 );
and ( n11366 , n11337 , n11365 );
xor ( n11367 , n11336 , n11366 );
and ( n11368 , n11367 , n11333 );
or ( n11369 , n11335 , n11368 );
buf ( n11370 , n11369 );
buf ( n11371 , n11370 );
buf ( n11372 , n10613 );
buf ( n11373 , n10613 );
buf ( n11374 , RI2107a660_489);
buf ( n11375 , n11374 );
not ( n11376 , n11375 );
buf ( n11377 , RI2107a6d8_488);
buf ( n11378 , n11377 );
not ( n11379 , n11378 );
buf ( n11380 , RI2107b218_486);
buf ( n11381 , n11380 );
not ( n11382 , n11381 );
buf ( n11383 , RI2107b290_485);
buf ( n11384 , n11383 );
not ( n11385 , n11384 );
buf ( n11386 , RI2107b308_484);
buf ( n11387 , n11386 );
not ( n11388 , n11387 );
buf ( n11389 , RI2107b380_483);
buf ( n11390 , n11389 );
not ( n11391 , n11390 );
buf ( n11392 , RI2107b3f8_482);
buf ( n11393 , n11392 );
not ( n11394 , n11393 );
buf ( n11395 , RI2107bec0_481);
buf ( n11396 , n11395 );
not ( n11397 , n11396 );
buf ( n11398 , RI2107bf38_480);
buf ( n11399 , n11398 );
not ( n11400 , n11399 );
buf ( n11401 , RI2107bfb0_479);
buf ( n11402 , n11401 );
not ( n11403 , n11402 );
buf ( n11404 , RI2107c028_478);
buf ( n11405 , n11404 );
not ( n11406 , n11405 );
buf ( n11407 , RI2107c0a0_477);
buf ( n11408 , n11407 );
not ( n11409 , n11408 );
buf ( n11410 , RI2107cbe0_475);
buf ( n11411 , n11410 );
not ( n11412 , n11411 );
buf ( n11413 , RI2107cc58_474);
buf ( n11414 , n11413 );
not ( n11415 , n11414 );
buf ( n11416 , RI2107ccd0_473);
buf ( n11417 , n11416 );
not ( n11418 , n11417 );
buf ( n11419 , RI2107cd48_472);
buf ( n11420 , n11419 );
not ( n11421 , n11420 );
buf ( n11422 , RI2107cdc0_471);
buf ( n11423 , n11422 );
not ( n11424 , n11423 );
buf ( n11425 , RI2107ce38_470);
buf ( n11426 , n11425 );
not ( n11427 , n11426 );
buf ( n11428 , RI2107d900_469);
buf ( n11429 , n11428 );
not ( n11430 , n11429 );
buf ( n11431 , RI2107d978_468);
buf ( n11432 , n11431 );
not ( n11433 , n11432 );
buf ( n11434 , RI2107d9f0_467);
buf ( n11435 , n11434 );
not ( n11436 , n11435 );
buf ( n11437 , RI2107da68_466);
buf ( n11438 , n11437 );
not ( n11439 , n11438 );
buf ( n11440 , RI210798c8_496);
buf ( n11441 , n11440 );
not ( n11442 , n11441 );
buf ( n11443 , RI21079940_495);
buf ( n11444 , n11443 );
not ( n11445 , n11444 );
buf ( n11446 , RI210799b8_494);
buf ( n11447 , n11446 );
not ( n11448 , n11447 );
buf ( n11449 , RI2107a480_493);
buf ( n11450 , n11449 );
not ( n11451 , n11450 );
buf ( n11452 , RI2107a4f8_492);
buf ( n11453 , n11452 );
not ( n11454 , n11453 );
buf ( n11455 , RI2107a570_491);
buf ( n11456 , n11455 );
not ( n11457 , n11456 );
buf ( n11458 , RI2107a5e8_490);
buf ( n11459 , n11458 );
not ( n11460 , n11459 );
buf ( n11461 , RI2107b1a0_487);
buf ( n11462 , n11461 );
not ( n11463 , n11462 );
buf ( n11464 , RI2107c118_476);
buf ( n11465 , n11464 );
not ( n11466 , n11465 );
buf ( n11467 , RI2106bde0_608);
buf ( n11468 , n11467 );
not ( n11469 , n11468 );
and ( n11470 , n11466 , n11469 );
and ( n11471 , n11463 , n11470 );
and ( n11472 , n11460 , n11471 );
and ( n11473 , n11457 , n11472 );
and ( n11474 , n11454 , n11473 );
and ( n11475 , n11451 , n11474 );
and ( n11476 , n11448 , n11475 );
and ( n11477 , n11445 , n11476 );
and ( n11478 , n11442 , n11477 );
and ( n11479 , n11439 , n11478 );
and ( n11480 , n11436 , n11479 );
and ( n11481 , n11433 , n11480 );
and ( n11482 , n11430 , n11481 );
and ( n11483 , n11427 , n11482 );
and ( n11484 , n11424 , n11483 );
and ( n11485 , n11421 , n11484 );
and ( n11486 , n11418 , n11485 );
and ( n11487 , n11415 , n11486 );
and ( n11488 , n11412 , n11487 );
and ( n11489 , n11409 , n11488 );
and ( n11490 , n11406 , n11489 );
and ( n11491 , n11403 , n11490 );
and ( n11492 , n11400 , n11491 );
and ( n11493 , n11397 , n11492 );
and ( n11494 , n11394 , n11493 );
and ( n11495 , n11391 , n11494 );
and ( n11496 , n11388 , n11495 );
and ( n11497 , n11385 , n11496 );
and ( n11498 , n11382 , n11497 );
and ( n11499 , n11379 , n11498 );
xor ( n11500 , n11376 , n11499 );
buf ( n11501 , n11500 );
buf ( n11502 , n11374 );
and ( n11503 , n11501 , n11502 );
or ( n11504 , C0 , n11503 );
buf ( n11505 , n11504 );
not ( n11506 , n11505 );
not ( n11507 , n11502 );
and ( n11508 , n11507 , n11398 );
xor ( n11509 , n11400 , n11491 );
buf ( n11510 , n11509 );
and ( n11511 , n11510 , n11502 );
or ( n11512 , n11508 , n11511 );
buf ( n11513 , n11512 );
and ( n11514 , n11506 , n11513 );
not ( n11515 , n11513 );
not ( n11516 , n11502 );
and ( n11517 , n11516 , n11401 );
xor ( n11518 , n11403 , n11490 );
buf ( n11519 , n11518 );
and ( n11520 , n11519 , n11502 );
or ( n11521 , n11517 , n11520 );
buf ( n11522 , n11521 );
not ( n11523 , n11522 );
not ( n11524 , n11502 );
and ( n11525 , n11524 , n11404 );
xor ( n11526 , n11406 , n11489 );
buf ( n11527 , n11526 );
and ( n11528 , n11527 , n11502 );
or ( n11529 , n11525 , n11528 );
buf ( n11530 , n11529 );
not ( n11531 , n11530 );
not ( n11532 , n11502 );
and ( n11533 , n11532 , n11407 );
xor ( n11534 , n11409 , n11488 );
buf ( n11535 , n11534 );
and ( n11536 , n11535 , n11502 );
or ( n11537 , n11533 , n11536 );
buf ( n11538 , n11537 );
not ( n11539 , n11538 );
not ( n11540 , n11502 );
and ( n11541 , n11540 , n11410 );
xor ( n11542 , n11412 , n11487 );
buf ( n11543 , n11542 );
and ( n11544 , n11543 , n11502 );
or ( n11545 , n11541 , n11544 );
buf ( n11546 , n11545 );
not ( n11547 , n11546 );
not ( n11548 , n11502 );
and ( n11549 , n11548 , n11413 );
xor ( n11550 , n11415 , n11486 );
buf ( n11551 , n11550 );
and ( n11552 , n11551 , n11502 );
or ( n11553 , n11549 , n11552 );
buf ( n11554 , n11553 );
not ( n11555 , n11554 );
not ( n11556 , n11502 );
and ( n11557 , n11556 , n11416 );
xor ( n11558 , n11418 , n11485 );
buf ( n11559 , n11558 );
and ( n11560 , n11559 , n11502 );
or ( n11561 , n11557 , n11560 );
buf ( n11562 , n11561 );
not ( n11563 , n11562 );
not ( n11564 , n11502 );
and ( n11565 , n11564 , n11419 );
xor ( n11566 , n11421 , n11484 );
buf ( n11567 , n11566 );
and ( n11568 , n11567 , n11502 );
or ( n11569 , n11565 , n11568 );
buf ( n11570 , n11569 );
not ( n11571 , n11570 );
not ( n11572 , n11502 );
and ( n11573 , n11572 , n11422 );
xor ( n11574 , n11424 , n11483 );
buf ( n11575 , n11574 );
and ( n11576 , n11575 , n11502 );
or ( n11577 , n11573 , n11576 );
buf ( n11578 , n11577 );
not ( n11579 , n11578 );
not ( n11580 , n11502 );
and ( n11581 , n11580 , n11425 );
xor ( n11582 , n11427 , n11482 );
buf ( n11583 , n11582 );
and ( n11584 , n11583 , n11502 );
or ( n11585 , n11581 , n11584 );
buf ( n11586 , n11585 );
not ( n11587 , n11586 );
not ( n11588 , n11502 );
and ( n11589 , n11588 , n11428 );
xor ( n11590 , n11430 , n11481 );
buf ( n11591 , n11590 );
and ( n11592 , n11591 , n11502 );
or ( n11593 , n11589 , n11592 );
buf ( n11594 , n11593 );
not ( n11595 , n11594 );
not ( n11596 , n11502 );
and ( n11597 , n11596 , n11431 );
xor ( n11598 , n11433 , n11480 );
buf ( n11599 , n11598 );
and ( n11600 , n11599 , n11502 );
or ( n11601 , n11597 , n11600 );
buf ( n11602 , n11601 );
not ( n11603 , n11602 );
not ( n11604 , n11502 );
and ( n11605 , n11604 , n11434 );
xor ( n11606 , n11436 , n11479 );
buf ( n11607 , n11606 );
and ( n11608 , n11607 , n11502 );
or ( n11609 , n11605 , n11608 );
buf ( n11610 , n11609 );
not ( n11611 , n11610 );
not ( n11612 , n11502 );
and ( n11613 , n11612 , n11437 );
xor ( n11614 , n11439 , n11478 );
buf ( n11615 , n11614 );
and ( n11616 , n11615 , n11502 );
or ( n11617 , n11613 , n11616 );
buf ( n11618 , n11617 );
not ( n11619 , n11618 );
not ( n11620 , n11502 );
and ( n11621 , n11620 , n11440 );
xor ( n11622 , n11442 , n11477 );
buf ( n11623 , n11622 );
and ( n11624 , n11623 , n11502 );
or ( n11625 , n11621 , n11624 );
buf ( n11626 , n11625 );
not ( n11627 , n11626 );
not ( n11628 , n11502 );
and ( n11629 , n11628 , n11443 );
xor ( n11630 , n11445 , n11476 );
buf ( n11631 , n11630 );
and ( n11632 , n11631 , n11502 );
or ( n11633 , n11629 , n11632 );
buf ( n11634 , n11633 );
not ( n11635 , n11634 );
not ( n11636 , n11502 );
and ( n11637 , n11636 , n11446 );
xor ( n11638 , n11448 , n11475 );
buf ( n11639 , n11638 );
and ( n11640 , n11639 , n11502 );
or ( n11641 , n11637 , n11640 );
buf ( n11642 , n11641 );
not ( n11643 , n11642 );
not ( n11644 , n11502 );
and ( n11645 , n11644 , n11449 );
xor ( n11646 , n11451 , n11474 );
buf ( n11647 , n11646 );
and ( n11648 , n11647 , n11502 );
or ( n11649 , n11645 , n11648 );
buf ( n11650 , n11649 );
not ( n11651 , n11650 );
not ( n11652 , n11502 );
and ( n11653 , n11652 , n11452 );
xor ( n11654 , n11454 , n11473 );
buf ( n11655 , n11654 );
and ( n11656 , n11655 , n11502 );
or ( n11657 , n11653 , n11656 );
buf ( n11658 , n11657 );
not ( n11659 , n11658 );
not ( n11660 , n11502 );
and ( n11661 , n11660 , n11455 );
xor ( n11662 , n11457 , n11472 );
buf ( n11663 , n11662 );
and ( n11664 , n11663 , n11502 );
or ( n11665 , n11661 , n11664 );
buf ( n11666 , n11665 );
not ( n11667 , n11666 );
not ( n11668 , n11502 );
and ( n11669 , n11668 , n11458 );
xor ( n11670 , n11460 , n11471 );
buf ( n11671 , n11670 );
and ( n11672 , n11671 , n11502 );
or ( n11673 , n11669 , n11672 );
buf ( n11674 , n11673 );
not ( n11675 , n11674 );
not ( n11676 , n11502 );
and ( n11677 , n11676 , n11461 );
xor ( n11678 , n11463 , n11470 );
buf ( n11679 , n11678 );
and ( n11680 , n11679 , n11502 );
or ( n11681 , n11677 , n11680 );
buf ( n11682 , n11681 );
not ( n11683 , n11682 );
not ( n11684 , n11502 );
and ( n11685 , n11684 , n11464 );
xor ( n11686 , n11466 , n11469 );
buf ( n11687 , n11686 );
and ( n11688 , n11687 , n11502 );
or ( n11689 , n11685 , n11688 );
buf ( n11690 , n11689 );
not ( n11691 , n11690 );
buf ( n11692 , n11467 );
buf ( n11693 , n11692 );
not ( n11694 , n11693 );
and ( n11695 , n11691 , n11694 );
and ( n11696 , n11683 , n11695 );
and ( n11697 , n11675 , n11696 );
and ( n11698 , n11667 , n11697 );
and ( n11699 , n11659 , n11698 );
and ( n11700 , n11651 , n11699 );
and ( n11701 , n11643 , n11700 );
and ( n11702 , n11635 , n11701 );
and ( n11703 , n11627 , n11702 );
and ( n11704 , n11619 , n11703 );
and ( n11705 , n11611 , n11704 );
and ( n11706 , n11603 , n11705 );
and ( n11707 , n11595 , n11706 );
and ( n11708 , n11587 , n11707 );
and ( n11709 , n11579 , n11708 );
and ( n11710 , n11571 , n11709 );
and ( n11711 , n11563 , n11710 );
and ( n11712 , n11555 , n11711 );
and ( n11713 , n11547 , n11712 );
and ( n11714 , n11539 , n11713 );
and ( n11715 , n11531 , n11714 );
and ( n11716 , n11523 , n11715 );
xor ( n11717 , n11515 , n11716 );
and ( n11718 , n11717 , n11505 );
or ( n11719 , n11514 , n11718 );
buf ( n11720 , n11719 );
not ( n11721 , n11720 );
buf ( n11722 , n11721 );
buf ( n11723 , n11722 );
not ( n11724 , n11723 );
buf ( n11725 , n11724 );
buf ( n11726 , n11725 );
not ( n11727 , n11726 );
buf ( n11728 , n11727 );
buf ( n11729 , n11728 );
not ( n11730 , n11729 );
or ( n11731 , n11730 , C0 );
or ( n11732 , n11731 , C0 );
or ( n11733 , n11732 , C0 );
or ( n11734 , n11733 , C0 );
or ( n11735 , n11734 , C0 );
or ( n11736 , n11735 , C0 );
or ( n11737 , n11736 , C0 );
or ( n11738 , n11737 , C0 );
or ( n11739 , n11738 , C0 );
or ( n11740 , n11739 , C0 );
or ( n11741 , n11740 , C0 );
or ( n11742 , n11741 , C0 );
or ( n11743 , n11742 , C0 );
or ( n11744 , n11743 , C0 );
or ( n11745 , n11744 , C0 );
or ( n11746 , n11745 , C0 );
or ( n11747 , n11746 , C0 );
or ( n11748 , n11747 , C0 );
or ( n11749 , n11748 , C0 );
or ( n11750 , n11749 , C0 );
or ( n11751 , n11750 , C0 );
or ( n11752 , n11751 , C0 );
or ( n11753 , n11752 , C0 );
or ( n11754 , n11753 , C0 );
or ( n11755 , n11754 , C0 );
or ( n11756 , n11755 , C0 );
or ( n11757 , n11756 , C0 );
or ( n11758 , n11757 , C0 );
or ( n11759 , n11758 , C0 );
or ( n11760 , n11759 , C0 );
buf ( n11761 , n11760 );
not ( n11762 , n11505 );
not ( n11763 , n11502 );
and ( n11764 , n11763 , n11377 );
xor ( n11765 , n11379 , n11498 );
buf ( n11766 , n11765 );
and ( n11767 , n11766 , n11502 );
or ( n11768 , n11764 , n11767 );
buf ( n11769 , n11768 );
not ( n11770 , n11769 );
not ( n11771 , n11502 );
and ( n11772 , n11771 , n11380 );
xor ( n11773 , n11382 , n11497 );
buf ( n11774 , n11773 );
and ( n11775 , n11774 , n11502 );
or ( n11776 , n11772 , n11775 );
buf ( n11777 , n11776 );
not ( n11778 , n11777 );
not ( n11779 , n11502 );
and ( n11780 , n11779 , n11383 );
xor ( n11781 , n11385 , n11496 );
buf ( n11782 , n11781 );
and ( n11783 , n11782 , n11502 );
or ( n11784 , n11780 , n11783 );
buf ( n11785 , n11784 );
not ( n11786 , n11785 );
not ( n11787 , n11502 );
and ( n11788 , n11787 , n11386 );
xor ( n11789 , n11388 , n11495 );
buf ( n11790 , n11789 );
and ( n11791 , n11790 , n11502 );
or ( n11792 , n11788 , n11791 );
buf ( n11793 , n11792 );
not ( n11794 , n11793 );
not ( n11795 , n11502 );
and ( n11796 , n11795 , n11389 );
xor ( n11797 , n11391 , n11494 );
buf ( n11798 , n11797 );
and ( n11799 , n11798 , n11502 );
or ( n11800 , n11796 , n11799 );
buf ( n11801 , n11800 );
not ( n11802 , n11801 );
not ( n11803 , n11502 );
and ( n11804 , n11803 , n11392 );
xor ( n11805 , n11394 , n11493 );
buf ( n11806 , n11805 );
and ( n11807 , n11806 , n11502 );
or ( n11808 , n11804 , n11807 );
buf ( n11809 , n11808 );
not ( n11810 , n11809 );
not ( n11811 , n11502 );
and ( n11812 , n11811 , n11395 );
xor ( n11813 , n11397 , n11492 );
buf ( n11814 , n11813 );
and ( n11815 , n11814 , n11502 );
or ( n11816 , n11812 , n11815 );
buf ( n11817 , n11816 );
not ( n11818 , n11817 );
and ( n11819 , n11515 , n11716 );
and ( n11820 , n11818 , n11819 );
and ( n11821 , n11810 , n11820 );
and ( n11822 , n11802 , n11821 );
and ( n11823 , n11794 , n11822 );
and ( n11824 , n11786 , n11823 );
and ( n11825 , n11778 , n11824 );
and ( n11826 , n11770 , n11825 );
xor ( n11827 , n11762 , n11826 );
buf ( n11828 , n11505 );
and ( n11829 , n11827 , n11828 );
or ( n11830 , C0 , n11829 );
buf ( n11831 , n11830 );
not ( n11832 , n11831 );
buf ( n11833 , n11832 );
buf ( n11834 , n11833 );
not ( n11835 , n11834 );
buf ( n11836 , n11835 );
not ( n11837 , n11836 );
buf ( n11838 , n11837 );
not ( n11839 , n11505 );
and ( n11840 , n11839 , n11769 );
xor ( n11841 , n11770 , n11825 );
and ( n11842 , n11841 , n11505 );
or ( n11843 , n11840 , n11842 );
buf ( n11844 , n11843 );
not ( n11845 , n11844 );
buf ( n11846 , n11845 );
buf ( n11847 , n11846 );
not ( n11848 , n11847 );
buf ( n11849 , n11848 );
not ( n11850 , n11849 );
buf ( n11851 , n11850 );
not ( n11852 , n11505 );
and ( n11853 , n11852 , n11777 );
xor ( n11854 , n11778 , n11824 );
and ( n11855 , n11854 , n11505 );
or ( n11856 , n11853 , n11855 );
buf ( n11857 , n11856 );
not ( n11858 , n11857 );
buf ( n11859 , n11858 );
buf ( n11860 , n11859 );
not ( n11861 , n11860 );
buf ( n11862 , n11861 );
not ( n11863 , n11862 );
buf ( n11864 , n11863 );
not ( n11865 , n11505 );
and ( n11866 , n11865 , n11785 );
xor ( n11867 , n11786 , n11823 );
and ( n11868 , n11867 , n11505 );
or ( n11869 , n11866 , n11868 );
buf ( n11870 , n11869 );
not ( n11871 , n11870 );
buf ( n11872 , n11871 );
buf ( n11873 , n11872 );
not ( n11874 , n11873 );
buf ( n11875 , n11874 );
not ( n11876 , n11875 );
buf ( n11877 , n11876 );
not ( n11878 , n11505 );
and ( n11879 , n11878 , n11793 );
xor ( n11880 , n11794 , n11822 );
and ( n11881 , n11880 , n11505 );
or ( n11882 , n11879 , n11881 );
buf ( n11883 , n11882 );
not ( n11884 , n11883 );
buf ( n11885 , n11884 );
buf ( n11886 , n11885 );
not ( n11887 , n11886 );
buf ( n11888 , n11887 );
not ( n11889 , n11888 );
buf ( n11890 , n11889 );
not ( n11891 , n11505 );
and ( n11892 , n11891 , n11801 );
xor ( n11893 , n11802 , n11821 );
and ( n11894 , n11893 , n11505 );
or ( n11895 , n11892 , n11894 );
buf ( n11896 , n11895 );
not ( n11897 , n11896 );
buf ( n11898 , n11897 );
buf ( n11899 , n11898 );
not ( n11900 , n11899 );
buf ( n11901 , n11900 );
not ( n11902 , n11901 );
buf ( n11903 , n11902 );
not ( n11904 , n11505 );
and ( n11905 , n11904 , n11809 );
xor ( n11906 , n11810 , n11820 );
and ( n11907 , n11906 , n11505 );
or ( n11908 , n11905 , n11907 );
buf ( n11909 , n11908 );
not ( n11910 , n11909 );
buf ( n11911 , n11910 );
buf ( n11912 , n11911 );
not ( n11913 , n11912 );
buf ( n11914 , n11913 );
not ( n11915 , n11914 );
buf ( n11916 , n11915 );
not ( n11917 , n11505 );
and ( n11918 , n11917 , n11817 );
xor ( n11919 , n11818 , n11819 );
and ( n11920 , n11919 , n11505 );
or ( n11921 , n11918 , n11920 );
buf ( n11922 , n11921 );
not ( n11923 , n11922 );
buf ( n11924 , n11923 );
buf ( n11925 , n11924 );
not ( n11926 , n11925 );
buf ( n11927 , n11926 );
not ( n11928 , n11927 );
buf ( n11929 , n11928 );
not ( n11930 , n11725 );
buf ( n11931 , n11930 );
and ( n11932 , n11929 , n11931 );
and ( n11933 , n11916 , n11932 );
and ( n11934 , n11903 , n11933 );
and ( n11935 , n11890 , n11934 );
and ( n11936 , n11877 , n11935 );
and ( n11937 , n11864 , n11936 );
and ( n11938 , n11851 , n11937 );
and ( n11939 , n11838 , n11938 );
not ( n11940 , n11939 );
buf ( n11941 , n11940 );
buf ( n11942 , n11505 );
and ( n11943 , n11941 , n11942 );
or ( n11944 , C0 , n11943 );
buf ( n11945 , n11944 );
buf ( n11946 , n11945 );
and ( n11947 , n11761 , n11946 );
not ( n11948 , n11947 );
and ( n11949 , n11948 , n11730 );
xor ( n11950 , n11730 , n11946 );
xor ( n11951 , n11950 , n11946 );
and ( n11952 , n11951 , n11947 );
or ( n11953 , n11949 , n11952 );
buf ( n11954 , n11953 );
not ( n11955 , n11954 );
buf ( n11956 , n11504 );
not ( n11957 , n11956 );
buf ( n11958 , n11816 );
and ( n11959 , n11957 , n11958 );
not ( n11960 , n11958 );
buf ( n11961 , n11512 );
not ( n11962 , n11961 );
buf ( n11963 , n11521 );
not ( n11964 , n11963 );
buf ( n11965 , n11529 );
not ( n11966 , n11965 );
buf ( n11967 , n11537 );
not ( n11968 , n11967 );
buf ( n11969 , n11545 );
not ( n11970 , n11969 );
buf ( n11971 , n11553 );
not ( n11972 , n11971 );
buf ( n11973 , n11561 );
not ( n11974 , n11973 );
buf ( n11975 , n11569 );
not ( n11976 , n11975 );
buf ( n11977 , n11577 );
not ( n11978 , n11977 );
buf ( n11979 , n11585 );
not ( n11980 , n11979 );
buf ( n11981 , n11593 );
not ( n11982 , n11981 );
buf ( n11983 , n11601 );
not ( n11984 , n11983 );
buf ( n11985 , n11609 );
not ( n11986 , n11985 );
buf ( n11987 , n11617 );
not ( n11988 , n11987 );
buf ( n11989 , n11625 );
not ( n11990 , n11989 );
buf ( n11991 , n11633 );
not ( n11992 , n11991 );
buf ( n11993 , n11641 );
not ( n11994 , n11993 );
buf ( n11995 , n11649 );
not ( n11996 , n11995 );
buf ( n11997 , n11657 );
not ( n11998 , n11997 );
buf ( n11999 , n11665 );
not ( n12000 , n11999 );
buf ( n12001 , n11673 );
not ( n12002 , n12001 );
buf ( n12003 , n11681 );
not ( n12004 , n12003 );
buf ( n12005 , n11689 );
not ( n12006 , n12005 );
buf ( n12007 , n11692 );
not ( n12008 , n12007 );
and ( n12009 , n12006 , n12008 );
and ( n12010 , n12004 , n12009 );
and ( n12011 , n12002 , n12010 );
and ( n12012 , n12000 , n12011 );
and ( n12013 , n11998 , n12012 );
and ( n12014 , n11996 , n12013 );
and ( n12015 , n11994 , n12014 );
and ( n12016 , n11992 , n12015 );
and ( n12017 , n11990 , n12016 );
and ( n12018 , n11988 , n12017 );
and ( n12019 , n11986 , n12018 );
and ( n12020 , n11984 , n12019 );
and ( n12021 , n11982 , n12020 );
and ( n12022 , n11980 , n12021 );
and ( n12023 , n11978 , n12022 );
and ( n12024 , n11976 , n12023 );
and ( n12025 , n11974 , n12024 );
and ( n12026 , n11972 , n12025 );
and ( n12027 , n11970 , n12026 );
and ( n12028 , n11968 , n12027 );
and ( n12029 , n11966 , n12028 );
and ( n12030 , n11964 , n12029 );
and ( n12031 , n11962 , n12030 );
xor ( n12032 , n11960 , n12031 );
and ( n12033 , n12032 , n11956 );
or ( n12034 , n11959 , n12033 );
buf ( n12035 , n12034 );
not ( n12036 , n12035 );
buf ( n12037 , n12036 );
buf ( n12038 , n12037 );
not ( n12039 , n12038 );
buf ( n12040 , n12039 );
buf ( n12041 , n12040 );
buf ( n12042 , n12041 );
not ( n12043 , n12042 );
buf ( n12044 , n12043 );
buf ( n12045 , n12044 );
not ( n12046 , n12045 );
not ( n12047 , n11956 );
buf ( n12048 , n11768 );
not ( n12049 , n12048 );
buf ( n12050 , n11776 );
not ( n12051 , n12050 );
buf ( n12052 , n11784 );
not ( n12053 , n12052 );
buf ( n12054 , n11792 );
not ( n12055 , n12054 );
buf ( n12056 , n11800 );
not ( n12057 , n12056 );
buf ( n12058 , n11808 );
not ( n12059 , n12058 );
and ( n12060 , n11960 , n12031 );
and ( n12061 , n12059 , n12060 );
and ( n12062 , n12057 , n12061 );
and ( n12063 , n12055 , n12062 );
and ( n12064 , n12053 , n12063 );
and ( n12065 , n12051 , n12064 );
and ( n12066 , n12049 , n12065 );
xor ( n12067 , n12047 , n12066 );
buf ( n12068 , n11956 );
and ( n12069 , n12067 , n12068 );
or ( n12070 , C0 , n12069 );
buf ( n12071 , n12070 );
not ( n12072 , n12071 );
buf ( n12073 , n12072 );
buf ( n12074 , n12073 );
not ( n12075 , n12074 );
buf ( n12076 , n12075 );
not ( n12077 , n12076 );
buf ( n12078 , n12077 );
not ( n12079 , n11956 );
and ( n12080 , n12079 , n12048 );
xor ( n12081 , n12049 , n12065 );
and ( n12082 , n12081 , n11956 );
or ( n12083 , n12080 , n12082 );
buf ( n12084 , n12083 );
not ( n12085 , n12084 );
buf ( n12086 , n12085 );
buf ( n12087 , n12086 );
not ( n12088 , n12087 );
buf ( n12089 , n12088 );
not ( n12090 , n12089 );
buf ( n12091 , n12090 );
not ( n12092 , n11956 );
and ( n12093 , n12092 , n12050 );
xor ( n12094 , n12051 , n12064 );
and ( n12095 , n12094 , n11956 );
or ( n12096 , n12093 , n12095 );
buf ( n12097 , n12096 );
not ( n12098 , n12097 );
buf ( n12099 , n12098 );
buf ( n12100 , n12099 );
not ( n12101 , n12100 );
buf ( n12102 , n12101 );
not ( n12103 , n12102 );
buf ( n12104 , n12103 );
not ( n12105 , n11956 );
and ( n12106 , n12105 , n12052 );
xor ( n12107 , n12053 , n12063 );
and ( n12108 , n12107 , n11956 );
or ( n12109 , n12106 , n12108 );
buf ( n12110 , n12109 );
not ( n12111 , n12110 );
buf ( n12112 , n12111 );
buf ( n12113 , n12112 );
not ( n12114 , n12113 );
buf ( n12115 , n12114 );
not ( n12116 , n12115 );
buf ( n12117 , n12116 );
not ( n12118 , n11956 );
and ( n12119 , n12118 , n12054 );
xor ( n12120 , n12055 , n12062 );
and ( n12121 , n12120 , n11956 );
or ( n12122 , n12119 , n12121 );
buf ( n12123 , n12122 );
not ( n12124 , n12123 );
buf ( n12125 , n12124 );
buf ( n12126 , n12125 );
not ( n12127 , n12126 );
buf ( n12128 , n12127 );
not ( n12129 , n12128 );
buf ( n12130 , n12129 );
not ( n12131 , n11956 );
and ( n12132 , n12131 , n12056 );
xor ( n12133 , n12057 , n12061 );
and ( n12134 , n12133 , n11956 );
or ( n12135 , n12132 , n12134 );
buf ( n12136 , n12135 );
not ( n12137 , n12136 );
buf ( n12138 , n12137 );
buf ( n12139 , n12138 );
not ( n12140 , n12139 );
buf ( n12141 , n12140 );
not ( n12142 , n12141 );
buf ( n12143 , n12142 );
not ( n12144 , n11956 );
and ( n12145 , n12144 , n12058 );
xor ( n12146 , n12059 , n12060 );
and ( n12147 , n12146 , n11956 );
or ( n12148 , n12145 , n12147 );
buf ( n12149 , n12148 );
not ( n12150 , n12149 );
buf ( n12151 , n12150 );
buf ( n12152 , n12151 );
not ( n12153 , n12152 );
buf ( n12154 , n12153 );
not ( n12155 , n12154 );
buf ( n12156 , n12155 );
not ( n12157 , n12040 );
buf ( n12158 , n12157 );
and ( n12159 , n12156 , n12158 );
and ( n12160 , n12143 , n12159 );
and ( n12161 , n12130 , n12160 );
and ( n12162 , n12117 , n12161 );
and ( n12163 , n12104 , n12162 );
and ( n12164 , n12091 , n12163 );
and ( n12165 , n12078 , n12164 );
not ( n12166 , n12165 );
buf ( n12167 , n12166 );
buf ( n12168 , n11956 );
and ( n12169 , n12167 , n12168 );
or ( n12170 , C0 , n12169 );
buf ( n12171 , n12170 );
buf ( n12172 , n12171 );
not ( n12173 , n12172 );
not ( n12174 , n12168 );
buf ( n12175 , n12154 );
and ( n12176 , n12174 , n12175 );
xor ( n12177 , n12156 , n12158 );
buf ( n12178 , n12177 );
and ( n12179 , n12178 , n12168 );
or ( n12180 , n12176 , n12179 );
buf ( n12181 , n12180 );
buf ( n12182 , n12181 );
and ( n12183 , n12173 , n12182 );
not ( n12184 , n12182 );
not ( n12185 , n12041 );
xor ( n12186 , n12184 , n12185 );
and ( n12187 , n12186 , n12172 );
or ( n12188 , n12183 , n12187 );
buf ( n12189 , n12188 );
not ( n12190 , n12189 );
buf ( n12191 , n12190 );
buf ( n12192 , n12191 );
not ( n12193 , n12192 );
or ( n12194 , n12046 , n12193 );
not ( n12195 , n12172 );
not ( n12196 , n12168 );
buf ( n12197 , n12141 );
and ( n12198 , n12196 , n12197 );
xor ( n12199 , n12143 , n12159 );
buf ( n12200 , n12199 );
and ( n12201 , n12200 , n12168 );
or ( n12202 , n12198 , n12201 );
buf ( n12203 , n12202 );
buf ( n12204 , n12203 );
and ( n12205 , n12195 , n12204 );
not ( n12206 , n12204 );
and ( n12207 , n12184 , n12185 );
xor ( n12208 , n12206 , n12207 );
and ( n12209 , n12208 , n12172 );
or ( n12210 , n12205 , n12209 );
buf ( n12211 , n12210 );
not ( n12212 , n12211 );
buf ( n12213 , n12212 );
buf ( n12214 , n12213 );
not ( n12215 , n12214 );
or ( n12216 , n12194 , n12215 );
buf ( n12217 , n12216 );
buf ( n12218 , n12217 );
and ( n12219 , n12218 , n12172 );
not ( n12220 , n12219 );
and ( n12221 , n12220 , n12046 );
xor ( n12222 , n12046 , n12172 );
xor ( n12223 , n12222 , n12172 );
and ( n12224 , n12223 , n12219 );
or ( n12225 , n12221 , n12224 );
buf ( n12226 , n12225 );
not ( n12227 , n12219 );
and ( n12228 , n12227 , n12193 );
xor ( n12229 , n12193 , n12172 );
and ( n12230 , n12222 , n12172 );
xor ( n12231 , n12229 , n12230 );
and ( n12232 , n12231 , n12219 );
or ( n12233 , n12228 , n12232 );
buf ( n12234 , n12233 );
not ( n12235 , n12219 );
and ( n12236 , n12235 , n12215 );
xor ( n12237 , n12215 , n12172 );
and ( n12238 , n12229 , n12230 );
xor ( n12239 , n12237 , n12238 );
and ( n12240 , n12239 , n12219 );
or ( n12241 , n12236 , n12240 );
buf ( n12242 , n12241 );
and ( n12243 , n12226 , n12234 , n12242 );
not ( n12244 , n12243 );
buf ( n12245 , GI20478f00_682);
buf ( n12246 , n12245 );
not ( n12247 , n12246 );
buf ( n12248 , RI2106c0b0_602);
buf ( n12249 , n12248 );
and ( n12250 , n12247 , n12249 );
not ( n12251 , n12249 );
buf ( n12252 , RI2106c128_601);
buf ( n12253 , n12252 );
not ( n12254 , n12253 );
buf ( n12255 , RI2106c1a0_600);
buf ( n12256 , n12255 );
not ( n12257 , n12256 );
buf ( n12258 , RI2106c218_599);
buf ( n12259 , n12258 );
not ( n12260 , n12259 );
buf ( n12261 , RI2106c290_598);
buf ( n12262 , n12261 );
not ( n12263 , n12262 );
buf ( n12264 , RI2106a238_641);
buf ( n12265 , n12264 );
not ( n12266 , n12265 );
buf ( n12267 , RI2106a2b0_640);
buf ( n12268 , n12267 );
not ( n12269 , n12268 );
buf ( n12270 , RI2106a328_639);
buf ( n12271 , n12270 );
not ( n12272 , n12271 );
buf ( n12273 , RI2106a3a0_638);
buf ( n12274 , n12273 );
not ( n12275 , n12274 );
buf ( n12276 , RI2106a490_636);
buf ( n12277 , n12276 );
not ( n12278 , n12277 );
buf ( n12279 , RI2106a508_635);
buf ( n12280 , n12279 );
not ( n12281 , n12280 );
buf ( n12282 , RI2106a580_634);
buf ( n12283 , n12282 );
not ( n12284 , n12283 );
buf ( n12285 , RI2106c308_597);
buf ( n12286 , n12285 );
not ( n12287 , n12286 );
buf ( n12288 , RI2106a5f8_633);
buf ( n12289 , n12288 );
not ( n12290 , n12289 );
buf ( n12291 , RI2106a670_632);
buf ( n12292 , n12291 );
not ( n12293 , n12292 );
buf ( n12294 , RI2106a6e8_631);
buf ( n12295 , n12294 );
not ( n12296 , n12295 );
buf ( n12297 , RI2106a760_630);
buf ( n12298 , n12297 );
not ( n12299 , n12298 );
buf ( n12300 , RI2106a7d8_629);
buf ( n12301 , n12300 );
not ( n12302 , n12301 );
buf ( n12303 , RI2106ae68_628);
buf ( n12304 , n12303 );
not ( n12305 , n12304 );
buf ( n12306 , RI21069a40_645);
buf ( n12307 , n12306 );
not ( n12308 , n12307 );
buf ( n12309 , RI2106bed0_606);
buf ( n12310 , n12309 );
not ( n12311 , n12310 );
buf ( n12312 , RI21069ab8_644);
buf ( n12313 , n12312 );
not ( n12314 , n12313 );
buf ( n12315 , RI2106bf48_605);
buf ( n12316 , n12315 );
not ( n12317 , n12316 );
buf ( n12318 , RI2106bfc0_604);
buf ( n12319 , n12318 );
not ( n12320 , n12319 );
buf ( n12321 , RI2106c038_603);
buf ( n12322 , n12321 );
not ( n12323 , n12322 );
buf ( n12324 , RI2106a148_643);
buf ( n12325 , n12324 );
not ( n12326 , n12325 );
buf ( n12327 , RI2106a1c0_642);
buf ( n12328 , n12327 );
not ( n12329 , n12328 );
buf ( n12330 , RI2106a418_637);
buf ( n12331 , n12330 );
not ( n12332 , n12331 );
buf ( n12333 , RI2106c380_596);
buf ( n12334 , n12333 );
not ( n12335 , n12334 );
and ( n12336 , n12332 , n12335 );
and ( n12337 , n12329 , n12336 );
and ( n12338 , n12326 , n12337 );
and ( n12339 , n12323 , n12338 );
and ( n12340 , n12320 , n12339 );
and ( n12341 , n12317 , n12340 );
and ( n12342 , n12314 , n12341 );
and ( n12343 , n12311 , n12342 );
and ( n12344 , n12308 , n12343 );
and ( n12345 , n12305 , n12344 );
and ( n12346 , n12302 , n12345 );
and ( n12347 , n12299 , n12346 );
and ( n12348 , n12296 , n12347 );
and ( n12349 , n12293 , n12348 );
and ( n12350 , n12290 , n12349 );
and ( n12351 , n12287 , n12350 );
and ( n12352 , n12284 , n12351 );
and ( n12353 , n12281 , n12352 );
and ( n12354 , n12278 , n12353 );
and ( n12355 , n12275 , n12354 );
and ( n12356 , n12272 , n12355 );
and ( n12357 , n12269 , n12356 );
and ( n12358 , n12266 , n12357 );
and ( n12359 , n12263 , n12358 );
and ( n12360 , n12260 , n12359 );
and ( n12361 , n12257 , n12360 );
and ( n12362 , n12254 , n12361 );
xor ( n12363 , n12251 , n12362 );
and ( n12364 , n12363 , n12246 );
or ( n12365 , n12250 , n12364 );
buf ( n12366 , n12365 );
not ( n12367 , n12366 );
buf ( n12368 , n12367 );
buf ( n12369 , n12368 );
not ( n12370 , n12369 );
xor ( n12371 , n12370 , n12246 );
not ( n12372 , n12246 );
and ( n12373 , n12372 , n12253 );
xor ( n12374 , n12254 , n12361 );
and ( n12375 , n12374 , n12246 );
or ( n12376 , n12373 , n12375 );
buf ( n12377 , n12376 );
not ( n12378 , n12377 );
buf ( n12379 , n12378 );
buf ( n12380 , n12379 );
not ( n12381 , n12380 );
xor ( n12382 , n12381 , n12246 );
not ( n12383 , n12246 );
and ( n12384 , n12383 , n12256 );
xor ( n12385 , n12257 , n12360 );
and ( n12386 , n12385 , n12246 );
or ( n12387 , n12384 , n12386 );
buf ( n12388 , n12387 );
not ( n12389 , n12388 );
buf ( n12390 , n12389 );
buf ( n12391 , n12390 );
not ( n12392 , n12391 );
xor ( n12393 , n12392 , n12246 );
not ( n12394 , n12246 );
and ( n12395 , n12394 , n12259 );
xor ( n12396 , n12260 , n12359 );
and ( n12397 , n12396 , n12246 );
or ( n12398 , n12395 , n12397 );
buf ( n12399 , n12398 );
not ( n12400 , n12399 );
buf ( n12401 , n12400 );
buf ( n12402 , n12401 );
not ( n12403 , n12402 );
xor ( n12404 , n12403 , n12246 );
not ( n12405 , n12246 );
and ( n12406 , n12405 , n12262 );
xor ( n12407 , n12263 , n12358 );
and ( n12408 , n12407 , n12246 );
or ( n12409 , n12406 , n12408 );
buf ( n12410 , n12409 );
not ( n12411 , n12410 );
buf ( n12412 , n12411 );
buf ( n12413 , n12412 );
not ( n12414 , n12413 );
xor ( n12415 , n12414 , n12246 );
not ( n12416 , n12246 );
and ( n12417 , n12416 , n12265 );
xor ( n12418 , n12266 , n12357 );
and ( n12419 , n12418 , n12246 );
or ( n12420 , n12417 , n12419 );
buf ( n12421 , n12420 );
not ( n12422 , n12421 );
buf ( n12423 , n12422 );
buf ( n12424 , n12423 );
not ( n12425 , n12424 );
xor ( n12426 , n12425 , n12246 );
not ( n12427 , n12246 );
and ( n12428 , n12427 , n12268 );
xor ( n12429 , n12269 , n12356 );
and ( n12430 , n12429 , n12246 );
or ( n12431 , n12428 , n12430 );
buf ( n12432 , n12431 );
not ( n12433 , n12432 );
buf ( n12434 , n12433 );
buf ( n12435 , n12434 );
not ( n12436 , n12435 );
xor ( n12437 , n12436 , n12246 );
not ( n12438 , n12246 );
and ( n12439 , n12438 , n12271 );
xor ( n12440 , n12272 , n12355 );
and ( n12441 , n12440 , n12246 );
or ( n12442 , n12439 , n12441 );
buf ( n12443 , n12442 );
not ( n12444 , n12443 );
buf ( n12445 , n12444 );
buf ( n12446 , n12445 );
not ( n12447 , n12446 );
xor ( n12448 , n12447 , n12246 );
not ( n12449 , n12246 );
and ( n12450 , n12449 , n12274 );
xor ( n12451 , n12275 , n12354 );
and ( n12452 , n12451 , n12246 );
or ( n12453 , n12450 , n12452 );
buf ( n12454 , n12453 );
not ( n12455 , n12454 );
buf ( n12456 , n12455 );
buf ( n12457 , n12456 );
not ( n12458 , n12457 );
xor ( n12459 , n12458 , n12246 );
not ( n12460 , n12246 );
and ( n12461 , n12460 , n12277 );
xor ( n12462 , n12278 , n12353 );
and ( n12463 , n12462 , n12246 );
or ( n12464 , n12461 , n12463 );
buf ( n12465 , n12464 );
not ( n12466 , n12465 );
buf ( n12467 , n12466 );
buf ( n12468 , n12467 );
not ( n12469 , n12468 );
xor ( n12470 , n12469 , n12246 );
not ( n12471 , n12246 );
and ( n12472 , n12471 , n12280 );
xor ( n12473 , n12281 , n12352 );
and ( n12474 , n12473 , n12246 );
or ( n12475 , n12472 , n12474 );
buf ( n12476 , n12475 );
not ( n12477 , n12476 );
buf ( n12478 , n12477 );
buf ( n12479 , n12478 );
not ( n12480 , n12479 );
xor ( n12481 , n12480 , n12246 );
not ( n12482 , n12246 );
and ( n12483 , n12482 , n12283 );
xor ( n12484 , n12284 , n12351 );
and ( n12485 , n12484 , n12246 );
or ( n12486 , n12483 , n12485 );
buf ( n12487 , n12486 );
not ( n12488 , n12487 );
buf ( n12489 , n12488 );
buf ( n12490 , n12489 );
not ( n12491 , n12490 );
xor ( n12492 , n12491 , n12246 );
not ( n12493 , n12246 );
and ( n12494 , n12493 , n12286 );
xor ( n12495 , n12287 , n12350 );
and ( n12496 , n12495 , n12246 );
or ( n12497 , n12494 , n12496 );
buf ( n12498 , n12497 );
not ( n12499 , n12498 );
buf ( n12500 , n12499 );
buf ( n12501 , n12500 );
not ( n12502 , n12501 );
xor ( n12503 , n12502 , n12246 );
not ( n12504 , n12246 );
and ( n12505 , n12504 , n12289 );
xor ( n12506 , n12290 , n12349 );
and ( n12507 , n12506 , n12246 );
or ( n12508 , n12505 , n12507 );
buf ( n12509 , n12508 );
not ( n12510 , n12509 );
buf ( n12511 , n12510 );
buf ( n12512 , n12511 );
not ( n12513 , n12512 );
xor ( n12514 , n12513 , n12246 );
not ( n12515 , n12246 );
and ( n12516 , n12515 , n12292 );
xor ( n12517 , n12293 , n12348 );
and ( n12518 , n12517 , n12246 );
or ( n12519 , n12516 , n12518 );
buf ( n12520 , n12519 );
not ( n12521 , n12520 );
buf ( n12522 , n12521 );
buf ( n12523 , n12522 );
not ( n12524 , n12523 );
xor ( n12525 , n12524 , n12246 );
not ( n12526 , n12246 );
and ( n12527 , n12526 , n12295 );
xor ( n12528 , n12296 , n12347 );
and ( n12529 , n12528 , n12246 );
or ( n12530 , n12527 , n12529 );
buf ( n12531 , n12530 );
not ( n12532 , n12531 );
buf ( n12533 , n12532 );
buf ( n12534 , n12533 );
not ( n12535 , n12534 );
xor ( n12536 , n12535 , n12246 );
not ( n12537 , n12246 );
and ( n12538 , n12537 , n12298 );
xor ( n12539 , n12299 , n12346 );
and ( n12540 , n12539 , n12246 );
or ( n12541 , n12538 , n12540 );
buf ( n12542 , n12541 );
not ( n12543 , n12542 );
buf ( n12544 , n12543 );
buf ( n12545 , n12544 );
not ( n12546 , n12545 );
xor ( n12547 , n12546 , n12246 );
not ( n12548 , n12246 );
and ( n12549 , n12548 , n12301 );
xor ( n12550 , n12302 , n12345 );
and ( n12551 , n12550 , n12246 );
or ( n12552 , n12549 , n12551 );
buf ( n12553 , n12552 );
not ( n12554 , n12553 );
buf ( n12555 , n12554 );
buf ( n12556 , n12555 );
not ( n12557 , n12556 );
xor ( n12558 , n12557 , n12246 );
not ( n12559 , n12246 );
and ( n12560 , n12559 , n12304 );
xor ( n12561 , n12305 , n12344 );
and ( n12562 , n12561 , n12246 );
or ( n12563 , n12560 , n12562 );
buf ( n12564 , n12563 );
not ( n12565 , n12564 );
buf ( n12566 , n12565 );
buf ( n12567 , n12566 );
not ( n12568 , n12567 );
xor ( n12569 , n12568 , n12246 );
not ( n12570 , n12246 );
and ( n12571 , n12570 , n12307 );
xor ( n12572 , n12308 , n12343 );
and ( n12573 , n12572 , n12246 );
or ( n12574 , n12571 , n12573 );
buf ( n12575 , n12574 );
not ( n12576 , n12575 );
buf ( n12577 , n12576 );
buf ( n12578 , n12577 );
not ( n12579 , n12578 );
xor ( n12580 , n12579 , n12246 );
not ( n12581 , n12246 );
and ( n12582 , n12581 , n12310 );
xor ( n12583 , n12311 , n12342 );
and ( n12584 , n12583 , n12246 );
or ( n12585 , n12582 , n12584 );
buf ( n12586 , n12585 );
not ( n12587 , n12586 );
buf ( n12588 , n12587 );
buf ( n12589 , n12588 );
not ( n12590 , n12589 );
xor ( n12591 , n12590 , n12246 );
not ( n12592 , n12246 );
and ( n12593 , n12592 , n12313 );
xor ( n12594 , n12314 , n12341 );
and ( n12595 , n12594 , n12246 );
or ( n12596 , n12593 , n12595 );
buf ( n12597 , n12596 );
not ( n12598 , n12597 );
buf ( n12599 , n12598 );
buf ( n12600 , n12599 );
not ( n12601 , n12600 );
xor ( n12602 , n12601 , n12246 );
not ( n12603 , n12246 );
and ( n12604 , n12603 , n12316 );
xor ( n12605 , n12317 , n12340 );
and ( n12606 , n12605 , n12246 );
or ( n12607 , n12604 , n12606 );
buf ( n12608 , n12607 );
not ( n12609 , n12608 );
buf ( n12610 , n12609 );
buf ( n12611 , n12610 );
not ( n12612 , n12611 );
xor ( n12613 , n12612 , n12246 );
not ( n12614 , n12246 );
and ( n12615 , n12614 , n12319 );
xor ( n12616 , n12320 , n12339 );
and ( n12617 , n12616 , n12246 );
or ( n12618 , n12615 , n12617 );
buf ( n12619 , n12618 );
not ( n12620 , n12619 );
buf ( n12621 , n12620 );
buf ( n12622 , n12621 );
not ( n12623 , n12622 );
xor ( n12624 , n12623 , n12246 );
not ( n12625 , n12246 );
and ( n12626 , n12625 , n12322 );
xor ( n12627 , n12323 , n12338 );
and ( n12628 , n12627 , n12246 );
or ( n12629 , n12626 , n12628 );
buf ( n12630 , n12629 );
not ( n12631 , n12630 );
buf ( n12632 , n12631 );
buf ( n12633 , n12632 );
not ( n12634 , n12633 );
xor ( n12635 , n12634 , n12246 );
not ( n12636 , n12246 );
and ( n12637 , n12636 , n12325 );
xor ( n12638 , n12326 , n12337 );
and ( n12639 , n12638 , n12246 );
or ( n12640 , n12637 , n12639 );
buf ( n12641 , n12640 );
not ( n12642 , n12641 );
buf ( n12643 , n12642 );
buf ( n12644 , n12643 );
not ( n12645 , n12644 );
xor ( n12646 , n12645 , n12246 );
not ( n12647 , n12246 );
and ( n12648 , n12647 , n12328 );
xor ( n12649 , n12329 , n12336 );
and ( n12650 , n12649 , n12246 );
or ( n12651 , n12648 , n12650 );
buf ( n12652 , n12651 );
not ( n12653 , n12652 );
buf ( n12654 , n12653 );
buf ( n12655 , n12654 );
not ( n12656 , n12655 );
xor ( n12657 , n12656 , n12246 );
not ( n12658 , n12246 );
and ( n12659 , n12658 , n12331 );
xor ( n12660 , n12332 , n12335 );
and ( n12661 , n12660 , n12246 );
or ( n12662 , n12659 , n12661 );
buf ( n12663 , n12662 );
not ( n12664 , n12663 );
buf ( n12665 , n12664 );
buf ( n12666 , n12665 );
not ( n12667 , n12666 );
xor ( n12668 , n12667 , n12246 );
buf ( n12669 , n12334 );
not ( n12670 , n12669 );
buf ( n12671 , n12670 );
buf ( n12672 , n12671 );
not ( n12673 , n12672 );
xor ( n12674 , n12673 , n12246 );
and ( n12675 , n12674 , n12246 );
and ( n12676 , n12668 , n12675 );
and ( n12677 , n12657 , n12676 );
and ( n12678 , n12646 , n12677 );
and ( n12679 , n12635 , n12678 );
and ( n12680 , n12624 , n12679 );
and ( n12681 , n12613 , n12680 );
and ( n12682 , n12602 , n12681 );
and ( n12683 , n12591 , n12682 );
and ( n12684 , n12580 , n12683 );
and ( n12685 , n12569 , n12684 );
and ( n12686 , n12558 , n12685 );
and ( n12687 , n12547 , n12686 );
and ( n12688 , n12536 , n12687 );
and ( n12689 , n12525 , n12688 );
and ( n12690 , n12514 , n12689 );
and ( n12691 , n12503 , n12690 );
and ( n12692 , n12492 , n12691 );
and ( n12693 , n12481 , n12692 );
and ( n12694 , n12470 , n12693 );
and ( n12695 , n12459 , n12694 );
and ( n12696 , n12448 , n12695 );
and ( n12697 , n12437 , n12696 );
and ( n12698 , n12426 , n12697 );
and ( n12699 , n12415 , n12698 );
and ( n12700 , n12404 , n12699 );
and ( n12701 , n12393 , n12700 );
and ( n12702 , n12382 , n12701 );
and ( n12703 , n12371 , n12702 );
buf ( n12704 , n12703 );
or ( n12705 , n12673 , n12667 );
or ( n12706 , n12705 , n12656 );
or ( n12707 , n12706 , n12645 );
or ( n12708 , n12707 , n12634 );
or ( n12709 , n12708 , n12623 );
or ( n12710 , n12709 , n12612 );
or ( n12711 , n12710 , n12601 );
or ( n12712 , n12711 , n12590 );
or ( n12713 , n12712 , n12579 );
or ( n12714 , n12713 , n12568 );
or ( n12715 , n12714 , n12557 );
or ( n12716 , n12715 , n12546 );
or ( n12717 , n12716 , n12535 );
or ( n12718 , n12717 , n12524 );
or ( n12719 , n12718 , n12513 );
or ( n12720 , n12719 , n12502 );
or ( n12721 , n12720 , n12491 );
or ( n12722 , n12721 , n12480 );
or ( n12723 , n12722 , n12469 );
or ( n12724 , n12723 , n12458 );
or ( n12725 , n12724 , n12447 );
or ( n12726 , n12725 , n12436 );
or ( n12727 , n12726 , n12425 );
or ( n12728 , n12727 , n12414 );
or ( n12729 , n12728 , n12403 );
or ( n12730 , n12729 , n12392 );
or ( n12731 , n12730 , n12381 );
or ( n12732 , n12731 , n12370 );
buf ( n12733 , n12732 );
buf ( n12734 , n12733 );
and ( n12735 , n12734 , n12246 );
and ( n12736 , n12704 , n12735 );
or ( n12737 , C0 , n12736 );
buf ( n12738 , n12737 );
buf ( n12739 , n12738 );
not ( n12740 , n12735 );
and ( n12741 , n12740 , n12370 );
xor ( n12742 , n12371 , n12702 );
and ( n12743 , n12742 , n12735 );
or ( n12744 , n12741 , n12743 );
buf ( n12745 , n12744 );
buf ( n12746 , n12745 );
not ( n12747 , n12735 );
and ( n12748 , n12747 , n12381 );
xor ( n12749 , n12382 , n12701 );
and ( n12750 , n12749 , n12735 );
or ( n12751 , n12748 , n12750 );
buf ( n12752 , n12751 );
buf ( n12753 , n12752 );
not ( n12754 , n12735 );
and ( n12755 , n12754 , n12392 );
xor ( n12756 , n12393 , n12700 );
and ( n12757 , n12756 , n12735 );
or ( n12758 , n12755 , n12757 );
buf ( n12759 , n12758 );
buf ( n12760 , n12759 );
not ( n12761 , n12735 );
and ( n12762 , n12761 , n12403 );
xor ( n12763 , n12404 , n12699 );
and ( n12764 , n12763 , n12735 );
or ( n12765 , n12762 , n12764 );
buf ( n12766 , n12765 );
buf ( n12767 , n12766 );
not ( n12768 , n12735 );
and ( n12769 , n12768 , n12414 );
xor ( n12770 , n12415 , n12698 );
and ( n12771 , n12770 , n12735 );
or ( n12772 , n12769 , n12771 );
buf ( n12773 , n12772 );
buf ( n12774 , n12773 );
not ( n12775 , n12735 );
and ( n12776 , n12775 , n12425 );
xor ( n12777 , n12426 , n12697 );
and ( n12778 , n12777 , n12735 );
or ( n12779 , n12776 , n12778 );
buf ( n12780 , n12779 );
buf ( n12781 , n12780 );
not ( n12782 , n12735 );
and ( n12783 , n12782 , n12436 );
xor ( n12784 , n12437 , n12696 );
and ( n12785 , n12784 , n12735 );
or ( n12786 , n12783 , n12785 );
buf ( n12787 , n12786 );
buf ( n12788 , n12787 );
not ( n12789 , n12735 );
and ( n12790 , n12789 , n12447 );
xor ( n12791 , n12448 , n12695 );
and ( n12792 , n12791 , n12735 );
or ( n12793 , n12790 , n12792 );
buf ( n12794 , n12793 );
buf ( n12795 , n12794 );
not ( n12796 , n12735 );
and ( n12797 , n12796 , n12458 );
xor ( n12798 , n12459 , n12694 );
and ( n12799 , n12798 , n12735 );
or ( n12800 , n12797 , n12799 );
buf ( n12801 , n12800 );
buf ( n12802 , n12801 );
not ( n12803 , n12735 );
and ( n12804 , n12803 , n12469 );
xor ( n12805 , n12470 , n12693 );
and ( n12806 , n12805 , n12735 );
or ( n12807 , n12804 , n12806 );
buf ( n12808 , n12807 );
buf ( n12809 , n12808 );
not ( n12810 , n12735 );
and ( n12811 , n12810 , n12480 );
xor ( n12812 , n12481 , n12692 );
and ( n12813 , n12812 , n12735 );
or ( n12814 , n12811 , n12813 );
buf ( n12815 , n12814 );
buf ( n12816 , n12815 );
not ( n12817 , n12735 );
and ( n12818 , n12817 , n12491 );
xor ( n12819 , n12492 , n12691 );
and ( n12820 , n12819 , n12735 );
or ( n12821 , n12818 , n12820 );
buf ( n12822 , n12821 );
buf ( n12823 , n12822 );
not ( n12824 , n12735 );
and ( n12825 , n12824 , n12502 );
xor ( n12826 , n12503 , n12690 );
and ( n12827 , n12826 , n12735 );
or ( n12828 , n12825 , n12827 );
buf ( n12829 , n12828 );
buf ( n12830 , n12829 );
not ( n12831 , n12735 );
and ( n12832 , n12831 , n12513 );
xor ( n12833 , n12514 , n12689 );
and ( n12834 , n12833 , n12735 );
or ( n12835 , n12832 , n12834 );
buf ( n12836 , n12835 );
buf ( n12837 , n12836 );
not ( n12838 , n12735 );
and ( n12839 , n12838 , n12524 );
xor ( n12840 , n12525 , n12688 );
and ( n12841 , n12840 , n12735 );
or ( n12842 , n12839 , n12841 );
buf ( n12843 , n12842 );
buf ( n12844 , n12843 );
not ( n12845 , n12735 );
and ( n12846 , n12845 , n12535 );
xor ( n12847 , n12536 , n12687 );
and ( n12848 , n12847 , n12735 );
or ( n12849 , n12846 , n12848 );
buf ( n12850 , n12849 );
buf ( n12851 , n12850 );
not ( n12852 , n12735 );
and ( n12853 , n12852 , n12546 );
xor ( n12854 , n12547 , n12686 );
and ( n12855 , n12854 , n12735 );
or ( n12856 , n12853 , n12855 );
buf ( n12857 , n12856 );
buf ( n12858 , n12857 );
not ( n12859 , n12735 );
and ( n12860 , n12859 , n12557 );
xor ( n12861 , n12558 , n12685 );
and ( n12862 , n12861 , n12735 );
or ( n12863 , n12860 , n12862 );
buf ( n12864 , n12863 );
buf ( n12865 , n12864 );
not ( n12866 , n12735 );
and ( n12867 , n12866 , n12568 );
xor ( n12868 , n12569 , n12684 );
and ( n12869 , n12868 , n12735 );
or ( n12870 , n12867 , n12869 );
buf ( n12871 , n12870 );
buf ( n12872 , n12871 );
not ( n12873 , n12735 );
and ( n12874 , n12873 , n12579 );
xor ( n12875 , n12580 , n12683 );
and ( n12876 , n12875 , n12735 );
or ( n12877 , n12874 , n12876 );
buf ( n12878 , n12877 );
buf ( n12879 , n12878 );
not ( n12880 , n12735 );
and ( n12881 , n12880 , n12590 );
xor ( n12882 , n12591 , n12682 );
and ( n12883 , n12882 , n12735 );
or ( n12884 , n12881 , n12883 );
buf ( n12885 , n12884 );
buf ( n12886 , n12885 );
not ( n12887 , n12735 );
and ( n12888 , n12887 , n12601 );
xor ( n12889 , n12602 , n12681 );
and ( n12890 , n12889 , n12735 );
or ( n12891 , n12888 , n12890 );
buf ( n12892 , n12891 );
buf ( n12893 , n12892 );
not ( n12894 , n12735 );
and ( n12895 , n12894 , n12612 );
xor ( n12896 , n12613 , n12680 );
and ( n12897 , n12896 , n12735 );
or ( n12898 , n12895 , n12897 );
buf ( n12899 , n12898 );
buf ( n12900 , n12899 );
not ( n12901 , n12735 );
and ( n12902 , n12901 , n12623 );
xor ( n12903 , n12624 , n12679 );
and ( n12904 , n12903 , n12735 );
or ( n12905 , n12902 , n12904 );
buf ( n12906 , n12905 );
buf ( n12907 , n12906 );
not ( n12908 , n12735 );
and ( n12909 , n12908 , n12634 );
xor ( n12910 , n12635 , n12678 );
and ( n12911 , n12910 , n12735 );
or ( n12912 , n12909 , n12911 );
buf ( n12913 , n12912 );
buf ( n12914 , n12913 );
not ( n12915 , n12735 );
and ( n12916 , n12915 , n12645 );
xor ( n12917 , n12646 , n12677 );
and ( n12918 , n12917 , n12735 );
or ( n12919 , n12916 , n12918 );
buf ( n12920 , n12919 );
buf ( n12921 , n12920 );
or ( n12922 , n12914 , n12921 );
or ( n12923 , n12907 , n12922 );
or ( n12924 , n12900 , n12923 );
or ( n12925 , n12893 , n12924 );
or ( n12926 , n12886 , n12925 );
or ( n12927 , n12879 , n12926 );
or ( n12928 , n12872 , n12927 );
or ( n12929 , n12865 , n12928 );
or ( n12930 , n12858 , n12929 );
or ( n12931 , n12851 , n12930 );
or ( n12932 , n12844 , n12931 );
or ( n12933 , n12837 , n12932 );
or ( n12934 , n12830 , n12933 );
or ( n12935 , n12823 , n12934 );
or ( n12936 , n12816 , n12935 );
or ( n12937 , n12809 , n12936 );
or ( n12938 , n12802 , n12937 );
or ( n12939 , n12795 , n12938 );
or ( n12940 , n12788 , n12939 );
or ( n12941 , n12781 , n12940 );
or ( n12942 , n12774 , n12941 );
or ( n12943 , n12767 , n12942 );
or ( n12944 , n12760 , n12943 );
or ( n12945 , n12753 , n12944 );
or ( n12946 , n12746 , n12945 );
or ( n12947 , n12739 , n12946 );
buf ( n12948 , n12947 );
not ( n12949 , n12948 );
buf ( n12950 , n12949 );
buf ( n12951 , n11504 );
not ( n12952 , n12951 );
buf ( n12953 , n11776 );
and ( n12954 , n12952 , n12953 );
not ( n12955 , n12953 );
buf ( n12956 , n11784 );
not ( n12957 , n12956 );
buf ( n12958 , n11792 );
not ( n12959 , n12958 );
buf ( n12960 , n11800 );
not ( n12961 , n12960 );
buf ( n12962 , n11808 );
not ( n12963 , n12962 );
buf ( n12964 , n11816 );
not ( n12965 , n12964 );
buf ( n12966 , n11512 );
not ( n12967 , n12966 );
buf ( n12968 , n11521 );
not ( n12969 , n12968 );
buf ( n12970 , n11529 );
not ( n12971 , n12970 );
buf ( n12972 , n11537 );
not ( n12973 , n12972 );
buf ( n12974 , n11545 );
not ( n12975 , n12974 );
buf ( n12976 , n11553 );
not ( n12977 , n12976 );
buf ( n12978 , n11561 );
not ( n12979 , n12978 );
buf ( n12980 , n11569 );
not ( n12981 , n12980 );
buf ( n12982 , n11577 );
not ( n12983 , n12982 );
buf ( n12984 , n11585 );
not ( n12985 , n12984 );
buf ( n12986 , n11593 );
not ( n12987 , n12986 );
buf ( n12988 , n11601 );
not ( n12989 , n12988 );
buf ( n12990 , n11609 );
not ( n12991 , n12990 );
buf ( n12992 , n11617 );
not ( n12993 , n12992 );
buf ( n12994 , n11625 );
not ( n12995 , n12994 );
buf ( n12996 , n11633 );
not ( n12997 , n12996 );
buf ( n12998 , n11641 );
not ( n12999 , n12998 );
buf ( n13000 , n11649 );
not ( n13001 , n13000 );
buf ( n13002 , n11657 );
not ( n13003 , n13002 );
buf ( n13004 , n11665 );
not ( n13005 , n13004 );
buf ( n13006 , n11673 );
not ( n13007 , n13006 );
buf ( n13008 , n11681 );
not ( n13009 , n13008 );
buf ( n13010 , n11689 );
not ( n13011 , n13010 );
buf ( n13012 , n11692 );
not ( n13013 , n13012 );
and ( n13014 , n13011 , n13013 );
and ( n13015 , n13009 , n13014 );
and ( n13016 , n13007 , n13015 );
and ( n13017 , n13005 , n13016 );
and ( n13018 , n13003 , n13017 );
and ( n13019 , n13001 , n13018 );
and ( n13020 , n12999 , n13019 );
and ( n13021 , n12997 , n13020 );
and ( n13022 , n12995 , n13021 );
and ( n13023 , n12993 , n13022 );
and ( n13024 , n12991 , n13023 );
and ( n13025 , n12989 , n13024 );
and ( n13026 , n12987 , n13025 );
and ( n13027 , n12985 , n13026 );
and ( n13028 , n12983 , n13027 );
and ( n13029 , n12981 , n13028 );
and ( n13030 , n12979 , n13029 );
and ( n13031 , n12977 , n13030 );
and ( n13032 , n12975 , n13031 );
and ( n13033 , n12973 , n13032 );
and ( n13034 , n12971 , n13033 );
and ( n13035 , n12969 , n13034 );
and ( n13036 , n12967 , n13035 );
and ( n13037 , n12965 , n13036 );
and ( n13038 , n12963 , n13037 );
and ( n13039 , n12961 , n13038 );
and ( n13040 , n12959 , n13039 );
and ( n13041 , n12957 , n13040 );
xor ( n13042 , n12955 , n13041 );
and ( n13043 , n13042 , n12951 );
or ( n13044 , n12954 , n13043 );
buf ( n13045 , n13044 );
not ( n13046 , n13045 );
buf ( n13047 , n13046 );
buf ( n13048 , n13047 );
not ( n13049 , n13048 );
buf ( n13050 , n13049 );
buf ( n13051 , n13050 );
buf ( n13052 , n13051 );
not ( n13053 , n13052 );
buf ( n13054 , n13053 );
buf ( n13055 , n13054 );
not ( n13056 , n13055 );
not ( n13057 , n12951 );
buf ( n13058 , n11768 );
not ( n13059 , n13058 );
and ( n13060 , n12955 , n13041 );
and ( n13061 , n13059 , n13060 );
xor ( n13062 , n13057 , n13061 );
buf ( n13063 , n12951 );
and ( n13064 , n13062 , n13063 );
or ( n13065 , C0 , n13064 );
buf ( n13066 , n13065 );
not ( n13067 , n13066 );
buf ( n13068 , n13067 );
buf ( n13069 , n13068 );
not ( n13070 , n13069 );
buf ( n13071 , n13070 );
not ( n13072 , n13071 );
buf ( n13073 , n13072 );
not ( n13074 , n12951 );
and ( n13075 , n13074 , n13058 );
xor ( n13076 , n13059 , n13060 );
and ( n13077 , n13076 , n12951 );
or ( n13078 , n13075 , n13077 );
buf ( n13079 , n13078 );
not ( n13080 , n13079 );
buf ( n13081 , n13080 );
buf ( n13082 , n13081 );
not ( n13083 , n13082 );
buf ( n13084 , n13083 );
not ( n13085 , n13084 );
buf ( n13086 , n13085 );
not ( n13087 , n13050 );
buf ( n13088 , n13087 );
and ( n13089 , n13086 , n13088 );
and ( n13090 , n13073 , n13089 );
not ( n13091 , n13090 );
buf ( n13092 , n13091 );
buf ( n13093 , n12951 );
and ( n13094 , n13092 , n13093 );
or ( n13095 , C0 , n13094 );
buf ( n13096 , n13095 );
buf ( n13097 , n13096 );
not ( n13098 , n13097 );
not ( n13099 , n13093 );
buf ( n13100 , n13084 );
and ( n13101 , n13099 , n13100 );
xor ( n13102 , n13086 , n13088 );
buf ( n13103 , n13102 );
and ( n13104 , n13103 , n13093 );
or ( n13105 , n13101 , n13104 );
buf ( n13106 , n13105 );
buf ( n13107 , n13106 );
and ( n13108 , n13098 , n13107 );
not ( n13109 , n13107 );
not ( n13110 , n13051 );
xor ( n13111 , n13109 , n13110 );
and ( n13112 , n13111 , n13097 );
or ( n13113 , n13108 , n13112 );
buf ( n13114 , n13113 );
not ( n13115 , n13114 );
buf ( n13116 , n13115 );
buf ( n13117 , n13116 );
not ( n13118 , n13117 );
or ( n13119 , n13056 , n13118 );
buf ( n13120 , n13119 );
buf ( n13121 , n13120 );
and ( n13122 , n13121 , n13097 );
not ( n13123 , n13122 );
and ( n13124 , n13123 , n13056 );
xor ( n13125 , n13056 , n13097 );
xor ( n13126 , n13125 , n13097 );
and ( n13127 , n13126 , n13122 );
or ( n13128 , n13124 , n13127 );
buf ( n13129 , n13128 );
not ( n13130 , n13122 );
and ( n13131 , n13130 , n13118 );
xor ( n13132 , n13118 , n13097 );
and ( n13133 , n13125 , n13097 );
xor ( n13134 , n13132 , n13133 );
and ( n13135 , n13134 , n13122 );
or ( n13136 , n13131 , n13135 );
buf ( n13137 , n13136 );
and ( n13138 , n13129 , n13137 );
and ( n13139 , n12950 , n13138 );
buf ( n13140 , RI2106cbf0_591);
not ( n13141 , n13129 );
and ( n13142 , n13141 , n13137 );
and ( n13143 , n13140 , n13142 );
buf ( n13144 , RI2106dd48_567);
nor ( n13145 , n13141 , n13137 );
and ( n13146 , n13144 , n13145 );
buf ( n13147 , RI21073040_543);
nor ( n13148 , n13129 , n13137 );
and ( n13149 , n13147 , n13148 );
or ( n13150 , n13139 , n13143 , n13146 , n13149 );
buf ( n13151 , n13150 );
not ( n13152 , n13151 );
xnor ( n13153 , n12746 , n12945 );
buf ( n13154 , n13153 );
and ( n13155 , n13154 , n13138 );
buf ( n13156 , RI2106cd58_588);
and ( n13157 , n13156 , n13142 );
buf ( n13158 , RI2106deb0_564);
and ( n13159 , n13158 , n13145 );
buf ( n13160 , RI21073c70_539);
and ( n13161 , n13160 , n13148 );
or ( n13162 , n13155 , n13157 , n13159 , n13161 );
buf ( n13163 , n13162 );
and ( n13164 , n13152 , n13163 );
not ( n13165 , n13163 );
xnor ( n13166 , n12753 , n12944 );
buf ( n13167 , n13166 );
and ( n13168 , n13167 , n13138 );
buf ( n13169 , RI2106cdd0_587);
and ( n13170 , n13169 , n13142 );
buf ( n13171 , RI2106df28_563);
and ( n13172 , n13171 , n13145 );
buf ( n13173 , RI21073ce8_538);
and ( n13174 , n13173 , n13148 );
or ( n13175 , n13168 , n13170 , n13172 , n13174 );
buf ( n13176 , n13175 );
not ( n13177 , n13176 );
xnor ( n13178 , n12760 , n12943 );
buf ( n13179 , n13178 );
and ( n13180 , n13179 , n13138 );
buf ( n13181 , RI2106ce48_586);
and ( n13182 , n13181 , n13142 );
buf ( n13183 , RI2106dfa0_562);
and ( n13184 , n13183 , n13145 );
buf ( n13185 , RI21073d60_537);
and ( n13186 , n13185 , n13148 );
or ( n13187 , n13180 , n13182 , n13184 , n13186 );
buf ( n13188 , n13187 );
not ( n13189 , n13188 );
xnor ( n13190 , n12767 , n12942 );
buf ( n13191 , n13190 );
and ( n13192 , n13191 , n13138 );
buf ( n13193 , RI2106cec0_585);
and ( n13194 , n13193 , n13142 );
buf ( n13195 , RI2106e018_561);
and ( n13196 , n13195 , n13145 );
buf ( n13197 , RI21073dd8_536);
and ( n13198 , n13197 , n13148 );
or ( n13199 , n13192 , n13194 , n13196 , n13198 );
buf ( n13200 , n13199 );
not ( n13201 , n13200 );
xnor ( n13202 , n12774 , n12941 );
buf ( n13203 , n13202 );
and ( n13204 , n13203 , n13138 );
buf ( n13205 , RI2106cf38_584);
and ( n13206 , n13205 , n13142 );
buf ( n13207 , RI2106e090_560);
and ( n13208 , n13207 , n13145 );
buf ( n13209 , RI210748a0_535);
and ( n13210 , n13209 , n13148 );
or ( n13211 , n13204 , n13206 , n13208 , n13210 );
buf ( n13212 , n13211 );
not ( n13213 , n13212 );
xnor ( n13214 , n12781 , n12940 );
buf ( n13215 , n13214 );
and ( n13216 , n13215 , n13138 );
buf ( n13217 , RI2106cfb0_583);
and ( n13218 , n13217 , n13142 );
buf ( n13219 , RI2106e108_559);
and ( n13220 , n13219 , n13145 );
buf ( n13221 , RI21074918_534);
and ( n13222 , n13221 , n13148 );
or ( n13223 , n13216 , n13218 , n13220 , n13222 );
buf ( n13224 , n13223 );
not ( n13225 , n13224 );
xnor ( n13226 , n12788 , n12939 );
buf ( n13227 , n13226 );
and ( n13228 , n13227 , n13138 );
buf ( n13229 , RI2106d028_582);
and ( n13230 , n13229 , n13142 );
buf ( n13231 , RI21070a48_558);
and ( n13232 , n13231 , n13145 );
buf ( n13233 , RI21074990_533);
and ( n13234 , n13233 , n13148 );
or ( n13235 , n13228 , n13230 , n13232 , n13234 );
buf ( n13236 , n13235 );
not ( n13237 , n13236 );
xnor ( n13238 , n12795 , n12938 );
buf ( n13239 , n13238 );
and ( n13240 , n13239 , n13138 );
buf ( n13241 , RI2106d0a0_581);
and ( n13242 , n13241 , n13142 );
buf ( n13243 , RI21070ac0_557);
and ( n13244 , n13243 , n13145 );
buf ( n13245 , RI21074a08_532);
and ( n13246 , n13245 , n13148 );
or ( n13247 , n13240 , n13242 , n13244 , n13246 );
buf ( n13248 , n13247 );
not ( n13249 , n13248 );
xnor ( n13250 , n12802 , n12937 );
buf ( n13251 , n13250 );
and ( n13252 , n13251 , n13138 );
buf ( n13253 , RI2106d118_580);
and ( n13254 , n13253 , n13142 );
buf ( n13255 , RI21071588_556);
and ( n13256 , n13255 , n13145 );
buf ( n13257 , RI21074a80_531);
and ( n13258 , n13257 , n13148 );
or ( n13259 , n13252 , n13254 , n13256 , n13258 );
buf ( n13260 , n13259 );
not ( n13261 , n13260 );
xnor ( n13262 , n12809 , n12936 );
buf ( n13263 , n13262 );
and ( n13264 , n13263 , n13138 );
buf ( n13265 , RI2106b138_622);
and ( n13266 , n13265 , n13142 );
buf ( n13267 , RI2106b4f8_614);
and ( n13268 , n13267 , n13145 );
buf ( n13269 , RI210755c0_529);
and ( n13270 , n13269 , n13148 );
or ( n13271 , n13264 , n13266 , n13268 , n13270 );
buf ( n13272 , n13271 );
not ( n13273 , n13272 );
xnor ( n13274 , n12816 , n12935 );
buf ( n13275 , n13274 );
and ( n13276 , n13275 , n13138 );
buf ( n13277 , RI2106b1b0_621);
and ( n13278 , n13277 , n13142 );
buf ( n13279 , RI2106b570_613);
and ( n13280 , n13279 , n13145 );
buf ( n13281 , RI21075638_528);
and ( n13282 , n13281 , n13148 );
or ( n13283 , n13276 , n13278 , n13280 , n13282 );
buf ( n13284 , n13283 );
not ( n13285 , n13284 );
xnor ( n13286 , n12823 , n12934 );
buf ( n13287 , n13286 );
and ( n13288 , n13287 , n13138 );
buf ( n13289 , RI2106b228_620);
and ( n13290 , n13289 , n13142 );
buf ( n13291 , RI2106bc00_612);
and ( n13292 , n13291 , n13145 );
buf ( n13293 , RI210756b0_527);
and ( n13294 , n13293 , n13148 );
or ( n13295 , n13288 , n13290 , n13292 , n13294 );
buf ( n13296 , n13295 );
not ( n13297 , n13296 );
xnor ( n13298 , n12830 , n12933 );
buf ( n13299 , n13298 );
and ( n13300 , n13299 , n13138 );
buf ( n13301 , RI2106d190_579);
and ( n13302 , n13301 , n13142 );
buf ( n13303 , RI21071600_555);
and ( n13304 , n13303 , n13145 );
buf ( n13305 , RI21075728_526);
and ( n13306 , n13305 , n13148 );
or ( n13307 , n13300 , n13302 , n13304 , n13306 );
buf ( n13308 , n13307 );
not ( n13309 , n13308 );
xnor ( n13310 , n12837 , n12932 );
buf ( n13311 , n13310 );
and ( n13312 , n13311 , n13138 );
buf ( n13313 , RI2106d208_578);
and ( n13314 , n13313 , n13142 );
buf ( n13315 , RI21071678_554);
and ( n13316 , n13315 , n13145 );
buf ( n13317 , RI210757a0_525);
and ( n13318 , n13317 , n13148 );
or ( n13319 , n13312 , n13314 , n13316 , n13318 );
buf ( n13320 , n13319 );
not ( n13321 , n13320 );
xnor ( n13322 , n12844 , n12931 );
buf ( n13323 , n13322 );
and ( n13324 , n13323 , n13138 );
buf ( n13325 , RI2106d898_577);
and ( n13326 , n13325 , n13142 );
buf ( n13327 , RI2106bc78_611);
and ( n13328 , n13327 , n13145 );
buf ( n13329 , RI21075818_524);
and ( n13330 , n13329 , n13148 );
or ( n13331 , n13324 , n13326 , n13328 , n13330 );
buf ( n13332 , n13331 );
not ( n13333 , n13332 );
xnor ( n13334 , n12851 , n12930 );
buf ( n13335 , n13334 );
and ( n13336 , n13335 , n13138 );
buf ( n13337 , RI2106d910_576);
and ( n13338 , n13337 , n13142 );
buf ( n13339 , RI2106bcf0_610);
and ( n13340 , n13339 , n13145 );
buf ( n13341 , RI210762e0_523);
and ( n13342 , n13341 , n13148 );
or ( n13343 , n13336 , n13338 , n13340 , n13342 );
buf ( n13344 , n13343 );
not ( n13345 , n13344 );
xnor ( n13346 , n12858 , n12929 );
buf ( n13347 , n13346 );
and ( n13348 , n13347 , n13138 );
buf ( n13349 , RI2106d988_575);
and ( n13350 , n13349 , n13142 );
buf ( n13351 , RI210716f0_553);
and ( n13352 , n13351 , n13145 );
buf ( n13353 , RI21076358_522);
and ( n13354 , n13353 , n13148 );
or ( n13355 , n13348 , n13350 , n13352 , n13354 );
buf ( n13356 , n13355 );
not ( n13357 , n13356 );
xnor ( n13358 , n12865 , n12928 );
buf ( n13359 , n13358 );
and ( n13360 , n13359 , n13138 );
buf ( n13361 , RI2106da00_574);
and ( n13362 , n13361 , n13142 );
buf ( n13363 , RI210721b8_552);
and ( n13364 , n13363 , n13145 );
buf ( n13365 , RI210763d0_521);
and ( n13366 , n13365 , n13148 );
or ( n13367 , n13360 , n13362 , n13364 , n13366 );
buf ( n13368 , n13367 );
not ( n13369 , n13368 );
xnor ( n13370 , n12872 , n12927 );
buf ( n13371 , n13370 );
and ( n13372 , n13371 , n13138 );
buf ( n13373 , RI2106da78_573);
and ( n13374 , n13373 , n13142 );
buf ( n13375 , RI2106bd68_609);
and ( n13376 , n13375 , n13145 );
buf ( n13377 , RI21076448_520);
and ( n13378 , n13377 , n13148 );
or ( n13379 , n13372 , n13374 , n13376 , n13378 );
buf ( n13380 , n13379 );
not ( n13381 , n13380 );
xnor ( n13382 , n12879 , n12926 );
buf ( n13383 , n13382 );
and ( n13384 , n13383 , n13138 );
buf ( n13385 , RI2106ca10_595);
and ( n13386 , n13385 , n13142 );
buf ( n13387 , RI2106db68_571);
and ( n13388 , n13387 , n13145 );
buf ( n13389 , RI210722a8_550);
and ( n13390 , n13389 , n13148 );
or ( n13391 , n13384 , n13386 , n13388 , n13390 );
buf ( n13392 , n13391 );
not ( n13393 , n13392 );
xnor ( n13394 , n12886 , n12925 );
buf ( n13395 , n13394 );
and ( n13396 , n13395 , n13138 );
buf ( n13397 , RI2106ca88_594);
and ( n13398 , n13397 , n13142 );
buf ( n13399 , RI2106dbe0_570);
and ( n13400 , n13399 , n13145 );
buf ( n13401 , RI21072320_549);
and ( n13402 , n13401 , n13148 );
or ( n13403 , n13396 , n13398 , n13400 , n13402 );
buf ( n13404 , n13403 );
not ( n13405 , n13404 );
xnor ( n13406 , n12893 , n12924 );
buf ( n13407 , n13406 );
and ( n13408 , n13407 , n13138 );
buf ( n13409 , RI2106aee0_627);
and ( n13410 , n13409 , n13142 );
buf ( n13411 , RI2106dc58_569);
and ( n13412 , n13411 , n13145 );
buf ( n13413 , RI21072398_548);
and ( n13414 , n13413 , n13148 );
or ( n13415 , n13408 , n13410 , n13412 , n13414 );
buf ( n13416 , n13415 );
not ( n13417 , n13416 );
xnor ( n13418 , n12900 , n12923 );
buf ( n13419 , n13418 );
and ( n13420 , n13419 , n13138 );
buf ( n13421 , RI2106af58_626);
and ( n13422 , n13421 , n13142 );
buf ( n13423 , RI2106dcd0_568);
and ( n13424 , n13423 , n13145 );
buf ( n13425 , RI21072e60_547);
and ( n13426 , n13425 , n13148 );
or ( n13427 , n13420 , n13422 , n13424 , n13426 );
buf ( n13428 , n13427 );
not ( n13429 , n13428 );
xnor ( n13430 , n12907 , n12922 );
buf ( n13431 , n13430 );
and ( n13432 , n13431 , n13138 );
buf ( n13433 , RI2106cb00_593);
and ( n13434 , n13433 , n13142 );
buf ( n13435 , RI2106b2a0_619);
and ( n13436 , n13435 , n13145 );
buf ( n13437 , RI21072ed8_546);
and ( n13438 , n13437 , n13148 );
or ( n13439 , n13432 , n13434 , n13436 , n13438 );
buf ( n13440 , n13439 );
not ( n13441 , n13440 );
xnor ( n13442 , n12914 , n12921 );
buf ( n13443 , n13442 );
and ( n13444 , n13443 , n13138 );
buf ( n13445 , RI2106afd0_625);
and ( n13446 , n13445 , n13142 );
buf ( n13447 , RI2106b318_618);
and ( n13448 , n13447 , n13145 );
buf ( n13449 , RI21072f50_545);
and ( n13450 , n13449 , n13148 );
or ( n13451 , n13444 , n13446 , n13448 , n13450 );
buf ( n13452 , n13451 );
not ( n13453 , n13452 );
not ( n13454 , n12921 );
buf ( n13455 , n13454 );
and ( n13456 , n13455 , n13138 );
buf ( n13457 , RI2106cb78_592);
and ( n13458 , n13457 , n13142 );
buf ( n13459 , RI2106b390_617);
and ( n13460 , n13459 , n13145 );
buf ( n13461 , RI21072fc8_544);
and ( n13462 , n13461 , n13148 );
or ( n13463 , n13456 , n13458 , n13460 , n13462 );
buf ( n13464 , n13463 );
not ( n13465 , n13464 );
not ( n13466 , n12735 );
and ( n13467 , n13466 , n12656 );
xor ( n13468 , n12657 , n12676 );
and ( n13469 , n13468 , n12735 );
or ( n13470 , n13467 , n13469 );
buf ( n13471 , n13470 );
buf ( n13472 , n13471 );
and ( n13473 , n13472 , n13138 );
buf ( n13474 , RI2106b048_624);
and ( n13475 , n13474 , n13142 );
buf ( n13476 , RI2106b408_616);
and ( n13477 , n13476 , n13145 );
buf ( n13478 , RI21073b80_541);
and ( n13479 , n13478 , n13148 );
or ( n13480 , n13473 , n13475 , n13477 , n13479 );
buf ( n13481 , n13480 );
not ( n13482 , n13481 );
not ( n13483 , n12735 );
and ( n13484 , n13483 , n12667 );
xor ( n13485 , n12668 , n12675 );
and ( n13486 , n13485 , n12735 );
or ( n13487 , n13484 , n13486 );
buf ( n13488 , n13487 );
buf ( n13489 , n13488 );
and ( n13490 , n13489 , n13138 );
buf ( n13491 , RI2106b0c0_623);
and ( n13492 , n13491 , n13142 );
buf ( n13493 , RI2106b480_615);
and ( n13494 , n13493 , n13145 );
buf ( n13495 , RI21074af8_530);
and ( n13496 , n13495 , n13148 );
or ( n13497 , n13490 , n13492 , n13494 , n13496 );
buf ( n13498 , n13497 );
not ( n13499 , n13498 );
not ( n13500 , n12735 );
and ( n13501 , n13500 , n12673 );
xor ( n13502 , n12674 , n12246 );
and ( n13503 , n13502 , n12735 );
or ( n13504 , n13501 , n13503 );
buf ( n13505 , n13504 );
buf ( n13506 , n13505 );
and ( n13507 , n13506 , n13138 );
buf ( n13508 , RI2106daf0_572);
and ( n13509 , n13508 , n13142 );
buf ( n13510 , RI21072230_551);
and ( n13511 , n13510 , n13145 );
buf ( n13512 , RI210764c0_519);
and ( n13513 , n13512 , n13148 );
or ( n13514 , n13507 , n13509 , n13511 , n13513 );
buf ( n13515 , n13514 );
not ( n13516 , n13515 );
and ( n13517 , n13499 , n13516 );
and ( n13518 , n13482 , n13517 );
and ( n13519 , n13465 , n13518 );
and ( n13520 , n13453 , n13519 );
and ( n13521 , n13441 , n13520 );
and ( n13522 , n13429 , n13521 );
and ( n13523 , n13417 , n13522 );
and ( n13524 , n13405 , n13523 );
and ( n13525 , n13393 , n13524 );
and ( n13526 , n13381 , n13525 );
and ( n13527 , n13369 , n13526 );
and ( n13528 , n13357 , n13527 );
and ( n13529 , n13345 , n13528 );
and ( n13530 , n13333 , n13529 );
and ( n13531 , n13321 , n13530 );
and ( n13532 , n13309 , n13531 );
and ( n13533 , n13297 , n13532 );
and ( n13534 , n13285 , n13533 );
and ( n13535 , n13273 , n13534 );
and ( n13536 , n13261 , n13535 );
and ( n13537 , n13249 , n13536 );
and ( n13538 , n13237 , n13537 );
and ( n13539 , n13225 , n13538 );
and ( n13540 , n13213 , n13539 );
and ( n13541 , n13201 , n13540 );
and ( n13542 , n13189 , n13541 );
and ( n13543 , n13177 , n13542 );
xor ( n13544 , n13165 , n13543 );
and ( n13545 , n13544 , n13151 );
or ( n13546 , n13164 , n13545 );
buf ( n13547 , n13546 );
not ( n13548 , n13547 );
buf ( n13549 , n13548 );
buf ( n13550 , n13549 );
not ( n13551 , n13550 );
xor ( n13552 , n13551 , n13151 );
not ( n13553 , n13151 );
and ( n13554 , n13553 , n13176 );
xor ( n13555 , n13177 , n13542 );
and ( n13556 , n13555 , n13151 );
or ( n13557 , n13554 , n13556 );
buf ( n13558 , n13557 );
not ( n13559 , n13558 );
buf ( n13560 , n13559 );
buf ( n13561 , n13560 );
not ( n13562 , n13561 );
xor ( n13563 , n13562 , n13151 );
not ( n13564 , n13151 );
and ( n13565 , n13564 , n13188 );
xor ( n13566 , n13189 , n13541 );
and ( n13567 , n13566 , n13151 );
or ( n13568 , n13565 , n13567 );
buf ( n13569 , n13568 );
not ( n13570 , n13569 );
buf ( n13571 , n13570 );
buf ( n13572 , n13571 );
not ( n13573 , n13572 );
xor ( n13574 , n13573 , n13151 );
not ( n13575 , n13151 );
and ( n13576 , n13575 , n13200 );
xor ( n13577 , n13201 , n13540 );
and ( n13578 , n13577 , n13151 );
or ( n13579 , n13576 , n13578 );
buf ( n13580 , n13579 );
not ( n13581 , n13580 );
buf ( n13582 , n13581 );
buf ( n13583 , n13582 );
not ( n13584 , n13583 );
xor ( n13585 , n13584 , n13151 );
not ( n13586 , n13151 );
and ( n13587 , n13586 , n13212 );
xor ( n13588 , n13213 , n13539 );
and ( n13589 , n13588 , n13151 );
or ( n13590 , n13587 , n13589 );
buf ( n13591 , n13590 );
not ( n13592 , n13591 );
buf ( n13593 , n13592 );
buf ( n13594 , n13593 );
not ( n13595 , n13594 );
xor ( n13596 , n13595 , n13151 );
not ( n13597 , n13151 );
and ( n13598 , n13597 , n13224 );
xor ( n13599 , n13225 , n13538 );
and ( n13600 , n13599 , n13151 );
or ( n13601 , n13598 , n13600 );
buf ( n13602 , n13601 );
not ( n13603 , n13602 );
buf ( n13604 , n13603 );
buf ( n13605 , n13604 );
not ( n13606 , n13605 );
xor ( n13607 , n13606 , n13151 );
not ( n13608 , n13151 );
and ( n13609 , n13608 , n13236 );
xor ( n13610 , n13237 , n13537 );
and ( n13611 , n13610 , n13151 );
or ( n13612 , n13609 , n13611 );
buf ( n13613 , n13612 );
not ( n13614 , n13613 );
buf ( n13615 , n13614 );
buf ( n13616 , n13615 );
not ( n13617 , n13616 );
xor ( n13618 , n13617 , n13151 );
not ( n13619 , n13151 );
and ( n13620 , n13619 , n13248 );
xor ( n13621 , n13249 , n13536 );
and ( n13622 , n13621 , n13151 );
or ( n13623 , n13620 , n13622 );
buf ( n13624 , n13623 );
not ( n13625 , n13624 );
buf ( n13626 , n13625 );
buf ( n13627 , n13626 );
not ( n13628 , n13627 );
xor ( n13629 , n13628 , n13151 );
not ( n13630 , n13151 );
and ( n13631 , n13630 , n13260 );
xor ( n13632 , n13261 , n13535 );
and ( n13633 , n13632 , n13151 );
or ( n13634 , n13631 , n13633 );
buf ( n13635 , n13634 );
not ( n13636 , n13635 );
buf ( n13637 , n13636 );
buf ( n13638 , n13637 );
not ( n13639 , n13638 );
xor ( n13640 , n13639 , n13151 );
not ( n13641 , n13151 );
and ( n13642 , n13641 , n13272 );
xor ( n13643 , n13273 , n13534 );
and ( n13644 , n13643 , n13151 );
or ( n13645 , n13642 , n13644 );
buf ( n13646 , n13645 );
not ( n13647 , n13646 );
buf ( n13648 , n13647 );
buf ( n13649 , n13648 );
not ( n13650 , n13649 );
xor ( n13651 , n13650 , n13151 );
not ( n13652 , n13151 );
and ( n13653 , n13652 , n13284 );
xor ( n13654 , n13285 , n13533 );
and ( n13655 , n13654 , n13151 );
or ( n13656 , n13653 , n13655 );
buf ( n13657 , n13656 );
not ( n13658 , n13657 );
buf ( n13659 , n13658 );
buf ( n13660 , n13659 );
not ( n13661 , n13660 );
xor ( n13662 , n13661 , n13151 );
not ( n13663 , n13151 );
and ( n13664 , n13663 , n13296 );
xor ( n13665 , n13297 , n13532 );
and ( n13666 , n13665 , n13151 );
or ( n13667 , n13664 , n13666 );
buf ( n13668 , n13667 );
not ( n13669 , n13668 );
buf ( n13670 , n13669 );
buf ( n13671 , n13670 );
not ( n13672 , n13671 );
xor ( n13673 , n13672 , n13151 );
not ( n13674 , n13151 );
and ( n13675 , n13674 , n13308 );
xor ( n13676 , n13309 , n13531 );
and ( n13677 , n13676 , n13151 );
or ( n13678 , n13675 , n13677 );
buf ( n13679 , n13678 );
not ( n13680 , n13679 );
buf ( n13681 , n13680 );
buf ( n13682 , n13681 );
not ( n13683 , n13682 );
xor ( n13684 , n13683 , n13151 );
not ( n13685 , n13151 );
and ( n13686 , n13685 , n13320 );
xor ( n13687 , n13321 , n13530 );
and ( n13688 , n13687 , n13151 );
or ( n13689 , n13686 , n13688 );
buf ( n13690 , n13689 );
not ( n13691 , n13690 );
buf ( n13692 , n13691 );
buf ( n13693 , n13692 );
not ( n13694 , n13693 );
xor ( n13695 , n13694 , n13151 );
not ( n13696 , n13151 );
and ( n13697 , n13696 , n13332 );
xor ( n13698 , n13333 , n13529 );
and ( n13699 , n13698 , n13151 );
or ( n13700 , n13697 , n13699 );
buf ( n13701 , n13700 );
not ( n13702 , n13701 );
buf ( n13703 , n13702 );
buf ( n13704 , n13703 );
not ( n13705 , n13704 );
xor ( n13706 , n13705 , n13151 );
not ( n13707 , n13151 );
and ( n13708 , n13707 , n13344 );
xor ( n13709 , n13345 , n13528 );
and ( n13710 , n13709 , n13151 );
or ( n13711 , n13708 , n13710 );
buf ( n13712 , n13711 );
not ( n13713 , n13712 );
buf ( n13714 , n13713 );
buf ( n13715 , n13714 );
not ( n13716 , n13715 );
xor ( n13717 , n13716 , n13151 );
not ( n13718 , n13151 );
and ( n13719 , n13718 , n13356 );
xor ( n13720 , n13357 , n13527 );
and ( n13721 , n13720 , n13151 );
or ( n13722 , n13719 , n13721 );
buf ( n13723 , n13722 );
not ( n13724 , n13723 );
buf ( n13725 , n13724 );
buf ( n13726 , n13725 );
not ( n13727 , n13726 );
xor ( n13728 , n13727 , n13151 );
not ( n13729 , n13151 );
and ( n13730 , n13729 , n13368 );
xor ( n13731 , n13369 , n13526 );
and ( n13732 , n13731 , n13151 );
or ( n13733 , n13730 , n13732 );
buf ( n13734 , n13733 );
not ( n13735 , n13734 );
buf ( n13736 , n13735 );
buf ( n13737 , n13736 );
not ( n13738 , n13737 );
xor ( n13739 , n13738 , n13151 );
not ( n13740 , n13151 );
and ( n13741 , n13740 , n13380 );
xor ( n13742 , n13381 , n13525 );
and ( n13743 , n13742 , n13151 );
or ( n13744 , n13741 , n13743 );
buf ( n13745 , n13744 );
not ( n13746 , n13745 );
buf ( n13747 , n13746 );
buf ( n13748 , n13747 );
not ( n13749 , n13748 );
xor ( n13750 , n13749 , n13151 );
not ( n13751 , n13151 );
and ( n13752 , n13751 , n13392 );
xor ( n13753 , n13393 , n13524 );
and ( n13754 , n13753 , n13151 );
or ( n13755 , n13752 , n13754 );
buf ( n13756 , n13755 );
not ( n13757 , n13756 );
buf ( n13758 , n13757 );
buf ( n13759 , n13758 );
not ( n13760 , n13759 );
xor ( n13761 , n13760 , n13151 );
not ( n13762 , n13151 );
and ( n13763 , n13762 , n13404 );
xor ( n13764 , n13405 , n13523 );
and ( n13765 , n13764 , n13151 );
or ( n13766 , n13763 , n13765 );
buf ( n13767 , n13766 );
not ( n13768 , n13767 );
buf ( n13769 , n13768 );
buf ( n13770 , n13769 );
not ( n13771 , n13770 );
xor ( n13772 , n13771 , n13151 );
not ( n13773 , n13151 );
and ( n13774 , n13773 , n13416 );
xor ( n13775 , n13417 , n13522 );
and ( n13776 , n13775 , n13151 );
or ( n13777 , n13774 , n13776 );
buf ( n13778 , n13777 );
not ( n13779 , n13778 );
buf ( n13780 , n13779 );
buf ( n13781 , n13780 );
not ( n13782 , n13781 );
xor ( n13783 , n13782 , n13151 );
not ( n13784 , n13151 );
and ( n13785 , n13784 , n13428 );
xor ( n13786 , n13429 , n13521 );
and ( n13787 , n13786 , n13151 );
or ( n13788 , n13785 , n13787 );
buf ( n13789 , n13788 );
not ( n13790 , n13789 );
buf ( n13791 , n13790 );
buf ( n13792 , n13791 );
not ( n13793 , n13792 );
xor ( n13794 , n13793 , n13151 );
not ( n13795 , n13151 );
and ( n13796 , n13795 , n13440 );
xor ( n13797 , n13441 , n13520 );
and ( n13798 , n13797 , n13151 );
or ( n13799 , n13796 , n13798 );
buf ( n13800 , n13799 );
not ( n13801 , n13800 );
buf ( n13802 , n13801 );
buf ( n13803 , n13802 );
not ( n13804 , n13803 );
xor ( n13805 , n13804 , n13151 );
not ( n13806 , n13151 );
and ( n13807 , n13806 , n13452 );
xor ( n13808 , n13453 , n13519 );
and ( n13809 , n13808 , n13151 );
or ( n13810 , n13807 , n13809 );
buf ( n13811 , n13810 );
not ( n13812 , n13811 );
buf ( n13813 , n13812 );
buf ( n13814 , n13813 );
not ( n13815 , n13814 );
xor ( n13816 , n13815 , n13151 );
not ( n13817 , n13151 );
and ( n13818 , n13817 , n13464 );
xor ( n13819 , n13465 , n13518 );
and ( n13820 , n13819 , n13151 );
or ( n13821 , n13818 , n13820 );
buf ( n13822 , n13821 );
not ( n13823 , n13822 );
buf ( n13824 , n13823 );
buf ( n13825 , n13824 );
not ( n13826 , n13825 );
xor ( n13827 , n13826 , n13151 );
not ( n13828 , n13151 );
and ( n13829 , n13828 , n13481 );
xor ( n13830 , n13482 , n13517 );
and ( n13831 , n13830 , n13151 );
or ( n13832 , n13829 , n13831 );
buf ( n13833 , n13832 );
not ( n13834 , n13833 );
buf ( n13835 , n13834 );
buf ( n13836 , n13835 );
not ( n13837 , n13836 );
xor ( n13838 , n13837 , n13151 );
not ( n13839 , n13151 );
and ( n13840 , n13839 , n13498 );
xor ( n13841 , n13499 , n13516 );
and ( n13842 , n13841 , n13151 );
or ( n13843 , n13840 , n13842 );
buf ( n13844 , n13843 );
not ( n13845 , n13844 );
buf ( n13846 , n13845 );
buf ( n13847 , n13846 );
not ( n13848 , n13847 );
xor ( n13849 , n13848 , n13151 );
buf ( n13850 , n13515 );
not ( n13851 , n13850 );
buf ( n13852 , n13851 );
buf ( n13853 , n13852 );
not ( n13854 , n13853 );
xor ( n13855 , n13854 , n13151 );
and ( n13856 , n13855 , n13151 );
and ( n13857 , n13849 , n13856 );
and ( n13858 , n13838 , n13857 );
and ( n13859 , n13827 , n13858 );
and ( n13860 , n13816 , n13859 );
and ( n13861 , n13805 , n13860 );
and ( n13862 , n13794 , n13861 );
and ( n13863 , n13783 , n13862 );
and ( n13864 , n13772 , n13863 );
and ( n13865 , n13761 , n13864 );
and ( n13866 , n13750 , n13865 );
and ( n13867 , n13739 , n13866 );
and ( n13868 , n13728 , n13867 );
and ( n13869 , n13717 , n13868 );
and ( n13870 , n13706 , n13869 );
and ( n13871 , n13695 , n13870 );
and ( n13872 , n13684 , n13871 );
and ( n13873 , n13673 , n13872 );
and ( n13874 , n13662 , n13873 );
and ( n13875 , n13651 , n13874 );
and ( n13876 , n13640 , n13875 );
and ( n13877 , n13629 , n13876 );
and ( n13878 , n13618 , n13877 );
and ( n13879 , n13607 , n13878 );
and ( n13880 , n13596 , n13879 );
and ( n13881 , n13585 , n13880 );
and ( n13882 , n13574 , n13881 );
and ( n13883 , n13563 , n13882 );
and ( n13884 , n13552 , n13883 );
buf ( n13885 , n13884 );
or ( n13886 , n13854 , n13848 );
or ( n13887 , n13886 , n13837 );
or ( n13888 , n13887 , n13826 );
or ( n13889 , n13888 , n13815 );
or ( n13890 , n13889 , n13804 );
or ( n13891 , n13890 , n13793 );
or ( n13892 , n13891 , n13782 );
or ( n13893 , n13892 , n13771 );
or ( n13894 , n13893 , n13760 );
or ( n13895 , n13894 , n13749 );
or ( n13896 , n13895 , n13738 );
or ( n13897 , n13896 , n13727 );
or ( n13898 , n13897 , n13716 );
or ( n13899 , n13898 , n13705 );
or ( n13900 , n13899 , n13694 );
or ( n13901 , n13900 , n13683 );
or ( n13902 , n13901 , n13672 );
or ( n13903 , n13902 , n13661 );
or ( n13904 , n13903 , n13650 );
or ( n13905 , n13904 , n13639 );
or ( n13906 , n13905 , n13628 );
or ( n13907 , n13906 , n13617 );
or ( n13908 , n13907 , n13606 );
or ( n13909 , n13908 , n13595 );
or ( n13910 , n13909 , n13584 );
or ( n13911 , n13910 , n13573 );
or ( n13912 , n13911 , n13562 );
or ( n13913 , n13912 , n13551 );
buf ( n13914 , n13913 );
buf ( n13915 , n13914 );
and ( n13916 , n13915 , n13151 );
and ( n13917 , n13885 , n13916 );
or ( n13918 , C0 , n13917 );
buf ( n13919 , n13918 );
buf ( n13920 , n13919 );
buf ( n13921 , n11504 );
not ( n13922 , n13921 );
buf ( n13923 , n11792 );
and ( n13924 , n13922 , n13923 );
not ( n13925 , n13923 );
buf ( n13926 , n11800 );
not ( n13927 , n13926 );
buf ( n13928 , n11808 );
not ( n13929 , n13928 );
buf ( n13930 , n11816 );
not ( n13931 , n13930 );
buf ( n13932 , n11512 );
not ( n13933 , n13932 );
buf ( n13934 , n11521 );
not ( n13935 , n13934 );
buf ( n13936 , n11529 );
not ( n13937 , n13936 );
buf ( n13938 , n11537 );
not ( n13939 , n13938 );
buf ( n13940 , n11545 );
not ( n13941 , n13940 );
buf ( n13942 , n11553 );
not ( n13943 , n13942 );
buf ( n13944 , n11561 );
not ( n13945 , n13944 );
buf ( n13946 , n11569 );
not ( n13947 , n13946 );
buf ( n13948 , n11577 );
not ( n13949 , n13948 );
buf ( n13950 , n11585 );
not ( n13951 , n13950 );
buf ( n13952 , n11593 );
not ( n13953 , n13952 );
buf ( n13954 , n11601 );
not ( n13955 , n13954 );
buf ( n13956 , n11609 );
not ( n13957 , n13956 );
buf ( n13958 , n11617 );
not ( n13959 , n13958 );
buf ( n13960 , n11625 );
not ( n13961 , n13960 );
buf ( n13962 , n11633 );
not ( n13963 , n13962 );
buf ( n13964 , n11641 );
not ( n13965 , n13964 );
buf ( n13966 , n11649 );
not ( n13967 , n13966 );
buf ( n13968 , n11657 );
not ( n13969 , n13968 );
buf ( n13970 , n11665 );
not ( n13971 , n13970 );
buf ( n13972 , n11673 );
not ( n13973 , n13972 );
buf ( n13974 , n11681 );
not ( n13975 , n13974 );
buf ( n13976 , n11689 );
not ( n13977 , n13976 );
buf ( n13978 , n11692 );
not ( n13979 , n13978 );
and ( n13980 , n13977 , n13979 );
and ( n13981 , n13975 , n13980 );
and ( n13982 , n13973 , n13981 );
and ( n13983 , n13971 , n13982 );
and ( n13984 , n13969 , n13983 );
and ( n13985 , n13967 , n13984 );
and ( n13986 , n13965 , n13985 );
and ( n13987 , n13963 , n13986 );
and ( n13988 , n13961 , n13987 );
and ( n13989 , n13959 , n13988 );
and ( n13990 , n13957 , n13989 );
and ( n13991 , n13955 , n13990 );
and ( n13992 , n13953 , n13991 );
and ( n13993 , n13951 , n13992 );
and ( n13994 , n13949 , n13993 );
and ( n13995 , n13947 , n13994 );
and ( n13996 , n13945 , n13995 );
and ( n13997 , n13943 , n13996 );
and ( n13998 , n13941 , n13997 );
and ( n13999 , n13939 , n13998 );
and ( n14000 , n13937 , n13999 );
and ( n14001 , n13935 , n14000 );
and ( n14002 , n13933 , n14001 );
and ( n14003 , n13931 , n14002 );
and ( n14004 , n13929 , n14003 );
and ( n14005 , n13927 , n14004 );
xor ( n14006 , n13925 , n14005 );
and ( n14007 , n14006 , n13921 );
or ( n14008 , n13924 , n14007 );
buf ( n14009 , n14008 );
not ( n14010 , n14009 );
buf ( n14011 , n14010 );
buf ( n14012 , n14011 );
not ( n14013 , n14012 );
buf ( n14014 , n14013 );
buf ( n14015 , n14014 );
buf ( n14016 , n14015 );
not ( n14017 , n14016 );
buf ( n14018 , n14017 );
buf ( n14019 , n14018 );
not ( n14020 , n14019 );
not ( n14021 , n13921 );
buf ( n14022 , n11768 );
not ( n14023 , n14022 );
buf ( n14024 , n11776 );
not ( n14025 , n14024 );
buf ( n14026 , n11784 );
not ( n14027 , n14026 );
and ( n14028 , n13925 , n14005 );
and ( n14029 , n14027 , n14028 );
and ( n14030 , n14025 , n14029 );
and ( n14031 , n14023 , n14030 );
xor ( n14032 , n14021 , n14031 );
buf ( n14033 , n13921 );
and ( n14034 , n14032 , n14033 );
or ( n14035 , C0 , n14034 );
buf ( n14036 , n14035 );
not ( n14037 , n14036 );
buf ( n14038 , n14037 );
buf ( n14039 , n14038 );
not ( n14040 , n14039 );
buf ( n14041 , n14040 );
not ( n14042 , n14041 );
buf ( n14043 , n14042 );
not ( n14044 , n13921 );
and ( n14045 , n14044 , n14022 );
xor ( n14046 , n14023 , n14030 );
and ( n14047 , n14046 , n13921 );
or ( n14048 , n14045 , n14047 );
buf ( n14049 , n14048 );
not ( n14050 , n14049 );
buf ( n14051 , n14050 );
buf ( n14052 , n14051 );
not ( n14053 , n14052 );
buf ( n14054 , n14053 );
not ( n14055 , n14054 );
buf ( n14056 , n14055 );
not ( n14057 , n13921 );
and ( n14058 , n14057 , n14024 );
xor ( n14059 , n14025 , n14029 );
and ( n14060 , n14059 , n13921 );
or ( n14061 , n14058 , n14060 );
buf ( n14062 , n14061 );
not ( n14063 , n14062 );
buf ( n14064 , n14063 );
buf ( n14065 , n14064 );
not ( n14066 , n14065 );
buf ( n14067 , n14066 );
not ( n14068 , n14067 );
buf ( n14069 , n14068 );
not ( n14070 , n13921 );
and ( n14071 , n14070 , n14026 );
xor ( n14072 , n14027 , n14028 );
and ( n14073 , n14072 , n13921 );
or ( n14074 , n14071 , n14073 );
buf ( n14075 , n14074 );
not ( n14076 , n14075 );
buf ( n14077 , n14076 );
buf ( n14078 , n14077 );
not ( n14079 , n14078 );
buf ( n14080 , n14079 );
not ( n14081 , n14080 );
buf ( n14082 , n14081 );
not ( n14083 , n14014 );
buf ( n14084 , n14083 );
and ( n14085 , n14082 , n14084 );
and ( n14086 , n14069 , n14085 );
and ( n14087 , n14056 , n14086 );
and ( n14088 , n14043 , n14087 );
not ( n14089 , n14088 );
buf ( n14090 , n14089 );
buf ( n14091 , n13921 );
and ( n14092 , n14090 , n14091 );
or ( n14093 , C0 , n14092 );
buf ( n14094 , n14093 );
buf ( n14095 , n14094 );
not ( n14096 , n14095 );
not ( n14097 , n14091 );
buf ( n14098 , n14080 );
and ( n14099 , n14097 , n14098 );
xor ( n14100 , n14082 , n14084 );
buf ( n14101 , n14100 );
and ( n14102 , n14101 , n14091 );
or ( n14103 , n14099 , n14102 );
buf ( n14104 , n14103 );
buf ( n14105 , n14104 );
and ( n14106 , n14096 , n14105 );
not ( n14107 , n14105 );
not ( n14108 , n14015 );
xor ( n14109 , n14107 , n14108 );
and ( n14110 , n14109 , n14095 );
or ( n14111 , n14106 , n14110 );
buf ( n14112 , n14111 );
not ( n14113 , n14112 );
buf ( n14114 , n14113 );
buf ( n14115 , n14114 );
not ( n14116 , n14115 );
or ( n14117 , n14020 , n14116 );
buf ( n14118 , n14117 );
buf ( n14119 , n14118 );
and ( n14120 , n14119 , n14095 );
not ( n14121 , n14120 );
and ( n14122 , n14121 , n14020 );
xor ( n14123 , n14020 , n14095 );
xor ( n14124 , n14123 , n14095 );
and ( n14125 , n14124 , n14120 );
or ( n14126 , n14122 , n14125 );
buf ( n14127 , n14126 );
not ( n14128 , n14127 );
not ( n14129 , n14120 );
and ( n14130 , n14129 , n14116 );
xor ( n14131 , n14116 , n14095 );
and ( n14132 , n14123 , n14095 );
xor ( n14133 , n14131 , n14132 );
and ( n14134 , n14133 , n14120 );
or ( n14135 , n14130 , n14134 );
buf ( n14136 , n14135 );
and ( n14137 , n14128 , n14136 );
and ( n14138 , n13920 , n14137 );
buf ( n14139 , RI2107dae0_465);
and ( n14140 , n14127 , n14136 );
nor ( n14141 , n14127 , n14136 );
or ( n14142 , n14140 , n14141 );
nor ( n14143 , n14128 , n14136 );
or ( n14144 , n14142 , n14143 );
and ( n14145 , n14139 , n14144 );
or ( n14146 , n14138 , n14145 );
buf ( n14147 , n11504 );
not ( n14148 , n14147 );
buf ( n14149 , n11545 );
and ( n14150 , n14148 , n14149 );
not ( n14151 , n14149 );
buf ( n14152 , n11553 );
not ( n14153 , n14152 );
buf ( n14154 , n11561 );
not ( n14155 , n14154 );
buf ( n14156 , n11569 );
not ( n14157 , n14156 );
buf ( n14158 , n11577 );
not ( n14159 , n14158 );
buf ( n14160 , n11585 );
not ( n14161 , n14160 );
buf ( n14162 , n11593 );
not ( n14163 , n14162 );
buf ( n14164 , n11601 );
not ( n14165 , n14164 );
buf ( n14166 , n11609 );
not ( n14167 , n14166 );
buf ( n14168 , n11617 );
not ( n14169 , n14168 );
buf ( n14170 , n11625 );
not ( n14171 , n14170 );
buf ( n14172 , n11633 );
not ( n14173 , n14172 );
buf ( n14174 , n11641 );
not ( n14175 , n14174 );
buf ( n14176 , n11649 );
not ( n14177 , n14176 );
buf ( n14178 , n11657 );
not ( n14179 , n14178 );
buf ( n14180 , n11665 );
not ( n14181 , n14180 );
buf ( n14182 , n11673 );
not ( n14183 , n14182 );
buf ( n14184 , n11681 );
not ( n14185 , n14184 );
buf ( n14186 , n11689 );
not ( n14187 , n14186 );
buf ( n14188 , n11692 );
not ( n14189 , n14188 );
and ( n14190 , n14187 , n14189 );
and ( n14191 , n14185 , n14190 );
and ( n14192 , n14183 , n14191 );
and ( n14193 , n14181 , n14192 );
and ( n14194 , n14179 , n14193 );
and ( n14195 , n14177 , n14194 );
and ( n14196 , n14175 , n14195 );
and ( n14197 , n14173 , n14196 );
and ( n14198 , n14171 , n14197 );
and ( n14199 , n14169 , n14198 );
and ( n14200 , n14167 , n14199 );
and ( n14201 , n14165 , n14200 );
and ( n14202 , n14163 , n14201 );
and ( n14203 , n14161 , n14202 );
and ( n14204 , n14159 , n14203 );
and ( n14205 , n14157 , n14204 );
and ( n14206 , n14155 , n14205 );
and ( n14207 , n14153 , n14206 );
xor ( n14208 , n14151 , n14207 );
and ( n14209 , n14208 , n14147 );
or ( n14210 , n14150 , n14209 );
buf ( n14211 , n14210 );
not ( n14212 , n14211 );
buf ( n14213 , n14212 );
buf ( n14214 , n14213 );
not ( n14215 , n14214 );
buf ( n14216 , n14215 );
buf ( n14217 , n14216 );
buf ( n14218 , n14217 );
not ( n14219 , n14218 );
buf ( n14220 , n14219 );
buf ( n14221 , n14220 );
not ( n14222 , n14221 );
not ( n14223 , n14147 );
buf ( n14224 , n11768 );
not ( n14225 , n14224 );
buf ( n14226 , n11776 );
not ( n14227 , n14226 );
buf ( n14228 , n11784 );
not ( n14229 , n14228 );
buf ( n14230 , n11792 );
not ( n14231 , n14230 );
buf ( n14232 , n11800 );
not ( n14233 , n14232 );
buf ( n14234 , n11808 );
not ( n14235 , n14234 );
buf ( n14236 , n11816 );
not ( n14237 , n14236 );
buf ( n14238 , n11512 );
not ( n14239 , n14238 );
buf ( n14240 , n11521 );
not ( n14241 , n14240 );
buf ( n14242 , n11529 );
not ( n14243 , n14242 );
buf ( n14244 , n11537 );
not ( n14245 , n14244 );
and ( n14246 , n14151 , n14207 );
and ( n14247 , n14245 , n14246 );
and ( n14248 , n14243 , n14247 );
and ( n14249 , n14241 , n14248 );
and ( n14250 , n14239 , n14249 );
and ( n14251 , n14237 , n14250 );
and ( n14252 , n14235 , n14251 );
and ( n14253 , n14233 , n14252 );
and ( n14254 , n14231 , n14253 );
and ( n14255 , n14229 , n14254 );
and ( n14256 , n14227 , n14255 );
and ( n14257 , n14225 , n14256 );
xor ( n14258 , n14223 , n14257 );
buf ( n14259 , n14147 );
and ( n14260 , n14258 , n14259 );
or ( n14261 , C0 , n14260 );
buf ( n14262 , n14261 );
not ( n14263 , n14262 );
buf ( n14264 , n14263 );
buf ( n14265 , n14264 );
not ( n14266 , n14265 );
buf ( n14267 , n14266 );
not ( n14268 , n14267 );
buf ( n14269 , n14268 );
not ( n14270 , n14147 );
and ( n14271 , n14270 , n14224 );
xor ( n14272 , n14225 , n14256 );
and ( n14273 , n14272 , n14147 );
or ( n14274 , n14271 , n14273 );
buf ( n14275 , n14274 );
not ( n14276 , n14275 );
buf ( n14277 , n14276 );
buf ( n14278 , n14277 );
not ( n14279 , n14278 );
buf ( n14280 , n14279 );
not ( n14281 , n14280 );
buf ( n14282 , n14281 );
not ( n14283 , n14147 );
and ( n14284 , n14283 , n14226 );
xor ( n14285 , n14227 , n14255 );
and ( n14286 , n14285 , n14147 );
or ( n14287 , n14284 , n14286 );
buf ( n14288 , n14287 );
not ( n14289 , n14288 );
buf ( n14290 , n14289 );
buf ( n14291 , n14290 );
not ( n14292 , n14291 );
buf ( n14293 , n14292 );
not ( n14294 , n14293 );
buf ( n14295 , n14294 );
not ( n14296 , n14147 );
and ( n14297 , n14296 , n14228 );
xor ( n14298 , n14229 , n14254 );
and ( n14299 , n14298 , n14147 );
or ( n14300 , n14297 , n14299 );
buf ( n14301 , n14300 );
not ( n14302 , n14301 );
buf ( n14303 , n14302 );
buf ( n14304 , n14303 );
not ( n14305 , n14304 );
buf ( n14306 , n14305 );
not ( n14307 , n14306 );
buf ( n14308 , n14307 );
not ( n14309 , n14147 );
and ( n14310 , n14309 , n14230 );
xor ( n14311 , n14231 , n14253 );
and ( n14312 , n14311 , n14147 );
or ( n14313 , n14310 , n14312 );
buf ( n14314 , n14313 );
not ( n14315 , n14314 );
buf ( n14316 , n14315 );
buf ( n14317 , n14316 );
not ( n14318 , n14317 );
buf ( n14319 , n14318 );
not ( n14320 , n14319 );
buf ( n14321 , n14320 );
not ( n14322 , n14147 );
and ( n14323 , n14322 , n14232 );
xor ( n14324 , n14233 , n14252 );
and ( n14325 , n14324 , n14147 );
or ( n14326 , n14323 , n14325 );
buf ( n14327 , n14326 );
not ( n14328 , n14327 );
buf ( n14329 , n14328 );
buf ( n14330 , n14329 );
not ( n14331 , n14330 );
buf ( n14332 , n14331 );
not ( n14333 , n14332 );
buf ( n14334 , n14333 );
not ( n14335 , n14147 );
and ( n14336 , n14335 , n14234 );
xor ( n14337 , n14235 , n14251 );
and ( n14338 , n14337 , n14147 );
or ( n14339 , n14336 , n14338 );
buf ( n14340 , n14339 );
not ( n14341 , n14340 );
buf ( n14342 , n14341 );
buf ( n14343 , n14342 );
not ( n14344 , n14343 );
buf ( n14345 , n14344 );
not ( n14346 , n14345 );
buf ( n14347 , n14346 );
not ( n14348 , n14147 );
and ( n14349 , n14348 , n14236 );
xor ( n14350 , n14237 , n14250 );
and ( n14351 , n14350 , n14147 );
or ( n14352 , n14349 , n14351 );
buf ( n14353 , n14352 );
not ( n14354 , n14353 );
buf ( n14355 , n14354 );
buf ( n14356 , n14355 );
not ( n14357 , n14356 );
buf ( n14358 , n14357 );
not ( n14359 , n14358 );
buf ( n14360 , n14359 );
not ( n14361 , n14147 );
and ( n14362 , n14361 , n14238 );
xor ( n14363 , n14239 , n14249 );
and ( n14364 , n14363 , n14147 );
or ( n14365 , n14362 , n14364 );
buf ( n14366 , n14365 );
not ( n14367 , n14366 );
buf ( n14368 , n14367 );
buf ( n14369 , n14368 );
not ( n14370 , n14369 );
buf ( n14371 , n14370 );
not ( n14372 , n14371 );
buf ( n14373 , n14372 );
not ( n14374 , n14147 );
and ( n14375 , n14374 , n14240 );
xor ( n14376 , n14241 , n14248 );
and ( n14377 , n14376 , n14147 );
or ( n14378 , n14375 , n14377 );
buf ( n14379 , n14378 );
not ( n14380 , n14379 );
buf ( n14381 , n14380 );
buf ( n14382 , n14381 );
not ( n14383 , n14382 );
buf ( n14384 , n14383 );
not ( n14385 , n14384 );
buf ( n14386 , n14385 );
not ( n14387 , n14147 );
and ( n14388 , n14387 , n14242 );
xor ( n14389 , n14243 , n14247 );
and ( n14390 , n14389 , n14147 );
or ( n14391 , n14388 , n14390 );
buf ( n14392 , n14391 );
not ( n14393 , n14392 );
buf ( n14394 , n14393 );
buf ( n14395 , n14394 );
not ( n14396 , n14395 );
buf ( n14397 , n14396 );
not ( n14398 , n14397 );
buf ( n14399 , n14398 );
not ( n14400 , n14147 );
and ( n14401 , n14400 , n14244 );
xor ( n14402 , n14245 , n14246 );
and ( n14403 , n14402 , n14147 );
or ( n14404 , n14401 , n14403 );
buf ( n14405 , n14404 );
not ( n14406 , n14405 );
buf ( n14407 , n14406 );
buf ( n14408 , n14407 );
not ( n14409 , n14408 );
buf ( n14410 , n14409 );
not ( n14411 , n14410 );
buf ( n14412 , n14411 );
not ( n14413 , n14216 );
buf ( n14414 , n14413 );
and ( n14415 , n14412 , n14414 );
and ( n14416 , n14399 , n14415 );
and ( n14417 , n14386 , n14416 );
and ( n14418 , n14373 , n14417 );
and ( n14419 , n14360 , n14418 );
and ( n14420 , n14347 , n14419 );
and ( n14421 , n14334 , n14420 );
and ( n14422 , n14321 , n14421 );
and ( n14423 , n14308 , n14422 );
and ( n14424 , n14295 , n14423 );
and ( n14425 , n14282 , n14424 );
and ( n14426 , n14269 , n14425 );
not ( n14427 , n14426 );
buf ( n14428 , n14427 );
buf ( n14429 , n14147 );
and ( n14430 , n14428 , n14429 );
or ( n14431 , C0 , n14430 );
buf ( n14432 , n14431 );
buf ( n14433 , n14432 );
not ( n14434 , n14433 );
not ( n14435 , n14429 );
buf ( n14436 , n14410 );
and ( n14437 , n14435 , n14436 );
xor ( n14438 , n14412 , n14414 );
buf ( n14439 , n14438 );
and ( n14440 , n14439 , n14429 );
or ( n14441 , n14437 , n14440 );
buf ( n14442 , n14441 );
buf ( n14443 , n14442 );
and ( n14444 , n14434 , n14443 );
not ( n14445 , n14443 );
not ( n14446 , n14217 );
xor ( n14447 , n14445 , n14446 );
and ( n14448 , n14447 , n14433 );
or ( n14449 , n14444 , n14448 );
buf ( n14450 , n14449 );
not ( n14451 , n14450 );
buf ( n14452 , n14451 );
buf ( n14453 , n14452 );
not ( n14454 , n14453 );
or ( n14455 , n14222 , n14454 );
not ( n14456 , n14433 );
not ( n14457 , n14429 );
buf ( n14458 , n14397 );
and ( n14459 , n14457 , n14458 );
xor ( n14460 , n14399 , n14415 );
buf ( n14461 , n14460 );
and ( n14462 , n14461 , n14429 );
or ( n14463 , n14459 , n14462 );
buf ( n14464 , n14463 );
buf ( n14465 , n14464 );
and ( n14466 , n14456 , n14465 );
not ( n14467 , n14465 );
and ( n14468 , n14445 , n14446 );
xor ( n14469 , n14467 , n14468 );
and ( n14470 , n14469 , n14433 );
or ( n14471 , n14466 , n14470 );
buf ( n14472 , n14471 );
not ( n14473 , n14472 );
buf ( n14474 , n14473 );
buf ( n14475 , n14474 );
not ( n14476 , n14475 );
or ( n14477 , n14455 , n14476 );
not ( n14478 , n14433 );
not ( n14479 , n14429 );
buf ( n14480 , n14384 );
and ( n14481 , n14479 , n14480 );
xor ( n14482 , n14386 , n14416 );
buf ( n14483 , n14482 );
and ( n14484 , n14483 , n14429 );
or ( n14485 , n14481 , n14484 );
buf ( n14486 , n14485 );
buf ( n14487 , n14486 );
and ( n14488 , n14478 , n14487 );
not ( n14489 , n14487 );
and ( n14490 , n14467 , n14468 );
xor ( n14491 , n14489 , n14490 );
and ( n14492 , n14491 , n14433 );
or ( n14493 , n14488 , n14492 );
buf ( n14494 , n14493 );
not ( n14495 , n14494 );
buf ( n14496 , n14495 );
buf ( n14497 , n14496 );
not ( n14498 , n14497 );
or ( n14499 , n14477 , n14498 );
or ( n14500 , n14499 , C0 );
or ( n14501 , n14500 , C0 );
or ( n14502 , n14501 , C0 );
or ( n14503 , n14502 , C0 );
or ( n14504 , n14503 , C0 );
or ( n14505 , n14504 , C0 );
or ( n14506 , n14505 , C0 );
or ( n14507 , n14506 , C0 );
or ( n14508 , n14507 , C0 );
or ( n14509 , n14508 , C0 );
or ( n14510 , n14509 , C0 );
or ( n14511 , n14510 , C0 );
or ( n14512 , n14511 , C0 );
or ( n14513 , n14512 , C0 );
or ( n14514 , n14513 , C0 );
or ( n14515 , n14514 , C0 );
or ( n14516 , n14515 , C0 );
or ( n14517 , n14516 , C0 );
or ( n14518 , n14517 , C0 );
or ( n14519 , n14518 , C0 );
or ( n14520 , n14519 , C0 );
or ( n14521 , n14520 , C0 );
or ( n14522 , n14521 , C0 );
or ( n14523 , n14522 , C0 );
or ( n14524 , n14523 , C0 );
or ( n14525 , n14524 , C0 );
or ( n14526 , n14525 , C0 );
buf ( n14527 , n14526 );
and ( n14528 , n14527 , n14433 );
not ( n14529 , n14528 );
and ( n14530 , n14529 , n14222 );
xor ( n14531 , n14222 , n14433 );
xor ( n14532 , n14531 , n14433 );
and ( n14533 , n14532 , n14528 );
or ( n14534 , n14530 , n14533 );
buf ( n14535 , n14534 );
not ( n14536 , n14535 );
not ( n14537 , n14528 );
and ( n14538 , n14537 , n14454 );
xor ( n14539 , n14454 , n14433 );
and ( n14540 , n14531 , n14433 );
xor ( n14541 , n14539 , n14540 );
and ( n14542 , n14541 , n14528 );
or ( n14543 , n14538 , n14542 );
buf ( n14544 , n14543 );
not ( n14545 , n14544 );
not ( n14546 , n14528 );
and ( n14547 , n14546 , n14476 );
xor ( n14548 , n14476 , n14433 );
and ( n14549 , n14539 , n14540 );
xor ( n14550 , n14548 , n14549 );
and ( n14551 , n14550 , n14528 );
or ( n14552 , n14547 , n14551 );
buf ( n14553 , n14552 );
not ( n14554 , n14528 );
and ( n14555 , n14554 , n14498 );
xor ( n14556 , n14498 , n14433 );
and ( n14557 , n14548 , n14549 );
xor ( n14558 , n14556 , n14557 );
and ( n14559 , n14558 , n14528 );
or ( n14560 , n14555 , n14559 );
buf ( n14561 , n14560 );
and ( n14562 , n14536 , n14545 , n14553 , n14561 );
and ( n14563 , n14146 , n14562 );
nor ( n14564 , n14536 , n14544 , n14553 , n14561 );
nor ( n14565 , n14535 , n14544 , n14553 , n14561 );
or ( n14566 , n14564 , n14565 );
nor ( n14567 , n14535 , n14545 , n14553 , n14561 );
or ( n14568 , n14566 , n14567 );
nor ( n14569 , n14536 , n14545 , n14553 , n14561 );
or ( n14570 , n14568 , n14569 );
not ( n14571 , n14561 );
and ( n14572 , n14536 , n14545 , n14553 , n14571 );
or ( n14573 , n14570 , n14572 );
and ( n14574 , n14535 , n14545 , n14553 , n14571 );
or ( n14575 , n14573 , n14574 );
and ( n14576 , n14536 , n14544 , n14553 , n14571 );
or ( n14577 , n14575 , n14576 );
and ( n14578 , n14535 , n14544 , n14553 , n14571 );
or ( n14579 , n14577 , n14578 );
nor ( n14580 , n14535 , n14544 , n14553 , n14571 );
or ( n14581 , n14579 , n14580 );
nor ( n14582 , n14536 , n14544 , n14553 , n14571 );
or ( n14583 , n14581 , n14582 );
nor ( n14584 , n14535 , n14545 , n14553 , n14571 );
or ( n14585 , n14583 , n14584 );
nor ( n14586 , n14536 , n14545 , n14553 , n14571 );
or ( n14587 , n14585 , n14586 );
and ( n14588 , n14535 , n14545 , n14553 , n14561 );
and ( n14589 , n14536 , n14544 , n14553 , n14561 );
or ( n14590 , n14588 , n14589 );
and ( n14591 , n14535 , n14544 , n14553 , n14561 );
or ( n14592 , n14590 , n14591 );
or ( n14593 , n14587 , n14592 );
and ( n14594 , n14139 , n14593 );
or ( n14595 , n14563 , n14594 );
and ( n14596 , n12244 , n14595 );
and ( n14597 , n14139 , n12243 );
or ( n14598 , n14596 , n14597 );
and ( n14599 , n11955 , n14598 );
buf ( n14600 , n13150 );
not ( n14601 , n14600 );
not ( n14602 , n12947 );
buf ( n14603 , n14602 );
and ( n14604 , n14603 , n13138 );
buf ( n14605 , RI2106cc68_590);
and ( n14606 , n14605 , n13142 );
buf ( n14607 , RI2106ddc0_566);
and ( n14608 , n14607 , n13145 );
buf ( n14609 , RI210730b8_542);
and ( n14610 , n14609 , n13148 );
or ( n14611 , n14604 , n14606 , n14608 , n14610 );
buf ( n14612 , n14611 );
and ( n14613 , n14601 , n14612 );
buf ( n14614 , n14613 );
not ( n14615 , n14614 );
and ( n14616 , n14615 , n13150 );
or ( n14617 , n14616 , C0 );
buf ( n14618 , n14617 );
buf ( n14619 , n10638 );
not ( n14620 , n14619 );
buf ( n14621 , n14620 );
buf ( n14622 , n10640 );
not ( n14623 , n14622 );
buf ( n14624 , n14623 );
and ( n14625 , n14621 , n14624 );
buf ( n14626 , n10797 );
and ( n14627 , n14625 , n14626 );
buf ( n14628 , RI21a0e608_121);
not ( n14629 , n14628 );
and ( n14630 , n14627 , n14629 );
buf ( n14631 , n10638 );
buf ( n14632 , n10640 );
and ( n14633 , n14631 , n14632 );
buf ( n14634 , n10797 );
not ( n14635 , n14634 );
buf ( n14636 , n14635 );
and ( n14637 , n14633 , n14636 );
buf ( n14638 , RI210b87a8_334);
not ( n14639 , n14638 );
and ( n14640 , n14637 , n14639 );
or ( n14641 , n14630 , n14640 );
not ( n14642 , n14641 );
buf ( n14643 , RI21a19a08_3);
and ( n14644 , n14642 , n14643 );
buf ( n14645 , RI21a0f058_113);
buf ( n14646 , n14645 );
buf ( n14647 , RI210b9b58_326);
buf ( n14648 , n14647 );
not ( n14649 , n14648 );
xor ( n14650 , n14646 , n14649 );
buf ( n14651 , RI21a0f0d0_112);
buf ( n14652 , n14651 );
buf ( n14653 , RI210b9bd0_325);
buf ( n14654 , n14653 );
not ( n14655 , n14654 );
and ( n14656 , n14652 , n14655 );
buf ( n14657 , RI21a0f850_110);
buf ( n14658 , n14657 );
buf ( n14659 , RI210b9c48_324);
buf ( n14660 , n14659 );
not ( n14661 , n14660 );
and ( n14662 , n14658 , n14661 );
buf ( n14663 , RI21a0f8c8_109);
buf ( n14664 , n14663 );
buf ( n14665 , RI210b9cc0_323);
buf ( n14666 , n14665 );
not ( n14667 , n14666 );
and ( n14668 , n14664 , n14667 );
buf ( n14669 , RI21a0f940_108);
buf ( n14670 , n14669 );
buf ( n14671 , RI210ba530_322);
buf ( n14672 , n14671 );
not ( n14673 , n14672 );
and ( n14674 , n14670 , n14673 );
buf ( n14675 , RI21a0f9b8_107);
buf ( n14676 , n14675 );
buf ( n14677 , RI210ba5a8_321);
buf ( n14678 , n14677 );
not ( n14679 , n14678 );
and ( n14680 , n14676 , n14679 );
buf ( n14681 , RI21a0fa30_106);
buf ( n14682 , n14681 );
buf ( n14683 , RI210ba620_320);
buf ( n14684 , n14683 );
not ( n14685 , n14684 );
and ( n14686 , n14682 , n14685 );
buf ( n14687 , RI21a0faa8_105);
buf ( n14688 , n14687 );
buf ( n14689 , RI210ba698_319);
buf ( n14690 , n14689 );
not ( n14691 , n14690 );
and ( n14692 , n14688 , n14691 );
buf ( n14693 , RI21a101b0_104);
buf ( n14694 , n14693 );
buf ( n14695 , RI210baf08_318);
buf ( n14696 , n14695 );
not ( n14697 , n14696 );
and ( n14698 , n14694 , n14697 );
buf ( n14699 , RI21a10228_103);
buf ( n14700 , n14699 );
buf ( n14701 , RI210baf80_317);
buf ( n14702 , n14701 );
not ( n14703 , n14702 );
and ( n14704 , n14700 , n14703 );
buf ( n14705 , RI21a102a0_102);
buf ( n14706 , n14705 );
buf ( n14707 , RI210baff8_316);
buf ( n14708 , n14707 );
not ( n14709 , n14708 );
and ( n14710 , n14706 , n14709 );
buf ( n14711 , RI21a10318_101);
buf ( n14712 , n14711 );
buf ( n14713 , RI210bb070_315);
buf ( n14714 , n14713 );
not ( n14715 , n14714 );
and ( n14716 , n14712 , n14715 );
buf ( n14717 , RI21a10390_100);
buf ( n14718 , n14717 );
buf ( n14719 , RI210bb8e0_314);
buf ( n14720 , n14719 );
not ( n14721 , n14720 );
and ( n14722 , n14718 , n14721 );
buf ( n14723 , RI21a10408_99);
buf ( n14724 , n14723 );
buf ( n14725 , RI210bb958_313);
buf ( n14726 , n14725 );
not ( n14727 , n14726 );
and ( n14728 , n14724 , n14727 );
buf ( n14729 , RI21a10b10_98);
buf ( n14730 , n14729 );
buf ( n14731 , RI210bb9d0_312);
buf ( n14732 , n14731 );
not ( n14733 , n14732 );
and ( n14734 , n14730 , n14733 );
buf ( n14735 , RI21a10b88_97);
buf ( n14736 , n14735 );
buf ( n14737 , RI210bba48_311);
buf ( n14738 , n14737 );
not ( n14739 , n14738 );
and ( n14740 , n14736 , n14739 );
buf ( n14741 , RI21a10c00_96);
buf ( n14742 , n14741 );
buf ( n14743 , RI210bc2b8_310);
buf ( n14744 , n14743 );
not ( n14745 , n14744 );
and ( n14746 , n14742 , n14745 );
buf ( n14747 , RI21a10c78_95);
buf ( n14748 , n14747 );
buf ( n14749 , RI210bc330_309);
buf ( n14750 , n14749 );
not ( n14751 , n14750 );
and ( n14752 , n14748 , n14751 );
buf ( n14753 , RI21a10cf0_94);
buf ( n14754 , n14753 );
buf ( n14755 , RI210bc3a8_308);
buf ( n14756 , n14755 );
not ( n14757 , n14756 );
and ( n14758 , n14754 , n14757 );
buf ( n14759 , RI21a10d68_93);
buf ( n14760 , n14759 );
buf ( n14761 , RI210bc420_307);
buf ( n14762 , n14761 );
not ( n14763 , n14762 );
and ( n14764 , n14760 , n14763 );
buf ( n14765 , RI21a11470_92);
buf ( n14766 , n14765 );
buf ( n14767 , RI210bcc90_306);
buf ( n14768 , n14767 );
not ( n14769 , n14768 );
and ( n14770 , n14766 , n14769 );
buf ( n14771 , RI21a114e8_91);
buf ( n14772 , n14771 );
buf ( n14773 , RI210bcd08_305);
buf ( n14774 , n14773 );
not ( n14775 , n14774 );
and ( n14776 , n14772 , n14775 );
buf ( n14777 , RI21a0e680_120);
buf ( n14778 , n14777 );
buf ( n14779 , RI210b8820_333);
buf ( n14780 , n14779 );
not ( n14781 , n14780 );
and ( n14782 , n14778 , n14781 );
buf ( n14783 , RI21a0e6f8_119);
buf ( n14784 , n14783 );
buf ( n14785 , RI210b8898_332);
buf ( n14786 , n14785 );
not ( n14787 , n14786 );
and ( n14788 , n14784 , n14787 );
buf ( n14789 , RI21a0e770_118);
buf ( n14790 , n14789 );
buf ( n14791 , RI210b8910_331);
buf ( n14792 , n14791 );
not ( n14793 , n14792 );
and ( n14794 , n14790 , n14793 );
buf ( n14795 , RI21a0e7e8_117);
buf ( n14796 , n14795 );
buf ( n14797 , RI210b9180_330);
buf ( n14798 , n14797 );
not ( n14799 , n14798 );
and ( n14800 , n14796 , n14799 );
buf ( n14801 , RI21a0eef0_116);
buf ( n14802 , n14801 );
buf ( n14803 , RI210b91f8_329);
buf ( n14804 , n14803 );
not ( n14805 , n14804 );
and ( n14806 , n14802 , n14805 );
buf ( n14807 , RI21a0ef68_115);
buf ( n14808 , n14807 );
buf ( n14809 , RI210b9270_328);
buf ( n14810 , n14809 );
not ( n14811 , n14810 );
and ( n14812 , n14808 , n14811 );
buf ( n14813 , RI21a0efe0_114);
buf ( n14814 , n14813 );
buf ( n14815 , RI210b92e8_327);
buf ( n14816 , n14815 );
not ( n14817 , n14816 );
and ( n14818 , n14814 , n14817 );
buf ( n14819 , RI21a0f148_111);
buf ( n14820 , n14819 );
buf ( n14821 , RI21084278_420);
buf ( n14822 , n14821 );
not ( n14823 , n14822 );
and ( n14824 , n14820 , n14823 );
buf ( n14825 , RI210cfcc8_237);
buf ( n14826 , n14825 );
buf ( n14827 , RI210842f0_419);
buf ( n14828 , n14827 );
not ( n14829 , n14828 );
and ( n14830 , n14826 , n14829 );
buf ( n14831 , RI21a11560_90);
buf ( n14832 , n14831 );
buf ( n14833 , RI210bcd80_304);
buf ( n14834 , n14833 );
not ( n14835 , n14834 );
or ( n14836 , n14832 , n14835 );
and ( n14837 , n14829 , n14836 );
and ( n14838 , n14826 , n14836 );
or ( n14839 , n14830 , n14837 , n14838 );
and ( n14840 , n14823 , n14839 );
and ( n14841 , n14820 , n14839 );
or ( n14842 , n14824 , n14840 , n14841 );
and ( n14843 , n14817 , n14842 );
and ( n14844 , n14814 , n14842 );
or ( n14845 , n14818 , n14843 , n14844 );
and ( n14846 , n14811 , n14845 );
and ( n14847 , n14808 , n14845 );
or ( n14848 , n14812 , n14846 , n14847 );
and ( n14849 , n14805 , n14848 );
and ( n14850 , n14802 , n14848 );
or ( n14851 , n14806 , n14849 , n14850 );
and ( n14852 , n14799 , n14851 );
and ( n14853 , n14796 , n14851 );
or ( n14854 , n14800 , n14852 , n14853 );
and ( n14855 , n14793 , n14854 );
and ( n14856 , n14790 , n14854 );
or ( n14857 , n14794 , n14855 , n14856 );
and ( n14858 , n14787 , n14857 );
and ( n14859 , n14784 , n14857 );
or ( n14860 , n14788 , n14858 , n14859 );
and ( n14861 , n14781 , n14860 );
and ( n14862 , n14778 , n14860 );
or ( n14863 , n14782 , n14861 , n14862 );
and ( n14864 , n14775 , n14863 );
and ( n14865 , n14772 , n14863 );
or ( n14866 , n14776 , n14864 , n14865 );
and ( n14867 , n14769 , n14866 );
and ( n14868 , n14766 , n14866 );
or ( n14869 , n14770 , n14867 , n14868 );
and ( n14870 , n14763 , n14869 );
and ( n14871 , n14760 , n14869 );
or ( n14872 , n14764 , n14870 , n14871 );
and ( n14873 , n14757 , n14872 );
and ( n14874 , n14754 , n14872 );
or ( n14875 , n14758 , n14873 , n14874 );
and ( n14876 , n14751 , n14875 );
and ( n14877 , n14748 , n14875 );
or ( n14878 , n14752 , n14876 , n14877 );
and ( n14879 , n14745 , n14878 );
and ( n14880 , n14742 , n14878 );
or ( n14881 , n14746 , n14879 , n14880 );
and ( n14882 , n14739 , n14881 );
and ( n14883 , n14736 , n14881 );
or ( n14884 , n14740 , n14882 , n14883 );
and ( n14885 , n14733 , n14884 );
and ( n14886 , n14730 , n14884 );
or ( n14887 , n14734 , n14885 , n14886 );
and ( n14888 , n14727 , n14887 );
and ( n14889 , n14724 , n14887 );
or ( n14890 , n14728 , n14888 , n14889 );
and ( n14891 , n14721 , n14890 );
and ( n14892 , n14718 , n14890 );
or ( n14893 , n14722 , n14891 , n14892 );
and ( n14894 , n14715 , n14893 );
and ( n14895 , n14712 , n14893 );
or ( n14896 , n14716 , n14894 , n14895 );
and ( n14897 , n14709 , n14896 );
and ( n14898 , n14706 , n14896 );
or ( n14899 , n14710 , n14897 , n14898 );
and ( n14900 , n14703 , n14899 );
and ( n14901 , n14700 , n14899 );
or ( n14902 , n14704 , n14900 , n14901 );
and ( n14903 , n14697 , n14902 );
and ( n14904 , n14694 , n14902 );
or ( n14905 , n14698 , n14903 , n14904 );
and ( n14906 , n14691 , n14905 );
and ( n14907 , n14688 , n14905 );
or ( n14908 , n14692 , n14906 , n14907 );
and ( n14909 , n14685 , n14908 );
and ( n14910 , n14682 , n14908 );
or ( n14911 , n14686 , n14909 , n14910 );
and ( n14912 , n14679 , n14911 );
and ( n14913 , n14676 , n14911 );
or ( n14914 , n14680 , n14912 , n14913 );
and ( n14915 , n14673 , n14914 );
and ( n14916 , n14670 , n14914 );
or ( n14917 , n14674 , n14915 , n14916 );
and ( n14918 , n14667 , n14917 );
and ( n14919 , n14664 , n14917 );
or ( n14920 , n14668 , n14918 , n14919 );
and ( n14921 , n14661 , n14920 );
and ( n14922 , n14658 , n14920 );
or ( n14923 , n14662 , n14921 , n14922 );
and ( n14924 , n14655 , n14923 );
and ( n14925 , n14652 , n14923 );
or ( n14926 , n14656 , n14924 , n14925 );
xor ( n14927 , n14650 , n14926 );
buf ( n14928 , n14927 );
and ( n14929 , n14928 , n14641 );
or ( n14930 , n14644 , n14929 );
or ( n14931 , n14143 , n14137 );
or ( n14932 , n14931 , n14140 );
and ( n14933 , n14930 , n14932 );
buf ( n14934 , n14933 );
buf ( n14935 , n14934 );
xor ( n14936 , n14618 , n14935 );
not ( n14937 , n14936 );
not ( n14938 , n14614 );
and ( n14939 , n14938 , n14611 );
or ( n14940 , n14939 , C0 );
buf ( n14941 , n14940 );
not ( n14942 , n14941 );
not ( n14943 , n14641 );
buf ( n14944 , RI21a19990_4);
and ( n14945 , n14943 , n14944 );
xor ( n14946 , n14652 , n14655 );
xor ( n14947 , n14946 , n14923 );
buf ( n14948 , n14947 );
and ( n14949 , n14948 , n14641 );
or ( n14950 , n14945 , n14949 );
and ( n14951 , n14950 , n14932 );
buf ( n14952 , n14951 );
buf ( n14953 , n14952 );
and ( n14954 , n14942 , n14953 );
xnor ( n14955 , n12739 , n12946 );
buf ( n14956 , n14955 );
and ( n14957 , n14956 , n13138 );
buf ( n14958 , RI2106cce0_589);
and ( n14959 , n14958 , n13142 );
buf ( n14960 , RI2106de38_565);
and ( n14961 , n14960 , n13145 );
buf ( n14962 , RI21073bf8_540);
and ( n14963 , n14962 , n13148 );
or ( n14964 , n14957 , n14959 , n14961 , n14963 );
buf ( n14965 , n14964 );
buf ( n14966 , n14965 );
not ( n14967 , n14966 );
not ( n14968 , n14641 );
buf ( n14969 , RI21a19918_5);
and ( n14970 , n14968 , n14969 );
xor ( n14971 , n14658 , n14661 );
xor ( n14972 , n14971 , n14920 );
buf ( n14973 , n14972 );
and ( n14974 , n14973 , n14641 );
or ( n14975 , n14970 , n14974 );
and ( n14976 , n14975 , n14932 );
buf ( n14977 , n14976 );
buf ( n14978 , n14977 );
and ( n14979 , n14967 , n14978 );
buf ( n14980 , n13162 );
buf ( n14981 , n14980 );
not ( n14982 , n14981 );
not ( n14983 , n14641 );
buf ( n14984 , RI21a198a0_6);
and ( n14985 , n14983 , n14984 );
xor ( n14986 , n14664 , n14667 );
xor ( n14987 , n14986 , n14917 );
buf ( n14988 , n14987 );
and ( n14989 , n14988 , n14641 );
or ( n14990 , n14985 , n14989 );
and ( n14991 , n14990 , n14932 );
buf ( n14992 , n14991 );
buf ( n14993 , n14992 );
and ( n14994 , n14982 , n14993 );
buf ( n14995 , n13175 );
buf ( n14996 , n14995 );
not ( n14997 , n14996 );
not ( n14998 , n14641 );
buf ( n14999 , RI21a19828_7);
and ( n15000 , n14998 , n14999 );
xor ( n15001 , n14670 , n14673 );
xor ( n15002 , n15001 , n14914 );
buf ( n15003 , n15002 );
and ( n15004 , n15003 , n14641 );
or ( n15005 , n15000 , n15004 );
and ( n15006 , n15005 , n14932 );
buf ( n15007 , n15006 );
buf ( n15008 , n15007 );
and ( n15009 , n14997 , n15008 );
buf ( n15010 , n13187 );
buf ( n15011 , n15010 );
not ( n15012 , n15011 );
not ( n15013 , n14641 );
buf ( n15014 , RI21a197b0_8);
and ( n15015 , n15013 , n15014 );
xor ( n15016 , n14676 , n14679 );
xor ( n15017 , n15016 , n14911 );
buf ( n15018 , n15017 );
and ( n15019 , n15018 , n14641 );
or ( n15020 , n15015 , n15019 );
and ( n15021 , n15020 , n14932 );
buf ( n15022 , n15021 );
buf ( n15023 , n15022 );
and ( n15024 , n15012 , n15023 );
buf ( n15025 , n13199 );
buf ( n15026 , n15025 );
not ( n15027 , n15026 );
not ( n15028 , n14641 );
buf ( n15029 , RI21a190a8_9);
and ( n15030 , n15028 , n15029 );
xor ( n15031 , n14682 , n14685 );
xor ( n15032 , n15031 , n14908 );
buf ( n15033 , n15032 );
and ( n15034 , n15033 , n14641 );
or ( n15035 , n15030 , n15034 );
and ( n15036 , n15035 , n14932 );
buf ( n15037 , n15036 );
buf ( n15038 , n15037 );
and ( n15039 , n15027 , n15038 );
buf ( n15040 , n13211 );
buf ( n15041 , n15040 );
not ( n15042 , n15041 );
not ( n15043 , n14641 );
buf ( n15044 , RI21a19030_10);
and ( n15045 , n15043 , n15044 );
xor ( n15046 , n14688 , n14691 );
xor ( n15047 , n15046 , n14905 );
buf ( n15048 , n15047 );
and ( n15049 , n15048 , n14641 );
or ( n15050 , n15045 , n15049 );
and ( n15051 , n15050 , n14932 );
buf ( n15052 , n15051 );
buf ( n15053 , n15052 );
and ( n15054 , n15042 , n15053 );
buf ( n15055 , n13223 );
buf ( n15056 , n15055 );
not ( n15057 , n15056 );
not ( n15058 , n14641 );
buf ( n15059 , RI21a18fb8_11);
and ( n15060 , n15058 , n15059 );
xor ( n15061 , n14694 , n14697 );
xor ( n15062 , n15061 , n14902 );
buf ( n15063 , n15062 );
and ( n15064 , n15063 , n14641 );
or ( n15065 , n15060 , n15064 );
and ( n15066 , n15065 , n14932 );
buf ( n15067 , n15066 );
buf ( n15068 , n15067 );
and ( n15069 , n15057 , n15068 );
buf ( n15070 , n13235 );
buf ( n15071 , n15070 );
not ( n15072 , n15071 );
not ( n15073 , n14641 );
buf ( n15074 , RI21a18f40_12);
and ( n15075 , n15073 , n15074 );
xor ( n15076 , n14700 , n14703 );
xor ( n15077 , n15076 , n14899 );
buf ( n15078 , n15077 );
and ( n15079 , n15078 , n14641 );
or ( n15080 , n15075 , n15079 );
and ( n15081 , n15080 , n14932 );
buf ( n15082 , n15081 );
buf ( n15083 , n15082 );
and ( n15084 , n15072 , n15083 );
buf ( n15085 , n13247 );
buf ( n15086 , n15085 );
not ( n15087 , n15086 );
not ( n15088 , n14641 );
buf ( n15089 , RI21a18ec8_13);
and ( n15090 , n15088 , n15089 );
xor ( n15091 , n14706 , n14709 );
xor ( n15092 , n15091 , n14896 );
buf ( n15093 , n15092 );
and ( n15094 , n15093 , n14641 );
or ( n15095 , n15090 , n15094 );
and ( n15096 , n15095 , n14932 );
buf ( n15097 , n15096 );
buf ( n15098 , n15097 );
and ( n15099 , n15087 , n15098 );
buf ( n15100 , n13259 );
buf ( n15101 , n15100 );
not ( n15102 , n15101 );
not ( n15103 , n14641 );
buf ( n15104 , RI21a18e50_14);
and ( n15105 , n15103 , n15104 );
xor ( n15106 , n14712 , n14715 );
xor ( n15107 , n15106 , n14893 );
buf ( n15108 , n15107 );
and ( n15109 , n15108 , n14641 );
or ( n15110 , n15105 , n15109 );
and ( n15111 , n15110 , n14932 );
buf ( n15112 , n15111 );
buf ( n15113 , n15112 );
and ( n15114 , n15102 , n15113 );
buf ( n15115 , n13271 );
buf ( n15116 , n15115 );
not ( n15117 , n15116 );
not ( n15118 , n14641 );
buf ( n15119 , RI21a18748_15);
and ( n15120 , n15118 , n15119 );
xor ( n15121 , n14718 , n14721 );
xor ( n15122 , n15121 , n14890 );
buf ( n15123 , n15122 );
and ( n15124 , n15123 , n14641 );
or ( n15125 , n15120 , n15124 );
and ( n15126 , n15125 , n14932 );
buf ( n15127 , n11692 );
buf ( n15128 , n15127 );
not ( n15129 , n15128 );
buf ( n15130 , n15129 );
buf ( n15131 , n15130 );
not ( n15132 , n15131 );
buf ( n15133 , n11504 );
not ( n15134 , n15133 );
buf ( n15135 , n11689 );
and ( n15136 , n15134 , n15135 );
not ( n15137 , n15135 );
not ( n15138 , n15127 );
xor ( n15139 , n15137 , n15138 );
and ( n15140 , n15139 , n15133 );
or ( n15141 , n15136 , n15140 );
buf ( n15142 , n15141 );
not ( n15143 , n15142 );
buf ( n15144 , n15143 );
buf ( n15145 , n15144 );
not ( n15146 , n15145 );
or ( n15147 , n15132 , n15146 );
not ( n15148 , n15133 );
buf ( n15149 , n11681 );
and ( n15150 , n15148 , n15149 );
not ( n15151 , n15149 );
and ( n15152 , n15137 , n15138 );
xor ( n15153 , n15151 , n15152 );
and ( n15154 , n15153 , n15133 );
or ( n15155 , n15150 , n15154 );
buf ( n15156 , n15155 );
not ( n15157 , n15156 );
buf ( n15158 , n15157 );
buf ( n15159 , n15158 );
not ( n15160 , n15159 );
or ( n15161 , n15147 , n15160 );
not ( n15162 , n15133 );
buf ( n15163 , n11673 );
and ( n15164 , n15162 , n15163 );
not ( n15165 , n15163 );
and ( n15166 , n15151 , n15152 );
xor ( n15167 , n15165 , n15166 );
and ( n15168 , n15167 , n15133 );
or ( n15169 , n15164 , n15168 );
buf ( n15170 , n15169 );
not ( n15171 , n15170 );
buf ( n15172 , n15171 );
buf ( n15173 , n15172 );
not ( n15174 , n15173 );
or ( n15175 , n15161 , n15174 );
not ( n15176 , n15133 );
buf ( n15177 , n11665 );
and ( n15178 , n15176 , n15177 );
not ( n15179 , n15177 );
and ( n15180 , n15165 , n15166 );
xor ( n15181 , n15179 , n15180 );
and ( n15182 , n15181 , n15133 );
or ( n15183 , n15178 , n15182 );
buf ( n15184 , n15183 );
not ( n15185 , n15184 );
buf ( n15186 , n15185 );
buf ( n15187 , n15186 );
not ( n15188 , n15187 );
or ( n15189 , n15175 , n15188 );
not ( n15190 , n15133 );
buf ( n15191 , n11657 );
and ( n15192 , n15190 , n15191 );
not ( n15193 , n15191 );
and ( n15194 , n15179 , n15180 );
xor ( n15195 , n15193 , n15194 );
and ( n15196 , n15195 , n15133 );
or ( n15197 , n15192 , n15196 );
buf ( n15198 , n15197 );
not ( n15199 , n15198 );
buf ( n15200 , n15199 );
buf ( n15201 , n15200 );
not ( n15202 , n15201 );
or ( n15203 , n15189 , n15202 );
not ( n15204 , n15133 );
buf ( n15205 , n11649 );
and ( n15206 , n15204 , n15205 );
not ( n15207 , n15205 );
and ( n15208 , n15193 , n15194 );
xor ( n15209 , n15207 , n15208 );
and ( n15210 , n15209 , n15133 );
or ( n15211 , n15206 , n15210 );
buf ( n15212 , n15211 );
not ( n15213 , n15212 );
buf ( n15214 , n15213 );
buf ( n15215 , n15214 );
not ( n15216 , n15215 );
or ( n15217 , n15203 , n15216 );
not ( n15218 , n15133 );
buf ( n15219 , n11641 );
and ( n15220 , n15218 , n15219 );
not ( n15221 , n15219 );
and ( n15222 , n15207 , n15208 );
xor ( n15223 , n15221 , n15222 );
and ( n15224 , n15223 , n15133 );
or ( n15225 , n15220 , n15224 );
buf ( n15226 , n15225 );
not ( n15227 , n15226 );
buf ( n15228 , n15227 );
buf ( n15229 , n15228 );
not ( n15230 , n15229 );
or ( n15231 , n15217 , n15230 );
not ( n15232 , n15133 );
buf ( n15233 , n11633 );
and ( n15234 , n15232 , n15233 );
not ( n15235 , n15233 );
and ( n15236 , n15221 , n15222 );
xor ( n15237 , n15235 , n15236 );
and ( n15238 , n15237 , n15133 );
or ( n15239 , n15234 , n15238 );
buf ( n15240 , n15239 );
not ( n15241 , n15240 );
buf ( n15242 , n15241 );
buf ( n15243 , n15242 );
not ( n15244 , n15243 );
or ( n15245 , n15231 , n15244 );
not ( n15246 , n15133 );
buf ( n15247 , n11625 );
and ( n15248 , n15246 , n15247 );
not ( n15249 , n15247 );
and ( n15250 , n15235 , n15236 );
xor ( n15251 , n15249 , n15250 );
and ( n15252 , n15251 , n15133 );
or ( n15253 , n15248 , n15252 );
buf ( n15254 , n15253 );
not ( n15255 , n15254 );
buf ( n15256 , n15255 );
buf ( n15257 , n15256 );
not ( n15258 , n15257 );
or ( n15259 , n15245 , n15258 );
not ( n15260 , n15133 );
buf ( n15261 , n11617 );
and ( n15262 , n15260 , n15261 );
not ( n15263 , n15261 );
and ( n15264 , n15249 , n15250 );
xor ( n15265 , n15263 , n15264 );
and ( n15266 , n15265 , n15133 );
or ( n15267 , n15262 , n15266 );
buf ( n15268 , n15267 );
not ( n15269 , n15268 );
buf ( n15270 , n15269 );
buf ( n15271 , n15270 );
not ( n15272 , n15271 );
or ( n15273 , n15259 , n15272 );
not ( n15274 , n15133 );
buf ( n15275 , n11609 );
and ( n15276 , n15274 , n15275 );
not ( n15277 , n15275 );
and ( n15278 , n15263 , n15264 );
xor ( n15279 , n15277 , n15278 );
and ( n15280 , n15279 , n15133 );
or ( n15281 , n15276 , n15280 );
buf ( n15282 , n15281 );
not ( n15283 , n15282 );
buf ( n15284 , n15283 );
buf ( n15285 , n15284 );
not ( n15286 , n15285 );
or ( n15287 , n15273 , n15286 );
not ( n15288 , n15133 );
buf ( n15289 , n11601 );
and ( n15290 , n15288 , n15289 );
not ( n15291 , n15289 );
and ( n15292 , n15277 , n15278 );
xor ( n15293 , n15291 , n15292 );
and ( n15294 , n15293 , n15133 );
or ( n15295 , n15290 , n15294 );
buf ( n15296 , n15295 );
not ( n15297 , n15296 );
buf ( n15298 , n15297 );
buf ( n15299 , n15298 );
not ( n15300 , n15299 );
or ( n15301 , n15287 , n15300 );
not ( n15302 , n15133 );
buf ( n15303 , n11593 );
and ( n15304 , n15302 , n15303 );
not ( n15305 , n15303 );
and ( n15306 , n15291 , n15292 );
xor ( n15307 , n15305 , n15306 );
and ( n15308 , n15307 , n15133 );
or ( n15309 , n15304 , n15308 );
buf ( n15310 , n15309 );
not ( n15311 , n15310 );
buf ( n15312 , n15311 );
buf ( n15313 , n15312 );
not ( n15314 , n15313 );
or ( n15315 , n15301 , n15314 );
not ( n15316 , n15133 );
buf ( n15317 , n11585 );
and ( n15318 , n15316 , n15317 );
not ( n15319 , n15317 );
and ( n15320 , n15305 , n15306 );
xor ( n15321 , n15319 , n15320 );
and ( n15322 , n15321 , n15133 );
or ( n15323 , n15318 , n15322 );
buf ( n15324 , n15323 );
not ( n15325 , n15324 );
buf ( n15326 , n15325 );
buf ( n15327 , n15326 );
not ( n15328 , n15327 );
or ( n15329 , n15315 , n15328 );
not ( n15330 , n15133 );
buf ( n15331 , n11577 );
and ( n15332 , n15330 , n15331 );
not ( n15333 , n15331 );
and ( n15334 , n15319 , n15320 );
xor ( n15335 , n15333 , n15334 );
and ( n15336 , n15335 , n15133 );
or ( n15337 , n15332 , n15336 );
buf ( n15338 , n15337 );
not ( n15339 , n15338 );
buf ( n15340 , n15339 );
buf ( n15341 , n15340 );
not ( n15342 , n15341 );
or ( n15343 , n15329 , n15342 );
not ( n15344 , n15133 );
buf ( n15345 , n11569 );
and ( n15346 , n15344 , n15345 );
not ( n15347 , n15345 );
and ( n15348 , n15333 , n15334 );
xor ( n15349 , n15347 , n15348 );
and ( n15350 , n15349 , n15133 );
or ( n15351 , n15346 , n15350 );
buf ( n15352 , n15351 );
not ( n15353 , n15352 );
buf ( n15354 , n15353 );
buf ( n15355 , n15354 );
not ( n15356 , n15355 );
or ( n15357 , n15343 , n15356 );
not ( n15358 , n15133 );
buf ( n15359 , n11561 );
and ( n15360 , n15358 , n15359 );
not ( n15361 , n15359 );
and ( n15362 , n15347 , n15348 );
xor ( n15363 , n15361 , n15362 );
and ( n15364 , n15363 , n15133 );
or ( n15365 , n15360 , n15364 );
buf ( n15366 , n15365 );
not ( n15367 , n15366 );
buf ( n15368 , n15367 );
buf ( n15369 , n15368 );
not ( n15370 , n15369 );
or ( n15371 , n15357 , n15370 );
not ( n15372 , n15133 );
buf ( n15373 , n11553 );
and ( n15374 , n15372 , n15373 );
not ( n15375 , n15373 );
and ( n15376 , n15361 , n15362 );
xor ( n15377 , n15375 , n15376 );
and ( n15378 , n15377 , n15133 );
or ( n15379 , n15374 , n15378 );
buf ( n15380 , n15379 );
not ( n15381 , n15380 );
buf ( n15382 , n15381 );
buf ( n15383 , n15382 );
not ( n15384 , n15383 );
or ( n15385 , n15371 , n15384 );
not ( n15386 , n15133 );
buf ( n15387 , n11545 );
and ( n15388 , n15386 , n15387 );
not ( n15389 , n15387 );
and ( n15390 , n15375 , n15376 );
xor ( n15391 , n15389 , n15390 );
and ( n15392 , n15391 , n15133 );
or ( n15393 , n15388 , n15392 );
buf ( n15394 , n15393 );
not ( n15395 , n15394 );
buf ( n15396 , n15395 );
buf ( n15397 , n15396 );
not ( n15398 , n15397 );
or ( n15399 , n15385 , n15398 );
buf ( n15400 , n15399 );
buf ( n15401 , n15400 );
and ( n15402 , n15401 , n15133 );
not ( n15403 , n15402 );
and ( n15404 , n15403 , n15398 );
xor ( n15405 , n15398 , n15133 );
xor ( n15406 , n15384 , n15133 );
xor ( n15407 , n15370 , n15133 );
xor ( n15408 , n15356 , n15133 );
xor ( n15409 , n15342 , n15133 );
xor ( n15410 , n15328 , n15133 );
xor ( n15411 , n15314 , n15133 );
xor ( n15412 , n15300 , n15133 );
xor ( n15413 , n15286 , n15133 );
xor ( n15414 , n15272 , n15133 );
xor ( n15415 , n15258 , n15133 );
xor ( n15416 , n15244 , n15133 );
xor ( n15417 , n15230 , n15133 );
xor ( n15418 , n15216 , n15133 );
xor ( n15419 , n15202 , n15133 );
xor ( n15420 , n15188 , n15133 );
xor ( n15421 , n15174 , n15133 );
xor ( n15422 , n15160 , n15133 );
xor ( n15423 , n15146 , n15133 );
xor ( n15424 , n15132 , n15133 );
and ( n15425 , n15424 , n15133 );
and ( n15426 , n15423 , n15425 );
and ( n15427 , n15422 , n15426 );
and ( n15428 , n15421 , n15427 );
and ( n15429 , n15420 , n15428 );
and ( n15430 , n15419 , n15429 );
and ( n15431 , n15418 , n15430 );
and ( n15432 , n15417 , n15431 );
and ( n15433 , n15416 , n15432 );
and ( n15434 , n15415 , n15433 );
and ( n15435 , n15414 , n15434 );
and ( n15436 , n15413 , n15435 );
and ( n15437 , n15412 , n15436 );
and ( n15438 , n15411 , n15437 );
and ( n15439 , n15410 , n15438 );
and ( n15440 , n15409 , n15439 );
and ( n15441 , n15408 , n15440 );
and ( n15442 , n15407 , n15441 );
and ( n15443 , n15406 , n15442 );
xor ( n15444 , n15405 , n15443 );
and ( n15445 , n15444 , n15402 );
or ( n15446 , n15404 , n15445 );
buf ( n15447 , n15446 );
and ( n15448 , n15447 , n14141 );
or ( n15449 , n15126 , n15448 );
buf ( n15450 , n15449 );
and ( n15451 , n15117 , n15450 );
buf ( n15452 , n13283 );
buf ( n15453 , n15452 );
not ( n15454 , n15453 );
not ( n15455 , n14641 );
buf ( n15456 , RI21a186d0_16);
and ( n15457 , n15455 , n15456 );
xor ( n15458 , n14724 , n14727 );
xor ( n15459 , n15458 , n14887 );
buf ( n15460 , n15459 );
and ( n15461 , n15460 , n14641 );
or ( n15462 , n15457 , n15461 );
and ( n15463 , n15462 , n14932 );
not ( n15464 , n15402 );
and ( n15465 , n15464 , n15384 );
xor ( n15466 , n15406 , n15442 );
and ( n15467 , n15466 , n15402 );
or ( n15468 , n15465 , n15467 );
buf ( n15469 , n15468 );
and ( n15470 , n15469 , n14141 );
or ( n15471 , n15463 , n15470 );
buf ( n15472 , n15471 );
and ( n15473 , n15454 , n15472 );
buf ( n15474 , n13295 );
buf ( n15475 , n15474 );
not ( n15476 , n15475 );
not ( n15477 , n14641 );
buf ( n15478 , RI21a18658_17);
and ( n15479 , n15477 , n15478 );
xor ( n15480 , n14730 , n14733 );
xor ( n15481 , n15480 , n14884 );
buf ( n15482 , n15481 );
and ( n15483 , n15482 , n14641 );
or ( n15484 , n15479 , n15483 );
and ( n15485 , n15484 , n14932 );
not ( n15486 , n15402 );
and ( n15487 , n15486 , n15370 );
xor ( n15488 , n15407 , n15441 );
and ( n15489 , n15488 , n15402 );
or ( n15490 , n15487 , n15489 );
buf ( n15491 , n15490 );
and ( n15492 , n15491 , n14141 );
or ( n15493 , n15485 , n15492 );
buf ( n15494 , n15493 );
and ( n15495 , n15476 , n15494 );
buf ( n15496 , n13307 );
buf ( n15497 , n15496 );
not ( n15498 , n15497 );
not ( n15499 , n14641 );
buf ( n15500 , RI21a185e0_18);
and ( n15501 , n15499 , n15500 );
xor ( n15502 , n14736 , n14739 );
xor ( n15503 , n15502 , n14881 );
buf ( n15504 , n15503 );
and ( n15505 , n15504 , n14641 );
or ( n15506 , n15501 , n15505 );
and ( n15507 , n15506 , n14932 );
not ( n15508 , n15402 );
and ( n15509 , n15508 , n15356 );
xor ( n15510 , n15408 , n15440 );
and ( n15511 , n15510 , n15402 );
or ( n15512 , n15509 , n15511 );
buf ( n15513 , n15512 );
and ( n15514 , n15513 , n14141 );
or ( n15515 , n15507 , n15514 );
buf ( n15516 , n15515 );
and ( n15517 , n15498 , n15516 );
buf ( n15518 , n13319 );
buf ( n15519 , n15518 );
not ( n15520 , n15519 );
not ( n15521 , n14641 );
buf ( n15522 , RI21a18568_19);
and ( n15523 , n15521 , n15522 );
xor ( n15524 , n14742 , n14745 );
xor ( n15525 , n15524 , n14878 );
buf ( n15526 , n15525 );
and ( n15527 , n15526 , n14641 );
or ( n15528 , n15523 , n15527 );
and ( n15529 , n15528 , n14932 );
not ( n15530 , n15402 );
and ( n15531 , n15530 , n15342 );
xor ( n15532 , n15409 , n15439 );
and ( n15533 , n15532 , n15402 );
or ( n15534 , n15531 , n15533 );
buf ( n15535 , n15534 );
and ( n15536 , n15535 , n14141 );
or ( n15537 , n15529 , n15536 );
buf ( n15538 , n15537 );
and ( n15539 , n15520 , n15538 );
buf ( n15540 , n13331 );
buf ( n15541 , n15540 );
not ( n15542 , n15541 );
not ( n15543 , n14641 );
buf ( n15544 , RI21a184f0_20);
and ( n15545 , n15543 , n15544 );
xor ( n15546 , n14748 , n14751 );
xor ( n15547 , n15546 , n14875 );
buf ( n15548 , n15547 );
and ( n15549 , n15548 , n14641 );
or ( n15550 , n15545 , n15549 );
and ( n15551 , n15550 , n14932 );
not ( n15552 , n15402 );
and ( n15553 , n15552 , n15328 );
xor ( n15554 , n15410 , n15438 );
and ( n15555 , n15554 , n15402 );
or ( n15556 , n15553 , n15555 );
buf ( n15557 , n15556 );
and ( n15558 , n15557 , n14141 );
or ( n15559 , n15551 , n15558 );
buf ( n15560 , n15559 );
and ( n15561 , n15542 , n15560 );
buf ( n15562 , n13343 );
buf ( n15563 , n15562 );
not ( n15564 , n15563 );
not ( n15565 , n14641 );
buf ( n15566 , RI21a17de8_21);
and ( n15567 , n15565 , n15566 );
xor ( n15568 , n14754 , n14757 );
xor ( n15569 , n15568 , n14872 );
buf ( n15570 , n15569 );
and ( n15571 , n15570 , n14641 );
or ( n15572 , n15567 , n15571 );
and ( n15573 , n15572 , n14932 );
not ( n15574 , n15402 );
and ( n15575 , n15574 , n15314 );
xor ( n15576 , n15411 , n15437 );
and ( n15577 , n15576 , n15402 );
or ( n15578 , n15575 , n15577 );
buf ( n15579 , n15578 );
and ( n15580 , n15579 , n14141 );
or ( n15581 , n15573 , n15580 );
buf ( n15582 , n15581 );
and ( n15583 , n15564 , n15582 );
buf ( n15584 , n13355 );
buf ( n15585 , n15584 );
not ( n15586 , n15585 );
not ( n15587 , n14641 );
buf ( n15588 , RI21a17d70_22);
and ( n15589 , n15587 , n15588 );
xor ( n15590 , n14760 , n14763 );
xor ( n15591 , n15590 , n14869 );
buf ( n15592 , n15591 );
and ( n15593 , n15592 , n14641 );
or ( n15594 , n15589 , n15593 );
and ( n15595 , n15594 , n14932 );
not ( n15596 , n15402 );
and ( n15597 , n15596 , n15300 );
xor ( n15598 , n15412 , n15436 );
and ( n15599 , n15598 , n15402 );
or ( n15600 , n15597 , n15599 );
buf ( n15601 , n15600 );
and ( n15602 , n15601 , n14141 );
or ( n15603 , n15595 , n15602 );
buf ( n15604 , n15603 );
and ( n15605 , n15586 , n15604 );
buf ( n15606 , n13367 );
buf ( n15607 , n15606 );
not ( n15608 , n15607 );
not ( n15609 , n14641 );
buf ( n15610 , RI21a17cf8_23);
and ( n15611 , n15609 , n15610 );
xor ( n15612 , n14766 , n14769 );
xor ( n15613 , n15612 , n14866 );
buf ( n15614 , n15613 );
and ( n15615 , n15614 , n14641 );
or ( n15616 , n15611 , n15615 );
and ( n15617 , n15616 , n14932 );
not ( n15618 , n15402 );
and ( n15619 , n15618 , n15286 );
xor ( n15620 , n15413 , n15435 );
and ( n15621 , n15620 , n15402 );
or ( n15622 , n15619 , n15621 );
buf ( n15623 , n15622 );
and ( n15624 , n15623 , n14141 );
or ( n15625 , n15617 , n15624 );
buf ( n15626 , n15625 );
and ( n15627 , n15608 , n15626 );
buf ( n15628 , n13379 );
buf ( n15629 , n15628 );
not ( n15630 , n15629 );
not ( n15631 , n14641 );
buf ( n15632 , RI21a17c80_24);
and ( n15633 , n15631 , n15632 );
xor ( n15634 , n14772 , n14775 );
xor ( n15635 , n15634 , n14863 );
buf ( n15636 , n15635 );
and ( n15637 , n15636 , n14641 );
or ( n15638 , n15633 , n15637 );
and ( n15639 , n15638 , n14932 );
not ( n15640 , n15402 );
and ( n15641 , n15640 , n15272 );
xor ( n15642 , n15414 , n15434 );
and ( n15643 , n15642 , n15402 );
or ( n15644 , n15641 , n15643 );
buf ( n15645 , n15644 );
and ( n15646 , n15645 , n14141 );
or ( n15647 , n15639 , n15646 );
buf ( n15648 , n15647 );
and ( n15649 , n15630 , n15648 );
buf ( n15650 , n13391 );
buf ( n15651 , n15650 );
not ( n15652 , n15651 );
not ( n15653 , n14641 );
buf ( n15654 , RI21a17c08_25);
and ( n15655 , n15653 , n15654 );
xor ( n15656 , n14778 , n14781 );
xor ( n15657 , n15656 , n14860 );
buf ( n15658 , n15657 );
and ( n15659 , n15658 , n14641 );
or ( n15660 , n15655 , n15659 );
and ( n15661 , n15660 , n14932 );
not ( n15662 , n15402 );
and ( n15663 , n15662 , n15258 );
xor ( n15664 , n15415 , n15433 );
and ( n15665 , n15664 , n15402 );
or ( n15666 , n15663 , n15665 );
buf ( n15667 , n15666 );
and ( n15668 , n15667 , n14141 );
or ( n15669 , n15661 , n15668 );
buf ( n15670 , n15669 );
and ( n15671 , n15652 , n15670 );
buf ( n15672 , n13403 );
buf ( n15673 , n15672 );
not ( n15674 , n15673 );
not ( n15675 , n14641 );
buf ( n15676 , RI21a17b90_26);
and ( n15677 , n15675 , n15676 );
xor ( n15678 , n14784 , n14787 );
xor ( n15679 , n15678 , n14857 );
buf ( n15680 , n15679 );
and ( n15681 , n15680 , n14641 );
or ( n15682 , n15677 , n15681 );
and ( n15683 , n15682 , n14932 );
not ( n15684 , n15402 );
and ( n15685 , n15684 , n15244 );
xor ( n15686 , n15416 , n15432 );
and ( n15687 , n15686 , n15402 );
or ( n15688 , n15685 , n15687 );
buf ( n15689 , n15688 );
and ( n15690 , n15689 , n14141 );
or ( n15691 , n15683 , n15690 );
buf ( n15692 , n15691 );
and ( n15693 , n15674 , n15692 );
buf ( n15694 , n13415 );
buf ( n15695 , n15694 );
not ( n15696 , n15695 );
not ( n15697 , n14641 );
buf ( n15698 , RI21a17488_27);
and ( n15699 , n15697 , n15698 );
xor ( n15700 , n14790 , n14793 );
xor ( n15701 , n15700 , n14854 );
buf ( n15702 , n15701 );
and ( n15703 , n15702 , n14641 );
or ( n15704 , n15699 , n15703 );
and ( n15705 , n15704 , n14932 );
not ( n15706 , n15402 );
and ( n15707 , n15706 , n15230 );
xor ( n15708 , n15417 , n15431 );
and ( n15709 , n15708 , n15402 );
or ( n15710 , n15707 , n15709 );
buf ( n15711 , n15710 );
and ( n15712 , n15711 , n14141 );
or ( n15713 , n15705 , n15712 );
buf ( n15714 , n15713 );
and ( n15715 , n15696 , n15714 );
buf ( n15716 , n13427 );
buf ( n15717 , n15716 );
not ( n15718 , n15717 );
not ( n15719 , n14641 );
buf ( n15720 , RI21a17410_28);
and ( n15721 , n15719 , n15720 );
xor ( n15722 , n14796 , n14799 );
xor ( n15723 , n15722 , n14851 );
buf ( n15724 , n15723 );
and ( n15725 , n15724 , n14641 );
or ( n15726 , n15721 , n15725 );
and ( n15727 , n15726 , n14932 );
not ( n15728 , n15402 );
and ( n15729 , n15728 , n15216 );
xor ( n15730 , n15418 , n15430 );
and ( n15731 , n15730 , n15402 );
or ( n15732 , n15729 , n15731 );
buf ( n15733 , n15732 );
and ( n15734 , n15733 , n14141 );
or ( n15735 , n15727 , n15734 );
buf ( n15736 , n15735 );
and ( n15737 , n15718 , n15736 );
buf ( n15738 , n13439 );
buf ( n15739 , n15738 );
not ( n15740 , n15739 );
not ( n15741 , n14641 );
buf ( n15742 , RI21a17398_29);
and ( n15743 , n15741 , n15742 );
xor ( n15744 , n14802 , n14805 );
xor ( n15745 , n15744 , n14848 );
buf ( n15746 , n15745 );
and ( n15747 , n15746 , n14641 );
or ( n15748 , n15743 , n15747 );
and ( n15749 , n15748 , n14932 );
not ( n15750 , n15402 );
and ( n15751 , n15750 , n15202 );
xor ( n15752 , n15419 , n15429 );
and ( n15753 , n15752 , n15402 );
or ( n15754 , n15751 , n15753 );
buf ( n15755 , n15754 );
and ( n15756 , n15755 , n14141 );
or ( n15757 , n15749 , n15756 );
buf ( n15758 , n15757 );
and ( n15759 , n15740 , n15758 );
buf ( n15760 , n13451 );
buf ( n15761 , n15760 );
not ( n15762 , n15761 );
not ( n15763 , n14641 );
buf ( n15764 , RI21a17320_30);
and ( n15765 , n15763 , n15764 );
xor ( n15766 , n14808 , n14811 );
xor ( n15767 , n15766 , n14845 );
buf ( n15768 , n15767 );
and ( n15769 , n15768 , n14641 );
or ( n15770 , n15765 , n15769 );
and ( n15771 , n15770 , n14932 );
not ( n15772 , n15402 );
and ( n15773 , n15772 , n15188 );
xor ( n15774 , n15420 , n15428 );
and ( n15775 , n15774 , n15402 );
or ( n15776 , n15773 , n15775 );
buf ( n15777 , n15776 );
and ( n15778 , n15777 , n14141 );
or ( n15779 , n15771 , n15778 );
buf ( n15780 , n15779 );
and ( n15781 , n15762 , n15780 );
buf ( n15782 , n13463 );
buf ( n15783 , n15782 );
not ( n15784 , n15783 );
not ( n15785 , n14641 );
buf ( n15786 , RI21a172a8_31);
and ( n15787 , n15785 , n15786 );
xor ( n15788 , n14814 , n14817 );
xor ( n15789 , n15788 , n14842 );
buf ( n15790 , n15789 );
and ( n15791 , n15790 , n14641 );
or ( n15792 , n15787 , n15791 );
and ( n15793 , n15792 , n14932 );
not ( n15794 , n15402 );
and ( n15795 , n15794 , n15174 );
xor ( n15796 , n15421 , n15427 );
and ( n15797 , n15796 , n15402 );
or ( n15798 , n15795 , n15797 );
buf ( n15799 , n15798 );
and ( n15800 , n15799 , n14141 );
or ( n15801 , n15793 , n15800 );
buf ( n15802 , n15801 );
and ( n15803 , n15784 , n15802 );
buf ( n15804 , n13480 );
buf ( n15805 , n15804 );
not ( n15806 , n15805 );
not ( n15807 , n14641 );
buf ( n15808 , RI21a17230_32);
and ( n15809 , n15807 , n15808 );
xor ( n15810 , n14820 , n14823 );
xor ( n15811 , n15810 , n14839 );
buf ( n15812 , n15811 );
and ( n15813 , n15812 , n14641 );
or ( n15814 , n15809 , n15813 );
and ( n15815 , n15814 , n14932 );
not ( n15816 , n15402 );
and ( n15817 , n15816 , n15160 );
xor ( n15818 , n15422 , n15426 );
and ( n15819 , n15818 , n15402 );
or ( n15820 , n15817 , n15819 );
buf ( n15821 , n15820 );
and ( n15822 , n15821 , n14141 );
or ( n15823 , n15815 , n15822 );
buf ( n15824 , n15823 );
and ( n15825 , n15806 , n15824 );
buf ( n15826 , n13497 );
buf ( n15827 , n15826 );
not ( n15828 , n15827 );
not ( n15829 , n14641 );
buf ( n15830 , RI21a16b28_33);
and ( n15831 , n15829 , n15830 );
xor ( n15832 , n14826 , n14829 );
xor ( n15833 , n15832 , n14836 );
buf ( n15834 , n15833 );
and ( n15835 , n15834 , n14641 );
or ( n15836 , n15831 , n15835 );
and ( n15837 , n15836 , n14932 );
not ( n15838 , n15402 );
and ( n15839 , n15838 , n15146 );
xor ( n15840 , n15423 , n15425 );
and ( n15841 , n15840 , n15402 );
or ( n15842 , n15839 , n15841 );
buf ( n15843 , n15842 );
and ( n15844 , n15843 , n14141 );
or ( n15845 , n15837 , n15844 );
buf ( n15846 , n15845 );
and ( n15847 , n15828 , n15846 );
buf ( n15848 , n13514 );
buf ( n15849 , n15848 );
not ( n15850 , n15849 );
not ( n15851 , n14641 );
buf ( n15852 , RI21a16ab0_34);
and ( n15853 , n15851 , n15852 );
xor ( n15854 , n14832 , n14834 );
buf ( n15855 , n15854 );
and ( n15856 , n15855 , n14641 );
or ( n15857 , n15853 , n15856 );
and ( n15858 , n15857 , n14932 );
not ( n15859 , n15402 );
and ( n15860 , n15859 , n15132 );
xor ( n15861 , n15424 , n15133 );
and ( n15862 , n15861 , n15402 );
or ( n15863 , n15860 , n15862 );
buf ( n15864 , n15863 );
and ( n15865 , n15864 , n14141 );
or ( n15866 , n15858 , n15865 );
buf ( n15867 , n15866 );
and ( n15868 , n15850 , n15867 );
xnor ( n15869 , n15827 , n15846 );
and ( n15870 , n15868 , n15869 );
or ( n15871 , n15847 , n15870 );
xnor ( n15872 , n15805 , n15824 );
and ( n15873 , n15871 , n15872 );
or ( n15874 , n15825 , n15873 );
xnor ( n15875 , n15783 , n15802 );
and ( n15876 , n15874 , n15875 );
or ( n15877 , n15803 , n15876 );
xnor ( n15878 , n15761 , n15780 );
and ( n15879 , n15877 , n15878 );
or ( n15880 , n15781 , n15879 );
xnor ( n15881 , n15739 , n15758 );
and ( n15882 , n15880 , n15881 );
or ( n15883 , n15759 , n15882 );
xnor ( n15884 , n15717 , n15736 );
and ( n15885 , n15883 , n15884 );
or ( n15886 , n15737 , n15885 );
xnor ( n15887 , n15695 , n15714 );
and ( n15888 , n15886 , n15887 );
or ( n15889 , n15715 , n15888 );
xnor ( n15890 , n15673 , n15692 );
and ( n15891 , n15889 , n15890 );
or ( n15892 , n15693 , n15891 );
xnor ( n15893 , n15651 , n15670 );
and ( n15894 , n15892 , n15893 );
or ( n15895 , n15671 , n15894 );
xnor ( n15896 , n15629 , n15648 );
and ( n15897 , n15895 , n15896 );
or ( n15898 , n15649 , n15897 );
xnor ( n15899 , n15607 , n15626 );
and ( n15900 , n15898 , n15899 );
or ( n15901 , n15627 , n15900 );
xnor ( n15902 , n15585 , n15604 );
and ( n15903 , n15901 , n15902 );
or ( n15904 , n15605 , n15903 );
xnor ( n15905 , n15563 , n15582 );
and ( n15906 , n15904 , n15905 );
or ( n15907 , n15583 , n15906 );
xnor ( n15908 , n15541 , n15560 );
and ( n15909 , n15907 , n15908 );
or ( n15910 , n15561 , n15909 );
xnor ( n15911 , n15519 , n15538 );
and ( n15912 , n15910 , n15911 );
or ( n15913 , n15539 , n15912 );
xnor ( n15914 , n15497 , n15516 );
and ( n15915 , n15913 , n15914 );
or ( n15916 , n15517 , n15915 );
xnor ( n15917 , n15475 , n15494 );
and ( n15918 , n15916 , n15917 );
or ( n15919 , n15495 , n15918 );
xnor ( n15920 , n15453 , n15472 );
and ( n15921 , n15919 , n15920 );
or ( n15922 , n15473 , n15921 );
xnor ( n15923 , n15116 , n15450 );
and ( n15924 , n15922 , n15923 );
or ( n15925 , n15451 , n15924 );
xnor ( n15926 , n15101 , n15113 );
and ( n15927 , n15925 , n15926 );
or ( n15928 , n15114 , n15927 );
xnor ( n15929 , n15086 , n15098 );
and ( n15930 , n15928 , n15929 );
or ( n15931 , n15099 , n15930 );
xnor ( n15932 , n15071 , n15083 );
and ( n15933 , n15931 , n15932 );
or ( n15934 , n15084 , n15933 );
xnor ( n15935 , n15056 , n15068 );
and ( n15936 , n15934 , n15935 );
or ( n15937 , n15069 , n15936 );
xnor ( n15938 , n15041 , n15053 );
and ( n15939 , n15937 , n15938 );
or ( n15940 , n15054 , n15939 );
xnor ( n15941 , n15026 , n15038 );
and ( n15942 , n15940 , n15941 );
or ( n15943 , n15039 , n15942 );
xnor ( n15944 , n15011 , n15023 );
and ( n15945 , n15943 , n15944 );
or ( n15946 , n15024 , n15945 );
xnor ( n15947 , n14996 , n15008 );
and ( n15948 , n15946 , n15947 );
or ( n15949 , n15009 , n15948 );
xnor ( n15950 , n14981 , n14993 );
and ( n15951 , n15949 , n15950 );
or ( n15952 , n14994 , n15951 );
xnor ( n15953 , n14966 , n14978 );
and ( n15954 , n15952 , n15953 );
or ( n15955 , n14979 , n15954 );
xnor ( n15956 , n14941 , n14953 );
and ( n15957 , n15955 , n15956 );
or ( n15958 , n14954 , n15957 );
and ( n15959 , n14937 , n15958 );
not ( n15960 , n14935 );
and ( n15961 , n15960 , n14618 );
and ( n15962 , n15961 , n14936 );
or ( n15963 , n15959 , n15962 );
buf ( n15964 , n15963 );
not ( n15965 , n15964 );
or ( n15966 , n15965 , n14139 );
and ( n15967 , n15966 , n14591 );
or ( n15968 , n15964 , n14139 );
and ( n15969 , n15968 , n14589 );
buf ( n15970 , n13150 );
buf ( n15971 , n14934 );
xor ( n15972 , n15970 , n15971 );
not ( n15973 , n15972 );
buf ( n15974 , n14952 );
not ( n15975 , n15974 );
buf ( n15976 , n14611 );
and ( n15977 , n15975 , n15976 );
buf ( n15978 , n14977 );
not ( n15979 , n15978 );
buf ( n15980 , n14964 );
and ( n15981 , n15979 , n15980 );
buf ( n15982 , n14992 );
not ( n15983 , n15982 );
buf ( n15984 , n13162 );
and ( n15985 , n15983 , n15984 );
buf ( n15986 , n15007 );
not ( n15987 , n15986 );
buf ( n15988 , n13175 );
and ( n15989 , n15987 , n15988 );
buf ( n15990 , n15022 );
not ( n15991 , n15990 );
buf ( n15992 , n13187 );
and ( n15993 , n15991 , n15992 );
buf ( n15994 , n15037 );
not ( n15995 , n15994 );
buf ( n15996 , n13199 );
and ( n15997 , n15995 , n15996 );
buf ( n15998 , n15052 );
not ( n15999 , n15998 );
buf ( n16000 , n13211 );
and ( n16001 , n15999 , n16000 );
buf ( n16002 , n15067 );
not ( n16003 , n16002 );
buf ( n16004 , n13223 );
and ( n16005 , n16003 , n16004 );
buf ( n16006 , n15082 );
not ( n16007 , n16006 );
buf ( n16008 , n13235 );
and ( n16009 , n16007 , n16008 );
buf ( n16010 , n15097 );
not ( n16011 , n16010 );
buf ( n16012 , n13247 );
and ( n16013 , n16011 , n16012 );
buf ( n16014 , n15112 );
not ( n16015 , n16014 );
buf ( n16016 , n13259 );
and ( n16017 , n16015 , n16016 );
buf ( n16018 , n15449 );
not ( n16019 , n16018 );
buf ( n16020 , n13271 );
and ( n16021 , n16019 , n16020 );
buf ( n16022 , n15471 );
not ( n16023 , n16022 );
buf ( n16024 , n13283 );
and ( n16025 , n16023 , n16024 );
buf ( n16026 , n15493 );
not ( n16027 , n16026 );
buf ( n16028 , n13295 );
and ( n16029 , n16027 , n16028 );
buf ( n16030 , n15515 );
not ( n16031 , n16030 );
buf ( n16032 , n13307 );
and ( n16033 , n16031 , n16032 );
buf ( n16034 , n15537 );
not ( n16035 , n16034 );
buf ( n16036 , n13319 );
and ( n16037 , n16035 , n16036 );
buf ( n16038 , n15559 );
not ( n16039 , n16038 );
buf ( n16040 , n13331 );
and ( n16041 , n16039 , n16040 );
buf ( n16042 , n15581 );
not ( n16043 , n16042 );
buf ( n16044 , n13343 );
and ( n16045 , n16043 , n16044 );
buf ( n16046 , n15603 );
not ( n16047 , n16046 );
buf ( n16048 , n13355 );
and ( n16049 , n16047 , n16048 );
buf ( n16050 , n15625 );
not ( n16051 , n16050 );
buf ( n16052 , n13367 );
and ( n16053 , n16051 , n16052 );
buf ( n16054 , n15647 );
not ( n16055 , n16054 );
buf ( n16056 , n13379 );
and ( n16057 , n16055 , n16056 );
buf ( n16058 , n15669 );
not ( n16059 , n16058 );
buf ( n16060 , n13391 );
and ( n16061 , n16059 , n16060 );
buf ( n16062 , n15691 );
not ( n16063 , n16062 );
buf ( n16064 , n13403 );
and ( n16065 , n16063 , n16064 );
buf ( n16066 , n15713 );
not ( n16067 , n16066 );
buf ( n16068 , n13415 );
and ( n16069 , n16067 , n16068 );
buf ( n16070 , n15735 );
not ( n16071 , n16070 );
buf ( n16072 , n13427 );
and ( n16073 , n16071 , n16072 );
buf ( n16074 , n15757 );
not ( n16075 , n16074 );
buf ( n16076 , n13439 );
and ( n16077 , n16075 , n16076 );
buf ( n16078 , n15779 );
not ( n16079 , n16078 );
buf ( n16080 , n13451 );
and ( n16081 , n16079 , n16080 );
buf ( n16082 , n15801 );
not ( n16083 , n16082 );
buf ( n16084 , n13463 );
and ( n16085 , n16083 , n16084 );
buf ( n16086 , n15823 );
not ( n16087 , n16086 );
buf ( n16088 , n13480 );
and ( n16089 , n16087 , n16088 );
buf ( n16090 , n15845 );
not ( n16091 , n16090 );
buf ( n16092 , n13497 );
and ( n16093 , n16091 , n16092 );
buf ( n16094 , n15866 );
not ( n16095 , n16094 );
buf ( n16096 , n13514 );
and ( n16097 , n16095 , n16096 );
xnor ( n16098 , n16092 , n16090 );
and ( n16099 , n16097 , n16098 );
or ( n16100 , n16093 , n16099 );
xnor ( n16101 , n16088 , n16086 );
and ( n16102 , n16100 , n16101 );
or ( n16103 , n16089 , n16102 );
xnor ( n16104 , n16084 , n16082 );
and ( n16105 , n16103 , n16104 );
or ( n16106 , n16085 , n16105 );
xnor ( n16107 , n16080 , n16078 );
and ( n16108 , n16106 , n16107 );
or ( n16109 , n16081 , n16108 );
xnor ( n16110 , n16076 , n16074 );
and ( n16111 , n16109 , n16110 );
or ( n16112 , n16077 , n16111 );
xnor ( n16113 , n16072 , n16070 );
and ( n16114 , n16112 , n16113 );
or ( n16115 , n16073 , n16114 );
xnor ( n16116 , n16068 , n16066 );
and ( n16117 , n16115 , n16116 );
or ( n16118 , n16069 , n16117 );
xnor ( n16119 , n16064 , n16062 );
and ( n16120 , n16118 , n16119 );
or ( n16121 , n16065 , n16120 );
xnor ( n16122 , n16060 , n16058 );
and ( n16123 , n16121 , n16122 );
or ( n16124 , n16061 , n16123 );
xnor ( n16125 , n16056 , n16054 );
and ( n16126 , n16124 , n16125 );
or ( n16127 , n16057 , n16126 );
xnor ( n16128 , n16052 , n16050 );
and ( n16129 , n16127 , n16128 );
or ( n16130 , n16053 , n16129 );
xnor ( n16131 , n16048 , n16046 );
and ( n16132 , n16130 , n16131 );
or ( n16133 , n16049 , n16132 );
xnor ( n16134 , n16044 , n16042 );
and ( n16135 , n16133 , n16134 );
or ( n16136 , n16045 , n16135 );
xnor ( n16137 , n16040 , n16038 );
and ( n16138 , n16136 , n16137 );
or ( n16139 , n16041 , n16138 );
xnor ( n16140 , n16036 , n16034 );
and ( n16141 , n16139 , n16140 );
or ( n16142 , n16037 , n16141 );
xnor ( n16143 , n16032 , n16030 );
and ( n16144 , n16142 , n16143 );
or ( n16145 , n16033 , n16144 );
xnor ( n16146 , n16028 , n16026 );
and ( n16147 , n16145 , n16146 );
or ( n16148 , n16029 , n16147 );
xnor ( n16149 , n16024 , n16022 );
and ( n16150 , n16148 , n16149 );
or ( n16151 , n16025 , n16150 );
xnor ( n16152 , n16020 , n16018 );
and ( n16153 , n16151 , n16152 );
or ( n16154 , n16021 , n16153 );
xnor ( n16155 , n16016 , n16014 );
and ( n16156 , n16154 , n16155 );
or ( n16157 , n16017 , n16156 );
xnor ( n16158 , n16012 , n16010 );
and ( n16159 , n16157 , n16158 );
or ( n16160 , n16013 , n16159 );
xnor ( n16161 , n16008 , n16006 );
and ( n16162 , n16160 , n16161 );
or ( n16163 , n16009 , n16162 );
xnor ( n16164 , n16004 , n16002 );
and ( n16165 , n16163 , n16164 );
or ( n16166 , n16005 , n16165 );
xnor ( n16167 , n16000 , n15998 );
and ( n16168 , n16166 , n16167 );
or ( n16169 , n16001 , n16168 );
xnor ( n16170 , n15996 , n15994 );
and ( n16171 , n16169 , n16170 );
or ( n16172 , n15997 , n16171 );
xnor ( n16173 , n15992 , n15990 );
and ( n16174 , n16172 , n16173 );
or ( n16175 , n15993 , n16174 );
xnor ( n16176 , n15988 , n15986 );
and ( n16177 , n16175 , n16176 );
or ( n16178 , n15989 , n16177 );
xnor ( n16179 , n15984 , n15982 );
and ( n16180 , n16178 , n16179 );
or ( n16181 , n15985 , n16180 );
xnor ( n16182 , n15980 , n15978 );
and ( n16183 , n16181 , n16182 );
or ( n16184 , n15981 , n16183 );
xnor ( n16185 , n15976 , n15974 );
and ( n16186 , n16184 , n16185 );
or ( n16187 , n15977 , n16186 );
and ( n16188 , n15973 , n16187 );
not ( n16189 , n15970 );
and ( n16190 , n16189 , n15971 );
and ( n16191 , n16190 , n15972 );
or ( n16192 , n16188 , n16191 );
buf ( n16193 , n16192 );
or ( n16194 , n16193 , n14139 );
and ( n16195 , n16194 , n14588 );
not ( n16196 , n16193 );
or ( n16197 , n16196 , n14139 );
and ( n16198 , n16197 , n14562 );
buf ( n16199 , n13150 );
buf ( n16200 , n14934 );
xor ( n16201 , n16199 , n16200 );
buf ( n16202 , n14611 );
buf ( n16203 , n14952 );
xor ( n16204 , n16202 , n16203 );
or ( n16205 , n16201 , n16204 );
buf ( n16206 , n14964 );
buf ( n16207 , n14977 );
xor ( n16208 , n16206 , n16207 );
or ( n16209 , n16205 , n16208 );
buf ( n16210 , n13162 );
buf ( n16211 , n14992 );
xor ( n16212 , n16210 , n16211 );
or ( n16213 , n16209 , n16212 );
buf ( n16214 , n13175 );
buf ( n16215 , n15007 );
xor ( n16216 , n16214 , n16215 );
or ( n16217 , n16213 , n16216 );
buf ( n16218 , n13187 );
buf ( n16219 , n15022 );
xor ( n16220 , n16218 , n16219 );
or ( n16221 , n16217 , n16220 );
buf ( n16222 , n13199 );
buf ( n16223 , n15037 );
xor ( n16224 , n16222 , n16223 );
or ( n16225 , n16221 , n16224 );
buf ( n16226 , n13211 );
buf ( n16227 , n15052 );
xor ( n16228 , n16226 , n16227 );
or ( n16229 , n16225 , n16228 );
buf ( n16230 , n13223 );
buf ( n16231 , n15067 );
xor ( n16232 , n16230 , n16231 );
or ( n16233 , n16229 , n16232 );
buf ( n16234 , n13235 );
buf ( n16235 , n15082 );
xor ( n16236 , n16234 , n16235 );
or ( n16237 , n16233 , n16236 );
buf ( n16238 , n13247 );
buf ( n16239 , n15097 );
xor ( n16240 , n16238 , n16239 );
or ( n16241 , n16237 , n16240 );
buf ( n16242 , n13259 );
buf ( n16243 , n15112 );
xor ( n16244 , n16242 , n16243 );
or ( n16245 , n16241 , n16244 );
buf ( n16246 , n13271 );
buf ( n16247 , n15449 );
xor ( n16248 , n16246 , n16247 );
or ( n16249 , n16245 , n16248 );
buf ( n16250 , n13283 );
buf ( n16251 , n15471 );
xor ( n16252 , n16250 , n16251 );
or ( n16253 , n16249 , n16252 );
buf ( n16254 , n13295 );
buf ( n16255 , n15493 );
xor ( n16256 , n16254 , n16255 );
or ( n16257 , n16253 , n16256 );
buf ( n16258 , n13307 );
buf ( n16259 , n15515 );
xor ( n16260 , n16258 , n16259 );
or ( n16261 , n16257 , n16260 );
buf ( n16262 , n13319 );
buf ( n16263 , n15537 );
xor ( n16264 , n16262 , n16263 );
or ( n16265 , n16261 , n16264 );
buf ( n16266 , n13331 );
buf ( n16267 , n15559 );
xor ( n16268 , n16266 , n16267 );
or ( n16269 , n16265 , n16268 );
buf ( n16270 , n13343 );
buf ( n16271 , n15581 );
xor ( n16272 , n16270 , n16271 );
or ( n16273 , n16269 , n16272 );
buf ( n16274 , n13355 );
buf ( n16275 , n15603 );
xor ( n16276 , n16274 , n16275 );
or ( n16277 , n16273 , n16276 );
buf ( n16278 , n13367 );
buf ( n16279 , n15625 );
xor ( n16280 , n16278 , n16279 );
or ( n16281 , n16277 , n16280 );
buf ( n16282 , n13379 );
buf ( n16283 , n15647 );
xor ( n16284 , n16282 , n16283 );
or ( n16285 , n16281 , n16284 );
buf ( n16286 , n13391 );
buf ( n16287 , n15669 );
xor ( n16288 , n16286 , n16287 );
or ( n16289 , n16285 , n16288 );
buf ( n16290 , n13403 );
buf ( n16291 , n15691 );
xor ( n16292 , n16290 , n16291 );
or ( n16293 , n16289 , n16292 );
buf ( n16294 , n13415 );
buf ( n16295 , n15713 );
xor ( n16296 , n16294 , n16295 );
or ( n16297 , n16293 , n16296 );
buf ( n16298 , n13427 );
buf ( n16299 , n15735 );
xor ( n16300 , n16298 , n16299 );
or ( n16301 , n16297 , n16300 );
buf ( n16302 , n13439 );
buf ( n16303 , n15757 );
xor ( n16304 , n16302 , n16303 );
or ( n16305 , n16301 , n16304 );
buf ( n16306 , n13451 );
buf ( n16307 , n15779 );
xor ( n16308 , n16306 , n16307 );
or ( n16309 , n16305 , n16308 );
buf ( n16310 , n13463 );
buf ( n16311 , n15801 );
xor ( n16312 , n16310 , n16311 );
or ( n16313 , n16309 , n16312 );
buf ( n16314 , n13480 );
buf ( n16315 , n15823 );
xor ( n16316 , n16314 , n16315 );
or ( n16317 , n16313 , n16316 );
buf ( n16318 , n13497 );
buf ( n16319 , n15845 );
xor ( n16320 , n16318 , n16319 );
or ( n16321 , n16317 , n16320 );
buf ( n16322 , n13514 );
buf ( n16323 , n15866 );
xor ( n16324 , n16322 , n16323 );
or ( n16325 , n16321 , n16324 );
not ( n16326 , n16325 );
buf ( n16327 , n16326 );
not ( n16328 , n16327 );
or ( n16329 , n16328 , n14139 );
and ( n16330 , n16329 , n14586 );
or ( n16331 , n16327 , n14139 );
and ( n16332 , n16331 , n14584 );
buf ( n16333 , n13150 );
buf ( n16334 , n14934 );
xor ( n16335 , n16333 , n16334 );
not ( n16336 , n16335 );
buf ( n16337 , n14611 );
not ( n16338 , n16337 );
buf ( n16339 , n14952 );
and ( n16340 , n16338 , n16339 );
buf ( n16341 , n14964 );
not ( n16342 , n16341 );
buf ( n16343 , n14977 );
and ( n16344 , n16342 , n16343 );
buf ( n16345 , n13162 );
not ( n16346 , n16345 );
buf ( n16347 , n14992 );
and ( n16348 , n16346 , n16347 );
buf ( n16349 , n13175 );
not ( n16350 , n16349 );
buf ( n16351 , n15007 );
and ( n16352 , n16350 , n16351 );
buf ( n16353 , n13187 );
not ( n16354 , n16353 );
buf ( n16355 , n15022 );
and ( n16356 , n16354 , n16355 );
buf ( n16357 , n13199 );
not ( n16358 , n16357 );
buf ( n16359 , n15037 );
and ( n16360 , n16358 , n16359 );
buf ( n16361 , n13211 );
not ( n16362 , n16361 );
buf ( n16363 , n15052 );
and ( n16364 , n16362 , n16363 );
buf ( n16365 , n13223 );
not ( n16366 , n16365 );
buf ( n16367 , n15067 );
and ( n16368 , n16366 , n16367 );
buf ( n16369 , n13235 );
not ( n16370 , n16369 );
buf ( n16371 , n15082 );
and ( n16372 , n16370 , n16371 );
buf ( n16373 , n13247 );
not ( n16374 , n16373 );
buf ( n16375 , n15097 );
and ( n16376 , n16374 , n16375 );
buf ( n16377 , n13259 );
not ( n16378 , n16377 );
buf ( n16379 , n15112 );
and ( n16380 , n16378 , n16379 );
buf ( n16381 , n13271 );
not ( n16382 , n16381 );
buf ( n16383 , n15449 );
and ( n16384 , n16382 , n16383 );
buf ( n16385 , n13283 );
not ( n16386 , n16385 );
buf ( n16387 , n15471 );
and ( n16388 , n16386 , n16387 );
buf ( n16389 , n13295 );
not ( n16390 , n16389 );
buf ( n16391 , n15493 );
and ( n16392 , n16390 , n16391 );
buf ( n16393 , n13307 );
not ( n16394 , n16393 );
buf ( n16395 , n15515 );
and ( n16396 , n16394 , n16395 );
buf ( n16397 , n13319 );
not ( n16398 , n16397 );
buf ( n16399 , n15537 );
and ( n16400 , n16398 , n16399 );
buf ( n16401 , n13331 );
not ( n16402 , n16401 );
buf ( n16403 , n15559 );
and ( n16404 , n16402 , n16403 );
buf ( n16405 , n13343 );
not ( n16406 , n16405 );
buf ( n16407 , n15581 );
and ( n16408 , n16406 , n16407 );
buf ( n16409 , n13355 );
not ( n16410 , n16409 );
buf ( n16411 , n15603 );
and ( n16412 , n16410 , n16411 );
buf ( n16413 , n13367 );
not ( n16414 , n16413 );
buf ( n16415 , n15625 );
and ( n16416 , n16414 , n16415 );
buf ( n16417 , n13379 );
not ( n16418 , n16417 );
buf ( n16419 , n15647 );
and ( n16420 , n16418 , n16419 );
buf ( n16421 , n13391 );
not ( n16422 , n16421 );
buf ( n16423 , n15669 );
and ( n16424 , n16422 , n16423 );
buf ( n16425 , n13403 );
not ( n16426 , n16425 );
buf ( n16427 , n15691 );
and ( n16428 , n16426 , n16427 );
buf ( n16429 , n13415 );
not ( n16430 , n16429 );
buf ( n16431 , n15713 );
and ( n16432 , n16430 , n16431 );
buf ( n16433 , n13427 );
not ( n16434 , n16433 );
buf ( n16435 , n15735 );
and ( n16436 , n16434 , n16435 );
buf ( n16437 , n13439 );
not ( n16438 , n16437 );
buf ( n16439 , n15757 );
and ( n16440 , n16438 , n16439 );
buf ( n16441 , n13451 );
not ( n16442 , n16441 );
buf ( n16443 , n15779 );
and ( n16444 , n16442 , n16443 );
buf ( n16445 , n13463 );
not ( n16446 , n16445 );
buf ( n16447 , n15801 );
and ( n16448 , n16446 , n16447 );
buf ( n16449 , n13480 );
not ( n16450 , n16449 );
buf ( n16451 , n15823 );
and ( n16452 , n16450 , n16451 );
buf ( n16453 , n13497 );
not ( n16454 , n16453 );
buf ( n16455 , n15845 );
and ( n16456 , n16454 , n16455 );
buf ( n16457 , n13514 );
not ( n16458 , n16457 );
buf ( n16459 , n15866 );
and ( n16460 , n16458 , n16459 );
xnor ( n16461 , n16453 , n16455 );
and ( n16462 , n16460 , n16461 );
or ( n16463 , n16456 , n16462 );
xnor ( n16464 , n16449 , n16451 );
and ( n16465 , n16463 , n16464 );
or ( n16466 , n16452 , n16465 );
xnor ( n16467 , n16445 , n16447 );
and ( n16468 , n16466 , n16467 );
or ( n16469 , n16448 , n16468 );
xnor ( n16470 , n16441 , n16443 );
and ( n16471 , n16469 , n16470 );
or ( n16472 , n16444 , n16471 );
xnor ( n16473 , n16437 , n16439 );
and ( n16474 , n16472 , n16473 );
or ( n16475 , n16440 , n16474 );
xnor ( n16476 , n16433 , n16435 );
and ( n16477 , n16475 , n16476 );
or ( n16478 , n16436 , n16477 );
xnor ( n16479 , n16429 , n16431 );
and ( n16480 , n16478 , n16479 );
or ( n16481 , n16432 , n16480 );
xnor ( n16482 , n16425 , n16427 );
and ( n16483 , n16481 , n16482 );
or ( n16484 , n16428 , n16483 );
xnor ( n16485 , n16421 , n16423 );
and ( n16486 , n16484 , n16485 );
or ( n16487 , n16424 , n16486 );
xnor ( n16488 , n16417 , n16419 );
and ( n16489 , n16487 , n16488 );
or ( n16490 , n16420 , n16489 );
xnor ( n16491 , n16413 , n16415 );
and ( n16492 , n16490 , n16491 );
or ( n16493 , n16416 , n16492 );
xnor ( n16494 , n16409 , n16411 );
and ( n16495 , n16493 , n16494 );
or ( n16496 , n16412 , n16495 );
xnor ( n16497 , n16405 , n16407 );
and ( n16498 , n16496 , n16497 );
or ( n16499 , n16408 , n16498 );
xnor ( n16500 , n16401 , n16403 );
and ( n16501 , n16499 , n16500 );
or ( n16502 , n16404 , n16501 );
xnor ( n16503 , n16397 , n16399 );
and ( n16504 , n16502 , n16503 );
or ( n16505 , n16400 , n16504 );
xnor ( n16506 , n16393 , n16395 );
and ( n16507 , n16505 , n16506 );
or ( n16508 , n16396 , n16507 );
xnor ( n16509 , n16389 , n16391 );
and ( n16510 , n16508 , n16509 );
or ( n16511 , n16392 , n16510 );
xnor ( n16512 , n16385 , n16387 );
and ( n16513 , n16511 , n16512 );
or ( n16514 , n16388 , n16513 );
xnor ( n16515 , n16381 , n16383 );
and ( n16516 , n16514 , n16515 );
or ( n16517 , n16384 , n16516 );
xnor ( n16518 , n16377 , n16379 );
and ( n16519 , n16517 , n16518 );
or ( n16520 , n16380 , n16519 );
xnor ( n16521 , n16373 , n16375 );
and ( n16522 , n16520 , n16521 );
or ( n16523 , n16376 , n16522 );
xnor ( n16524 , n16369 , n16371 );
and ( n16525 , n16523 , n16524 );
or ( n16526 , n16372 , n16525 );
xnor ( n16527 , n16365 , n16367 );
and ( n16528 , n16526 , n16527 );
or ( n16529 , n16368 , n16528 );
xnor ( n16530 , n16361 , n16363 );
and ( n16531 , n16529 , n16530 );
or ( n16532 , n16364 , n16531 );
xnor ( n16533 , n16357 , n16359 );
and ( n16534 , n16532 , n16533 );
or ( n16535 , n16360 , n16534 );
xnor ( n16536 , n16353 , n16355 );
and ( n16537 , n16535 , n16536 );
or ( n16538 , n16356 , n16537 );
xnor ( n16539 , n16349 , n16351 );
and ( n16540 , n16538 , n16539 );
or ( n16541 , n16352 , n16540 );
xnor ( n16542 , n16345 , n16347 );
and ( n16543 , n16541 , n16542 );
or ( n16544 , n16348 , n16543 );
xnor ( n16545 , n16341 , n16343 );
and ( n16546 , n16544 , n16545 );
or ( n16547 , n16344 , n16546 );
xnor ( n16548 , n16337 , n16339 );
and ( n16549 , n16547 , n16548 );
or ( n16550 , n16340 , n16549 );
and ( n16551 , n16336 , n16550 );
not ( n16552 , n16334 );
and ( n16553 , n16552 , n16333 );
and ( n16554 , n16553 , n16335 );
or ( n16555 , n16551 , n16554 );
buf ( n16556 , n16555 );
not ( n16557 , n16556 );
or ( n16558 , n16557 , n14139 );
and ( n16559 , n16558 , n14582 );
or ( n16560 , n16556 , n14139 );
and ( n16561 , n16560 , n14580 );
and ( n16562 , n15965 , n14578 );
and ( n16563 , n15964 , n14576 );
and ( n16564 , n16193 , n14574 );
and ( n16565 , n16196 , n14572 );
and ( n16566 , n16328 , n14569 );
and ( n16567 , n16327 , n14567 );
and ( n16568 , n16557 , n14564 );
and ( n16569 , n16556 , n14565 );
or ( n16570 , n15967 , n15969 , n16195 , n16198 , n16330 , n16332 , n16559 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 );
and ( n16571 , n16570 , n11954 );
or ( n16572 , n14599 , n16571 );
buf ( n16573 , RI2106be58_607);
buf ( n16574 , n16573 );
and ( n16575 , n16572 , n16574 );
not ( n16576 , n16573 );
and ( n16577 , n14139 , n16576 );
or ( n16578 , n16575 , n16577 );
buf ( n16579 , n16578 );
buf ( n16580 , n16579 );
buf ( n16581 , n10613 );
buf ( n16582 , RI21a14440_60);
buf ( n16583 , n16582 );
not ( n16584 , n16583 );
buf ( n16585 , RI21a144b8_59);
buf ( n16586 , n16585 );
not ( n16587 , n16586 );
buf ( n16588 , RI21a145a8_57);
buf ( n16589 , n16588 );
not ( n16590 , n16589 );
buf ( n16591 , RI21a14cb0_56);
buf ( n16592 , n16591 );
not ( n16593 , n16592 );
buf ( n16594 , RI21a14d28_55);
buf ( n16595 , n16594 );
not ( n16596 , n16595 );
buf ( n16597 , RI21a14da0_54);
buf ( n16598 , n16597 );
not ( n16599 , n16598 );
buf ( n16600 , RI21a14e18_53);
buf ( n16601 , n16600 );
not ( n16602 , n16601 );
buf ( n16603 , RI21a14e90_52);
buf ( n16604 , n16603 );
not ( n16605 , n16604 );
buf ( n16606 , RI21a14f08_51);
buf ( n16607 , n16606 );
not ( n16608 , n16607 );
buf ( n16609 , RI21a15610_50);
buf ( n16610 , n16609 );
not ( n16611 , n16610 );
buf ( n16612 , RI21a15688_49);
buf ( n16613 , n16612 );
not ( n16614 , n16613 );
buf ( n16615 , RI21a15700_48);
buf ( n16616 , n16615 );
not ( n16617 , n16616 );
buf ( n16618 , RI21a157f0_46);
buf ( n16619 , n16618 );
not ( n16620 , n16619 );
buf ( n16621 , RI21a15868_45);
buf ( n16622 , n16621 );
not ( n16623 , n16622 );
buf ( n16624 , RI21a15f70_44);
buf ( n16625 , n16624 );
not ( n16626 , n16625 );
buf ( n16627 , RI21a15fe8_43);
buf ( n16628 , n16627 );
not ( n16629 , n16628 );
buf ( n16630 , RI21a16060_42);
buf ( n16631 , n16630 );
not ( n16632 , n16631 );
buf ( n16633 , RI21a160d8_41);
buf ( n16634 , n16633 );
not ( n16635 , n16634 );
buf ( n16636 , RI21a16150_40);
buf ( n16637 , n16636 );
not ( n16638 , n16637 );
buf ( n16639 , RI21a161c8_39);
buf ( n16640 , n16639 );
not ( n16641 , n16640 );
buf ( n16642 , RI21a168d0_38);
buf ( n16643 , n16642 );
not ( n16644 , n16643 );
buf ( n16645 , RI21a16948_37);
buf ( n16646 , n16645 );
not ( n16647 , n16646 );
buf ( n16648 , RI21a13a68_67);
buf ( n16649 , n16648 );
not ( n16650 , n16649 );
buf ( n16651 , RI21a13ae0_66);
buf ( n16652 , n16651 );
not ( n16653 , n16652 );
buf ( n16654 , RI21a13b58_65);
buf ( n16655 , n16654 );
not ( n16656 , n16655 );
buf ( n16657 , RI21a13bd0_64);
buf ( n16658 , n16657 );
not ( n16659 , n16658 );
buf ( n16660 , RI21a13c48_63);
buf ( n16661 , n16660 );
not ( n16662 , n16661 );
buf ( n16663 , RI21a14350_62);
buf ( n16664 , n16663 );
not ( n16665 , n16664 );
buf ( n16666 , RI21a143c8_61);
buf ( n16667 , n16666 );
not ( n16668 , n16667 );
buf ( n16669 , RI21a14530_58);
buf ( n16670 , n16669 );
not ( n16671 , n16670 );
buf ( n16672 , RI21a15778_47);
buf ( n16673 , n16672 );
not ( n16674 , n16673 );
buf ( n16675 , RI21a169c0_36);
buf ( n16676 , n16675 );
not ( n16677 , n16676 );
and ( n16678 , n16674 , n16677 );
and ( n16679 , n16671 , n16678 );
and ( n16680 , n16668 , n16679 );
and ( n16681 , n16665 , n16680 );
and ( n16682 , n16662 , n16681 );
and ( n16683 , n16659 , n16682 );
and ( n16684 , n16656 , n16683 );
and ( n16685 , n16653 , n16684 );
and ( n16686 , n16650 , n16685 );
and ( n16687 , n16647 , n16686 );
and ( n16688 , n16644 , n16687 );
and ( n16689 , n16641 , n16688 );
and ( n16690 , n16638 , n16689 );
and ( n16691 , n16635 , n16690 );
and ( n16692 , n16632 , n16691 );
and ( n16693 , n16629 , n16692 );
and ( n16694 , n16626 , n16693 );
and ( n16695 , n16623 , n16694 );
and ( n16696 , n16620 , n16695 );
and ( n16697 , n16617 , n16696 );
and ( n16698 , n16614 , n16697 );
and ( n16699 , n16611 , n16698 );
and ( n16700 , n16608 , n16699 );
and ( n16701 , n16605 , n16700 );
and ( n16702 , n16602 , n16701 );
and ( n16703 , n16599 , n16702 );
and ( n16704 , n16596 , n16703 );
and ( n16705 , n16593 , n16704 );
and ( n16706 , n16590 , n16705 );
and ( n16707 , n16587 , n16706 );
xor ( n16708 , n16584 , n16707 );
buf ( n16709 , n16708 );
buf ( n16710 , n16582 );
and ( n16711 , n16709 , n16710 );
or ( n16712 , C0 , n16711 );
buf ( n16713 , n16712 );
not ( n16714 , n16713 );
not ( n16715 , n16710 );
and ( n16716 , n16715 , n16606 );
xor ( n16717 , n16608 , n16699 );
buf ( n16718 , n16717 );
and ( n16719 , n16718 , n16710 );
or ( n16720 , n16716 , n16719 );
buf ( n16721 , n16720 );
and ( n16722 , n16714 , n16721 );
not ( n16723 , n16721 );
not ( n16724 , n16710 );
and ( n16725 , n16724 , n16609 );
xor ( n16726 , n16611 , n16698 );
buf ( n16727 , n16726 );
and ( n16728 , n16727 , n16710 );
or ( n16729 , n16725 , n16728 );
buf ( n16730 , n16729 );
not ( n16731 , n16730 );
not ( n16732 , n16710 );
and ( n16733 , n16732 , n16612 );
xor ( n16734 , n16614 , n16697 );
buf ( n16735 , n16734 );
and ( n16736 , n16735 , n16710 );
or ( n16737 , n16733 , n16736 );
buf ( n16738 , n16737 );
not ( n16739 , n16738 );
not ( n16740 , n16710 );
and ( n16741 , n16740 , n16615 );
xor ( n16742 , n16617 , n16696 );
buf ( n16743 , n16742 );
and ( n16744 , n16743 , n16710 );
or ( n16745 , n16741 , n16744 );
buf ( n16746 , n16745 );
not ( n16747 , n16746 );
not ( n16748 , n16710 );
and ( n16749 , n16748 , n16618 );
xor ( n16750 , n16620 , n16695 );
buf ( n16751 , n16750 );
and ( n16752 , n16751 , n16710 );
or ( n16753 , n16749 , n16752 );
buf ( n16754 , n16753 );
not ( n16755 , n16754 );
not ( n16756 , n16710 );
and ( n16757 , n16756 , n16621 );
xor ( n16758 , n16623 , n16694 );
buf ( n16759 , n16758 );
and ( n16760 , n16759 , n16710 );
or ( n16761 , n16757 , n16760 );
buf ( n16762 , n16761 );
not ( n16763 , n16762 );
not ( n16764 , n16710 );
and ( n16765 , n16764 , n16624 );
xor ( n16766 , n16626 , n16693 );
buf ( n16767 , n16766 );
and ( n16768 , n16767 , n16710 );
or ( n16769 , n16765 , n16768 );
buf ( n16770 , n16769 );
not ( n16771 , n16770 );
not ( n16772 , n16710 );
and ( n16773 , n16772 , n16627 );
xor ( n16774 , n16629 , n16692 );
buf ( n16775 , n16774 );
and ( n16776 , n16775 , n16710 );
or ( n16777 , n16773 , n16776 );
buf ( n16778 , n16777 );
not ( n16779 , n16778 );
not ( n16780 , n16710 );
and ( n16781 , n16780 , n16630 );
xor ( n16782 , n16632 , n16691 );
buf ( n16783 , n16782 );
and ( n16784 , n16783 , n16710 );
or ( n16785 , n16781 , n16784 );
buf ( n16786 , n16785 );
not ( n16787 , n16786 );
not ( n16788 , n16710 );
and ( n16789 , n16788 , n16633 );
xor ( n16790 , n16635 , n16690 );
buf ( n16791 , n16790 );
and ( n16792 , n16791 , n16710 );
or ( n16793 , n16789 , n16792 );
buf ( n16794 , n16793 );
not ( n16795 , n16794 );
not ( n16796 , n16710 );
and ( n16797 , n16796 , n16636 );
xor ( n16798 , n16638 , n16689 );
buf ( n16799 , n16798 );
and ( n16800 , n16799 , n16710 );
or ( n16801 , n16797 , n16800 );
buf ( n16802 , n16801 );
not ( n16803 , n16802 );
not ( n16804 , n16710 );
and ( n16805 , n16804 , n16639 );
xor ( n16806 , n16641 , n16688 );
buf ( n16807 , n16806 );
and ( n16808 , n16807 , n16710 );
or ( n16809 , n16805 , n16808 );
buf ( n16810 , n16809 );
not ( n16811 , n16810 );
not ( n16812 , n16710 );
and ( n16813 , n16812 , n16642 );
xor ( n16814 , n16644 , n16687 );
buf ( n16815 , n16814 );
and ( n16816 , n16815 , n16710 );
or ( n16817 , n16813 , n16816 );
buf ( n16818 , n16817 );
not ( n16819 , n16818 );
not ( n16820 , n16710 );
and ( n16821 , n16820 , n16645 );
xor ( n16822 , n16647 , n16686 );
buf ( n16823 , n16822 );
and ( n16824 , n16823 , n16710 );
or ( n16825 , n16821 , n16824 );
buf ( n16826 , n16825 );
not ( n16827 , n16826 );
not ( n16828 , n16710 );
and ( n16829 , n16828 , n16648 );
xor ( n16830 , n16650 , n16685 );
buf ( n16831 , n16830 );
and ( n16832 , n16831 , n16710 );
or ( n16833 , n16829 , n16832 );
buf ( n16834 , n16833 );
not ( n16835 , n16834 );
not ( n16836 , n16710 );
and ( n16837 , n16836 , n16651 );
xor ( n16838 , n16653 , n16684 );
buf ( n16839 , n16838 );
and ( n16840 , n16839 , n16710 );
or ( n16841 , n16837 , n16840 );
buf ( n16842 , n16841 );
not ( n16843 , n16842 );
not ( n16844 , n16710 );
and ( n16845 , n16844 , n16654 );
xor ( n16846 , n16656 , n16683 );
buf ( n16847 , n16846 );
and ( n16848 , n16847 , n16710 );
or ( n16849 , n16845 , n16848 );
buf ( n16850 , n16849 );
not ( n16851 , n16850 );
not ( n16852 , n16710 );
and ( n16853 , n16852 , n16657 );
xor ( n16854 , n16659 , n16682 );
buf ( n16855 , n16854 );
and ( n16856 , n16855 , n16710 );
or ( n16857 , n16853 , n16856 );
buf ( n16858 , n16857 );
not ( n16859 , n16858 );
not ( n16860 , n16710 );
and ( n16861 , n16860 , n16660 );
xor ( n16862 , n16662 , n16681 );
buf ( n16863 , n16862 );
and ( n16864 , n16863 , n16710 );
or ( n16865 , n16861 , n16864 );
buf ( n16866 , n16865 );
not ( n16867 , n16866 );
not ( n16868 , n16710 );
and ( n16869 , n16868 , n16663 );
xor ( n16870 , n16665 , n16680 );
buf ( n16871 , n16870 );
and ( n16872 , n16871 , n16710 );
or ( n16873 , n16869 , n16872 );
buf ( n16874 , n16873 );
not ( n16875 , n16874 );
not ( n16876 , n16710 );
and ( n16877 , n16876 , n16666 );
xor ( n16878 , n16668 , n16679 );
buf ( n16879 , n16878 );
and ( n16880 , n16879 , n16710 );
or ( n16881 , n16877 , n16880 );
buf ( n16882 , n16881 );
not ( n16883 , n16882 );
not ( n16884 , n16710 );
and ( n16885 , n16884 , n16669 );
xor ( n16886 , n16671 , n16678 );
buf ( n16887 , n16886 );
and ( n16888 , n16887 , n16710 );
or ( n16889 , n16885 , n16888 );
buf ( n16890 , n16889 );
not ( n16891 , n16890 );
not ( n16892 , n16710 );
and ( n16893 , n16892 , n16672 );
xor ( n16894 , n16674 , n16677 );
buf ( n16895 , n16894 );
and ( n16896 , n16895 , n16710 );
or ( n16897 , n16893 , n16896 );
buf ( n16898 , n16897 );
not ( n16899 , n16898 );
buf ( n16900 , n16675 );
buf ( n16901 , n16900 );
not ( n16902 , n16901 );
and ( n16903 , n16899 , n16902 );
and ( n16904 , n16891 , n16903 );
and ( n16905 , n16883 , n16904 );
and ( n16906 , n16875 , n16905 );
and ( n16907 , n16867 , n16906 );
and ( n16908 , n16859 , n16907 );
and ( n16909 , n16851 , n16908 );
and ( n16910 , n16843 , n16909 );
and ( n16911 , n16835 , n16910 );
and ( n16912 , n16827 , n16911 );
and ( n16913 , n16819 , n16912 );
and ( n16914 , n16811 , n16913 );
and ( n16915 , n16803 , n16914 );
and ( n16916 , n16795 , n16915 );
and ( n16917 , n16787 , n16916 );
and ( n16918 , n16779 , n16917 );
and ( n16919 , n16771 , n16918 );
and ( n16920 , n16763 , n16919 );
and ( n16921 , n16755 , n16920 );
and ( n16922 , n16747 , n16921 );
and ( n16923 , n16739 , n16922 );
and ( n16924 , n16731 , n16923 );
xor ( n16925 , n16723 , n16924 );
and ( n16926 , n16925 , n16713 );
or ( n16927 , n16722 , n16926 );
buf ( n16928 , n16927 );
not ( n16929 , n16928 );
buf ( n16930 , n16929 );
buf ( n16931 , n16930 );
not ( n16932 , n16931 );
buf ( n16933 , n16932 );
buf ( n16934 , n16933 );
not ( n16935 , n16934 );
buf ( n16936 , n16935 );
buf ( n16937 , n16936 );
not ( n16938 , n16937 );
or ( n16939 , n16938 , C0 );
or ( n16940 , n16939 , C0 );
or ( n16941 , n16940 , C0 );
or ( n16942 , n16941 , C0 );
or ( n16943 , n16942 , C0 );
or ( n16944 , n16943 , C0 );
or ( n16945 , n16944 , C0 );
or ( n16946 , n16945 , C0 );
or ( n16947 , n16946 , C0 );
or ( n16948 , n16947 , C0 );
or ( n16949 , n16948 , C0 );
or ( n16950 , n16949 , C0 );
or ( n16951 , n16950 , C0 );
or ( n16952 , n16951 , C0 );
or ( n16953 , n16952 , C0 );
or ( n16954 , n16953 , C0 );
or ( n16955 , n16954 , C0 );
or ( n16956 , n16955 , C0 );
or ( n16957 , n16956 , C0 );
or ( n16958 , n16957 , C0 );
or ( n16959 , n16958 , C0 );
or ( n16960 , n16959 , C0 );
or ( n16961 , n16960 , C0 );
or ( n16962 , n16961 , C0 );
or ( n16963 , n16962 , C0 );
or ( n16964 , n16963 , C0 );
or ( n16965 , n16964 , C0 );
or ( n16966 , n16965 , C0 );
or ( n16967 , n16966 , C0 );
or ( n16968 , n16967 , C0 );
buf ( n16969 , n16968 );
not ( n16970 , n16713 );
not ( n16971 , n16710 );
and ( n16972 , n16971 , n16585 );
xor ( n16973 , n16587 , n16706 );
buf ( n16974 , n16973 );
and ( n16975 , n16974 , n16710 );
or ( n16976 , n16972 , n16975 );
buf ( n16977 , n16976 );
not ( n16978 , n16977 );
not ( n16979 , n16710 );
and ( n16980 , n16979 , n16588 );
xor ( n16981 , n16590 , n16705 );
buf ( n16982 , n16981 );
and ( n16983 , n16982 , n16710 );
or ( n16984 , n16980 , n16983 );
buf ( n16985 , n16984 );
not ( n16986 , n16985 );
not ( n16987 , n16710 );
and ( n16988 , n16987 , n16591 );
xor ( n16989 , n16593 , n16704 );
buf ( n16990 , n16989 );
and ( n16991 , n16990 , n16710 );
or ( n16992 , n16988 , n16991 );
buf ( n16993 , n16992 );
not ( n16994 , n16993 );
not ( n16995 , n16710 );
and ( n16996 , n16995 , n16594 );
xor ( n16997 , n16596 , n16703 );
buf ( n16998 , n16997 );
and ( n16999 , n16998 , n16710 );
or ( n17000 , n16996 , n16999 );
buf ( n17001 , n17000 );
not ( n17002 , n17001 );
not ( n17003 , n16710 );
and ( n17004 , n17003 , n16597 );
xor ( n17005 , n16599 , n16702 );
buf ( n17006 , n17005 );
and ( n17007 , n17006 , n16710 );
or ( n17008 , n17004 , n17007 );
buf ( n17009 , n17008 );
not ( n17010 , n17009 );
not ( n17011 , n16710 );
and ( n17012 , n17011 , n16600 );
xor ( n17013 , n16602 , n16701 );
buf ( n17014 , n17013 );
and ( n17015 , n17014 , n16710 );
or ( n17016 , n17012 , n17015 );
buf ( n17017 , n17016 );
not ( n17018 , n17017 );
not ( n17019 , n16710 );
and ( n17020 , n17019 , n16603 );
xor ( n17021 , n16605 , n16700 );
buf ( n17022 , n17021 );
and ( n17023 , n17022 , n16710 );
or ( n17024 , n17020 , n17023 );
buf ( n17025 , n17024 );
not ( n17026 , n17025 );
and ( n17027 , n16723 , n16924 );
and ( n17028 , n17026 , n17027 );
and ( n17029 , n17018 , n17028 );
and ( n17030 , n17010 , n17029 );
and ( n17031 , n17002 , n17030 );
and ( n17032 , n16994 , n17031 );
and ( n17033 , n16986 , n17032 );
and ( n17034 , n16978 , n17033 );
xor ( n17035 , n16970 , n17034 );
buf ( n17036 , n16713 );
and ( n17037 , n17035 , n17036 );
or ( n17038 , C0 , n17037 );
buf ( n17039 , n17038 );
not ( n17040 , n17039 );
buf ( n17041 , n17040 );
buf ( n17042 , n17041 );
not ( n17043 , n17042 );
buf ( n17044 , n17043 );
not ( n17045 , n17044 );
buf ( n17046 , n17045 );
not ( n17047 , n16713 );
and ( n17048 , n17047 , n16977 );
xor ( n17049 , n16978 , n17033 );
and ( n17050 , n17049 , n16713 );
or ( n17051 , n17048 , n17050 );
buf ( n17052 , n17051 );
not ( n17053 , n17052 );
buf ( n17054 , n17053 );
buf ( n17055 , n17054 );
not ( n17056 , n17055 );
buf ( n17057 , n17056 );
not ( n17058 , n17057 );
buf ( n17059 , n17058 );
not ( n17060 , n16713 );
and ( n17061 , n17060 , n16985 );
xor ( n17062 , n16986 , n17032 );
and ( n17063 , n17062 , n16713 );
or ( n17064 , n17061 , n17063 );
buf ( n17065 , n17064 );
not ( n17066 , n17065 );
buf ( n17067 , n17066 );
buf ( n17068 , n17067 );
not ( n17069 , n17068 );
buf ( n17070 , n17069 );
not ( n17071 , n17070 );
buf ( n17072 , n17071 );
not ( n17073 , n16713 );
and ( n17074 , n17073 , n16993 );
xor ( n17075 , n16994 , n17031 );
and ( n17076 , n17075 , n16713 );
or ( n17077 , n17074 , n17076 );
buf ( n17078 , n17077 );
not ( n17079 , n17078 );
buf ( n17080 , n17079 );
buf ( n17081 , n17080 );
not ( n17082 , n17081 );
buf ( n17083 , n17082 );
not ( n17084 , n17083 );
buf ( n17085 , n17084 );
not ( n17086 , n16713 );
and ( n17087 , n17086 , n17001 );
xor ( n17088 , n17002 , n17030 );
and ( n17089 , n17088 , n16713 );
or ( n17090 , n17087 , n17089 );
buf ( n17091 , n17090 );
not ( n17092 , n17091 );
buf ( n17093 , n17092 );
buf ( n17094 , n17093 );
not ( n17095 , n17094 );
buf ( n17096 , n17095 );
not ( n17097 , n17096 );
buf ( n17098 , n17097 );
not ( n17099 , n16713 );
and ( n17100 , n17099 , n17009 );
xor ( n17101 , n17010 , n17029 );
and ( n17102 , n17101 , n16713 );
or ( n17103 , n17100 , n17102 );
buf ( n17104 , n17103 );
not ( n17105 , n17104 );
buf ( n17106 , n17105 );
buf ( n17107 , n17106 );
not ( n17108 , n17107 );
buf ( n17109 , n17108 );
not ( n17110 , n17109 );
buf ( n17111 , n17110 );
not ( n17112 , n16713 );
and ( n17113 , n17112 , n17017 );
xor ( n17114 , n17018 , n17028 );
and ( n17115 , n17114 , n16713 );
or ( n17116 , n17113 , n17115 );
buf ( n17117 , n17116 );
not ( n17118 , n17117 );
buf ( n17119 , n17118 );
buf ( n17120 , n17119 );
not ( n17121 , n17120 );
buf ( n17122 , n17121 );
not ( n17123 , n17122 );
buf ( n17124 , n17123 );
not ( n17125 , n16713 );
and ( n17126 , n17125 , n17025 );
xor ( n17127 , n17026 , n17027 );
and ( n17128 , n17127 , n16713 );
or ( n17129 , n17126 , n17128 );
buf ( n17130 , n17129 );
not ( n17131 , n17130 );
buf ( n17132 , n17131 );
buf ( n17133 , n17132 );
not ( n17134 , n17133 );
buf ( n17135 , n17134 );
not ( n17136 , n17135 );
buf ( n17137 , n17136 );
not ( n17138 , n16933 );
buf ( n17139 , n17138 );
and ( n17140 , n17137 , n17139 );
and ( n17141 , n17124 , n17140 );
and ( n17142 , n17111 , n17141 );
and ( n17143 , n17098 , n17142 );
and ( n17144 , n17085 , n17143 );
and ( n17145 , n17072 , n17144 );
and ( n17146 , n17059 , n17145 );
and ( n17147 , n17046 , n17146 );
not ( n17148 , n17147 );
buf ( n17149 , n17148 );
buf ( n17150 , n16713 );
and ( n17151 , n17149 , n17150 );
or ( n17152 , C0 , n17151 );
buf ( n17153 , n17152 );
buf ( n17154 , n17153 );
and ( n17155 , n16969 , n17154 );
not ( n17156 , n17155 );
and ( n17157 , n17156 , n16938 );
xor ( n17158 , n16938 , n17154 );
xor ( n17159 , n17158 , n17154 );
and ( n17160 , n17159 , n17155 );
or ( n17161 , n17157 , n17160 );
buf ( n17162 , n17161 );
buf ( n17163 , n16712 );
not ( n17164 , n17163 );
buf ( n17165 , n17024 );
and ( n17166 , n17164 , n17165 );
not ( n17167 , n17165 );
buf ( n17168 , n16720 );
not ( n17169 , n17168 );
buf ( n17170 , n16729 );
not ( n17171 , n17170 );
buf ( n17172 , n16737 );
not ( n17173 , n17172 );
buf ( n17174 , n16745 );
not ( n17175 , n17174 );
buf ( n17176 , n16753 );
not ( n17177 , n17176 );
buf ( n17178 , n16761 );
not ( n17179 , n17178 );
buf ( n17180 , n16769 );
not ( n17181 , n17180 );
buf ( n17182 , n16777 );
not ( n17183 , n17182 );
buf ( n17184 , n16785 );
not ( n17185 , n17184 );
buf ( n17186 , n16793 );
not ( n17187 , n17186 );
buf ( n17188 , n16801 );
not ( n17189 , n17188 );
buf ( n17190 , n16809 );
not ( n17191 , n17190 );
buf ( n17192 , n16817 );
not ( n17193 , n17192 );
buf ( n17194 , n16825 );
not ( n17195 , n17194 );
buf ( n17196 , n16833 );
not ( n17197 , n17196 );
buf ( n17198 , n16841 );
not ( n17199 , n17198 );
buf ( n17200 , n16849 );
not ( n17201 , n17200 );
buf ( n17202 , n16857 );
not ( n17203 , n17202 );
buf ( n17204 , n16865 );
not ( n17205 , n17204 );
buf ( n17206 , n16873 );
not ( n17207 , n17206 );
buf ( n17208 , n16881 );
not ( n17209 , n17208 );
buf ( n17210 , n16889 );
not ( n17211 , n17210 );
buf ( n17212 , n16897 );
not ( n17213 , n17212 );
buf ( n17214 , n16900 );
not ( n17215 , n17214 );
and ( n17216 , n17213 , n17215 );
and ( n17217 , n17211 , n17216 );
and ( n17218 , n17209 , n17217 );
and ( n17219 , n17207 , n17218 );
and ( n17220 , n17205 , n17219 );
and ( n17221 , n17203 , n17220 );
and ( n17222 , n17201 , n17221 );
and ( n17223 , n17199 , n17222 );
and ( n17224 , n17197 , n17223 );
and ( n17225 , n17195 , n17224 );
and ( n17226 , n17193 , n17225 );
and ( n17227 , n17191 , n17226 );
and ( n17228 , n17189 , n17227 );
and ( n17229 , n17187 , n17228 );
and ( n17230 , n17185 , n17229 );
and ( n17231 , n17183 , n17230 );
and ( n17232 , n17181 , n17231 );
and ( n17233 , n17179 , n17232 );
and ( n17234 , n17177 , n17233 );
and ( n17235 , n17175 , n17234 );
and ( n17236 , n17173 , n17235 );
and ( n17237 , n17171 , n17236 );
and ( n17238 , n17169 , n17237 );
xor ( n17239 , n17167 , n17238 );
and ( n17240 , n17239 , n17163 );
or ( n17241 , n17166 , n17240 );
buf ( n17242 , n17241 );
not ( n17243 , n17242 );
buf ( n17244 , n17243 );
buf ( n17245 , n17244 );
not ( n17246 , n17245 );
buf ( n17247 , n17246 );
buf ( n17248 , n17247 );
buf ( n17249 , n17248 );
not ( n17250 , n17249 );
buf ( n17251 , n17250 );
buf ( n17252 , n17251 );
not ( n17253 , n17252 );
not ( n17254 , n17163 );
buf ( n17255 , n16976 );
not ( n17256 , n17255 );
buf ( n17257 , n16984 );
not ( n17258 , n17257 );
buf ( n17259 , n16992 );
not ( n17260 , n17259 );
buf ( n17261 , n17000 );
not ( n17262 , n17261 );
buf ( n17263 , n17008 );
not ( n17264 , n17263 );
buf ( n17265 , n17016 );
not ( n17266 , n17265 );
and ( n17267 , n17167 , n17238 );
and ( n17268 , n17266 , n17267 );
and ( n17269 , n17264 , n17268 );
and ( n17270 , n17262 , n17269 );
and ( n17271 , n17260 , n17270 );
and ( n17272 , n17258 , n17271 );
and ( n17273 , n17256 , n17272 );
xor ( n17274 , n17254 , n17273 );
buf ( n17275 , n17163 );
and ( n17276 , n17274 , n17275 );
or ( n17277 , C0 , n17276 );
buf ( n17278 , n17277 );
not ( n17279 , n17278 );
buf ( n17280 , n17279 );
buf ( n17281 , n17280 );
not ( n17282 , n17281 );
buf ( n17283 , n17282 );
not ( n17284 , n17283 );
buf ( n17285 , n17284 );
not ( n17286 , n17163 );
and ( n17287 , n17286 , n17255 );
xor ( n17288 , n17256 , n17272 );
and ( n17289 , n17288 , n17163 );
or ( n17290 , n17287 , n17289 );
buf ( n17291 , n17290 );
not ( n17292 , n17291 );
buf ( n17293 , n17292 );
buf ( n17294 , n17293 );
not ( n17295 , n17294 );
buf ( n17296 , n17295 );
not ( n17297 , n17296 );
buf ( n17298 , n17297 );
not ( n17299 , n17163 );
and ( n17300 , n17299 , n17257 );
xor ( n17301 , n17258 , n17271 );
and ( n17302 , n17301 , n17163 );
or ( n17303 , n17300 , n17302 );
buf ( n17304 , n17303 );
not ( n17305 , n17304 );
buf ( n17306 , n17305 );
buf ( n17307 , n17306 );
not ( n17308 , n17307 );
buf ( n17309 , n17308 );
not ( n17310 , n17309 );
buf ( n17311 , n17310 );
not ( n17312 , n17163 );
and ( n17313 , n17312 , n17259 );
xor ( n17314 , n17260 , n17270 );
and ( n17315 , n17314 , n17163 );
or ( n17316 , n17313 , n17315 );
buf ( n17317 , n17316 );
not ( n17318 , n17317 );
buf ( n17319 , n17318 );
buf ( n17320 , n17319 );
not ( n17321 , n17320 );
buf ( n17322 , n17321 );
not ( n17323 , n17322 );
buf ( n17324 , n17323 );
not ( n17325 , n17163 );
and ( n17326 , n17325 , n17261 );
xor ( n17327 , n17262 , n17269 );
and ( n17328 , n17327 , n17163 );
or ( n17329 , n17326 , n17328 );
buf ( n17330 , n17329 );
not ( n17331 , n17330 );
buf ( n17332 , n17331 );
buf ( n17333 , n17332 );
not ( n17334 , n17333 );
buf ( n17335 , n17334 );
not ( n17336 , n17335 );
buf ( n17337 , n17336 );
not ( n17338 , n17163 );
and ( n17339 , n17338 , n17263 );
xor ( n17340 , n17264 , n17268 );
and ( n17341 , n17340 , n17163 );
or ( n17342 , n17339 , n17341 );
buf ( n17343 , n17342 );
not ( n17344 , n17343 );
buf ( n17345 , n17344 );
buf ( n17346 , n17345 );
not ( n17347 , n17346 );
buf ( n17348 , n17347 );
not ( n17349 , n17348 );
buf ( n17350 , n17349 );
not ( n17351 , n17163 );
and ( n17352 , n17351 , n17265 );
xor ( n17353 , n17266 , n17267 );
and ( n17354 , n17353 , n17163 );
or ( n17355 , n17352 , n17354 );
buf ( n17356 , n17355 );
not ( n17357 , n17356 );
buf ( n17358 , n17357 );
buf ( n17359 , n17358 );
not ( n17360 , n17359 );
buf ( n17361 , n17360 );
not ( n17362 , n17361 );
buf ( n17363 , n17362 );
not ( n17364 , n17247 );
buf ( n17365 , n17364 );
and ( n17366 , n17363 , n17365 );
and ( n17367 , n17350 , n17366 );
and ( n17368 , n17337 , n17367 );
and ( n17369 , n17324 , n17368 );
and ( n17370 , n17311 , n17369 );
and ( n17371 , n17298 , n17370 );
and ( n17372 , n17285 , n17371 );
not ( n17373 , n17372 );
buf ( n17374 , n17373 );
buf ( n17375 , n17163 );
and ( n17376 , n17374 , n17375 );
or ( n17377 , C0 , n17376 );
buf ( n17378 , n17377 );
buf ( n17379 , n17378 );
not ( n17380 , n17379 );
not ( n17381 , n17375 );
buf ( n17382 , n17361 );
and ( n17383 , n17381 , n17382 );
xor ( n17384 , n17363 , n17365 );
buf ( n17385 , n17384 );
and ( n17386 , n17385 , n17375 );
or ( n17387 , n17383 , n17386 );
buf ( n17388 , n17387 );
buf ( n17389 , n17388 );
and ( n17390 , n17380 , n17389 );
not ( n17391 , n17389 );
not ( n17392 , n17248 );
xor ( n17393 , n17391 , n17392 );
and ( n17394 , n17393 , n17379 );
or ( n17395 , n17390 , n17394 );
buf ( n17396 , n17395 );
not ( n17397 , n17396 );
buf ( n17398 , n17397 );
buf ( n17399 , n17398 );
not ( n17400 , n17399 );
or ( n17401 , n17253 , n17400 );
not ( n17402 , n17379 );
not ( n17403 , n17375 );
buf ( n17404 , n17348 );
and ( n17405 , n17403 , n17404 );
xor ( n17406 , n17350 , n17366 );
buf ( n17407 , n17406 );
and ( n17408 , n17407 , n17375 );
or ( n17409 , n17405 , n17408 );
buf ( n17410 , n17409 );
buf ( n17411 , n17410 );
and ( n17412 , n17402 , n17411 );
not ( n17413 , n17411 );
and ( n17414 , n17391 , n17392 );
xor ( n17415 , n17413 , n17414 );
and ( n17416 , n17415 , n17379 );
or ( n17417 , n17412 , n17416 );
buf ( n17418 , n17417 );
not ( n17419 , n17418 );
buf ( n17420 , n17419 );
buf ( n17421 , n17420 );
not ( n17422 , n17421 );
or ( n17423 , n17401 , n17422 );
buf ( n17424 , n17423 );
buf ( n17425 , n17424 );
and ( n17426 , n17425 , n17379 );
not ( n17427 , n17426 );
and ( n17428 , n17427 , n17253 );
xor ( n17429 , n17253 , n17379 );
xor ( n17430 , n17429 , n17379 );
and ( n17431 , n17430 , n17426 );
or ( n17432 , n17428 , n17431 );
buf ( n17433 , n17432 );
not ( n17434 , n17426 );
and ( n17435 , n17434 , n17400 );
xor ( n17436 , n17400 , n17379 );
and ( n17437 , n17429 , n17379 );
xor ( n17438 , n17436 , n17437 );
and ( n17439 , n17438 , n17426 );
or ( n17440 , n17435 , n17439 );
buf ( n17441 , n17440 );
not ( n17442 , n17426 );
and ( n17443 , n17442 , n17422 );
xor ( n17444 , n17422 , n17379 );
and ( n17445 , n17436 , n17437 );
xor ( n17446 , n17444 , n17445 );
and ( n17447 , n17446 , n17426 );
or ( n17448 , n17443 , n17447 );
buf ( n17449 , n17448 );
and ( n17450 , n17433 , n17441 , n17449 );
or ( n17451 , n17162 , n17450 );
not ( n17452 , n17451 );
buf ( n17453 , RI210d6910_193);
buf ( n17454 , n16712 );
not ( n17455 , n17454 );
buf ( n17456 , n16753 );
and ( n17457 , n17455 , n17456 );
not ( n17458 , n17456 );
buf ( n17459 , n16761 );
not ( n17460 , n17459 );
buf ( n17461 , n16769 );
not ( n17462 , n17461 );
buf ( n17463 , n16777 );
not ( n17464 , n17463 );
buf ( n17465 , n16785 );
not ( n17466 , n17465 );
buf ( n17467 , n16793 );
not ( n17468 , n17467 );
buf ( n17469 , n16801 );
not ( n17470 , n17469 );
buf ( n17471 , n16809 );
not ( n17472 , n17471 );
buf ( n17473 , n16817 );
not ( n17474 , n17473 );
buf ( n17475 , n16825 );
not ( n17476 , n17475 );
buf ( n17477 , n16833 );
not ( n17478 , n17477 );
buf ( n17479 , n16841 );
not ( n17480 , n17479 );
buf ( n17481 , n16849 );
not ( n17482 , n17481 );
buf ( n17483 , n16857 );
not ( n17484 , n17483 );
buf ( n17485 , n16865 );
not ( n17486 , n17485 );
buf ( n17487 , n16873 );
not ( n17488 , n17487 );
buf ( n17489 , n16881 );
not ( n17490 , n17489 );
buf ( n17491 , n16889 );
not ( n17492 , n17491 );
buf ( n17493 , n16897 );
not ( n17494 , n17493 );
buf ( n17495 , n16900 );
not ( n17496 , n17495 );
and ( n17497 , n17494 , n17496 );
and ( n17498 , n17492 , n17497 );
and ( n17499 , n17490 , n17498 );
and ( n17500 , n17488 , n17499 );
and ( n17501 , n17486 , n17500 );
and ( n17502 , n17484 , n17501 );
and ( n17503 , n17482 , n17502 );
and ( n17504 , n17480 , n17503 );
and ( n17505 , n17478 , n17504 );
and ( n17506 , n17476 , n17505 );
and ( n17507 , n17474 , n17506 );
and ( n17508 , n17472 , n17507 );
and ( n17509 , n17470 , n17508 );
and ( n17510 , n17468 , n17509 );
and ( n17511 , n17466 , n17510 );
and ( n17512 , n17464 , n17511 );
and ( n17513 , n17462 , n17512 );
and ( n17514 , n17460 , n17513 );
xor ( n17515 , n17458 , n17514 );
and ( n17516 , n17515 , n17454 );
or ( n17517 , n17457 , n17516 );
buf ( n17518 , n17517 );
not ( n17519 , n17518 );
buf ( n17520 , n17519 );
buf ( n17521 , n17520 );
not ( n17522 , n17521 );
buf ( n17523 , n17522 );
buf ( n17524 , n17523 );
buf ( n17525 , n17524 );
not ( n17526 , n17525 );
buf ( n17527 , n17526 );
buf ( n17528 , n17527 );
not ( n17529 , n17528 );
not ( n17530 , n17454 );
buf ( n17531 , n16976 );
not ( n17532 , n17531 );
buf ( n17533 , n16984 );
not ( n17534 , n17533 );
buf ( n17535 , n16992 );
not ( n17536 , n17535 );
buf ( n17537 , n17000 );
not ( n17538 , n17537 );
buf ( n17539 , n17008 );
not ( n17540 , n17539 );
buf ( n17541 , n17016 );
not ( n17542 , n17541 );
buf ( n17543 , n17024 );
not ( n17544 , n17543 );
buf ( n17545 , n16720 );
not ( n17546 , n17545 );
buf ( n17547 , n16729 );
not ( n17548 , n17547 );
buf ( n17549 , n16737 );
not ( n17550 , n17549 );
buf ( n17551 , n16745 );
not ( n17552 , n17551 );
and ( n17553 , n17458 , n17514 );
and ( n17554 , n17552 , n17553 );
and ( n17555 , n17550 , n17554 );
and ( n17556 , n17548 , n17555 );
and ( n17557 , n17546 , n17556 );
and ( n17558 , n17544 , n17557 );
and ( n17559 , n17542 , n17558 );
and ( n17560 , n17540 , n17559 );
and ( n17561 , n17538 , n17560 );
and ( n17562 , n17536 , n17561 );
and ( n17563 , n17534 , n17562 );
and ( n17564 , n17532 , n17563 );
xor ( n17565 , n17530 , n17564 );
buf ( n17566 , n17454 );
and ( n17567 , n17565 , n17566 );
or ( n17568 , C0 , n17567 );
buf ( n17569 , n17568 );
not ( n17570 , n17569 );
buf ( n17571 , n17570 );
buf ( n17572 , n17571 );
not ( n17573 , n17572 );
buf ( n17574 , n17573 );
not ( n17575 , n17574 );
buf ( n17576 , n17575 );
not ( n17577 , n17454 );
and ( n17578 , n17577 , n17531 );
xor ( n17579 , n17532 , n17563 );
and ( n17580 , n17579 , n17454 );
or ( n17581 , n17578 , n17580 );
buf ( n17582 , n17581 );
not ( n17583 , n17582 );
buf ( n17584 , n17583 );
buf ( n17585 , n17584 );
not ( n17586 , n17585 );
buf ( n17587 , n17586 );
not ( n17588 , n17587 );
buf ( n17589 , n17588 );
not ( n17590 , n17454 );
and ( n17591 , n17590 , n17533 );
xor ( n17592 , n17534 , n17562 );
and ( n17593 , n17592 , n17454 );
or ( n17594 , n17591 , n17593 );
buf ( n17595 , n17594 );
not ( n17596 , n17595 );
buf ( n17597 , n17596 );
buf ( n17598 , n17597 );
not ( n17599 , n17598 );
buf ( n17600 , n17599 );
not ( n17601 , n17600 );
buf ( n17602 , n17601 );
not ( n17603 , n17454 );
and ( n17604 , n17603 , n17535 );
xor ( n17605 , n17536 , n17561 );
and ( n17606 , n17605 , n17454 );
or ( n17607 , n17604 , n17606 );
buf ( n17608 , n17607 );
not ( n17609 , n17608 );
buf ( n17610 , n17609 );
buf ( n17611 , n17610 );
not ( n17612 , n17611 );
buf ( n17613 , n17612 );
not ( n17614 , n17613 );
buf ( n17615 , n17614 );
not ( n17616 , n17454 );
and ( n17617 , n17616 , n17537 );
xor ( n17618 , n17538 , n17560 );
and ( n17619 , n17618 , n17454 );
or ( n17620 , n17617 , n17619 );
buf ( n17621 , n17620 );
not ( n17622 , n17621 );
buf ( n17623 , n17622 );
buf ( n17624 , n17623 );
not ( n17625 , n17624 );
buf ( n17626 , n17625 );
not ( n17627 , n17626 );
buf ( n17628 , n17627 );
not ( n17629 , n17454 );
and ( n17630 , n17629 , n17539 );
xor ( n17631 , n17540 , n17559 );
and ( n17632 , n17631 , n17454 );
or ( n17633 , n17630 , n17632 );
buf ( n17634 , n17633 );
not ( n17635 , n17634 );
buf ( n17636 , n17635 );
buf ( n17637 , n17636 );
not ( n17638 , n17637 );
buf ( n17639 , n17638 );
not ( n17640 , n17639 );
buf ( n17641 , n17640 );
not ( n17642 , n17454 );
and ( n17643 , n17642 , n17541 );
xor ( n17644 , n17542 , n17558 );
and ( n17645 , n17644 , n17454 );
or ( n17646 , n17643 , n17645 );
buf ( n17647 , n17646 );
not ( n17648 , n17647 );
buf ( n17649 , n17648 );
buf ( n17650 , n17649 );
not ( n17651 , n17650 );
buf ( n17652 , n17651 );
not ( n17653 , n17652 );
buf ( n17654 , n17653 );
not ( n17655 , n17454 );
and ( n17656 , n17655 , n17543 );
xor ( n17657 , n17544 , n17557 );
and ( n17658 , n17657 , n17454 );
or ( n17659 , n17656 , n17658 );
buf ( n17660 , n17659 );
not ( n17661 , n17660 );
buf ( n17662 , n17661 );
buf ( n17663 , n17662 );
not ( n17664 , n17663 );
buf ( n17665 , n17664 );
not ( n17666 , n17665 );
buf ( n17667 , n17666 );
not ( n17668 , n17454 );
and ( n17669 , n17668 , n17545 );
xor ( n17670 , n17546 , n17556 );
and ( n17671 , n17670 , n17454 );
or ( n17672 , n17669 , n17671 );
buf ( n17673 , n17672 );
not ( n17674 , n17673 );
buf ( n17675 , n17674 );
buf ( n17676 , n17675 );
not ( n17677 , n17676 );
buf ( n17678 , n17677 );
not ( n17679 , n17678 );
buf ( n17680 , n17679 );
not ( n17681 , n17454 );
and ( n17682 , n17681 , n17547 );
xor ( n17683 , n17548 , n17555 );
and ( n17684 , n17683 , n17454 );
or ( n17685 , n17682 , n17684 );
buf ( n17686 , n17685 );
not ( n17687 , n17686 );
buf ( n17688 , n17687 );
buf ( n17689 , n17688 );
not ( n17690 , n17689 );
buf ( n17691 , n17690 );
not ( n17692 , n17691 );
buf ( n17693 , n17692 );
not ( n17694 , n17454 );
and ( n17695 , n17694 , n17549 );
xor ( n17696 , n17550 , n17554 );
and ( n17697 , n17696 , n17454 );
or ( n17698 , n17695 , n17697 );
buf ( n17699 , n17698 );
not ( n17700 , n17699 );
buf ( n17701 , n17700 );
buf ( n17702 , n17701 );
not ( n17703 , n17702 );
buf ( n17704 , n17703 );
not ( n17705 , n17704 );
buf ( n17706 , n17705 );
not ( n17707 , n17454 );
and ( n17708 , n17707 , n17551 );
xor ( n17709 , n17552 , n17553 );
and ( n17710 , n17709 , n17454 );
or ( n17711 , n17708 , n17710 );
buf ( n17712 , n17711 );
not ( n17713 , n17712 );
buf ( n17714 , n17713 );
buf ( n17715 , n17714 );
not ( n17716 , n17715 );
buf ( n17717 , n17716 );
not ( n17718 , n17717 );
buf ( n17719 , n17718 );
not ( n17720 , n17523 );
buf ( n17721 , n17720 );
and ( n17722 , n17719 , n17721 );
and ( n17723 , n17706 , n17722 );
and ( n17724 , n17693 , n17723 );
and ( n17725 , n17680 , n17724 );
and ( n17726 , n17667 , n17725 );
and ( n17727 , n17654 , n17726 );
and ( n17728 , n17641 , n17727 );
and ( n17729 , n17628 , n17728 );
and ( n17730 , n17615 , n17729 );
and ( n17731 , n17602 , n17730 );
and ( n17732 , n17589 , n17731 );
and ( n17733 , n17576 , n17732 );
not ( n17734 , n17733 );
buf ( n17735 , n17734 );
buf ( n17736 , n17454 );
and ( n17737 , n17735 , n17736 );
or ( n17738 , C0 , n17737 );
buf ( n17739 , n17738 );
buf ( n17740 , n17739 );
not ( n17741 , n17740 );
not ( n17742 , n17736 );
buf ( n17743 , n17717 );
and ( n17744 , n17742 , n17743 );
xor ( n17745 , n17719 , n17721 );
buf ( n17746 , n17745 );
and ( n17747 , n17746 , n17736 );
or ( n17748 , n17744 , n17747 );
buf ( n17749 , n17748 );
buf ( n17750 , n17749 );
and ( n17751 , n17741 , n17750 );
not ( n17752 , n17750 );
not ( n17753 , n17524 );
xor ( n17754 , n17752 , n17753 );
and ( n17755 , n17754 , n17740 );
or ( n17756 , n17751 , n17755 );
buf ( n17757 , n17756 );
not ( n17758 , n17757 );
buf ( n17759 , n17758 );
buf ( n17760 , n17759 );
not ( n17761 , n17760 );
or ( n17762 , n17529 , n17761 );
not ( n17763 , n17740 );
not ( n17764 , n17736 );
buf ( n17765 , n17704 );
and ( n17766 , n17764 , n17765 );
xor ( n17767 , n17706 , n17722 );
buf ( n17768 , n17767 );
and ( n17769 , n17768 , n17736 );
or ( n17770 , n17766 , n17769 );
buf ( n17771 , n17770 );
buf ( n17772 , n17771 );
and ( n17773 , n17763 , n17772 );
not ( n17774 , n17772 );
and ( n17775 , n17752 , n17753 );
xor ( n17776 , n17774 , n17775 );
and ( n17777 , n17776 , n17740 );
or ( n17778 , n17773 , n17777 );
buf ( n17779 , n17778 );
not ( n17780 , n17779 );
buf ( n17781 , n17780 );
buf ( n17782 , n17781 );
not ( n17783 , n17782 );
or ( n17784 , n17762 , n17783 );
not ( n17785 , n17740 );
not ( n17786 , n17736 );
buf ( n17787 , n17691 );
and ( n17788 , n17786 , n17787 );
xor ( n17789 , n17693 , n17723 );
buf ( n17790 , n17789 );
and ( n17791 , n17790 , n17736 );
or ( n17792 , n17788 , n17791 );
buf ( n17793 , n17792 );
buf ( n17794 , n17793 );
and ( n17795 , n17785 , n17794 );
not ( n17796 , n17794 );
and ( n17797 , n17774 , n17775 );
xor ( n17798 , n17796 , n17797 );
and ( n17799 , n17798 , n17740 );
or ( n17800 , n17795 , n17799 );
buf ( n17801 , n17800 );
not ( n17802 , n17801 );
buf ( n17803 , n17802 );
buf ( n17804 , n17803 );
not ( n17805 , n17804 );
or ( n17806 , n17784 , n17805 );
or ( n17807 , n17806 , C0 );
or ( n17808 , n17807 , C0 );
or ( n17809 , n17808 , C0 );
or ( n17810 , n17809 , C0 );
or ( n17811 , n17810 , C0 );
or ( n17812 , n17811 , C0 );
or ( n17813 , n17812 , C0 );
or ( n17814 , n17813 , C0 );
or ( n17815 , n17814 , C0 );
or ( n17816 , n17815 , C0 );
or ( n17817 , n17816 , C0 );
or ( n17818 , n17817 , C0 );
or ( n17819 , n17818 , C0 );
or ( n17820 , n17819 , C0 );
or ( n17821 , n17820 , C0 );
or ( n17822 , n17821 , C0 );
or ( n17823 , n17822 , C0 );
or ( n17824 , n17823 , C0 );
or ( n17825 , n17824 , C0 );
or ( n17826 , n17825 , C0 );
or ( n17827 , n17826 , C0 );
or ( n17828 , n17827 , C0 );
or ( n17829 , n17828 , C0 );
or ( n17830 , n17829 , C0 );
or ( n17831 , n17830 , C0 );
or ( n17832 , n17831 , C0 );
or ( n17833 , n17832 , C0 );
buf ( n17834 , n17833 );
and ( n17835 , n17834 , n17740 );
not ( n17836 , n17835 );
and ( n17837 , n17836 , n17529 );
xor ( n17838 , n17529 , n17740 );
xor ( n17839 , n17838 , n17740 );
and ( n17840 , n17839 , n17835 );
or ( n17841 , n17837 , n17840 );
buf ( n17842 , n17841 );
not ( n17843 , n17835 );
and ( n17844 , n17843 , n17761 );
xor ( n17845 , n17761 , n17740 );
and ( n17846 , n17838 , n17740 );
xor ( n17847 , n17845 , n17846 );
and ( n17848 , n17847 , n17835 );
or ( n17849 , n17844 , n17848 );
buf ( n17850 , n17849 );
not ( n17851 , n17850 );
not ( n17852 , n17835 );
and ( n17853 , n17852 , n17783 );
xor ( n17854 , n17783 , n17740 );
and ( n17855 , n17845 , n17846 );
xor ( n17856 , n17854 , n17855 );
and ( n17857 , n17856 , n17835 );
or ( n17858 , n17853 , n17857 );
buf ( n17859 , n17858 );
not ( n17860 , n17835 );
and ( n17861 , n17860 , n17805 );
xor ( n17862 , n17805 , n17740 );
and ( n17863 , n17854 , n17855 );
xor ( n17864 , n17862 , n17863 );
and ( n17865 , n17864 , n17835 );
or ( n17866 , n17861 , n17865 );
buf ( n17867 , n17866 );
and ( n17868 , n17842 , n17851 , n17859 , n17867 );
not ( n17869 , n17842 );
and ( n17870 , n17869 , n17850 , n17859 , n17867 );
or ( n17871 , n17868 , n17870 );
and ( n17872 , n17842 , n17850 , n17859 , n17867 );
or ( n17873 , n17871 , n17872 );
and ( n17874 , n17453 , n17873 );
buf ( n17875 , RI210cdfb8_248);
buf ( n17876 , n17875 );
buf ( n17877 , n17876 );
not ( n17878 , n17877 );
buf ( n17879 , n17878 );
buf ( n17880 , n17879 );
not ( n17881 , n17880 );
buf ( n17882 , GI2046a680_186);
buf ( n17883 , n17882 );
not ( n17884 , n17883 );
buf ( n17885 , RI210d2d88_218);
buf ( n17886 , n17885 );
and ( n17887 , n17884 , n17886 );
not ( n17888 , n17886 );
not ( n17889 , n17876 );
xor ( n17890 , n17888 , n17889 );
and ( n17891 , n17890 , n17883 );
or ( n17892 , n17887 , n17891 );
buf ( n17893 , n17892 );
not ( n17894 , n17893 );
buf ( n17895 , n17894 );
buf ( n17896 , n17895 );
not ( n17897 , n17896 );
or ( n17898 , n17881 , n17897 );
not ( n17899 , n17883 );
buf ( n17900 , RI210d10f0_228);
buf ( n17901 , n17900 );
and ( n17902 , n17899 , n17901 );
not ( n17903 , n17901 );
and ( n17904 , n17888 , n17889 );
xor ( n17905 , n17903 , n17904 );
and ( n17906 , n17905 , n17883 );
or ( n17907 , n17902 , n17906 );
buf ( n17908 , n17907 );
not ( n17909 , n17908 );
buf ( n17910 , n17909 );
buf ( n17911 , n17910 );
not ( n17912 , n17911 );
or ( n17913 , n17898 , n17912 );
not ( n17914 , n17883 );
buf ( n17915 , RI210d1078_229);
buf ( n17916 , n17915 );
and ( n17917 , n17914 , n17916 );
not ( n17918 , n17916 );
and ( n17919 , n17903 , n17904 );
xor ( n17920 , n17918 , n17919 );
and ( n17921 , n17920 , n17883 );
or ( n17922 , n17917 , n17921 );
buf ( n17923 , n17922 );
not ( n17924 , n17923 );
buf ( n17925 , n17924 );
buf ( n17926 , n17925 );
not ( n17927 , n17926 );
or ( n17928 , n17913 , n17927 );
not ( n17929 , n17883 );
buf ( n17930 , RI210d1000_230);
buf ( n17931 , n17930 );
and ( n17932 , n17929 , n17931 );
not ( n17933 , n17931 );
and ( n17934 , n17918 , n17919 );
xor ( n17935 , n17933 , n17934 );
and ( n17936 , n17935 , n17883 );
or ( n17937 , n17932 , n17936 );
buf ( n17938 , n17937 );
not ( n17939 , n17938 );
buf ( n17940 , n17939 );
buf ( n17941 , n17940 );
not ( n17942 , n17941 );
or ( n17943 , n17928 , n17942 );
not ( n17944 , n17883 );
buf ( n17945 , RI210d0790_231);
buf ( n17946 , n17945 );
and ( n17947 , n17944 , n17946 );
not ( n17948 , n17946 );
and ( n17949 , n17933 , n17934 );
xor ( n17950 , n17948 , n17949 );
and ( n17951 , n17950 , n17883 );
or ( n17952 , n17947 , n17951 );
buf ( n17953 , n17952 );
not ( n17954 , n17953 );
buf ( n17955 , n17954 );
buf ( n17956 , n17955 );
not ( n17957 , n17956 );
or ( n17958 , n17943 , n17957 );
not ( n17959 , n17883 );
buf ( n17960 , RI210d0718_232);
buf ( n17961 , n17960 );
and ( n17962 , n17959 , n17961 );
not ( n17963 , n17961 );
and ( n17964 , n17948 , n17949 );
xor ( n17965 , n17963 , n17964 );
and ( n17966 , n17965 , n17883 );
or ( n17967 , n17962 , n17966 );
buf ( n17968 , n17967 );
not ( n17969 , n17968 );
buf ( n17970 , n17969 );
buf ( n17971 , n17970 );
not ( n17972 , n17971 );
or ( n17973 , n17958 , n17972 );
not ( n17974 , n17883 );
buf ( n17975 , RI210d06a0_233);
buf ( n17976 , n17975 );
and ( n17977 , n17974 , n17976 );
not ( n17978 , n17976 );
and ( n17979 , n17963 , n17964 );
xor ( n17980 , n17978 , n17979 );
and ( n17981 , n17980 , n17883 );
or ( n17982 , n17977 , n17981 );
buf ( n17983 , n17982 );
not ( n17984 , n17983 );
buf ( n17985 , n17984 );
buf ( n17986 , n17985 );
not ( n17987 , n17986 );
or ( n17988 , n17973 , n17987 );
not ( n17989 , n17883 );
buf ( n17990 , RI210d0628_234);
buf ( n17991 , n17990 );
and ( n17992 , n17989 , n17991 );
not ( n17993 , n17991 );
and ( n17994 , n17978 , n17979 );
xor ( n17995 , n17993 , n17994 );
and ( n17996 , n17995 , n17883 );
or ( n17997 , n17992 , n17996 );
buf ( n17998 , n17997 );
not ( n17999 , n17998 );
buf ( n18000 , n17999 );
buf ( n18001 , n18000 );
not ( n18002 , n18001 );
or ( n18003 , n17988 , n18002 );
not ( n18004 , n17883 );
buf ( n18005 , RI210cfdb8_235);
buf ( n18006 , n18005 );
and ( n18007 , n18004 , n18006 );
not ( n18008 , n18006 );
and ( n18009 , n17993 , n17994 );
xor ( n18010 , n18008 , n18009 );
and ( n18011 , n18010 , n17883 );
or ( n18012 , n18007 , n18011 );
buf ( n18013 , n18012 );
not ( n18014 , n18013 );
buf ( n18015 , n18014 );
buf ( n18016 , n18015 );
not ( n18017 , n18016 );
or ( n18018 , n18003 , n18017 );
not ( n18019 , n17883 );
buf ( n18020 , RI210d4228_208);
buf ( n18021 , n18020 );
and ( n18022 , n18019 , n18021 );
not ( n18023 , n18021 );
and ( n18024 , n18008 , n18009 );
xor ( n18025 , n18023 , n18024 );
and ( n18026 , n18025 , n17883 );
or ( n18027 , n18022 , n18026 );
buf ( n18028 , n18027 );
not ( n18029 , n18028 );
buf ( n18030 , n18029 );
buf ( n18031 , n18030 );
not ( n18032 , n18031 );
or ( n18033 , n18018 , n18032 );
not ( n18034 , n17883 );
buf ( n18035 , RI210d41b0_209);
buf ( n18036 , n18035 );
and ( n18037 , n18034 , n18036 );
not ( n18038 , n18036 );
and ( n18039 , n18023 , n18024 );
xor ( n18040 , n18038 , n18039 );
and ( n18041 , n18040 , n17883 );
or ( n18042 , n18037 , n18041 );
buf ( n18043 , n18042 );
not ( n18044 , n18043 );
buf ( n18045 , n18044 );
buf ( n18046 , n18045 );
not ( n18047 , n18046 );
or ( n18048 , n18033 , n18047 );
not ( n18049 , n17883 );
buf ( n18050 , RI210d4138_210);
buf ( n18051 , n18050 );
and ( n18052 , n18049 , n18051 );
not ( n18053 , n18051 );
and ( n18054 , n18038 , n18039 );
xor ( n18055 , n18053 , n18054 );
and ( n18056 , n18055 , n17883 );
or ( n18057 , n18052 , n18056 );
buf ( n18058 , n18057 );
not ( n18059 , n18058 );
buf ( n18060 , n18059 );
buf ( n18061 , n18060 );
not ( n18062 , n18061 );
or ( n18063 , n18048 , n18062 );
not ( n18064 , n17883 );
buf ( n18065 , RI210d38c8_211);
buf ( n18066 , n18065 );
and ( n18067 , n18064 , n18066 );
not ( n18068 , n18066 );
and ( n18069 , n18053 , n18054 );
xor ( n18070 , n18068 , n18069 );
and ( n18071 , n18070 , n17883 );
or ( n18072 , n18067 , n18071 );
buf ( n18073 , n18072 );
not ( n18074 , n18073 );
buf ( n18075 , n18074 );
buf ( n18076 , n18075 );
not ( n18077 , n18076 );
or ( n18078 , n18063 , n18077 );
not ( n18079 , n17883 );
buf ( n18080 , RI210d3850_212);
buf ( n18081 , n18080 );
and ( n18082 , n18079 , n18081 );
not ( n18083 , n18081 );
and ( n18084 , n18068 , n18069 );
xor ( n18085 , n18083 , n18084 );
and ( n18086 , n18085 , n17883 );
or ( n18087 , n18082 , n18086 );
buf ( n18088 , n18087 );
not ( n18089 , n18088 );
buf ( n18090 , n18089 );
buf ( n18091 , n18090 );
not ( n18092 , n18091 );
or ( n18093 , n18078 , n18092 );
not ( n18094 , n17883 );
buf ( n18095 , RI210d37d8_213);
buf ( n18096 , n18095 );
and ( n18097 , n18094 , n18096 );
not ( n18098 , n18096 );
and ( n18099 , n18083 , n18084 );
xor ( n18100 , n18098 , n18099 );
and ( n18101 , n18100 , n17883 );
or ( n18102 , n18097 , n18101 );
buf ( n18103 , n18102 );
not ( n18104 , n18103 );
buf ( n18105 , n18104 );
buf ( n18106 , n18105 );
not ( n18107 , n18106 );
or ( n18108 , n18093 , n18107 );
not ( n18109 , n17883 );
buf ( n18110 , RI210d3760_214);
buf ( n18111 , n18110 );
and ( n18112 , n18109 , n18111 );
not ( n18113 , n18111 );
and ( n18114 , n18098 , n18099 );
xor ( n18115 , n18113 , n18114 );
and ( n18116 , n18115 , n17883 );
or ( n18117 , n18112 , n18116 );
buf ( n18118 , n18117 );
not ( n18119 , n18118 );
buf ( n18120 , n18119 );
buf ( n18121 , n18120 );
not ( n18122 , n18121 );
or ( n18123 , n18108 , n18122 );
not ( n18124 , n17883 );
buf ( n18125 , RI210d2ef0_215);
buf ( n18126 , n18125 );
and ( n18127 , n18124 , n18126 );
not ( n18128 , n18126 );
and ( n18129 , n18113 , n18114 );
xor ( n18130 , n18128 , n18129 );
and ( n18131 , n18130 , n17883 );
or ( n18132 , n18127 , n18131 );
buf ( n18133 , n18132 );
not ( n18134 , n18133 );
buf ( n18135 , n18134 );
buf ( n18136 , n18135 );
not ( n18137 , n18136 );
or ( n18138 , n18123 , n18137 );
not ( n18139 , n17883 );
buf ( n18140 , RI210d2e78_216);
buf ( n18141 , n18140 );
and ( n18142 , n18139 , n18141 );
not ( n18143 , n18141 );
and ( n18144 , n18128 , n18129 );
xor ( n18145 , n18143 , n18144 );
and ( n18146 , n18145 , n17883 );
or ( n18147 , n18142 , n18146 );
buf ( n18148 , n18147 );
not ( n18149 , n18148 );
buf ( n18150 , n18149 );
buf ( n18151 , n18150 );
not ( n18152 , n18151 );
or ( n18153 , n18138 , n18152 );
not ( n18154 , n17883 );
buf ( n18155 , RI210d2e00_217);
buf ( n18156 , n18155 );
and ( n18157 , n18154 , n18156 );
not ( n18158 , n18156 );
and ( n18159 , n18143 , n18144 );
xor ( n18160 , n18158 , n18159 );
and ( n18161 , n18160 , n17883 );
or ( n18162 , n18157 , n18161 );
buf ( n18163 , n18162 );
not ( n18164 , n18163 );
buf ( n18165 , n18164 );
buf ( n18166 , n18165 );
not ( n18167 , n18166 );
or ( n18168 , n18153 , n18167 );
not ( n18169 , n17883 );
buf ( n18170 , RI210d2518_219);
buf ( n18171 , n18170 );
and ( n18172 , n18169 , n18171 );
not ( n18173 , n18171 );
and ( n18174 , n18158 , n18159 );
xor ( n18175 , n18173 , n18174 );
and ( n18176 , n18175 , n17883 );
or ( n18177 , n18172 , n18176 );
buf ( n18178 , n18177 );
not ( n18179 , n18178 );
buf ( n18180 , n18179 );
buf ( n18181 , n18180 );
not ( n18182 , n18181 );
or ( n18183 , n18168 , n18182 );
not ( n18184 , n17883 );
buf ( n18185 , RI210d24a0_220);
buf ( n18186 , n18185 );
and ( n18187 , n18184 , n18186 );
not ( n18188 , n18186 );
and ( n18189 , n18173 , n18174 );
xor ( n18190 , n18188 , n18189 );
and ( n18191 , n18190 , n17883 );
or ( n18192 , n18187 , n18191 );
buf ( n18193 , n18192 );
not ( n18194 , n18193 );
buf ( n18195 , n18194 );
buf ( n18196 , n18195 );
not ( n18197 , n18196 );
or ( n18198 , n18183 , n18197 );
not ( n18199 , n17883 );
buf ( n18200 , RI210d2428_221);
buf ( n18201 , n18200 );
and ( n18202 , n18199 , n18201 );
not ( n18203 , n18201 );
and ( n18204 , n18188 , n18189 );
xor ( n18205 , n18203 , n18204 );
and ( n18206 , n18205 , n17883 );
or ( n18207 , n18202 , n18206 );
buf ( n18208 , n18207 );
not ( n18209 , n18208 );
buf ( n18210 , n18209 );
buf ( n18211 , n18210 );
not ( n18212 , n18211 );
or ( n18213 , n18198 , n18212 );
not ( n18214 , n17883 );
buf ( n18215 , RI210d23b0_222);
buf ( n18216 , n18215 );
and ( n18217 , n18214 , n18216 );
not ( n18218 , n18216 );
and ( n18219 , n18203 , n18204 );
xor ( n18220 , n18218 , n18219 );
and ( n18221 , n18220 , n17883 );
or ( n18222 , n18217 , n18221 );
buf ( n18223 , n18222 );
not ( n18224 , n18223 );
buf ( n18225 , n18224 );
buf ( n18226 , n18225 );
not ( n18227 , n18226 );
or ( n18228 , n18213 , n18227 );
not ( n18229 , n17883 );
buf ( n18230 , RI210d1b40_223);
buf ( n18231 , n18230 );
and ( n18232 , n18229 , n18231 );
not ( n18233 , n18231 );
and ( n18234 , n18218 , n18219 );
xor ( n18235 , n18233 , n18234 );
and ( n18236 , n18235 , n17883 );
or ( n18237 , n18232 , n18236 );
buf ( n18238 , n18237 );
not ( n18239 , n18238 );
buf ( n18240 , n18239 );
buf ( n18241 , n18240 );
not ( n18242 , n18241 );
or ( n18243 , n18228 , n18242 );
not ( n18244 , n17883 );
buf ( n18245 , RI210d1ac8_224);
buf ( n18246 , n18245 );
and ( n18247 , n18244 , n18246 );
not ( n18248 , n18246 );
and ( n18249 , n18233 , n18234 );
xor ( n18250 , n18248 , n18249 );
and ( n18251 , n18250 , n17883 );
or ( n18252 , n18247 , n18251 );
buf ( n18253 , n18252 );
not ( n18254 , n18253 );
buf ( n18255 , n18254 );
buf ( n18256 , n18255 );
not ( n18257 , n18256 );
or ( n18258 , n18243 , n18257 );
not ( n18259 , n17883 );
buf ( n18260 , RI210d1a50_225);
buf ( n18261 , n18260 );
and ( n18262 , n18259 , n18261 );
not ( n18263 , n18261 );
and ( n18264 , n18248 , n18249 );
xor ( n18265 , n18263 , n18264 );
and ( n18266 , n18265 , n17883 );
or ( n18267 , n18262 , n18266 );
buf ( n18268 , n18267 );
not ( n18269 , n18268 );
buf ( n18270 , n18269 );
buf ( n18271 , n18270 );
not ( n18272 , n18271 );
or ( n18273 , n18258 , n18272 );
not ( n18274 , n17883 );
buf ( n18275 , RI210d19d8_226);
buf ( n18276 , n18275 );
and ( n18277 , n18274 , n18276 );
not ( n18278 , n18276 );
and ( n18279 , n18263 , n18264 );
xor ( n18280 , n18278 , n18279 );
and ( n18281 , n18280 , n17883 );
or ( n18282 , n18277 , n18281 );
buf ( n18283 , n18282 );
not ( n18284 , n18283 );
buf ( n18285 , n18284 );
buf ( n18286 , n18285 );
not ( n18287 , n18286 );
or ( n18288 , n18273 , n18287 );
not ( n18289 , n17883 );
buf ( n18290 , RI210d1168_227);
buf ( n18291 , n18290 );
and ( n18292 , n18289 , n18291 );
not ( n18293 , n18291 );
and ( n18294 , n18278 , n18279 );
xor ( n18295 , n18293 , n18294 );
and ( n18296 , n18295 , n17883 );
or ( n18297 , n18292 , n18296 );
buf ( n18298 , n18297 );
not ( n18299 , n18298 );
buf ( n18300 , n18299 );
buf ( n18301 , n18300 );
not ( n18302 , n18301 );
or ( n18303 , n18288 , n18302 );
buf ( n18304 , n18303 );
buf ( n18305 , n18304 );
and ( n18306 , n18305 , n17883 );
not ( n18307 , n18306 );
and ( n18308 , n18307 , n17881 );
xor ( n18309 , n17881 , n17883 );
xor ( n18310 , n18309 , n17883 );
and ( n18311 , n18310 , n18306 );
or ( n18312 , n18308 , n18311 );
buf ( n18313 , n18312 );
buf ( n18314 , n18313 );
buf ( n18315 , n16712 );
not ( n18316 , n18315 );
buf ( n18317 , n16984 );
and ( n18318 , n18316 , n18317 );
not ( n18319 , n18317 );
buf ( n18320 , n16992 );
not ( n18321 , n18320 );
buf ( n18322 , n17000 );
not ( n18323 , n18322 );
buf ( n18324 , n17008 );
not ( n18325 , n18324 );
buf ( n18326 , n17016 );
not ( n18327 , n18326 );
buf ( n18328 , n17024 );
not ( n18329 , n18328 );
buf ( n18330 , n16720 );
not ( n18331 , n18330 );
buf ( n18332 , n16729 );
not ( n18333 , n18332 );
buf ( n18334 , n16737 );
not ( n18335 , n18334 );
buf ( n18336 , n16745 );
not ( n18337 , n18336 );
buf ( n18338 , n16753 );
not ( n18339 , n18338 );
buf ( n18340 , n16761 );
not ( n18341 , n18340 );
buf ( n18342 , n16769 );
not ( n18343 , n18342 );
buf ( n18344 , n16777 );
not ( n18345 , n18344 );
buf ( n18346 , n16785 );
not ( n18347 , n18346 );
buf ( n18348 , n16793 );
not ( n18349 , n18348 );
buf ( n18350 , n16801 );
not ( n18351 , n18350 );
buf ( n18352 , n16809 );
not ( n18353 , n18352 );
buf ( n18354 , n16817 );
not ( n18355 , n18354 );
buf ( n18356 , n16825 );
not ( n18357 , n18356 );
buf ( n18358 , n16833 );
not ( n18359 , n18358 );
buf ( n18360 , n16841 );
not ( n18361 , n18360 );
buf ( n18362 , n16849 );
not ( n18363 , n18362 );
buf ( n18364 , n16857 );
not ( n18365 , n18364 );
buf ( n18366 , n16865 );
not ( n18367 , n18366 );
buf ( n18368 , n16873 );
not ( n18369 , n18368 );
buf ( n18370 , n16881 );
not ( n18371 , n18370 );
buf ( n18372 , n16889 );
not ( n18373 , n18372 );
buf ( n18374 , n16897 );
not ( n18375 , n18374 );
buf ( n18376 , n16900 );
not ( n18377 , n18376 );
and ( n18378 , n18375 , n18377 );
and ( n18379 , n18373 , n18378 );
and ( n18380 , n18371 , n18379 );
and ( n18381 , n18369 , n18380 );
and ( n18382 , n18367 , n18381 );
and ( n18383 , n18365 , n18382 );
and ( n18384 , n18363 , n18383 );
and ( n18385 , n18361 , n18384 );
and ( n18386 , n18359 , n18385 );
and ( n18387 , n18357 , n18386 );
and ( n18388 , n18355 , n18387 );
and ( n18389 , n18353 , n18388 );
and ( n18390 , n18351 , n18389 );
and ( n18391 , n18349 , n18390 );
and ( n18392 , n18347 , n18391 );
and ( n18393 , n18345 , n18392 );
and ( n18394 , n18343 , n18393 );
and ( n18395 , n18341 , n18394 );
and ( n18396 , n18339 , n18395 );
and ( n18397 , n18337 , n18396 );
and ( n18398 , n18335 , n18397 );
and ( n18399 , n18333 , n18398 );
and ( n18400 , n18331 , n18399 );
and ( n18401 , n18329 , n18400 );
and ( n18402 , n18327 , n18401 );
and ( n18403 , n18325 , n18402 );
and ( n18404 , n18323 , n18403 );
and ( n18405 , n18321 , n18404 );
xor ( n18406 , n18319 , n18405 );
and ( n18407 , n18406 , n18315 );
or ( n18408 , n18318 , n18407 );
buf ( n18409 , n18408 );
not ( n18410 , n18409 );
buf ( n18411 , n18410 );
buf ( n18412 , n18411 );
not ( n18413 , n18412 );
buf ( n18414 , n18413 );
buf ( n18415 , n18414 );
buf ( n18416 , n18415 );
not ( n18417 , n18416 );
buf ( n18418 , n18417 );
buf ( n18419 , n18418 );
not ( n18420 , n18419 );
not ( n18421 , n18315 );
buf ( n18422 , n16976 );
not ( n18423 , n18422 );
and ( n18424 , n18319 , n18405 );
and ( n18425 , n18423 , n18424 );
xor ( n18426 , n18421 , n18425 );
buf ( n18427 , n18315 );
and ( n18428 , n18426 , n18427 );
or ( n18429 , C0 , n18428 );
buf ( n18430 , n18429 );
not ( n18431 , n18430 );
buf ( n18432 , n18431 );
buf ( n18433 , n18432 );
not ( n18434 , n18433 );
buf ( n18435 , n18434 );
not ( n18436 , n18435 );
buf ( n18437 , n18436 );
not ( n18438 , n18315 );
and ( n18439 , n18438 , n18422 );
xor ( n18440 , n18423 , n18424 );
and ( n18441 , n18440 , n18315 );
or ( n18442 , n18439 , n18441 );
buf ( n18443 , n18442 );
not ( n18444 , n18443 );
buf ( n18445 , n18444 );
buf ( n18446 , n18445 );
not ( n18447 , n18446 );
buf ( n18448 , n18447 );
not ( n18449 , n18448 );
buf ( n18450 , n18449 );
not ( n18451 , n18414 );
buf ( n18452 , n18451 );
and ( n18453 , n18450 , n18452 );
and ( n18454 , n18437 , n18453 );
not ( n18455 , n18454 );
buf ( n18456 , n18455 );
buf ( n18457 , n18315 );
and ( n18458 , n18456 , n18457 );
or ( n18459 , C0 , n18458 );
buf ( n18460 , n18459 );
buf ( n18461 , n18460 );
not ( n18462 , n18461 );
not ( n18463 , n18457 );
buf ( n18464 , n18448 );
and ( n18465 , n18463 , n18464 );
xor ( n18466 , n18450 , n18452 );
buf ( n18467 , n18466 );
and ( n18468 , n18467 , n18457 );
or ( n18469 , n18465 , n18468 );
buf ( n18470 , n18469 );
buf ( n18471 , n18470 );
and ( n18472 , n18462 , n18471 );
not ( n18473 , n18471 );
not ( n18474 , n18415 );
xor ( n18475 , n18473 , n18474 );
and ( n18476 , n18475 , n18461 );
or ( n18477 , n18472 , n18476 );
buf ( n18478 , n18477 );
not ( n18479 , n18478 );
buf ( n18480 , n18479 );
buf ( n18481 , n18480 );
not ( n18482 , n18481 );
or ( n18483 , n18420 , n18482 );
buf ( n18484 , n18483 );
buf ( n18485 , n18484 );
and ( n18486 , n18485 , n18461 );
not ( n18487 , n18486 );
and ( n18488 , n18487 , n18420 );
xor ( n18489 , n18420 , n18461 );
xor ( n18490 , n18489 , n18461 );
and ( n18491 , n18490 , n18486 );
or ( n18492 , n18488 , n18491 );
buf ( n18493 , n18492 );
not ( n18494 , n18486 );
and ( n18495 , n18494 , n18482 );
xor ( n18496 , n18482 , n18461 );
and ( n18497 , n18489 , n18461 );
xor ( n18498 , n18496 , n18497 );
and ( n18499 , n18498 , n18486 );
or ( n18500 , n18495 , n18499 );
buf ( n18501 , n18500 );
and ( n18502 , n18493 , n18501 );
and ( n18503 , n18314 , n18502 );
buf ( n18504 , RI210d8ff8_178);
not ( n18505 , n18493 );
and ( n18506 , n18505 , n18501 );
and ( n18507 , n18504 , n18506 );
buf ( n18508 , RI21a0b7a0_150);
nor ( n18509 , n18505 , n18501 );
and ( n18510 , n18508 , n18509 );
buf ( n18511 , RI21a0e590_122);
nor ( n18512 , n18493 , n18501 );
and ( n18513 , n18511 , n18512 );
or ( n18514 , n18503 , n18507 , n18510 , n18513 );
buf ( n18515 , n18514 );
buf ( n18516 , n18515 );
not ( n18517 , n18516 );
buf ( n18518 , n18517 );
buf ( n18519 , n18518 );
not ( n18520 , n18519 );
buf ( n18521 , RI210d55d8_200);
and ( n18522 , n18521 , n18506 );
buf ( n18523 , RI210da3a8_170);
and ( n18524 , n18523 , n18509 );
buf ( n18525 , RI21a0c178_143);
and ( n18526 , n18525 , n18512 );
or ( n18527 , C0 , n18522 , n18524 , n18526 );
buf ( n18528 , n18527 );
not ( n18529 , n18528 );
not ( n18530 , n18306 );
and ( n18531 , n18530 , n17897 );
xor ( n18532 , n17897 , n17883 );
and ( n18533 , n18309 , n17883 );
xor ( n18534 , n18532 , n18533 );
and ( n18535 , n18534 , n18306 );
or ( n18536 , n18531 , n18535 );
buf ( n18537 , n18536 );
buf ( n18538 , n18537 );
and ( n18539 , n18538 , n18502 );
buf ( n18540 , RI210d73d8_187);
and ( n18541 , n18540 , n18506 );
buf ( n18542 , RI21a0a6c0_158);
and ( n18543 , n18542 , n18509 );
buf ( n18544 , RI21a0d438_131);
and ( n18545 , n18544 , n18512 );
or ( n18546 , n18539 , n18541 , n18543 , n18545 );
buf ( n18547 , n18546 );
and ( n18548 , n18529 , n18547 );
not ( n18549 , n18547 );
not ( n18550 , n18515 );
xor ( n18551 , n18549 , n18550 );
and ( n18552 , n18551 , n18528 );
or ( n18553 , n18548 , n18552 );
buf ( n18554 , n18553 );
not ( n18555 , n18554 );
buf ( n18556 , n18555 );
buf ( n18557 , n18556 );
not ( n18558 , n18557 );
or ( n18559 , n18520 , n18558 );
not ( n18560 , n18528 );
not ( n18561 , n18306 );
and ( n18562 , n18561 , n17912 );
xor ( n18563 , n17912 , n17883 );
and ( n18564 , n18532 , n18533 );
xor ( n18565 , n18563 , n18564 );
and ( n18566 , n18565 , n18306 );
or ( n18567 , n18562 , n18566 );
buf ( n18568 , n18567 );
buf ( n18569 , n18568 );
and ( n18570 , n18569 , n18502 );
buf ( n18571 , RI210d5ec0_198);
and ( n18572 , n18571 , n18506 );
buf ( n18573 , RI210da498_168);
and ( n18574 , n18573 , n18509 );
buf ( n18575 , RI21a0c268_141);
and ( n18576 , n18575 , n18512 );
or ( n18577 , n18570 , n18572 , n18574 , n18576 );
buf ( n18578 , n18577 );
and ( n18579 , n18560 , n18578 );
not ( n18580 , n18578 );
and ( n18581 , n18549 , n18550 );
xor ( n18582 , n18580 , n18581 );
and ( n18583 , n18582 , n18528 );
or ( n18584 , n18579 , n18583 );
buf ( n18585 , n18584 );
not ( n18586 , n18585 );
buf ( n18587 , n18586 );
buf ( n18588 , n18587 );
not ( n18589 , n18588 );
or ( n18590 , n18559 , n18589 );
not ( n18591 , n18528 );
not ( n18592 , n18306 );
and ( n18593 , n18592 , n17927 );
xor ( n18594 , n17927 , n17883 );
and ( n18595 , n18563 , n18564 );
xor ( n18596 , n18594 , n18595 );
and ( n18597 , n18596 , n18306 );
or ( n18598 , n18593 , n18597 );
buf ( n18599 , n18598 );
buf ( n18600 , n18599 );
not ( n18601 , n18600 );
buf ( n18602 , n18601 );
and ( n18603 , n18602 , n18502 );
buf ( n18604 , RI210d5560_201);
and ( n18605 , n18604 , n18506 );
buf ( n18606 , RI210d9b38_171);
and ( n18607 , n18606 , n18509 );
buf ( n18608 , RI21a0c100_144);
and ( n18609 , n18608 , n18512 );
or ( n18610 , n18603 , n18605 , n18607 , n18609 );
buf ( n18611 , n18610 );
and ( n18612 , n18591 , n18611 );
not ( n18613 , n18611 );
and ( n18614 , n18580 , n18581 );
xor ( n18615 , n18613 , n18614 );
and ( n18616 , n18615 , n18528 );
or ( n18617 , n18612 , n18616 );
buf ( n18618 , n18617 );
not ( n18619 , n18618 );
buf ( n18620 , n18619 );
buf ( n18621 , n18620 );
not ( n18622 , n18621 );
or ( n18623 , n18590 , n18622 );
not ( n18624 , n18528 );
not ( n18625 , n18306 );
and ( n18626 , n18625 , n17942 );
xor ( n18627 , n17942 , n17883 );
and ( n18628 , n18594 , n18595 );
xor ( n18629 , n18627 , n18628 );
and ( n18630 , n18629 , n18306 );
or ( n18631 , n18626 , n18630 );
buf ( n18632 , n18631 );
buf ( n18633 , n18632 );
xor ( n18634 , n18633 , n18600 );
buf ( n18635 , n18634 );
and ( n18636 , n18635 , n18502 );
buf ( n18637 , RI210d54e8_202);
and ( n18638 , n18637 , n18506 );
buf ( n18639 , RI210d9ac0_172);
and ( n18640 , n18639 , n18509 );
buf ( n18641 , RI210cf2f0_241);
and ( n18642 , n18641 , n18512 );
or ( n18643 , n18636 , n18638 , n18640 , n18642 );
buf ( n18644 , n18643 );
and ( n18645 , n18624 , n18644 );
not ( n18646 , n18644 );
and ( n18647 , n18613 , n18614 );
xor ( n18648 , n18646 , n18647 );
and ( n18649 , n18648 , n18528 );
or ( n18650 , n18645 , n18649 );
buf ( n18651 , n18650 );
not ( n18652 , n18651 );
buf ( n18653 , n18652 );
buf ( n18654 , n18653 );
not ( n18655 , n18654 );
or ( n18656 , n18623 , n18655 );
not ( n18657 , n18528 );
not ( n18658 , n18306 );
and ( n18659 , n18658 , n17957 );
xor ( n18660 , n17957 , n17883 );
and ( n18661 , n18627 , n18628 );
xor ( n18662 , n18660 , n18661 );
and ( n18663 , n18662 , n18306 );
or ( n18664 , n18659 , n18663 );
buf ( n18665 , n18664 );
buf ( n18666 , n18665 );
and ( n18667 , n18633 , n18600 );
xor ( n18668 , n18666 , n18667 );
buf ( n18669 , n18668 );
and ( n18670 , n18669 , n18502 );
buf ( n18671 , RI210d4c78_203);
and ( n18672 , n18671 , n18506 );
buf ( n18673 , RI210d9a48_173);
and ( n18674 , n18673 , n18509 );
buf ( n18675 , RI21a0c088_145);
and ( n18676 , n18675 , n18512 );
or ( n18677 , n18670 , n18672 , n18674 , n18676 );
buf ( n18678 , n18677 );
and ( n18679 , n18657 , n18678 );
not ( n18680 , n18678 );
and ( n18681 , n18646 , n18647 );
xor ( n18682 , n18680 , n18681 );
and ( n18683 , n18682 , n18528 );
or ( n18684 , n18679 , n18683 );
buf ( n18685 , n18684 );
not ( n18686 , n18685 );
buf ( n18687 , n18686 );
buf ( n18688 , n18687 );
not ( n18689 , n18688 );
or ( n18690 , n18656 , n18689 );
not ( n18691 , n18528 );
not ( n18692 , n18306 );
and ( n18693 , n18692 , n17972 );
xor ( n18694 , n17972 , n17883 );
and ( n18695 , n18660 , n18661 );
xor ( n18696 , n18694 , n18695 );
and ( n18697 , n18696 , n18306 );
or ( n18698 , n18693 , n18697 );
buf ( n18699 , n18698 );
buf ( n18700 , n18699 );
and ( n18701 , n18666 , n18667 );
xor ( n18702 , n18700 , n18701 );
buf ( n18703 , n18702 );
and ( n18704 , n18703 , n18502 );
buf ( n18705 , RI210d4c00_204);
and ( n18706 , n18705 , n18506 );
buf ( n18707 , RI210d99d0_174);
and ( n18708 , n18707 , n18509 );
buf ( n18709 , RI21a0c010_146);
and ( n18710 , n18709 , n18512 );
or ( n18711 , n18704 , n18706 , n18708 , n18710 );
buf ( n18712 , n18711 );
and ( n18713 , n18691 , n18712 );
not ( n18714 , n18712 );
and ( n18715 , n18680 , n18681 );
xor ( n18716 , n18714 , n18715 );
and ( n18717 , n18716 , n18528 );
or ( n18718 , n18713 , n18717 );
buf ( n18719 , n18718 );
not ( n18720 , n18719 );
buf ( n18721 , n18720 );
buf ( n18722 , n18721 );
not ( n18723 , n18722 );
or ( n18724 , n18690 , n18723 );
not ( n18725 , n18528 );
not ( n18726 , n18306 );
and ( n18727 , n18726 , n17987 );
xor ( n18728 , n17987 , n17883 );
and ( n18729 , n18694 , n18695 );
xor ( n18730 , n18728 , n18729 );
and ( n18731 , n18730 , n18306 );
or ( n18732 , n18727 , n18731 );
buf ( n18733 , n18732 );
buf ( n18734 , n18733 );
and ( n18735 , n18700 , n18701 );
xor ( n18736 , n18734 , n18735 );
buf ( n18737 , n18736 );
and ( n18738 , n18737 , n18502 );
buf ( n18739 , RI210d4b88_205);
and ( n18740 , n18739 , n18506 );
buf ( n18741 , RI210d9160_175);
and ( n18742 , n18741 , n18509 );
buf ( n18743 , RI21a0b908_147);
and ( n18744 , n18743 , n18512 );
or ( n18745 , n18738 , n18740 , n18742 , n18744 );
buf ( n18746 , n18745 );
and ( n18747 , n18725 , n18746 );
not ( n18748 , n18746 );
and ( n18749 , n18714 , n18715 );
xor ( n18750 , n18748 , n18749 );
and ( n18751 , n18750 , n18528 );
or ( n18752 , n18747 , n18751 );
buf ( n18753 , n18752 );
not ( n18754 , n18753 );
buf ( n18755 , n18754 );
buf ( n18756 , n18755 );
not ( n18757 , n18756 );
or ( n18758 , n18724 , n18757 );
not ( n18759 , n18528 );
not ( n18760 , n18306 );
and ( n18761 , n18760 , n18002 );
xor ( n18762 , n18002 , n17883 );
and ( n18763 , n18728 , n18729 );
xor ( n18764 , n18762 , n18763 );
and ( n18765 , n18764 , n18306 );
or ( n18766 , n18761 , n18765 );
buf ( n18767 , n18766 );
buf ( n18768 , n18767 );
and ( n18769 , n18734 , n18735 );
xor ( n18770 , n18768 , n18769 );
buf ( n18771 , n18770 );
and ( n18772 , n18771 , n18502 );
buf ( n18773 , RI210d4b10_206);
and ( n18774 , n18773 , n18506 );
buf ( n18775 , RI210d90e8_176);
and ( n18776 , n18775 , n18509 );
buf ( n18777 , RI21a0b890_148);
and ( n18778 , n18777 , n18512 );
or ( n18779 , n18772 , n18774 , n18776 , n18778 );
buf ( n18780 , n18779 );
and ( n18781 , n18759 , n18780 );
not ( n18782 , n18780 );
and ( n18783 , n18748 , n18749 );
xor ( n18784 , n18782 , n18783 );
and ( n18785 , n18784 , n18528 );
or ( n18786 , n18781 , n18785 );
buf ( n18787 , n18786 );
not ( n18788 , n18787 );
buf ( n18789 , n18788 );
buf ( n18790 , n18789 );
not ( n18791 , n18790 );
or ( n18792 , n18758 , n18791 );
not ( n18793 , n18528 );
not ( n18794 , n18306 );
and ( n18795 , n18794 , n18017 );
xor ( n18796 , n18017 , n17883 );
and ( n18797 , n18762 , n18763 );
xor ( n18798 , n18796 , n18797 );
and ( n18799 , n18798 , n18306 );
or ( n18800 , n18795 , n18799 );
buf ( n18801 , n18800 );
buf ( n18802 , n18801 );
and ( n18803 , n18768 , n18769 );
xor ( n18804 , n18802 , n18803 );
buf ( n18805 , n18804 );
and ( n18806 , n18805 , n18502 );
buf ( n18807 , RI210d42a0_207);
and ( n18808 , n18807 , n18506 );
buf ( n18809 , RI210d9070_177);
and ( n18810 , n18809 , n18509 );
buf ( n18811 , RI21a0b818_149);
and ( n18812 , n18811 , n18512 );
or ( n18813 , n18806 , n18808 , n18810 , n18812 );
buf ( n18814 , n18813 );
and ( n18815 , n18793 , n18814 );
not ( n18816 , n18814 );
and ( n18817 , n18782 , n18783 );
xor ( n18818 , n18816 , n18817 );
and ( n18819 , n18818 , n18528 );
or ( n18820 , n18815 , n18819 );
buf ( n18821 , n18820 );
not ( n18822 , n18821 );
buf ( n18823 , n18822 );
buf ( n18824 , n18823 );
not ( n18825 , n18824 );
or ( n18826 , n18792 , n18825 );
not ( n18827 , n18528 );
not ( n18828 , n18306 );
and ( n18829 , n18828 , n18032 );
xor ( n18830 , n18032 , n17883 );
and ( n18831 , n18796 , n18797 );
xor ( n18832 , n18830 , n18831 );
and ( n18833 , n18832 , n18306 );
or ( n18834 , n18829 , n18833 );
buf ( n18835 , n18834 );
buf ( n18836 , n18835 );
and ( n18837 , n18802 , n18803 );
xor ( n18838 , n18836 , n18837 );
buf ( n18839 , n18838 );
and ( n18840 , n18839 , n18502 );
buf ( n18841 , RI210d8788_179);
and ( n18842 , n18841 , n18506 );
buf ( n18843 , RI21a0b728_151);
and ( n18844 , n18843 , n18509 );
buf ( n18845 , RI21a0de88_123);
and ( n18846 , n18845 , n18512 );
or ( n18847 , n18840 , n18842 , n18844 , n18846 );
buf ( n18848 , n18847 );
and ( n18849 , n18827 , n18848 );
not ( n18850 , n18848 );
and ( n18851 , n18816 , n18817 );
xor ( n18852 , n18850 , n18851 );
and ( n18853 , n18852 , n18528 );
or ( n18854 , n18849 , n18853 );
buf ( n18855 , n18854 );
not ( n18856 , n18855 );
buf ( n18857 , n18856 );
buf ( n18858 , n18857 );
not ( n18859 , n18858 );
or ( n18860 , n18826 , n18859 );
not ( n18861 , n18528 );
not ( n18862 , n18306 );
and ( n18863 , n18862 , n18047 );
xor ( n18864 , n18047 , n17883 );
and ( n18865 , n18830 , n18831 );
xor ( n18866 , n18864 , n18865 );
and ( n18867 , n18866 , n18306 );
or ( n18868 , n18863 , n18867 );
buf ( n18869 , n18868 );
buf ( n18870 , n18869 );
and ( n18871 , n18836 , n18837 );
xor ( n18872 , n18870 , n18871 );
buf ( n18873 , n18872 );
and ( n18874 , n18873 , n18502 );
buf ( n18875 , RI210d8710_180);
and ( n18876 , n18875 , n18506 );
buf ( n18877 , RI21a0b6b0_152);
and ( n18878 , n18877 , n18509 );
buf ( n18879 , RI21a0de10_124);
and ( n18880 , n18879 , n18512 );
or ( n18881 , n18874 , n18876 , n18878 , n18880 );
buf ( n18882 , n18881 );
and ( n18883 , n18861 , n18882 );
not ( n18884 , n18882 );
and ( n18885 , n18850 , n18851 );
xor ( n18886 , n18884 , n18885 );
and ( n18887 , n18886 , n18528 );
or ( n18888 , n18883 , n18887 );
buf ( n18889 , n18888 );
not ( n18890 , n18889 );
buf ( n18891 , n18890 );
buf ( n18892 , n18891 );
not ( n18893 , n18892 );
or ( n18894 , n18860 , n18893 );
not ( n18895 , n18528 );
not ( n18896 , n18306 );
and ( n18897 , n18896 , n18062 );
xor ( n18898 , n18062 , n17883 );
and ( n18899 , n18864 , n18865 );
xor ( n18900 , n18898 , n18899 );
and ( n18901 , n18900 , n18306 );
or ( n18902 , n18897 , n18901 );
buf ( n18903 , n18902 );
buf ( n18904 , n18903 );
and ( n18905 , n18870 , n18871 );
xor ( n18906 , n18904 , n18905 );
buf ( n18907 , n18906 );
and ( n18908 , n18907 , n18502 );
buf ( n18909 , RI210d8698_181);
and ( n18910 , n18909 , n18506 );
buf ( n18911 , RI21a0afa8_153);
and ( n18912 , n18911 , n18509 );
buf ( n18913 , RI21a0dd98_125);
and ( n18914 , n18913 , n18512 );
or ( n18915 , n18908 , n18910 , n18912 , n18914 );
buf ( n18916 , n18915 );
and ( n18917 , n18895 , n18916 );
not ( n18918 , n18916 );
and ( n18919 , n18884 , n18885 );
xor ( n18920 , n18918 , n18919 );
and ( n18921 , n18920 , n18528 );
or ( n18922 , n18917 , n18921 );
buf ( n18923 , n18922 );
not ( n18924 , n18923 );
buf ( n18925 , n18924 );
buf ( n18926 , n18925 );
not ( n18927 , n18926 );
or ( n18928 , n18894 , n18927 );
not ( n18929 , n18528 );
not ( n18930 , n18306 );
and ( n18931 , n18930 , n18077 );
xor ( n18932 , n18077 , n17883 );
and ( n18933 , n18898 , n18899 );
xor ( n18934 , n18932 , n18933 );
and ( n18935 , n18934 , n18306 );
or ( n18936 , n18931 , n18935 );
buf ( n18937 , n18936 );
buf ( n18938 , n18937 );
and ( n18939 , n18904 , n18905 );
xor ( n18940 , n18938 , n18939 );
buf ( n18941 , n18940 );
and ( n18942 , n18941 , n18502 );
buf ( n18943 , RI210d8620_182);
and ( n18944 , n18943 , n18506 );
buf ( n18945 , RI21a0af30_154);
and ( n18946 , n18945 , n18509 );
buf ( n18947 , RI21a0dd20_126);
and ( n18948 , n18947 , n18512 );
or ( n18949 , n18942 , n18944 , n18946 , n18948 );
buf ( n18950 , n18949 );
and ( n18951 , n18929 , n18950 );
not ( n18952 , n18950 );
and ( n18953 , n18918 , n18919 );
xor ( n18954 , n18952 , n18953 );
and ( n18955 , n18954 , n18528 );
or ( n18956 , n18951 , n18955 );
buf ( n18957 , n18956 );
not ( n18958 , n18957 );
buf ( n18959 , n18958 );
buf ( n18960 , n18959 );
not ( n18961 , n18960 );
or ( n18962 , n18928 , n18961 );
not ( n18963 , n18528 );
not ( n18964 , n18306 );
and ( n18965 , n18964 , n18092 );
xor ( n18966 , n18092 , n17883 );
and ( n18967 , n18932 , n18933 );
xor ( n18968 , n18966 , n18967 );
and ( n18969 , n18968 , n18306 );
or ( n18970 , n18965 , n18969 );
buf ( n18971 , n18970 );
buf ( n18972 , n18971 );
and ( n18973 , n18938 , n18939 );
xor ( n18974 , n18972 , n18973 );
buf ( n18975 , n18974 );
and ( n18976 , n18975 , n18502 );
buf ( n18977 , RI210d7db0_183);
and ( n18978 , n18977 , n18506 );
buf ( n18979 , RI21a0aeb8_155);
and ( n18980 , n18979 , n18509 );
buf ( n18981 , RI21a0dca8_127);
and ( n18982 , n18981 , n18512 );
or ( n18983 , n18976 , n18978 , n18980 , n18982 );
buf ( n18984 , n18983 );
and ( n18985 , n18963 , n18984 );
not ( n18986 , n18984 );
and ( n18987 , n18952 , n18953 );
xor ( n18988 , n18986 , n18987 );
and ( n18989 , n18988 , n18528 );
or ( n18990 , n18985 , n18989 );
buf ( n18991 , n18990 );
not ( n18992 , n18991 );
buf ( n18993 , n18992 );
buf ( n18994 , n18993 );
not ( n18995 , n18994 );
or ( n18996 , n18962 , n18995 );
not ( n18997 , n18528 );
not ( n18998 , n18306 );
and ( n18999 , n18998 , n18107 );
xor ( n19000 , n18107 , n17883 );
and ( n19001 , n18966 , n18967 );
xor ( n19002 , n19000 , n19001 );
and ( n19003 , n19002 , n18306 );
or ( n19004 , n18999 , n19003 );
buf ( n19005 , n19004 );
buf ( n19006 , n19005 );
and ( n19007 , n18972 , n18973 );
xor ( n19008 , n19006 , n19007 );
buf ( n19009 , n19008 );
and ( n19010 , n19009 , n18502 );
buf ( n19011 , RI210d7d38_184);
and ( n19012 , n19011 , n18506 );
buf ( n19013 , RI21a0ae40_156);
and ( n19014 , n19013 , n18509 );
buf ( n19015 , RI21a0dc30_128);
and ( n19016 , n19015 , n18512 );
or ( n19017 , n19010 , n19012 , n19014 , n19016 );
buf ( n19018 , n19017 );
and ( n19019 , n18997 , n19018 );
not ( n19020 , n19018 );
and ( n19021 , n18986 , n18987 );
xor ( n19022 , n19020 , n19021 );
and ( n19023 , n19022 , n18528 );
or ( n19024 , n19019 , n19023 );
buf ( n19025 , n19024 );
not ( n19026 , n19025 );
buf ( n19027 , n19026 );
buf ( n19028 , n19027 );
not ( n19029 , n19028 );
or ( n19030 , n18996 , n19029 );
not ( n19031 , n18528 );
not ( n19032 , n18306 );
and ( n19033 , n19032 , n18122 );
xor ( n19034 , n18122 , n17883 );
and ( n19035 , n19000 , n19001 );
xor ( n19036 , n19034 , n19035 );
and ( n19037 , n19036 , n18306 );
or ( n19038 , n19033 , n19037 );
buf ( n19039 , n19038 );
buf ( n19040 , n19039 );
and ( n19041 , n19006 , n19007 );
xor ( n19042 , n19040 , n19041 );
buf ( n19043 , n19042 );
and ( n19044 , n19043 , n18502 );
buf ( n19045 , RI210ce8a0_246);
and ( n19046 , n19045 , n18506 );
buf ( n19047 , RI210cf278_242);
and ( n19048 , n19047 , n18509 );
buf ( n19049 , RI21a0d528_129);
and ( n19050 , n19049 , n18512 );
or ( n19051 , n19044 , n19046 , n19048 , n19050 );
buf ( n19052 , n19051 );
and ( n19053 , n19031 , n19052 );
not ( n19054 , n19052 );
and ( n19055 , n19020 , n19021 );
xor ( n19056 , n19054 , n19055 );
and ( n19057 , n19056 , n18528 );
or ( n19058 , n19053 , n19057 );
buf ( n19059 , n19058 );
not ( n19060 , n19059 );
buf ( n19061 , n19060 );
buf ( n19062 , n19061 );
not ( n19063 , n19062 );
or ( n19064 , n19030 , n19063 );
not ( n19065 , n18528 );
not ( n19066 , n18306 );
and ( n19067 , n19066 , n18137 );
xor ( n19068 , n18137 , n17883 );
and ( n19069 , n19034 , n19035 );
xor ( n19070 , n19068 , n19069 );
and ( n19071 , n19070 , n18306 );
or ( n19072 , n19067 , n19071 );
buf ( n19073 , n19072 );
buf ( n19074 , n19073 );
and ( n19075 , n19040 , n19041 );
xor ( n19076 , n19074 , n19075 );
buf ( n19077 , n19076 );
and ( n19078 , n19077 , n18502 );
buf ( n19079 , RI210d7cc0_185);
and ( n19080 , n19079 , n18506 );
buf ( n19081 , RI210cea08_243);
and ( n19082 , n19081 , n18509 );
buf ( n19083 , RI210cfc50_238);
and ( n19084 , n19083 , n18512 );
or ( n19085 , n19078 , n19080 , n19082 , n19084 );
buf ( n19086 , n19085 );
and ( n19087 , n19065 , n19086 );
not ( n19088 , n19086 );
and ( n19089 , n19054 , n19055 );
xor ( n19090 , n19088 , n19089 );
and ( n19091 , n19090 , n18528 );
or ( n19092 , n19087 , n19091 );
buf ( n19093 , n19092 );
not ( n19094 , n19093 );
buf ( n19095 , n19094 );
buf ( n19096 , n19095 );
not ( n19097 , n19096 );
or ( n19098 , n19064 , n19097 );
not ( n19099 , n18528 );
not ( n19100 , n18306 );
and ( n19101 , n19100 , n18152 );
xor ( n19102 , n18152 , n17883 );
and ( n19103 , n19068 , n19069 );
xor ( n19104 , n19102 , n19103 );
and ( n19105 , n19104 , n18306 );
or ( n19106 , n19101 , n19105 );
buf ( n19107 , n19106 );
buf ( n19108 , n19107 );
and ( n19109 , n19074 , n19075 );
xor ( n19110 , n19108 , n19109 );
buf ( n19111 , n19110 );
and ( n19112 , n19111 , n18502 );
buf ( n19113 , RI210ce030_247);
and ( n19114 , n19113 , n18506 );
buf ( n19115 , RI21a0adc8_157);
and ( n19116 , n19115 , n18509 );
buf ( n19117 , RI21a0d4b0_130);
and ( n19118 , n19117 , n18512 );
or ( n19119 , n19112 , n19114 , n19116 , n19118 );
buf ( n19120 , n19119 );
and ( n19121 , n19099 , n19120 );
not ( n19122 , n19120 );
and ( n19123 , n19088 , n19089 );
xor ( n19124 , n19122 , n19123 );
and ( n19125 , n19124 , n18528 );
or ( n19126 , n19121 , n19125 );
buf ( n19127 , n19126 );
not ( n19128 , n19127 );
buf ( n19129 , n19128 );
buf ( n19130 , n19129 );
not ( n19131 , n19130 );
or ( n19132 , n19098 , n19131 );
not ( n19133 , n18528 );
not ( n19134 , n18306 );
and ( n19135 , n19134 , n18167 );
xor ( n19136 , n18167 , n17883 );
and ( n19137 , n19102 , n19103 );
xor ( n19138 , n19136 , n19137 );
and ( n19139 , n19138 , n18306 );
or ( n19140 , n19135 , n19139 );
buf ( n19141 , n19140 );
buf ( n19142 , n19141 );
and ( n19143 , n19108 , n19109 );
xor ( n19144 , n19142 , n19143 );
buf ( n19145 , n19144 );
and ( n19146 , n19145 , n18502 );
buf ( n19147 , RI210d7c48_186);
and ( n19148 , n19147 , n18506 );
buf ( n19149 , RI210ce990_244);
and ( n19150 , n19149 , n18509 );
buf ( n19151 , RI210cf3e0_239);
and ( n19152 , n19151 , n18512 );
or ( n19153 , n19146 , n19148 , n19150 , n19152 );
buf ( n19154 , n19153 );
and ( n19155 , n19133 , n19154 );
not ( n19156 , n19154 );
and ( n19157 , n19122 , n19123 );
xor ( n19158 , n19156 , n19157 );
and ( n19159 , n19158 , n18528 );
or ( n19160 , n19155 , n19159 );
buf ( n19161 , n19160 );
not ( n19162 , n19161 );
buf ( n19163 , n19162 );
buf ( n19164 , n19163 );
not ( n19165 , n19164 );
or ( n19166 , n19132 , n19165 );
not ( n19167 , n18528 );
not ( n19168 , n18306 );
and ( n19169 , n19168 , n18182 );
xor ( n19170 , n18182 , n17883 );
and ( n19171 , n19136 , n19137 );
xor ( n19172 , n19170 , n19171 );
and ( n19173 , n19172 , n18306 );
or ( n19174 , n19169 , n19173 );
buf ( n19175 , n19174 );
buf ( n19176 , n19175 );
and ( n19177 , n19142 , n19143 );
xor ( n19178 , n19176 , n19177 );
buf ( n19179 , n19178 );
and ( n19180 , n19179 , n18502 );
buf ( n19181 , RI210d7360_188);
and ( n19182 , n19181 , n18506 );
buf ( n19183 , RI210ce918_245);
and ( n19184 , n19183 , n18509 );
buf ( n19185 , RI210cf368_240);
and ( n19186 , n19185 , n18512 );
or ( n19187 , n19180 , n19182 , n19184 , n19186 );
buf ( n19188 , n19187 );
and ( n19189 , n19167 , n19188 );
not ( n19190 , n19188 );
and ( n19191 , n19156 , n19157 );
xor ( n19192 , n19190 , n19191 );
and ( n19193 , n19192 , n18528 );
or ( n19194 , n19189 , n19193 );
buf ( n19195 , n19194 );
not ( n19196 , n19195 );
buf ( n19197 , n19196 );
buf ( n19198 , n19197 );
not ( n19199 , n19198 );
or ( n19200 , n19166 , n19199 );
not ( n19201 , n18528 );
not ( n19202 , n18306 );
and ( n19203 , n19202 , n18197 );
xor ( n19204 , n18197 , n17883 );
and ( n19205 , n19170 , n19171 );
xor ( n19206 , n19204 , n19205 );
and ( n19207 , n19206 , n18306 );
or ( n19208 , n19203 , n19207 );
buf ( n19209 , n19208 );
buf ( n19210 , n19209 );
and ( n19211 , n19176 , n19177 );
xor ( n19212 , n19210 , n19211 );
buf ( n19213 , n19212 );
and ( n19214 , n19213 , n18502 );
buf ( n19215 , RI210d72e8_189);
and ( n19216 , n19215 , n18506 );
buf ( n19217 , RI21a0a648_159);
and ( n19218 , n19217 , n18509 );
buf ( n19219 , RI21a0d3c0_132);
and ( n19220 , n19219 , n18512 );
or ( n19221 , n19214 , n19216 , n19218 , n19220 );
buf ( n19222 , n19221 );
and ( n19223 , n19201 , n19222 );
not ( n19224 , n19222 );
and ( n19225 , n19190 , n19191 );
xor ( n19226 , n19224 , n19225 );
and ( n19227 , n19226 , n18528 );
or ( n19228 , n19223 , n19227 );
buf ( n19229 , n19228 );
not ( n19230 , n19229 );
buf ( n19231 , n19230 );
buf ( n19232 , n19231 );
not ( n19233 , n19232 );
or ( n19234 , n19200 , n19233 );
not ( n19235 , n18528 );
not ( n19236 , n18306 );
and ( n19237 , n19236 , n18212 );
xor ( n19238 , n18212 , n17883 );
and ( n19239 , n19204 , n19205 );
xor ( n19240 , n19238 , n19239 );
and ( n19241 , n19240 , n18306 );
or ( n19242 , n19237 , n19241 );
buf ( n19243 , n19242 );
buf ( n19244 , n19243 );
and ( n19245 , n19210 , n19211 );
xor ( n19246 , n19244 , n19245 );
buf ( n19247 , n19246 );
and ( n19248 , n19247 , n18502 );
buf ( n19249 , RI210d7270_190);
and ( n19250 , n19249 , n18506 );
buf ( n19251 , RI21a0a5d0_160);
and ( n19252 , n19251 , n18509 );
buf ( n19253 , RI21a0d348_133);
and ( n19254 , n19253 , n18512 );
or ( n19255 , n19248 , n19250 , n19252 , n19254 );
buf ( n19256 , n19255 );
and ( n19257 , n19235 , n19256 );
not ( n19258 , n19256 );
and ( n19259 , n19224 , n19225 );
xor ( n19260 , n19258 , n19259 );
and ( n19261 , n19260 , n18528 );
or ( n19262 , n19257 , n19261 );
buf ( n19263 , n19262 );
not ( n19264 , n19263 );
buf ( n19265 , n19264 );
buf ( n19266 , n19265 );
not ( n19267 , n19266 );
or ( n19268 , n19234 , n19267 );
not ( n19269 , n18528 );
not ( n19270 , n18306 );
and ( n19271 , n19270 , n18227 );
xor ( n19272 , n18227 , n17883 );
and ( n19273 , n19238 , n19239 );
xor ( n19274 , n19272 , n19273 );
and ( n19275 , n19274 , n18306 );
or ( n19276 , n19271 , n19275 );
buf ( n19277 , n19276 );
buf ( n19278 , n19277 );
and ( n19279 , n19244 , n19245 );
xor ( n19280 , n19278 , n19279 );
buf ( n19281 , n19280 );
and ( n19282 , n19281 , n18502 );
buf ( n19283 , RI210d6a00_191);
and ( n19284 , n19283 , n18506 );
buf ( n19285 , RI21a0a558_161);
and ( n19286 , n19285 , n18509 );
buf ( n19287 , RI21a0d2d0_134);
and ( n19288 , n19287 , n18512 );
or ( n19289 , n19282 , n19284 , n19286 , n19288 );
buf ( n19290 , n19289 );
and ( n19291 , n19269 , n19290 );
not ( n19292 , n19290 );
and ( n19293 , n19258 , n19259 );
xor ( n19294 , n19292 , n19293 );
and ( n19295 , n19294 , n18528 );
or ( n19296 , n19291 , n19295 );
buf ( n19297 , n19296 );
not ( n19298 , n19297 );
buf ( n19299 , n19298 );
buf ( n19300 , n19299 );
not ( n19301 , n19300 );
or ( n19302 , n19268 , n19301 );
not ( n19303 , n18528 );
not ( n19304 , n18306 );
and ( n19305 , n19304 , n18242 );
xor ( n19306 , n18242 , n17883 );
and ( n19307 , n19272 , n19273 );
xor ( n19308 , n19306 , n19307 );
and ( n19309 , n19308 , n18306 );
or ( n19310 , n19305 , n19309 );
buf ( n19311 , n19310 );
buf ( n19312 , n19311 );
and ( n19313 , n19278 , n19279 );
xor ( n19314 , n19312 , n19313 );
buf ( n19315 , n19314 );
and ( n19316 , n19315 , n18502 );
buf ( n19317 , RI210d6988_192);
and ( n19318 , n19317 , n18506 );
buf ( n19319 , RI21a09e50_162);
and ( n19320 , n19319 , n18509 );
buf ( n19321 , RI21a0cbc8_135);
and ( n19322 , n19321 , n18512 );
or ( n19323 , n19316 , n19318 , n19320 , n19322 );
buf ( n19324 , n19323 );
and ( n19325 , n19303 , n19324 );
not ( n19326 , n19324 );
and ( n19327 , n19292 , n19293 );
xor ( n19328 , n19326 , n19327 );
and ( n19329 , n19328 , n18528 );
or ( n19330 , n19325 , n19329 );
buf ( n19331 , n19330 );
not ( n19332 , n19331 );
buf ( n19333 , n19332 );
buf ( n19334 , n19333 );
not ( n19335 , n19334 );
or ( n19336 , n19302 , n19335 );
not ( n19337 , n18528 );
not ( n19338 , n18306 );
and ( n19339 , n19338 , n18257 );
xor ( n19340 , n18257 , n17883 );
and ( n19341 , n19306 , n19307 );
xor ( n19342 , n19340 , n19341 );
and ( n19343 , n19342 , n18306 );
or ( n19344 , n19339 , n19343 );
buf ( n19345 , n19344 );
buf ( n19346 , n19345 );
and ( n19347 , n19312 , n19313 );
xor ( n19348 , n19346 , n19347 );
buf ( n19349 , n19348 );
and ( n19350 , n19349 , n18502 );
and ( n19351 , n17453 , n18506 );
buf ( n19352 , RI21a09dd8_163);
and ( n19353 , n19352 , n18509 );
buf ( n19354 , RI21a0cb50_136);
and ( n19355 , n19354 , n18512 );
or ( n19356 , n19350 , n19351 , n19353 , n19355 );
buf ( n19357 , n19356 );
and ( n19358 , n19337 , n19357 );
not ( n19359 , n19357 );
and ( n19360 , n19326 , n19327 );
xor ( n19361 , n19359 , n19360 );
and ( n19362 , n19361 , n18528 );
or ( n19363 , n19358 , n19362 );
buf ( n19364 , n19363 );
not ( n19365 , n19364 );
buf ( n19366 , n19365 );
buf ( n19367 , n19366 );
not ( n19368 , n19367 );
or ( n19369 , n19336 , n19368 );
not ( n19370 , n18528 );
not ( n19371 , n18306 );
and ( n19372 , n19371 , n18272 );
xor ( n19373 , n18272 , n17883 );
and ( n19374 , n19340 , n19341 );
xor ( n19375 , n19373 , n19374 );
and ( n19376 , n19375 , n18306 );
or ( n19377 , n19372 , n19376 );
buf ( n19378 , n19377 );
buf ( n19379 , n19378 );
and ( n19380 , n19346 , n19347 );
xor ( n19381 , n19379 , n19380 );
buf ( n19382 , n19381 );
and ( n19383 , n19382 , n18502 );
buf ( n19384 , RI210d6898_194);
and ( n19385 , n19384 , n18506 );
buf ( n19386 , RI21a09478_164);
and ( n19387 , n19386 , n18509 );
buf ( n19388 , RI21a0cad8_137);
and ( n19389 , n19388 , n18512 );
or ( n19390 , n19383 , n19385 , n19387 , n19389 );
buf ( n19391 , n19390 );
and ( n19392 , n19370 , n19391 );
not ( n19393 , n19391 );
and ( n19394 , n19359 , n19360 );
xor ( n19395 , n19393 , n19394 );
and ( n19396 , n19395 , n18528 );
or ( n19397 , n19392 , n19396 );
buf ( n19398 , n19397 );
not ( n19399 , n19398 );
buf ( n19400 , n19399 );
buf ( n19401 , n19400 );
not ( n19402 , n19401 );
or ( n19403 , n19369 , n19402 );
not ( n19404 , n18528 );
not ( n19405 , n18306 );
and ( n19406 , n19405 , n18287 );
xor ( n19407 , n18287 , n17883 );
and ( n19408 , n19373 , n19374 );
xor ( n19409 , n19407 , n19408 );
and ( n19410 , n19409 , n18306 );
or ( n19411 , n19406 , n19410 );
buf ( n19412 , n19411 );
buf ( n19413 , n19412 );
and ( n19414 , n19379 , n19380 );
xor ( n19415 , n19413 , n19414 );
buf ( n19416 , n19415 );
and ( n19417 , n19416 , n18502 );
buf ( n19418 , RI210d6028_195);
and ( n19419 , n19418 , n18506 );
buf ( n19420 , RI210dadf8_165);
and ( n19421 , n19420 , n18509 );
buf ( n19422 , RI21a0ca60_138);
and ( n19423 , n19422 , n18512 );
or ( n19424 , n19417 , n19419 , n19421 , n19423 );
buf ( n19425 , n19424 );
and ( n19426 , n19404 , n19425 );
not ( n19427 , n19425 );
and ( n19428 , n19393 , n19394 );
xor ( n19429 , n19427 , n19428 );
and ( n19430 , n19429 , n18528 );
or ( n19431 , n19426 , n19430 );
buf ( n19432 , n19431 );
not ( n19433 , n19432 );
buf ( n19434 , n19433 );
buf ( n19435 , n19434 );
not ( n19436 , n19435 );
or ( n19437 , n19403 , n19436 );
not ( n19438 , n18528 );
not ( n19439 , n18306 );
and ( n19440 , n19439 , n18302 );
xor ( n19441 , n18302 , n17883 );
and ( n19442 , n19407 , n19408 );
xor ( n19443 , n19441 , n19442 );
and ( n19444 , n19443 , n18306 );
or ( n19445 , n19440 , n19444 );
buf ( n19446 , n19445 );
buf ( n19447 , n19446 );
and ( n19448 , n19413 , n19414 );
xor ( n19449 , n19447 , n19448 );
buf ( n19450 , n19449 );
and ( n19451 , n19450 , n18502 );
buf ( n19452 , RI210d5fb0_196);
and ( n19453 , n19452 , n18506 );
buf ( n19454 , RI210dad80_166);
and ( n19455 , n19454 , n18509 );
buf ( n19456 , RI21a0c9e8_139);
and ( n19457 , n19456 , n18512 );
or ( n19458 , n19451 , n19453 , n19455 , n19457 );
buf ( n19459 , n19458 );
and ( n19460 , n19438 , n19459 );
not ( n19461 , n19459 );
and ( n19462 , n19427 , n19428 );
xor ( n19463 , n19461 , n19462 );
and ( n19464 , n19463 , n18528 );
or ( n19465 , n19460 , n19464 );
buf ( n19466 , n19465 );
not ( n19467 , n19466 );
buf ( n19468 , n19467 );
buf ( n19469 , n19468 );
not ( n19470 , n19469 );
or ( n19471 , n19437 , n19470 );
buf ( n19472 , n19471 );
buf ( n19473 , n19472 );
and ( n19474 , n19473 , n18528 );
not ( n19475 , n19474 );
and ( n19476 , n19475 , n19335 );
xor ( n19477 , n19335 , n18528 );
xor ( n19478 , n19301 , n18528 );
xor ( n19479 , n19267 , n18528 );
xor ( n19480 , n19233 , n18528 );
xor ( n19481 , n19199 , n18528 );
xor ( n19482 , n19165 , n18528 );
xor ( n19483 , n19131 , n18528 );
xor ( n19484 , n19097 , n18528 );
xor ( n19485 , n19063 , n18528 );
xor ( n19486 , n19029 , n18528 );
xor ( n19487 , n18995 , n18528 );
xor ( n19488 , n18961 , n18528 );
xor ( n19489 , n18927 , n18528 );
xor ( n19490 , n18893 , n18528 );
xor ( n19491 , n18859 , n18528 );
xor ( n19492 , n18825 , n18528 );
xor ( n19493 , n18791 , n18528 );
xor ( n19494 , n18757 , n18528 );
xor ( n19495 , n18723 , n18528 );
xor ( n19496 , n18689 , n18528 );
xor ( n19497 , n18655 , n18528 );
xor ( n19498 , n18622 , n18528 );
xor ( n19499 , n18589 , n18528 );
xor ( n19500 , n18558 , n18528 );
xor ( n19501 , n18520 , n18528 );
and ( n19502 , n19501 , n18528 );
and ( n19503 , n19500 , n19502 );
and ( n19504 , n19499 , n19503 );
and ( n19505 , n19498 , n19504 );
and ( n19506 , n19497 , n19505 );
and ( n19507 , n19496 , n19506 );
and ( n19508 , n19495 , n19507 );
and ( n19509 , n19494 , n19508 );
and ( n19510 , n19493 , n19509 );
and ( n19511 , n19492 , n19510 );
and ( n19512 , n19491 , n19511 );
and ( n19513 , n19490 , n19512 );
and ( n19514 , n19489 , n19513 );
and ( n19515 , n19488 , n19514 );
and ( n19516 , n19487 , n19515 );
and ( n19517 , n19486 , n19516 );
and ( n19518 , n19485 , n19517 );
and ( n19519 , n19484 , n19518 );
and ( n19520 , n19483 , n19519 );
and ( n19521 , n19482 , n19520 );
and ( n19522 , n19481 , n19521 );
and ( n19523 , n19480 , n19522 );
and ( n19524 , n19479 , n19523 );
and ( n19525 , n19478 , n19524 );
xor ( n19526 , n19477 , n19525 );
and ( n19527 , n19526 , n19474 );
or ( n19528 , n19476 , n19527 );
buf ( n19529 , n19528 );
buf ( n19530 , n16712 );
not ( n19531 , n19530 );
buf ( n19532 , n17000 );
and ( n19533 , n19531 , n19532 );
not ( n19534 , n19532 );
buf ( n19535 , n17008 );
not ( n19536 , n19535 );
buf ( n19537 , n17016 );
not ( n19538 , n19537 );
buf ( n19539 , n17024 );
not ( n19540 , n19539 );
buf ( n19541 , n16720 );
not ( n19542 , n19541 );
buf ( n19543 , n16729 );
not ( n19544 , n19543 );
buf ( n19545 , n16737 );
not ( n19546 , n19545 );
buf ( n19547 , n16745 );
not ( n19548 , n19547 );
buf ( n19549 , n16753 );
not ( n19550 , n19549 );
buf ( n19551 , n16761 );
not ( n19552 , n19551 );
buf ( n19553 , n16769 );
not ( n19554 , n19553 );
buf ( n19555 , n16777 );
not ( n19556 , n19555 );
buf ( n19557 , n16785 );
not ( n19558 , n19557 );
buf ( n19559 , n16793 );
not ( n19560 , n19559 );
buf ( n19561 , n16801 );
not ( n19562 , n19561 );
buf ( n19563 , n16809 );
not ( n19564 , n19563 );
buf ( n19565 , n16817 );
not ( n19566 , n19565 );
buf ( n19567 , n16825 );
not ( n19568 , n19567 );
buf ( n19569 , n16833 );
not ( n19570 , n19569 );
buf ( n19571 , n16841 );
not ( n19572 , n19571 );
buf ( n19573 , n16849 );
not ( n19574 , n19573 );
buf ( n19575 , n16857 );
not ( n19576 , n19575 );
buf ( n19577 , n16865 );
not ( n19578 , n19577 );
buf ( n19579 , n16873 );
not ( n19580 , n19579 );
buf ( n19581 , n16881 );
not ( n19582 , n19581 );
buf ( n19583 , n16889 );
not ( n19584 , n19583 );
buf ( n19585 , n16897 );
not ( n19586 , n19585 );
buf ( n19587 , n16900 );
not ( n19588 , n19587 );
and ( n19589 , n19586 , n19588 );
and ( n19590 , n19584 , n19589 );
and ( n19591 , n19582 , n19590 );
and ( n19592 , n19580 , n19591 );
and ( n19593 , n19578 , n19592 );
and ( n19594 , n19576 , n19593 );
and ( n19595 , n19574 , n19594 );
and ( n19596 , n19572 , n19595 );
and ( n19597 , n19570 , n19596 );
and ( n19598 , n19568 , n19597 );
and ( n19599 , n19566 , n19598 );
and ( n19600 , n19564 , n19599 );
and ( n19601 , n19562 , n19600 );
and ( n19602 , n19560 , n19601 );
and ( n19603 , n19558 , n19602 );
and ( n19604 , n19556 , n19603 );
and ( n19605 , n19554 , n19604 );
and ( n19606 , n19552 , n19605 );
and ( n19607 , n19550 , n19606 );
and ( n19608 , n19548 , n19607 );
and ( n19609 , n19546 , n19608 );
and ( n19610 , n19544 , n19609 );
and ( n19611 , n19542 , n19610 );
and ( n19612 , n19540 , n19611 );
and ( n19613 , n19538 , n19612 );
and ( n19614 , n19536 , n19613 );
xor ( n19615 , n19534 , n19614 );
and ( n19616 , n19615 , n19530 );
or ( n19617 , n19533 , n19616 );
buf ( n19618 , n19617 );
not ( n19619 , n19618 );
buf ( n19620 , n19619 );
buf ( n19621 , n19620 );
not ( n19622 , n19621 );
buf ( n19623 , n19622 );
buf ( n19624 , n19623 );
buf ( n19625 , n19624 );
not ( n19626 , n19625 );
buf ( n19627 , n19626 );
buf ( n19628 , n19627 );
not ( n19629 , n19628 );
not ( n19630 , n19530 );
buf ( n19631 , n16976 );
not ( n19632 , n19631 );
buf ( n19633 , n16984 );
not ( n19634 , n19633 );
buf ( n19635 , n16992 );
not ( n19636 , n19635 );
and ( n19637 , n19534 , n19614 );
and ( n19638 , n19636 , n19637 );
and ( n19639 , n19634 , n19638 );
and ( n19640 , n19632 , n19639 );
xor ( n19641 , n19630 , n19640 );
buf ( n19642 , n19530 );
and ( n19643 , n19641 , n19642 );
or ( n19644 , C0 , n19643 );
buf ( n19645 , n19644 );
not ( n19646 , n19645 );
buf ( n19647 , n19646 );
buf ( n19648 , n19647 );
not ( n19649 , n19648 );
buf ( n19650 , n19649 );
not ( n19651 , n19650 );
buf ( n19652 , n19651 );
not ( n19653 , n19530 );
and ( n19654 , n19653 , n19631 );
xor ( n19655 , n19632 , n19639 );
and ( n19656 , n19655 , n19530 );
or ( n19657 , n19654 , n19656 );
buf ( n19658 , n19657 );
not ( n19659 , n19658 );
buf ( n19660 , n19659 );
buf ( n19661 , n19660 );
not ( n19662 , n19661 );
buf ( n19663 , n19662 );
not ( n19664 , n19663 );
buf ( n19665 , n19664 );
not ( n19666 , n19530 );
and ( n19667 , n19666 , n19633 );
xor ( n19668 , n19634 , n19638 );
and ( n19669 , n19668 , n19530 );
or ( n19670 , n19667 , n19669 );
buf ( n19671 , n19670 );
not ( n19672 , n19671 );
buf ( n19673 , n19672 );
buf ( n19674 , n19673 );
not ( n19675 , n19674 );
buf ( n19676 , n19675 );
not ( n19677 , n19676 );
buf ( n19678 , n19677 );
not ( n19679 , n19530 );
and ( n19680 , n19679 , n19635 );
xor ( n19681 , n19636 , n19637 );
and ( n19682 , n19681 , n19530 );
or ( n19683 , n19680 , n19682 );
buf ( n19684 , n19683 );
not ( n19685 , n19684 );
buf ( n19686 , n19685 );
buf ( n19687 , n19686 );
not ( n19688 , n19687 );
buf ( n19689 , n19688 );
not ( n19690 , n19689 );
buf ( n19691 , n19690 );
not ( n19692 , n19623 );
buf ( n19693 , n19692 );
and ( n19694 , n19691 , n19693 );
and ( n19695 , n19678 , n19694 );
and ( n19696 , n19665 , n19695 );
and ( n19697 , n19652 , n19696 );
not ( n19698 , n19697 );
buf ( n19699 , n19698 );
buf ( n19700 , n19530 );
and ( n19701 , n19699 , n19700 );
or ( n19702 , C0 , n19701 );
buf ( n19703 , n19702 );
buf ( n19704 , n19703 );
not ( n19705 , n19704 );
not ( n19706 , n19700 );
buf ( n19707 , n19689 );
and ( n19708 , n19706 , n19707 );
xor ( n19709 , n19691 , n19693 );
buf ( n19710 , n19709 );
and ( n19711 , n19710 , n19700 );
or ( n19712 , n19708 , n19711 );
buf ( n19713 , n19712 );
buf ( n19714 , n19713 );
and ( n19715 , n19705 , n19714 );
not ( n19716 , n19714 );
not ( n19717 , n19624 );
xor ( n19718 , n19716 , n19717 );
and ( n19719 , n19718 , n19704 );
or ( n19720 , n19715 , n19719 );
buf ( n19721 , n19720 );
not ( n19722 , n19721 );
buf ( n19723 , n19722 );
buf ( n19724 , n19723 );
not ( n19725 , n19724 );
or ( n19726 , n19629 , n19725 );
buf ( n19727 , n19726 );
buf ( n19728 , n19727 );
and ( n19729 , n19728 , n19704 );
not ( n19730 , n19729 );
and ( n19731 , n19730 , n19629 );
xor ( n19732 , n19629 , n19704 );
xor ( n19733 , n19732 , n19704 );
and ( n19734 , n19733 , n19729 );
or ( n19735 , n19731 , n19734 );
buf ( n19736 , n19735 );
not ( n19737 , n19729 );
and ( n19738 , n19737 , n19725 );
xor ( n19739 , n19725 , n19704 );
and ( n19740 , n19732 , n19704 );
xor ( n19741 , n19739 , n19740 );
and ( n19742 , n19741 , n19729 );
or ( n19743 , n19738 , n19742 );
buf ( n19744 , n19743 );
and ( n19745 , n19736 , n19744 );
and ( n19746 , n19529 , n19745 );
not ( n19747 , n19736 );
and ( n19748 , n19747 , n19744 );
and ( n19749 , n19529 , n19748 );
buf ( n19750 , RI21a16a38_35);
not ( n19751 , n19750 );
buf ( n19752 , n18527 );
buf ( n19753 , n19752 );
not ( n19754 , n19753 );
not ( n19755 , n19752 );
buf ( n19756 , n19390 );
and ( n19757 , n19755 , n19756 );
not ( n19758 , n19756 );
buf ( n19759 , n19356 );
not ( n19760 , n19759 );
buf ( n19761 , n19323 );
not ( n19762 , n19761 );
buf ( n19763 , n19289 );
not ( n19764 , n19763 );
buf ( n19765 , n19255 );
not ( n19766 , n19765 );
buf ( n19767 , n19221 );
not ( n19768 , n19767 );
buf ( n19769 , n19187 );
not ( n19770 , n19769 );
buf ( n19771 , n19153 );
not ( n19772 , n19771 );
buf ( n19773 , n19119 );
not ( n19774 , n19773 );
buf ( n19775 , n19085 );
not ( n19776 , n19775 );
buf ( n19777 , n19051 );
not ( n19778 , n19777 );
buf ( n19779 , n19017 );
not ( n19780 , n19779 );
buf ( n19781 , n18983 );
not ( n19782 , n19781 );
buf ( n19783 , n18949 );
not ( n19784 , n19783 );
buf ( n19785 , n18915 );
not ( n19786 , n19785 );
buf ( n19787 , n18881 );
not ( n19788 , n19787 );
buf ( n19789 , n18847 );
not ( n19790 , n19789 );
buf ( n19791 , n18813 );
not ( n19792 , n19791 );
buf ( n19793 , n18779 );
not ( n19794 , n19793 );
buf ( n19795 , n18745 );
not ( n19796 , n19795 );
buf ( n19797 , n18711 );
not ( n19798 , n19797 );
buf ( n19799 , n18677 );
not ( n19800 , n19799 );
buf ( n19801 , n18643 );
not ( n19802 , n19801 );
buf ( n19803 , n18610 );
not ( n19804 , n19803 );
buf ( n19805 , n18577 );
not ( n19806 , n19805 );
buf ( n19807 , n18546 );
not ( n19808 , n19807 );
buf ( n19809 , n18514 );
not ( n19810 , n19809 );
and ( n19811 , n19808 , n19810 );
and ( n19812 , n19806 , n19811 );
and ( n19813 , n19804 , n19812 );
and ( n19814 , n19802 , n19813 );
and ( n19815 , n19800 , n19814 );
and ( n19816 , n19798 , n19815 );
and ( n19817 , n19796 , n19816 );
and ( n19818 , n19794 , n19817 );
and ( n19819 , n19792 , n19818 );
and ( n19820 , n19790 , n19819 );
and ( n19821 , n19788 , n19820 );
and ( n19822 , n19786 , n19821 );
and ( n19823 , n19784 , n19822 );
and ( n19824 , n19782 , n19823 );
and ( n19825 , n19780 , n19824 );
and ( n19826 , n19778 , n19825 );
and ( n19827 , n19776 , n19826 );
and ( n19828 , n19774 , n19827 );
and ( n19829 , n19772 , n19828 );
and ( n19830 , n19770 , n19829 );
and ( n19831 , n19768 , n19830 );
and ( n19832 , n19766 , n19831 );
and ( n19833 , n19764 , n19832 );
and ( n19834 , n19762 , n19833 );
and ( n19835 , n19760 , n19834 );
xor ( n19836 , n19758 , n19835 );
and ( n19837 , n19836 , n19752 );
or ( n19838 , n19757 , n19837 );
buf ( n19839 , n19838 );
not ( n19840 , n19839 );
buf ( n19841 , n19840 );
buf ( n19842 , n19841 );
not ( n19843 , n19842 );
buf ( n19844 , n19843 );
buf ( n19845 , n19844 );
and ( n19846 , n19754 , n19845 );
not ( n19847 , n19844 );
buf ( n19848 , n19847 );
not ( n19849 , n19752 );
and ( n19850 , n19849 , n19759 );
xor ( n19851 , n19760 , n19834 );
and ( n19852 , n19851 , n19752 );
or ( n19853 , n19850 , n19852 );
buf ( n19854 , n19853 );
not ( n19855 , n19854 );
buf ( n19856 , n19855 );
buf ( n19857 , n19856 );
not ( n19858 , n19857 );
buf ( n19859 , n19858 );
not ( n19860 , n19859 );
buf ( n19861 , n19860 );
not ( n19862 , n19752 );
and ( n19863 , n19862 , n19761 );
xor ( n19864 , n19762 , n19833 );
and ( n19865 , n19864 , n19752 );
or ( n19866 , n19863 , n19865 );
buf ( n19867 , n19866 );
not ( n19868 , n19867 );
buf ( n19869 , n19868 );
buf ( n19870 , n19869 );
not ( n19871 , n19870 );
buf ( n19872 , n19871 );
not ( n19873 , n19872 );
buf ( n19874 , n19873 );
not ( n19875 , n19752 );
and ( n19876 , n19875 , n19763 );
xor ( n19877 , n19764 , n19832 );
and ( n19878 , n19877 , n19752 );
or ( n19879 , n19876 , n19878 );
buf ( n19880 , n19879 );
not ( n19881 , n19880 );
buf ( n19882 , n19881 );
buf ( n19883 , n19882 );
not ( n19884 , n19883 );
buf ( n19885 , n19884 );
not ( n19886 , n19885 );
buf ( n19887 , n19886 );
not ( n19888 , n19752 );
and ( n19889 , n19888 , n19765 );
xor ( n19890 , n19766 , n19831 );
and ( n19891 , n19890 , n19752 );
or ( n19892 , n19889 , n19891 );
buf ( n19893 , n19892 );
not ( n19894 , n19893 );
buf ( n19895 , n19894 );
buf ( n19896 , n19895 );
not ( n19897 , n19896 );
buf ( n19898 , n19897 );
not ( n19899 , n19898 );
buf ( n19900 , n19899 );
not ( n19901 , n19752 );
and ( n19902 , n19901 , n19767 );
xor ( n19903 , n19768 , n19830 );
and ( n19904 , n19903 , n19752 );
or ( n19905 , n19902 , n19904 );
buf ( n19906 , n19905 );
not ( n19907 , n19906 );
buf ( n19908 , n19907 );
buf ( n19909 , n19908 );
not ( n19910 , n19909 );
buf ( n19911 , n19910 );
not ( n19912 , n19911 );
buf ( n19913 , n19912 );
not ( n19914 , n19752 );
and ( n19915 , n19914 , n19769 );
xor ( n19916 , n19770 , n19829 );
and ( n19917 , n19916 , n19752 );
or ( n19918 , n19915 , n19917 );
buf ( n19919 , n19918 );
not ( n19920 , n19919 );
buf ( n19921 , n19920 );
buf ( n19922 , n19921 );
not ( n19923 , n19922 );
buf ( n19924 , n19923 );
not ( n19925 , n19924 );
buf ( n19926 , n19925 );
not ( n19927 , n19752 );
and ( n19928 , n19927 , n19771 );
xor ( n19929 , n19772 , n19828 );
and ( n19930 , n19929 , n19752 );
or ( n19931 , n19928 , n19930 );
buf ( n19932 , n19931 );
not ( n19933 , n19932 );
buf ( n19934 , n19933 );
buf ( n19935 , n19934 );
not ( n19936 , n19935 );
buf ( n19937 , n19936 );
not ( n19938 , n19937 );
buf ( n19939 , n19938 );
not ( n19940 , n19752 );
and ( n19941 , n19940 , n19773 );
xor ( n19942 , n19774 , n19827 );
and ( n19943 , n19942 , n19752 );
or ( n19944 , n19941 , n19943 );
buf ( n19945 , n19944 );
not ( n19946 , n19945 );
buf ( n19947 , n19946 );
buf ( n19948 , n19947 );
not ( n19949 , n19948 );
buf ( n19950 , n19949 );
not ( n19951 , n19950 );
buf ( n19952 , n19951 );
not ( n19953 , n19752 );
and ( n19954 , n19953 , n19775 );
xor ( n19955 , n19776 , n19826 );
and ( n19956 , n19955 , n19752 );
or ( n19957 , n19954 , n19956 );
buf ( n19958 , n19957 );
not ( n19959 , n19958 );
buf ( n19960 , n19959 );
buf ( n19961 , n19960 );
not ( n19962 , n19961 );
buf ( n19963 , n19962 );
not ( n19964 , n19963 );
buf ( n19965 , n19964 );
not ( n19966 , n19752 );
and ( n19967 , n19966 , n19777 );
xor ( n19968 , n19778 , n19825 );
and ( n19969 , n19968 , n19752 );
or ( n19970 , n19967 , n19969 );
buf ( n19971 , n19970 );
not ( n19972 , n19971 );
buf ( n19973 , n19972 );
buf ( n19974 , n19973 );
not ( n19975 , n19974 );
buf ( n19976 , n19975 );
not ( n19977 , n19976 );
buf ( n19978 , n19977 );
not ( n19979 , n19752 );
and ( n19980 , n19979 , n19779 );
xor ( n19981 , n19780 , n19824 );
and ( n19982 , n19981 , n19752 );
or ( n19983 , n19980 , n19982 );
buf ( n19984 , n19983 );
not ( n19985 , n19984 );
buf ( n19986 , n19985 );
buf ( n19987 , n19986 );
not ( n19988 , n19987 );
buf ( n19989 , n19988 );
not ( n19990 , n19989 );
buf ( n19991 , n19990 );
not ( n19992 , n19752 );
and ( n19993 , n19992 , n19781 );
xor ( n19994 , n19782 , n19823 );
and ( n19995 , n19994 , n19752 );
or ( n19996 , n19993 , n19995 );
buf ( n19997 , n19996 );
not ( n19998 , n19997 );
buf ( n19999 , n19998 );
buf ( n20000 , n19999 );
not ( n20001 , n20000 );
buf ( n20002 , n20001 );
not ( n20003 , n20002 );
buf ( n20004 , n20003 );
not ( n20005 , n19752 );
and ( n20006 , n20005 , n19783 );
xor ( n20007 , n19784 , n19822 );
and ( n20008 , n20007 , n19752 );
or ( n20009 , n20006 , n20008 );
buf ( n20010 , n20009 );
not ( n20011 , n20010 );
buf ( n20012 , n20011 );
buf ( n20013 , n20012 );
not ( n20014 , n20013 );
buf ( n20015 , n20014 );
not ( n20016 , n20015 );
buf ( n20017 , n20016 );
not ( n20018 , n19752 );
and ( n20019 , n20018 , n19785 );
xor ( n20020 , n19786 , n19821 );
and ( n20021 , n20020 , n19752 );
or ( n20022 , n20019 , n20021 );
buf ( n20023 , n20022 );
not ( n20024 , n20023 );
buf ( n20025 , n20024 );
buf ( n20026 , n20025 );
not ( n20027 , n20026 );
buf ( n20028 , n20027 );
not ( n20029 , n20028 );
buf ( n20030 , n20029 );
not ( n20031 , n19752 );
and ( n20032 , n20031 , n19787 );
or ( n20033 , n19788 , n19820 );
and ( n20034 , n20033 , n19752 );
or ( n20035 , n20032 , n20034 );
buf ( n20036 , n20035 );
not ( n20037 , n20036 );
buf ( n20038 , n20037 );
buf ( n20039 , n20038 );
not ( n20040 , n20039 );
buf ( n20041 , n20040 );
not ( n20042 , n20041 );
buf ( n20043 , n20042 );
not ( n20044 , n19752 );
and ( n20045 , n20044 , n19789 );
xor ( n20046 , n19790 , n19819 );
and ( n20047 , n20046 , n19752 );
or ( n20048 , n20045 , n20047 );
buf ( n20049 , n20048 );
not ( n20050 , n20049 );
buf ( n20051 , n20050 );
buf ( n20052 , n20051 );
and ( n20053 , C1 , n20052 );
and ( n20054 , C1 , n20053 );
and ( n20055 , C1 , n20054 );
and ( n20056 , C1 , n20055 );
nand ( n20057 , C1 , n20056 );
and ( n20058 , C1 , n20057 );
and ( n20059 , C1 , n20058 );
and ( n20060 , C1 , n20059 );
and ( n20061 , C1 , n20060 );
and ( n20062 , C1 , n20061 );
and ( n20063 , C1 , n20062 );
and ( n20064 , C1 , n20063 );
and ( n20065 , C1 , n20064 );
and ( n20066 , C1 , n20065 );
and ( n20067 , C1 , n20066 );
and ( n20068 , C1 , n20067 );
and ( n20069 , C1 , n20068 );
and ( n20070 , C1 , n20069 );
and ( n20071 , C1 , n20070 );
and ( n20072 , C1 , n20071 );
and ( n20073 , C1 , n20072 );
not ( n20074 , n20073 );
buf ( n20075 , n20074 );
not ( n20076 , n20075 );
buf ( n20077 , n20076 );
not ( n20078 , n19752 );
and ( n20079 , n20078 , n19791 );
xor ( n20080 , n19792 , n19818 );
and ( n20081 , n20080 , n19752 );
or ( n20082 , n20079 , n20081 );
buf ( n20083 , n20082 );
not ( n20084 , n20083 );
buf ( n20085 , n20084 );
buf ( n20086 , n20085 );
and ( n20087 , C1 , n20086 );
and ( n20088 , C1 , n20087 );
and ( n20089 , C1 , n20088 );
and ( n20090 , C1 , n20089 );
and ( n20091 , C1 , n20090 );
and ( n20092 , C1 , n20091 );
and ( n20093 , C1 , n20092 );
and ( n20094 , C1 , n20093 );
and ( n20095 , C1 , n20094 );
and ( n20096 , C1 , n20095 );
and ( n20097 , C1 , n20096 );
and ( n20098 , C1 , n20097 );
and ( n20099 , C1 , n20098 );
and ( n20100 , C1 , n20099 );
and ( n20101 , C1 , n20100 );
and ( n20102 , C1 , n20101 );
and ( n20103 , C1 , n20102 );
and ( n20104 , C1 , n20103 );
and ( n20105 , C1 , n20104 );
and ( n20106 , C1 , n20105 );
and ( n20107 , C1 , n20106 );
buf ( n20108 , n20107 );
not ( n20109 , n20108 );
buf ( n20110 , n20109 );
not ( n20111 , n20110 );
buf ( n20112 , n20111 );
not ( n20113 , n19752 );
and ( n20114 , n20113 , n19793 );
xor ( n20115 , n19794 , n19817 );
and ( n20116 , n20115 , n19752 );
or ( n20117 , n20114 , n20116 );
buf ( n20118 , n20117 );
not ( n20119 , n20118 );
buf ( n20120 , n20119 );
buf ( n20121 , n20120 );
and ( n20122 , C1 , n20121 );
and ( n20123 , C1 , n20122 );
and ( n20124 , C1 , n20123 );
and ( n20125 , C1 , n20124 );
and ( n20126 , C1 , n20125 );
and ( n20127 , C1 , n20126 );
and ( n20128 , C1 , n20127 );
and ( n20129 , C1 , n20128 );
and ( n20130 , C1 , n20129 );
and ( n20131 , C1 , n20130 );
and ( n20132 , C1 , n20131 );
and ( n20133 , C1 , n20132 );
and ( n20134 , C1 , n20133 );
and ( n20135 , C1 , n20134 );
and ( n20136 , C1 , n20135 );
and ( n20137 , C1 , n20136 );
and ( n20138 , C1 , n20137 );
and ( n20139 , C1 , n20138 );
and ( n20140 , C1 , n20139 );
and ( n20141 , C1 , n20140 );
and ( n20142 , C1 , n20141 );
and ( n20143 , C1 , n20142 );
buf ( n20144 , n20143 );
not ( n20145 , n20144 );
buf ( n20146 , n20145 );
not ( n20147 , n20146 );
buf ( n20148 , n20147 );
not ( n20149 , n19752 );
and ( n20150 , n20149 , n19795 );
xor ( n20151 , n19796 , n19816 );
and ( n20152 , n20151 , n19752 );
or ( n20153 , n20150 , n20152 );
buf ( n20154 , n20153 );
not ( n20155 , n20154 );
buf ( n20156 , n20155 );
buf ( n20157 , n20156 );
and ( n20158 , C1 , n20157 );
and ( n20159 , C1 , n20158 );
and ( n20160 , C1 , n20159 );
and ( n20161 , C1 , n20160 );
and ( n20162 , C1 , n20161 );
and ( n20163 , C1 , n20162 );
and ( n20164 , C1 , n20163 );
and ( n20165 , C1 , n20164 );
and ( n20166 , C1 , n20165 );
and ( n20167 , C1 , n20166 );
and ( n20168 , C1 , n20167 );
and ( n20169 , C1 , n20168 );
and ( n20170 , C1 , n20169 );
and ( n20171 , C1 , n20170 );
and ( n20172 , C1 , n20171 );
and ( n20173 , C1 , n20172 );
and ( n20174 , C1 , n20173 );
and ( n20175 , C1 , n20174 );
and ( n20176 , C1 , n20175 );
and ( n20177 , C1 , n20176 );
and ( n20178 , C1 , n20177 );
and ( n20179 , C1 , n20178 );
and ( n20180 , C1 , n20179 );
buf ( n20181 , n20180 );
not ( n20182 , n20181 );
buf ( n20183 , n20182 );
not ( n20184 , n20183 );
buf ( n20185 , n20184 );
not ( n20186 , n19752 );
and ( n20187 , n20186 , n19797 );
xor ( n20188 , n19798 , n19815 );
and ( n20189 , n20188 , n19752 );
or ( n20190 , n20187 , n20189 );
buf ( n20191 , n20190 );
not ( n20192 , n20191 );
buf ( n20193 , n20192 );
buf ( n20194 , n20193 );
and ( n20195 , C1 , n20194 );
and ( n20196 , C1 , n20195 );
and ( n20197 , C1 , n20196 );
and ( n20198 , C1 , n20197 );
and ( n20199 , C1 , n20198 );
and ( n20200 , C1 , n20199 );
and ( n20201 , C1 , n20200 );
and ( n20202 , C1 , n20201 );
and ( n20203 , C1 , n20202 );
and ( n20204 , C1 , n20203 );
and ( n20205 , C1 , n20204 );
and ( n20206 , C1 , n20205 );
and ( n20207 , C1 , n20206 );
nand ( n20208 , C1 , n20207 );
and ( n20209 , C1 , n20208 );
and ( n20210 , C1 , n20209 );
and ( n20211 , C1 , n20210 );
and ( n20212 , C1 , n20211 );
and ( n20213 , C1 , n20212 );
and ( n20214 , C1 , n20213 );
and ( n20215 , C1 , n20214 );
and ( n20216 , C1 , n20215 );
and ( n20217 , C1 , n20216 );
and ( n20218 , C1 , n20217 );
buf ( n20219 , n20218 );
not ( n20220 , n20219 );
buf ( n20221 , n20220 );
not ( n20222 , n20221 );
buf ( n20223 , n20222 );
not ( n20224 , n19752 );
and ( n20225 , n20224 , n19799 );
xor ( n20226 , n19800 , n19814 );
and ( n20227 , n20226 , n19752 );
or ( n20228 , n20225 , n20227 );
buf ( n20229 , n20228 );
not ( n20230 , n20229 );
buf ( n20231 , n20230 );
buf ( n20232 , n20231 );
and ( n20233 , C1 , n20232 );
and ( n20234 , C1 , n20233 );
and ( n20235 , C1 , n20234 );
and ( n20236 , C1 , n20235 );
and ( n20237 , C1 , n20236 );
and ( n20238 , C1 , n20237 );
and ( n20239 , C1 , n20238 );
and ( n20240 , C1 , n20239 );
and ( n20241 , C1 , n20240 );
and ( n20242 , C1 , n20241 );
and ( n20243 , C1 , n20242 );
and ( n20244 , C1 , n20243 );
and ( n20245 , C1 , n20244 );
and ( n20246 , C1 , n20245 );
and ( n20247 , C1 , n20246 );
and ( n20248 , C1 , n20247 );
and ( n20249 , C1 , n20248 );
and ( n20250 , C1 , n20249 );
and ( n20251 , C1 , n20250 );
and ( n20252 , C1 , n20251 );
and ( n20253 , C1 , n20252 );
and ( n20254 , C1 , n20253 );
and ( n20255 , C1 , n20254 );
and ( n20256 , C1 , n20255 );
and ( n20257 , C1 , n20256 );
buf ( n20258 , n20257 );
not ( n20259 , n20258 );
buf ( n20260 , n20259 );
not ( n20261 , n20260 );
buf ( n20262 , n20261 );
not ( n20263 , n19752 );
and ( n20264 , n20263 , n19801 );
xor ( n20265 , n19802 , n19813 );
and ( n20266 , n20265 , n19752 );
or ( n20267 , n20264 , n20266 );
buf ( n20268 , n20267 );
not ( n20269 , n20268 );
buf ( n20270 , n20269 );
buf ( n20271 , n20270 );
and ( n20272 , C1 , n20271 );
and ( n20273 , C1 , n20272 );
and ( n20274 , C1 , n20273 );
and ( n20275 , C1 , n20274 );
and ( n20276 , C1 , n20275 );
and ( n20277 , C1 , n20276 );
and ( n20278 , C1 , n20277 );
and ( n20279 , C1 , n20278 );
and ( n20280 , C1 , n20279 );
and ( n20281 , C1 , n20280 );
and ( n20282 , C1 , n20281 );
and ( n20283 , C1 , n20282 );
and ( n20284 , C1 , n20283 );
and ( n20285 , C1 , n20284 );
and ( n20286 , C1 , n20285 );
and ( n20287 , C1 , n20286 );
and ( n20288 , C1 , n20287 );
and ( n20289 , C1 , n20288 );
and ( n20290 , C1 , n20289 );
and ( n20291 , C1 , n20290 );
and ( n20292 , C1 , n20291 );
and ( n20293 , C1 , n20292 );
and ( n20294 , C1 , n20293 );
and ( n20295 , C1 , n20294 );
and ( n20296 , C1 , n20295 );
and ( n20297 , C1 , n20296 );
buf ( n20298 , n20297 );
not ( n20299 , n20298 );
buf ( n20300 , n20299 );
not ( n20301 , n20300 );
buf ( n20302 , n20301 );
not ( n20303 , n19752 );
and ( n20304 , n20303 , n19803 );
xor ( n20305 , n19804 , n19812 );
and ( n20306 , n20305 , n19752 );
or ( n20307 , n20304 , n20306 );
buf ( n20308 , n20307 );
not ( n20309 , n20308 );
buf ( n20310 , n20309 );
buf ( n20311 , n20310 );
and ( n20312 , C1 , n20311 );
and ( n20313 , C1 , n20312 );
and ( n20314 , C1 , n20313 );
and ( n20315 , C1 , n20314 );
and ( n20316 , C1 , n20315 );
and ( n20317 , C1 , n20316 );
and ( n20318 , C1 , n20317 );
and ( n20319 , C1 , n20318 );
and ( n20320 , C1 , n20319 );
and ( n20321 , C1 , n20320 );
and ( n20322 , C1 , n20321 );
and ( n20323 , C1 , n20322 );
and ( n20324 , C1 , n20323 );
and ( n20325 , C1 , n20324 );
and ( n20326 , C1 , n20325 );
and ( n20327 , C1 , n20326 );
and ( n20328 , C1 , n20327 );
and ( n20329 , C1 , n20328 );
and ( n20330 , C1 , n20329 );
and ( n20331 , C1 , n20330 );
and ( n20332 , C1 , n20331 );
and ( n20333 , C1 , n20332 );
and ( n20334 , C1 , n20333 );
and ( n20335 , C1 , n20334 );
and ( n20336 , C1 , n20335 );
and ( n20337 , C1 , n20336 );
and ( n20338 , C1 , n20337 );
buf ( n20339 , n20338 );
not ( n20340 , n20339 );
buf ( n20341 , n20340 );
not ( n20342 , n20341 );
buf ( n20343 , n20342 );
not ( n20344 , n19752 );
and ( n20345 , n20344 , n19805 );
xor ( n20346 , n19806 , n19811 );
and ( n20347 , n20346 , n19752 );
or ( n20348 , n20345 , n20347 );
buf ( n20349 , n20348 );
not ( n20350 , n20349 );
buf ( n20351 , n20350 );
buf ( n20352 , n20351 );
and ( n20353 , C1 , n20352 );
and ( n20354 , C1 , n20353 );
and ( n20355 , C1 , n20354 );
and ( n20356 , C1 , n20355 );
and ( n20357 , C1 , n20356 );
and ( n20358 , C1 , n20357 );
and ( n20359 , C1 , n20358 );
and ( n20360 , C1 , n20359 );
and ( n20361 , C1 , n20360 );
and ( n20362 , C1 , n20361 );
and ( n20363 , C1 , n20362 );
and ( n20364 , C1 , n20363 );
and ( n20365 , C1 , n20364 );
and ( n20366 , C1 , n20365 );
and ( n20367 , C1 , n20366 );
and ( n20368 , C1 , n20367 );
and ( n20369 , C1 , n20368 );
and ( n20370 , C1 , n20369 );
and ( n20371 , C1 , n20370 );
and ( n20372 , C1 , n20371 );
and ( n20373 , C1 , n20372 );
and ( n20374 , C1 , n20373 );
and ( n20375 , C1 , n20374 );
and ( n20376 , C1 , n20375 );
and ( n20377 , C1 , n20376 );
and ( n20378 , C1 , n20377 );
and ( n20379 , C1 , n20378 );
and ( n20380 , C1 , n20379 );
buf ( n20381 , n20380 );
not ( n20382 , n20381 );
buf ( n20383 , n20382 );
not ( n20384 , n20383 );
buf ( n20385 , n20384 );
not ( n20386 , n19752 );
and ( n20387 , n20386 , n19807 );
xor ( n20388 , n19808 , n19810 );
and ( n20389 , n20388 , n19752 );
or ( n20390 , n20387 , n20389 );
buf ( n20391 , n20390 );
not ( n20392 , n20391 );
buf ( n20393 , n20392 );
buf ( n20394 , n20393 );
and ( n20395 , C1 , n20394 );
and ( n20396 , C1 , n20395 );
and ( n20397 , C1 , n20396 );
and ( n20398 , C1 , n20397 );
and ( n20399 , C1 , n20398 );
and ( n20400 , C1 , n20399 );
and ( n20401 , C1 , n20400 );
and ( n20402 , C1 , n20401 );
and ( n20403 , C1 , n20402 );
and ( n20404 , C1 , n20403 );
and ( n20405 , C1 , n20404 );
and ( n20406 , C1 , n20405 );
and ( n20407 , C1 , n20406 );
and ( n20408 , C1 , n20407 );
and ( n20409 , C1 , n20408 );
and ( n20410 , C1 , n20409 );
and ( n20411 , C1 , n20410 );
and ( n20412 , C1 , n20411 );
and ( n20413 , C1 , n20412 );
and ( n20414 , C1 , n20413 );
and ( n20415 , C1 , n20414 );
and ( n20416 , C1 , n20415 );
and ( n20417 , C1 , n20416 );
and ( n20418 , C1 , n20417 );
and ( n20419 , C1 , n20418 );
and ( n20420 , C1 , n20419 );
and ( n20421 , C1 , n20420 );
and ( n20422 , C1 , n20421 );
and ( n20423 , C1 , n20422 );
buf ( n20424 , n20423 );
not ( n20425 , n20424 );
buf ( n20426 , n20425 );
not ( n20427 , n20426 );
buf ( n20428 , n20427 );
and ( n20429 , n20385 , n20428 );
and ( n20430 , n20343 , n20429 );
and ( n20431 , n20302 , n20430 );
and ( n20432 , n20262 , n20431 );
and ( n20433 , n20223 , n20432 );
and ( n20434 , n20185 , n20433 );
and ( n20435 , n20148 , n20434 );
nand ( n20436 , n20112 , n20435 );
or ( n20437 , n20077 , n20436 );
and ( n20438 , n20043 , n20437 );
and ( n20439 , n20030 , n20438 );
and ( n20440 , n20017 , n20439 );
and ( n20441 , n20004 , n20440 );
and ( n20442 , n19991 , n20441 );
and ( n20443 , n19978 , n20442 );
and ( n20444 , n19965 , n20443 );
and ( n20445 , n19952 , n20444 );
and ( n20446 , n19939 , n20445 );
and ( n20447 , n19926 , n20446 );
and ( n20448 , n19913 , n20447 );
and ( n20449 , n19900 , n20448 );
and ( n20450 , n19887 , n20449 );
and ( n20451 , n19874 , n20450 );
and ( n20452 , n19861 , n20451 );
xor ( n20453 , n19848 , n20452 );
buf ( n20454 , n20453 );
and ( n20455 , n20454 , n19753 );
or ( n20456 , n19846 , n20455 );
buf ( n20457 , n20456 );
and ( n20458 , n19751 , n20457 );
buf ( n20459 , n20426 );
buf ( n20460 , n20459 );
buf ( n20461 , n20460 );
not ( n20462 , n20461 );
buf ( n20463 , n20462 );
buf ( n20464 , n20463 );
not ( n20465 , n20464 );
not ( n20466 , n19752 );
and ( n20467 , n19441 , n19442 );
buf ( n20468 , n20467 );
and ( n20469 , n20468 , n18306 );
or ( n20470 , C0 , n20469 );
buf ( n20471 , n20470 );
buf ( n20472 , n20471 );
and ( n20473 , n19447 , n19448 );
and ( n20474 , n20472 , n20473 );
buf ( n20475 , n20474 );
buf ( n20476 , n20475 );
and ( n20477 , n20476 , n18502 );
buf ( n20478 , RI210d5650_199);
and ( n20479 , n20478 , n18506 );
buf ( n20480 , RI210da420_169);
and ( n20481 , n20480 , n18509 );
buf ( n20482 , RI21a0c1f0_142);
and ( n20483 , n20482 , n18512 );
or ( n20484 , n20477 , n20479 , n20481 , n20483 );
buf ( n20485 , n20484 );
not ( n20486 , n20485 );
xor ( n20487 , n20472 , n20473 );
buf ( n20488 , n20487 );
and ( n20489 , n20488 , n18502 );
buf ( n20490 , RI210d5f38_197);
and ( n20491 , n20490 , n18506 );
buf ( n20492 , RI210da510_167);
and ( n20493 , n20492 , n18509 );
buf ( n20494 , RI21a0c970_140);
and ( n20495 , n20494 , n18512 );
or ( n20496 , n20489 , n20491 , n20493 , n20495 );
buf ( n20497 , n20496 );
not ( n20498 , n20497 );
buf ( n20499 , n19458 );
not ( n20500 , n20499 );
buf ( n20501 , n19424 );
not ( n20502 , n20501 );
and ( n20503 , n19758 , n19835 );
and ( n20504 , n20502 , n20503 );
and ( n20505 , n20500 , n20504 );
and ( n20506 , n20498 , n20505 );
and ( n20507 , n20486 , n20506 );
xor ( n20508 , n20466 , n20507 );
buf ( n20509 , n19752 );
and ( n20510 , n20508 , n20509 );
or ( n20511 , C0 , n20510 );
buf ( n20512 , n20511 );
not ( n20513 , n20512 );
buf ( n20514 , n20513 );
not ( n20515 , n20514 );
buf ( n20516 , n20515 );
not ( n20517 , n20516 );
buf ( n20518 , n20517 );
not ( n20519 , n19752 );
and ( n20520 , n20519 , n20485 );
xor ( n20521 , n20486 , n20506 );
and ( n20522 , n20521 , n19752 );
or ( n20523 , n20520 , n20522 );
buf ( n20524 , n20523 );
not ( n20525 , n20524 );
buf ( n20526 , n20525 );
buf ( n20527 , n20526 );
not ( n20528 , n20527 );
buf ( n20529 , n20528 );
not ( n20530 , n20529 );
buf ( n20531 , n20530 );
not ( n20532 , n19752 );
and ( n20533 , n20532 , n20497 );
xor ( n20534 , n20498 , n20505 );
and ( n20535 , n20534 , n19752 );
or ( n20536 , n20533 , n20535 );
buf ( n20537 , n20536 );
not ( n20538 , n20537 );
buf ( n20539 , n20538 );
buf ( n20540 , n20539 );
not ( n20541 , n20540 );
buf ( n20542 , n20541 );
not ( n20543 , n20542 );
buf ( n20544 , n20543 );
not ( n20545 , n19752 );
and ( n20546 , n20545 , n20499 );
xor ( n20547 , n20500 , n20504 );
and ( n20548 , n20547 , n19752 );
or ( n20549 , n20546 , n20548 );
buf ( n20550 , n20549 );
not ( n20551 , n20550 );
buf ( n20552 , n20551 );
buf ( n20553 , n20552 );
not ( n20554 , n20553 );
buf ( n20555 , n20554 );
not ( n20556 , n20555 );
buf ( n20557 , n20556 );
not ( n20558 , n19752 );
and ( n20559 , n20558 , n20501 );
xor ( n20560 , n20502 , n20503 );
and ( n20561 , n20560 , n19752 );
or ( n20562 , n20559 , n20561 );
buf ( n20563 , n20562 );
not ( n20564 , n20563 );
buf ( n20565 , n20564 );
buf ( n20566 , n20565 );
not ( n20567 , n20566 );
buf ( n20568 , n20567 );
not ( n20569 , n20568 );
buf ( n20570 , n20569 );
and ( n20571 , n19848 , n20452 );
and ( n20572 , n20570 , n20571 );
and ( n20573 , n20557 , n20572 );
and ( n20574 , n20544 , n20573 );
and ( n20575 , n20531 , n20574 );
and ( n20576 , n20518 , n20575 );
not ( n20577 , n20576 );
buf ( n20578 , n20577 );
and ( n20579 , n20578 , n19753 );
or ( n20580 , C0 , n20579 );
buf ( n20581 , n20580 );
buf ( n20582 , n20581 );
not ( n20583 , n20582 );
not ( n20584 , n19753 );
buf ( n20585 , n20383 );
and ( n20586 , n20584 , n20585 );
xor ( n20587 , n20385 , n20428 );
buf ( n20588 , n20587 );
and ( n20589 , n20588 , n19753 );
or ( n20590 , n20586 , n20589 );
buf ( n20591 , n20590 );
buf ( n20592 , n20591 );
and ( n20593 , n20583 , n20592 );
not ( n20594 , n20592 );
not ( n20595 , n20460 );
xor ( n20596 , n20594 , n20595 );
and ( n20597 , n20596 , n20582 );
or ( n20598 , n20593 , n20597 );
buf ( n20599 , n20598 );
not ( n20600 , n20599 );
buf ( n20601 , n20600 );
buf ( n20602 , n20601 );
not ( n20603 , n20602 );
or ( n20604 , n20465 , n20603 );
not ( n20605 , n20582 );
not ( n20606 , n19753 );
buf ( n20607 , n20341 );
and ( n20608 , n20606 , n20607 );
xor ( n20609 , n20343 , n20429 );
buf ( n20610 , n20609 );
and ( n20611 , n20610 , n19753 );
or ( n20612 , n20608 , n20611 );
buf ( n20613 , n20612 );
buf ( n20614 , n20613 );
and ( n20615 , n20605 , n20614 );
not ( n20616 , n20614 );
and ( n20617 , n20594 , n20595 );
xor ( n20618 , n20616 , n20617 );
and ( n20619 , n20618 , n20582 );
or ( n20620 , n20615 , n20619 );
buf ( n20621 , n20620 );
not ( n20622 , n20621 );
buf ( n20623 , n20622 );
buf ( n20624 , n20623 );
not ( n20625 , n20624 );
or ( n20626 , n20604 , n20625 );
not ( n20627 , n20582 );
not ( n20628 , n19753 );
buf ( n20629 , n20300 );
and ( n20630 , n20628 , n20629 );
xor ( n20631 , n20302 , n20430 );
buf ( n20632 , n20631 );
and ( n20633 , n20632 , n19753 );
or ( n20634 , n20630 , n20633 );
buf ( n20635 , n20634 );
buf ( n20636 , n20635 );
and ( n20637 , n20627 , n20636 );
not ( n20638 , n20636 );
and ( n20639 , n20616 , n20617 );
xor ( n20640 , n20638 , n20639 );
and ( n20641 , n20640 , n20582 );
or ( n20642 , n20637 , n20641 );
buf ( n20643 , n20642 );
not ( n20644 , n20643 );
buf ( n20645 , n20644 );
buf ( n20646 , n20645 );
not ( n20647 , n20646 );
or ( n20648 , n20626 , n20647 );
not ( n20649 , n20582 );
not ( n20650 , n19753 );
buf ( n20651 , n20260 );
and ( n20652 , n20650 , n20651 );
xor ( n20653 , n20262 , n20431 );
buf ( n20654 , n20653 );
and ( n20655 , n20654 , n19753 );
nor ( n20656 , n20652 , n20655 );
buf ( n20657 , n20656 );
buf ( n20658 , n20657 );
and ( n20659 , n20649 , n20658 );
not ( n20660 , n20658 );
and ( n20661 , n20638 , n20639 );
or ( n20662 , n20660 , n20661 );
nand ( n20663 , n20662 , n20582 );
nor ( n20664 , n20659 , n20663 );
buf ( n20665 , n20664 );
not ( n20666 , n20665 );
buf ( n20667 , n20666 );
buf ( n20668 , n20667 );
not ( n20669 , n20668 );
or ( n20670 , n20648 , n20669 );
not ( n20671 , n20582 );
not ( n20672 , n19753 );
buf ( n20673 , n20221 );
and ( n20674 , n20672 , n20673 );
xor ( n20675 , n20223 , n20432 );
buf ( n20676 , n20675 );
and ( n20677 , n20676 , n19753 );
or ( n20678 , n20674 , n20677 );
buf ( n20679 , n20678 );
buf ( n20680 , n20679 );
and ( n20681 , n20671 , n20680 );
not ( n20682 , n20680 );
and ( n20683 , n20660 , n20661 );
xor ( n20684 , n20682 , n20683 );
and ( n20685 , n20684 , n20582 );
or ( n20686 , n20681 , n20685 );
buf ( n20687 , n20686 );
not ( n20688 , n20687 );
buf ( n20689 , n20688 );
buf ( n20690 , n20689 );
not ( n20691 , n20690 );
or ( n20692 , n20670 , n20691 );
not ( n20693 , n20582 );
not ( n20694 , n19753 );
buf ( n20695 , n20183 );
and ( n20696 , n20694 , n20695 );
xor ( n20697 , n20185 , n20433 );
buf ( n20698 , n20697 );
and ( n20699 , n20698 , n19753 );
or ( n20700 , n20696 , n20699 );
buf ( n20701 , n20700 );
buf ( n20702 , n20701 );
and ( n20703 , n20693 , n20702 );
not ( n20704 , n20702 );
and ( n20705 , n20682 , n20683 );
xor ( n20706 , n20704 , n20705 );
and ( n20707 , n20706 , n20582 );
or ( n20708 , n20703 , n20707 );
buf ( n20709 , n20708 );
not ( n20710 , n20709 );
buf ( n20711 , n20710 );
buf ( n20712 , n20711 );
not ( n20713 , n20712 );
or ( n20714 , n20692 , n20713 );
not ( n20715 , n20582 );
not ( n20716 , n19753 );
buf ( n20717 , n20146 );
and ( n20718 , n20716 , n20717 );
xor ( n20719 , n20148 , n20434 );
buf ( n20720 , n20719 );
and ( n20721 , n20720 , n19753 );
or ( n20722 , n20718 , n20721 );
buf ( n20723 , n20722 );
buf ( n20724 , n20723 );
and ( n20725 , n20715 , n20724 );
not ( n20726 , n20724 );
and ( n20727 , n20704 , n20705 );
xor ( n20728 , n20726 , n20727 );
and ( n20729 , n20728 , n20582 );
or ( n20730 , n20725 , n20729 );
buf ( n20731 , n20730 );
not ( n20732 , n20731 );
buf ( n20733 , n20732 );
buf ( n20734 , n20733 );
not ( n20735 , n20734 );
or ( n20736 , n20714 , n20735 );
not ( n20737 , n20582 );
not ( n20738 , n19753 );
buf ( n20739 , n20110 );
and ( n20740 , n20738 , n20739 );
xor ( n20741 , n20112 , n20435 );
buf ( n20742 , n20741 );
and ( n20743 , n20742 , n19753 );
or ( n20744 , n20740 , n20743 );
buf ( n20745 , n20744 );
buf ( n20746 , n20745 );
and ( n20747 , n20737 , n20746 );
not ( n20748 , n20746 );
and ( n20749 , n20726 , n20727 );
xor ( n20750 , n20748 , n20749 );
and ( n20751 , n20750 , n20582 );
or ( n20752 , n20747 , n20751 );
buf ( n20753 , n20752 );
not ( n20754 , n20753 );
buf ( n20755 , n20754 );
buf ( n20756 , n20755 );
not ( n20757 , n20756 );
or ( n20758 , n20736 , n20757 );
not ( n20759 , n20582 );
not ( n20760 , n19753 );
buf ( n20761 , n20075 );
and ( n20762 , n20760 , n20761 );
xor ( n20763 , n20077 , n20436 );
buf ( n20764 , n20763 );
and ( n20765 , n20764 , n19753 );
or ( n20766 , n20762 , n20765 );
buf ( n20767 , n20766 );
buf ( n20768 , n20767 );
and ( n20769 , n20759 , n20768 );
not ( n20770 , n20768 );
and ( n20771 , n20748 , n20749 );
xor ( n20772 , n20770 , n20771 );
and ( n20773 , n20772 , n20582 );
or ( n20774 , n20769 , n20773 );
buf ( n20775 , n20774 );
not ( n20776 , n20775 );
buf ( n20777 , n20776 );
buf ( n20778 , n20777 );
not ( n20779 , n20778 );
or ( n20780 , n20758 , n20779 );
not ( n20781 , n20582 );
not ( n20782 , n19753 );
buf ( n20783 , n20041 );
and ( n20784 , n20782 , n20783 );
xor ( n20785 , n20043 , n20437 );
buf ( n20786 , n20785 );
and ( n20787 , n20786 , n19753 );
or ( n20788 , n20784 , n20787 );
buf ( n20789 , n20788 );
buf ( n20790 , n20789 );
and ( n20791 , n20781 , n20790 );
not ( n20792 , n20790 );
and ( n20793 , n20770 , n20771 );
xor ( n20794 , n20792 , n20793 );
and ( n20795 , n20794 , n20582 );
or ( n20796 , n20791 , n20795 );
buf ( n20797 , n20796 );
not ( n20798 , n20797 );
buf ( n20799 , n20798 );
buf ( n20800 , n20799 );
not ( n20801 , n20800 );
or ( n20802 , n20780 , n20801 );
not ( n20803 , n20582 );
not ( n20804 , n19753 );
buf ( n20805 , n20028 );
and ( n20806 , n20804 , n20805 );
xor ( n20807 , n20030 , n20438 );
buf ( n20808 , n20807 );
and ( n20809 , n20808 , n19753 );
or ( n20810 , n20806 , n20809 );
buf ( n20811 , n20810 );
buf ( n20812 , n20811 );
and ( n20813 , n20803 , n20812 );
not ( n20814 , n20812 );
and ( n20815 , n20792 , n20793 );
xor ( n20816 , n20814 , n20815 );
and ( n20817 , n20816 , n20582 );
or ( n20818 , n20813 , n20817 );
buf ( n20819 , n20818 );
not ( n20820 , n20819 );
buf ( n20821 , n20820 );
buf ( n20822 , n20821 );
not ( n20823 , n20822 );
or ( n20824 , n20802 , n20823 );
not ( n20825 , n20582 );
not ( n20826 , n19753 );
buf ( n20827 , n20015 );
and ( n20828 , n20826 , n20827 );
xor ( n20829 , n20017 , n20439 );
buf ( n20830 , n20829 );
and ( n20831 , n20830 , n19753 );
or ( n20832 , n20828 , n20831 );
buf ( n20833 , n20832 );
buf ( n20834 , n20833 );
and ( n20835 , n20825 , n20834 );
not ( n20836 , n20834 );
and ( n20837 , n20814 , n20815 );
xor ( n20838 , n20836 , n20837 );
and ( n20839 , n20838 , n20582 );
or ( n20840 , n20835 , n20839 );
buf ( n20841 , n20840 );
not ( n20842 , n20841 );
buf ( n20843 , n20842 );
buf ( n20844 , n20843 );
not ( n20845 , n20844 );
or ( n20846 , n20824 , n20845 );
not ( n20847 , n20582 );
not ( n20848 , n19753 );
buf ( n20849 , n20002 );
and ( n20850 , n20848 , n20849 );
xor ( n20851 , n20004 , n20440 );
buf ( n20852 , n20851 );
and ( n20853 , n20852 , n19753 );
or ( n20854 , n20850 , n20853 );
buf ( n20855 , n20854 );
buf ( n20856 , n20855 );
and ( n20857 , n20847 , n20856 );
not ( n20858 , n20856 );
and ( n20859 , n20836 , n20837 );
xor ( n20860 , n20858 , n20859 );
and ( n20861 , n20860 , n20582 );
or ( n20862 , n20857 , n20861 );
buf ( n20863 , n20862 );
not ( n20864 , n20863 );
buf ( n20865 , n20864 );
buf ( n20866 , n20865 );
not ( n20867 , n20866 );
or ( n20868 , n20846 , n20867 );
not ( n20869 , n20582 );
not ( n20870 , n19753 );
buf ( n20871 , n19989 );
and ( n20872 , n20870 , n20871 );
xor ( n20873 , n19991 , n20441 );
buf ( n20874 , n20873 );
and ( n20875 , n20874 , n19753 );
or ( n20876 , n20872 , n20875 );
not ( n20877 , n20876 );
buf ( n20878 , n20877 );
and ( n20879 , n20869 , n20878 );
not ( n20880 , n20878 );
or ( n20881 , n20858 , n20859 );
xor ( n20882 , n20880 , n20881 );
and ( n20883 , n20882 , n20582 );
or ( n20884 , n20879 , n20883 );
buf ( n20885 , n20884 );
not ( n20886 , n20885 );
buf ( n20887 , n20886 );
buf ( n20888 , n20887 );
not ( n20889 , n20888 );
or ( n20890 , n20868 , n20889 );
not ( n20891 , n20582 );
not ( n20892 , n19753 );
buf ( n20893 , n19976 );
and ( n20894 , n20892 , n20893 );
xor ( n20895 , n19978 , n20442 );
buf ( n20896 , n20895 );
and ( n20897 , n20896 , n19753 );
or ( n20898 , n20894 , n20897 );
buf ( n20899 , n20898 );
buf ( n20900 , n20899 );
and ( n20901 , n20891 , n20900 );
not ( n20902 , n20900 );
and ( n20903 , n20880 , n20881 );
xor ( n20904 , n20902 , n20903 );
and ( n20905 , n20904 , n20582 );
or ( n20906 , n20901 , n20905 );
buf ( n20907 , n20906 );
not ( n20908 , n20907 );
buf ( n20909 , n20908 );
buf ( n20910 , n20909 );
not ( n20911 , n20910 );
or ( n20912 , n20890 , n20911 );
not ( n20913 , n20582 );
not ( n20914 , n19753 );
buf ( n20915 , n19963 );
and ( n20916 , n20914 , n20915 );
xor ( n20917 , n19965 , n20443 );
buf ( n20918 , n20917 );
and ( n20919 , n20918 , n19753 );
or ( n20920 , n20916 , n20919 );
buf ( n20921 , n20920 );
buf ( n20922 , n20921 );
nand ( n20923 , n20913 , n20922 );
not ( n20924 , n20922 );
and ( n20925 , n20902 , n20903 );
xor ( n20926 , n20924 , n20925 );
and ( n20927 , n20926 , n20582 );
xor ( n20928 , n20923 , n20927 );
buf ( n20929 , n20928 );
not ( n20930 , n20929 );
buf ( n20931 , n20930 );
buf ( n20932 , n20931 );
not ( n20933 , n20932 );
or ( n20934 , n20912 , n20933 );
not ( n20935 , n20582 );
not ( n20936 , n19753 );
buf ( n20937 , n19950 );
and ( n20938 , n20936 , n20937 );
xor ( n20939 , n19952 , n20444 );
buf ( n20940 , n20939 );
and ( n20941 , n20940 , n19753 );
or ( n20942 , n20938 , n20941 );
buf ( n20943 , n20942 );
buf ( n20944 , n20943 );
and ( n20945 , n20935 , n20944 );
not ( n20946 , n20944 );
and ( n20947 , n20924 , n20925 );
xor ( n20948 , n20946 , n20947 );
and ( n20949 , n20948 , n20582 );
or ( n20950 , n20945 , n20949 );
buf ( n20951 , n20950 );
not ( n20952 , n20951 );
buf ( n20953 , n20952 );
buf ( n20954 , n20953 );
not ( n20955 , n20954 );
or ( n20956 , n20934 , n20955 );
not ( n20957 , n20582 );
not ( n20958 , n19753 );
buf ( n20959 , n19937 );
and ( n20960 , n20958 , n20959 );
xor ( n20961 , n19939 , n20445 );
buf ( n20962 , n20961 );
and ( n20963 , n20962 , n19753 );
or ( n20964 , n20960 , n20963 );
buf ( n20965 , n20964 );
buf ( n20966 , n20965 );
and ( n20967 , n20957 , n20966 );
not ( n20968 , n20966 );
and ( n20969 , n20946 , n20947 );
xor ( n20970 , n20968 , n20969 );
and ( n20971 , n20970 , n20582 );
or ( n20972 , n20967 , n20971 );
buf ( n20973 , n20972 );
not ( n20974 , n20973 );
buf ( n20975 , n20974 );
buf ( n20976 , n20975 );
not ( n20977 , n20976 );
or ( n20978 , n20956 , n20977 );
not ( n20979 , n20582 );
not ( n20980 , n19753 );
buf ( n20981 , n19924 );
and ( n20982 , n20980 , n20981 );
xor ( n20983 , n19926 , n20446 );
buf ( n20984 , n20983 );
and ( n20985 , n20984 , n19753 );
or ( n20986 , n20982 , n20985 );
buf ( n20987 , n20986 );
buf ( n20988 , n20987 );
and ( n20989 , n20979 , n20988 );
not ( n20990 , n20988 );
and ( n20991 , n20968 , n20969 );
xor ( n20992 , n20990 , n20991 );
and ( n20993 , n20992 , n20582 );
or ( n20994 , n20989 , n20993 );
buf ( n20995 , n20994 );
not ( n20996 , n20995 );
buf ( n20997 , n20996 );
buf ( n20998 , n20997 );
not ( n20999 , n20998 );
or ( n21000 , n20978 , n20999 );
not ( n21001 , n20582 );
not ( n21002 , n19753 );
buf ( n21003 , n19911 );
and ( n21004 , n21002 , n21003 );
xor ( n21005 , n19913 , n20447 );
buf ( n21006 , n21005 );
and ( n21007 , n21006 , n19753 );
or ( n21008 , n21004 , n21007 );
buf ( n21009 , n21008 );
buf ( n21010 , n21009 );
and ( n21011 , n21001 , n21010 );
not ( n21012 , n21010 );
and ( n21013 , n20990 , n20991 );
xor ( n21014 , n21012 , n21013 );
and ( n21015 , n21014 , n20582 );
or ( n21016 , n21011 , n21015 );
buf ( n21017 , n21016 );
not ( n21018 , n21017 );
buf ( n21019 , n21018 );
buf ( n21020 , n21019 );
not ( n21021 , n21020 );
or ( n21022 , n21000 , n21021 );
not ( n21023 , n20582 );
not ( n21024 , n19753 );
buf ( n21025 , n19898 );
and ( n21026 , n21024 , n21025 );
xor ( n21027 , n19900 , n20448 );
buf ( n21028 , n21027 );
and ( n21029 , n21028 , n19753 );
or ( n21030 , n21026 , n21029 );
buf ( n21031 , n21030 );
buf ( n21032 , n21031 );
and ( n21033 , n21023 , n21032 );
not ( n21034 , n21032 );
and ( n21035 , n21012 , n21013 );
xor ( n21036 , n21034 , n21035 );
and ( n21037 , n21036 , n20582 );
or ( n21038 , n21033 , n21037 );
buf ( n21039 , n21038 );
not ( n21040 , n21039 );
buf ( n21041 , n21040 );
buf ( n21042 , n21041 );
not ( n21043 , n21042 );
or ( n21044 , n21022 , n21043 );
not ( n21045 , n20582 );
not ( n21046 , n19753 );
buf ( n21047 , n19885 );
and ( n21048 , n21046 , n21047 );
xor ( n21049 , n19887 , n20449 );
buf ( n21050 , n21049 );
and ( n21051 , n21050 , n19753 );
or ( n21052 , n21048 , n21051 );
buf ( n21053 , n21052 );
buf ( n21054 , n21053 );
and ( n21055 , n21045 , n21054 );
not ( n21056 , n21054 );
and ( n21057 , n21034 , n21035 );
xor ( n21058 , n21056 , n21057 );
and ( n21059 , n21058 , n20582 );
or ( n21060 , n21055 , n21059 );
buf ( n21061 , n21060 );
not ( n21062 , n21061 );
buf ( n21063 , n21062 );
buf ( n21064 , n21063 );
not ( n21065 , n21064 );
or ( n21066 , n21044 , n21065 );
not ( n21067 , n20582 );
not ( n21068 , n19753 );
buf ( n21069 , n19872 );
and ( n21070 , n21068 , n21069 );
xor ( n21071 , n19874 , n20450 );
buf ( n21072 , n21071 );
and ( n21073 , n21072 , n19753 );
or ( n21074 , n21070 , n21073 );
buf ( n21075 , n21074 );
buf ( n21076 , n21075 );
and ( n21077 , n21067 , n21076 );
not ( n21078 , n21076 );
and ( n21079 , n21056 , n21057 );
xor ( n21080 , n21078 , n21079 );
and ( n21081 , n21080 , n20582 );
or ( n21082 , n21077 , n21081 );
buf ( n21083 , n21082 );
not ( n21084 , n21083 );
buf ( n21085 , n21084 );
buf ( n21086 , n21085 );
not ( n21087 , n21086 );
or ( n21088 , n21066 , n21087 );
not ( n21089 , n20582 );
not ( n21090 , n19753 );
buf ( n21091 , n19859 );
and ( n21092 , n21090 , n21091 );
xor ( n21093 , n19861 , n20451 );
buf ( n21094 , n21093 );
and ( n21095 , n21094 , n19753 );
or ( n21096 , n21092 , n21095 );
buf ( n21097 , n21096 );
buf ( n21098 , n21097 );
and ( n21099 , n21089 , n21098 );
not ( n21100 , n21098 );
and ( n21101 , n21078 , n21079 );
xor ( n21102 , n21100 , n21101 );
and ( n21103 , n21102 , n20582 );
or ( n21104 , n21099 , n21103 );
buf ( n21105 , n21104 );
not ( n21106 , n21105 );
buf ( n21107 , n21106 );
buf ( n21108 , n21107 );
not ( n21109 , n21108 );
or ( n21110 , n21088 , n21109 );
not ( n21111 , n20582 );
buf ( n21112 , n20457 );
and ( n21113 , n21111 , n21112 );
not ( n21114 , n21112 );
and ( n21115 , n21100 , n21101 );
xor ( n21116 , n21114 , n21115 );
and ( n21117 , n21116 , n20582 );
or ( n21118 , n21113 , n21117 );
buf ( n21119 , n21118 );
not ( n21120 , n21119 );
buf ( n21121 , n21120 );
buf ( n21122 , n21121 );
not ( n21123 , n21122 );
or ( n21124 , n21110 , n21123 );
not ( n21125 , n20582 );
not ( n21126 , n19753 );
buf ( n21127 , n20568 );
and ( n21128 , n21126 , n21127 );
xor ( n21129 , n20570 , n20571 );
buf ( n21130 , n21129 );
and ( n21131 , n21130 , n19753 );
or ( n21132 , n21128 , n21131 );
buf ( n21133 , n21132 );
buf ( n21134 , n21133 );
and ( n21135 , n21125 , n21134 );
not ( n21136 , n21134 );
and ( n21137 , n21114 , n21115 );
xor ( n21138 , n21136 , n21137 );
and ( n21139 , n21138 , n20582 );
or ( n21140 , n21135 , n21139 );
buf ( n21141 , n21140 );
not ( n21142 , n21141 );
buf ( n21143 , n21142 );
buf ( n21144 , n21143 );
not ( n21145 , n21144 );
or ( n21146 , n21124 , n21145 );
not ( n21147 , n20582 );
not ( n21148 , n19753 );
buf ( n21149 , n20555 );
and ( n21150 , n21148 , n21149 );
xor ( n21151 , n20557 , n20572 );
buf ( n21152 , n21151 );
and ( n21153 , n21152 , n19753 );
or ( n21154 , n21150 , n21153 );
buf ( n21155 , n21154 );
buf ( n21156 , n21155 );
and ( n21157 , n21147 , n21156 );
not ( n21158 , n21156 );
and ( n21159 , n21136 , n21137 );
xor ( n21160 , n21158 , n21159 );
and ( n21161 , n21160 , n20582 );
or ( n21162 , n21157 , n21161 );
buf ( n21163 , n21162 );
not ( n21164 , n21163 );
buf ( n21165 , n21164 );
buf ( n21166 , n21165 );
not ( n21167 , n21166 );
or ( n21168 , n21146 , n21167 );
not ( n21169 , n20582 );
not ( n21170 , n19753 );
buf ( n21171 , n20542 );
and ( n21172 , n21170 , n21171 );
xor ( n21173 , n20544 , n20573 );
buf ( n21174 , n21173 );
and ( n21175 , n21174 , n19753 );
or ( n21176 , n21172 , n21175 );
buf ( n21177 , n21176 );
buf ( n21178 , n21177 );
and ( n21179 , n21169 , n21178 );
not ( n21180 , n21178 );
and ( n21181 , n21158 , n21159 );
xor ( n21182 , n21180 , n21181 );
and ( n21183 , n21182 , n20582 );
or ( n21184 , n21179 , n21183 );
buf ( n21185 , n21184 );
not ( n21186 , n21185 );
buf ( n21187 , n21186 );
buf ( n21188 , n21187 );
not ( n21189 , n21188 );
or ( n21190 , n21168 , n21189 );
buf ( n21191 , n21190 );
buf ( n21192 , n21191 );
and ( n21193 , n21192 , n20582 );
not ( n21194 , n21193 );
and ( n21195 , n21194 , n21123 );
xor ( n21196 , n21123 , n20582 );
xor ( n21197 , n21109 , n20582 );
xor ( n21198 , n21087 , n20582 );
xor ( n21199 , n21065 , n20582 );
xor ( n21200 , n21043 , n20582 );
xor ( n21201 , n21021 , n20582 );
xor ( n21202 , n20999 , n20582 );
xor ( n21203 , n20977 , n20582 );
xor ( n21204 , n20955 , n20582 );
xor ( n21205 , n20933 , n20582 );
xor ( n21206 , n20911 , n20582 );
xor ( n21207 , n20889 , n20582 );
xor ( n21208 , n20867 , n20582 );
xor ( n21209 , n20845 , n20582 );
xor ( n21210 , n20823 , n20582 );
xor ( n21211 , n20801 , n20582 );
xor ( n21212 , n20779 , n20582 );
xor ( n21213 , n20757 , n20582 );
xor ( n21214 , n20735 , n20582 );
xor ( n21215 , n20713 , n20582 );
xor ( n21216 , n20691 , n20582 );
xor ( n21217 , n20669 , n20582 );
xor ( n21218 , n20647 , n20582 );
xor ( n21219 , n20625 , n20582 );
xor ( n21220 , n20603 , n20582 );
xor ( n21221 , n20465 , n20582 );
and ( n21222 , n21221 , n20582 );
and ( n21223 , n21220 , n21222 );
and ( n21224 , n21219 , n21223 );
and ( n21225 , n21218 , n21224 );
and ( n21226 , n21217 , n21225 );
and ( n21227 , n21216 , n21226 );
and ( n21228 , n21215 , n21227 );
and ( n21229 , n21214 , n21228 );
and ( n21230 , n21213 , n21229 );
and ( n21231 , n21212 , n21230 );
and ( n21232 , n21211 , n21231 );
and ( n21233 , n21210 , n21232 );
and ( n21234 , n21209 , n21233 );
and ( n21235 , n21208 , n21234 );
and ( n21236 , n21207 , n21235 );
and ( n21237 , n21206 , n21236 );
and ( n21238 , n21205 , n21237 );
and ( n21239 , n21204 , n21238 );
and ( n21240 , n21203 , n21239 );
and ( n21241 , n21202 , n21240 );
and ( n21242 , n21201 , n21241 );
and ( n21243 , n21200 , n21242 );
and ( n21244 , n21199 , n21243 );
and ( n21245 , n21198 , n21244 );
and ( n21246 , n21197 , n21245 );
xor ( n21247 , n21196 , n21246 );
and ( n21248 , n21247 , n21193 );
or ( n21249 , n21195 , n21248 );
buf ( n21250 , n21249 );
and ( n21251 , n21250 , n19750 );
or ( n21252 , n20458 , n21251 );
nor ( n21253 , n19747 , n19744 );
and ( n21254 , n21252 , n21253 );
nor ( n21255 , n19736 , n19744 );
and ( n21256 , n20457 , n21255 );
or ( n21257 , n19746 , n19749 , n21254 , n21256 );
not ( n21258 , n17433 );
not ( n21259 , n17449 );
nor ( n21260 , n21258 , n17441 , n21259 );
not ( n21261 , n21260 );
nor ( n21262 , n17433 , n17441 , n21259 );
not ( n21263 , n21262 );
and ( n21264 , n17433 , n17441 , n21259 );
not ( n21265 , n21264 );
and ( n21266 , n21258 , n17441 , n21259 );
not ( n21267 , n21266 );
nor ( n21268 , n21258 , n17441 , n17449 );
not ( n21269 , n21268 );
nor ( n21270 , n17433 , n17441 , n17449 );
not ( n21271 , n21270 );
buf ( n21272 , RI21a11650_88);
and ( n21273 , n21271 , n21272 );
or ( n21274 , n21273 , C0 );
and ( n21275 , n21269 , n21274 );
and ( n21276 , C1 , n21268 );
or ( n21277 , n21275 , n21276 );
and ( n21278 , n21267 , n21277 );
or ( n21279 , n21278 , C0 );
and ( n21280 , n21265 , n21279 );
and ( n21281 , C1 , n21264 );
or ( n21282 , n21280 , n21281 );
and ( n21283 , n21263 , n21282 );
not ( n21284 , n19750 );
and ( n21285 , n21284 , n21272 );
and ( n21286 , C1 , n19750 );
or ( n21287 , n21285 , n21286 );
and ( n21288 , n21287 , n21262 );
or ( n21289 , n21283 , n21288 );
and ( n21290 , n21261 , n21289 );
not ( n21291 , n19750 );
not ( n21292 , n21291 );
and ( n21293 , n21292 , n21272 );
and ( n21294 , C1 , n21291 );
or ( n21295 , n21293 , n21294 );
and ( n21296 , n21295 , n21260 );
or ( n21297 , n21290 , n21296 );
not ( n21298 , n21260 );
not ( n21299 , n21262 );
not ( n21300 , n21264 );
not ( n21301 , n21266 );
not ( n21302 , n21268 );
not ( n21303 , n21270 );
buf ( n21304 , RI21a115d8_89);
and ( n21305 , n21303 , n21304 );
or ( n21306 , n21305 , C0 );
and ( n21307 , n21302 , n21306 );
or ( n21308 , n21307 , C0 );
and ( n21309 , n21301 , n21308 );
and ( n21310 , C1 , n21266 );
or ( n21311 , n21309 , n21310 );
and ( n21312 , n21300 , n21311 );
and ( n21313 , C1 , n21264 );
or ( n21314 , n21312 , n21313 );
and ( n21315 , n21299 , n21314 );
not ( n21316 , n19750 );
and ( n21317 , n21316 , n21304 );
and ( n21318 , C1 , n19750 );
or ( n21319 , n21317 , n21318 );
and ( n21320 , n21319 , n21262 );
or ( n21321 , n21315 , n21320 );
and ( n21322 , n21298 , n21321 );
not ( n21323 , n21291 );
and ( n21324 , n21323 , n21304 );
and ( n21325 , C1 , n21291 );
or ( n21326 , n21324 , n21325 );
and ( n21327 , n21326 , n21260 );
or ( n21328 , n21322 , n21327 );
not ( n21329 , n21328 );
nor ( n21330 , n21297 , n21329 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n21331 , n21257 , n21330 );
not ( n21332 , n21297 );
nor ( n21333 , n21332 , n21328 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
nor ( n21334 , n21297 , n21328 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
or ( n21335 , n21333 , n21334 );
nor ( n21336 , n21332 , n21329 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
or ( n21337 , n21335 , n21336 );
or ( n21338 , n21337 , C0 );
and ( n21339 , n17453 , n21338 );
or ( n21340 , n21331 , n21339 );
and ( n21341 , n17869 , n17851 , n17859 , n17867 );
and ( n21342 , n21340 , n21341 );
buf ( n21343 , n18514 );
not ( n21344 , n14641 );
and ( n21345 , n21344 , n14833 );
buf ( n21346 , n14833 );
buf ( n21347 , n15852 );
xor ( n21348 , n21346 , n21347 );
buf ( n21349 , n21348 );
and ( n21350 , n21349 , n14641 );
or ( n21351 , n21345 , n21350 );
or ( n21352 , n21253 , n19748 );
or ( n21353 , n21352 , n19745 );
and ( n21354 , n21351 , n21353 );
buf ( n21355 , n16900 );
buf ( n21356 , n21355 );
not ( n21357 , n21356 );
buf ( n21358 , n21357 );
buf ( n21359 , n21358 );
not ( n21360 , n21359 );
buf ( n21361 , n16712 );
not ( n21362 , n21361 );
buf ( n21363 , n16897 );
and ( n21364 , n21362 , n21363 );
not ( n21365 , n21363 );
not ( n21366 , n21355 );
xor ( n21367 , n21365 , n21366 );
and ( n21368 , n21367 , n21361 );
or ( n21369 , n21364 , n21368 );
buf ( n21370 , n21369 );
not ( n21371 , n21370 );
buf ( n21372 , n21371 );
buf ( n21373 , n21372 );
not ( n21374 , n21373 );
or ( n21375 , n21360 , n21374 );
not ( n21376 , n21361 );
buf ( n21377 , n16889 );
and ( n21378 , n21376 , n21377 );
not ( n21379 , n21377 );
and ( n21380 , n21365 , n21366 );
xor ( n21381 , n21379 , n21380 );
and ( n21382 , n21381 , n21361 );
or ( n21383 , n21378 , n21382 );
buf ( n21384 , n21383 );
not ( n21385 , n21384 );
buf ( n21386 , n21385 );
buf ( n21387 , n21386 );
not ( n21388 , n21387 );
or ( n21389 , n21375 , n21388 );
not ( n21390 , n21361 );
buf ( n21391 , n16881 );
and ( n21392 , n21390 , n21391 );
not ( n21393 , n21391 );
and ( n21394 , n21379 , n21380 );
xor ( n21395 , n21393 , n21394 );
and ( n21396 , n21395 , n21361 );
or ( n21397 , n21392 , n21396 );
buf ( n21398 , n21397 );
not ( n21399 , n21398 );
buf ( n21400 , n21399 );
buf ( n21401 , n21400 );
not ( n21402 , n21401 );
or ( n21403 , n21389 , n21402 );
not ( n21404 , n21361 );
buf ( n21405 , n16873 );
and ( n21406 , n21404 , n21405 );
not ( n21407 , n21405 );
and ( n21408 , n21393 , n21394 );
xor ( n21409 , n21407 , n21408 );
and ( n21410 , n21409 , n21361 );
or ( n21411 , n21406 , n21410 );
buf ( n21412 , n21411 );
not ( n21413 , n21412 );
buf ( n21414 , n21413 );
buf ( n21415 , n21414 );
not ( n21416 , n21415 );
or ( n21417 , n21403 , n21416 );
not ( n21418 , n21361 );
buf ( n21419 , n16865 );
and ( n21420 , n21418 , n21419 );
not ( n21421 , n21419 );
and ( n21422 , n21407 , n21408 );
xor ( n21423 , n21421 , n21422 );
and ( n21424 , n21423 , n21361 );
or ( n21425 , n21420 , n21424 );
buf ( n21426 , n21425 );
not ( n21427 , n21426 );
buf ( n21428 , n21427 );
buf ( n21429 , n21428 );
not ( n21430 , n21429 );
or ( n21431 , n21417 , n21430 );
not ( n21432 , n21361 );
buf ( n21433 , n16857 );
and ( n21434 , n21432 , n21433 );
not ( n21435 , n21433 );
and ( n21436 , n21421 , n21422 );
xor ( n21437 , n21435 , n21436 );
and ( n21438 , n21437 , n21361 );
or ( n21439 , n21434 , n21438 );
buf ( n21440 , n21439 );
not ( n21441 , n21440 );
buf ( n21442 , n21441 );
buf ( n21443 , n21442 );
not ( n21444 , n21443 );
or ( n21445 , n21431 , n21444 );
not ( n21446 , n21361 );
buf ( n21447 , n16849 );
and ( n21448 , n21446 , n21447 );
not ( n21449 , n21447 );
and ( n21450 , n21435 , n21436 );
xor ( n21451 , n21449 , n21450 );
and ( n21452 , n21451 , n21361 );
or ( n21453 , n21448 , n21452 );
buf ( n21454 , n21453 );
not ( n21455 , n21454 );
buf ( n21456 , n21455 );
buf ( n21457 , n21456 );
not ( n21458 , n21457 );
or ( n21459 , n21445 , n21458 );
not ( n21460 , n21361 );
buf ( n21461 , n16841 );
and ( n21462 , n21460 , n21461 );
not ( n21463 , n21461 );
and ( n21464 , n21449 , n21450 );
xor ( n21465 , n21463 , n21464 );
and ( n21466 , n21465 , n21361 );
or ( n21467 , n21462 , n21466 );
buf ( n21468 , n21467 );
not ( n21469 , n21468 );
buf ( n21470 , n21469 );
buf ( n21471 , n21470 );
not ( n21472 , n21471 );
or ( n21473 , n21459 , n21472 );
not ( n21474 , n21361 );
buf ( n21475 , n16833 );
and ( n21476 , n21474 , n21475 );
not ( n21477 , n21475 );
and ( n21478 , n21463 , n21464 );
xor ( n21479 , n21477 , n21478 );
and ( n21480 , n21479 , n21361 );
or ( n21481 , n21476 , n21480 );
buf ( n21482 , n21481 );
not ( n21483 , n21482 );
buf ( n21484 , n21483 );
buf ( n21485 , n21484 );
not ( n21486 , n21485 );
or ( n21487 , n21473 , n21486 );
not ( n21488 , n21361 );
buf ( n21489 , n16825 );
and ( n21490 , n21488 , n21489 );
not ( n21491 , n21489 );
and ( n21492 , n21477 , n21478 );
xor ( n21493 , n21491 , n21492 );
and ( n21494 , n21493 , n21361 );
or ( n21495 , n21490 , n21494 );
buf ( n21496 , n21495 );
not ( n21497 , n21496 );
buf ( n21498 , n21497 );
buf ( n21499 , n21498 );
not ( n21500 , n21499 );
or ( n21501 , n21487 , n21500 );
not ( n21502 , n21361 );
buf ( n21503 , n16817 );
and ( n21504 , n21502 , n21503 );
not ( n21505 , n21503 );
and ( n21506 , n21491 , n21492 );
xor ( n21507 , n21505 , n21506 );
and ( n21508 , n21507 , n21361 );
or ( n21509 , n21504 , n21508 );
buf ( n21510 , n21509 );
not ( n21511 , n21510 );
buf ( n21512 , n21511 );
buf ( n21513 , n21512 );
not ( n21514 , n21513 );
or ( n21515 , n21501 , n21514 );
not ( n21516 , n21361 );
buf ( n21517 , n16809 );
and ( n21518 , n21516 , n21517 );
not ( n21519 , n21517 );
and ( n21520 , n21505 , n21506 );
xor ( n21521 , n21519 , n21520 );
and ( n21522 , n21521 , n21361 );
or ( n21523 , n21518 , n21522 );
buf ( n21524 , n21523 );
not ( n21525 , n21524 );
buf ( n21526 , n21525 );
buf ( n21527 , n21526 );
not ( n21528 , n21527 );
or ( n21529 , n21515 , n21528 );
not ( n21530 , n21361 );
buf ( n21531 , n16801 );
and ( n21532 , n21530 , n21531 );
not ( n21533 , n21531 );
and ( n21534 , n21519 , n21520 );
xor ( n21535 , n21533 , n21534 );
and ( n21536 , n21535 , n21361 );
or ( n21537 , n21532 , n21536 );
buf ( n21538 , n21537 );
not ( n21539 , n21538 );
buf ( n21540 , n21539 );
buf ( n21541 , n21540 );
not ( n21542 , n21541 );
or ( n21543 , n21529 , n21542 );
not ( n21544 , n21361 );
buf ( n21545 , n16793 );
and ( n21546 , n21544 , n21545 );
not ( n21547 , n21545 );
and ( n21548 , n21533 , n21534 );
xor ( n21549 , n21547 , n21548 );
and ( n21550 , n21549 , n21361 );
or ( n21551 , n21546 , n21550 );
buf ( n21552 , n21551 );
not ( n21553 , n21552 );
buf ( n21554 , n21553 );
buf ( n21555 , n21554 );
not ( n21556 , n21555 );
or ( n21557 , n21543 , n21556 );
not ( n21558 , n21361 );
buf ( n21559 , n16785 );
and ( n21560 , n21558 , n21559 );
not ( n21561 , n21559 );
and ( n21562 , n21547 , n21548 );
xor ( n21563 , n21561 , n21562 );
and ( n21564 , n21563 , n21361 );
or ( n21565 , n21560 , n21564 );
buf ( n21566 , n21565 );
not ( n21567 , n21566 );
buf ( n21568 , n21567 );
buf ( n21569 , n21568 );
not ( n21570 , n21569 );
or ( n21571 , n21557 , n21570 );
not ( n21572 , n21361 );
buf ( n21573 , n16777 );
and ( n21574 , n21572 , n21573 );
not ( n21575 , n21573 );
and ( n21576 , n21561 , n21562 );
xor ( n21577 , n21575 , n21576 );
and ( n21578 , n21577 , n21361 );
or ( n21579 , n21574 , n21578 );
buf ( n21580 , n21579 );
not ( n21581 , n21580 );
buf ( n21582 , n21581 );
buf ( n21583 , n21582 );
not ( n21584 , n21583 );
or ( n21585 , n21571 , n21584 );
not ( n21586 , n21361 );
buf ( n21587 , n16769 );
and ( n21588 , n21586 , n21587 );
not ( n21589 , n21587 );
and ( n21590 , n21575 , n21576 );
xor ( n21591 , n21589 , n21590 );
and ( n21592 , n21591 , n21361 );
or ( n21593 , n21588 , n21592 );
buf ( n21594 , n21593 );
not ( n21595 , n21594 );
buf ( n21596 , n21595 );
buf ( n21597 , n21596 );
not ( n21598 , n21597 );
or ( n21599 , n21585 , n21598 );
not ( n21600 , n21361 );
buf ( n21601 , n16761 );
and ( n21602 , n21600 , n21601 );
not ( n21603 , n21601 );
and ( n21604 , n21589 , n21590 );
xor ( n21605 , n21603 , n21604 );
and ( n21606 , n21605 , n21361 );
or ( n21607 , n21602 , n21606 );
buf ( n21608 , n21607 );
not ( n21609 , n21608 );
buf ( n21610 , n21609 );
buf ( n21611 , n21610 );
not ( n21612 , n21611 );
or ( n21613 , n21599 , n21612 );
not ( n21614 , n21361 );
buf ( n21615 , n16753 );
and ( n21616 , n21614 , n21615 );
not ( n21617 , n21615 );
and ( n21618 , n21603 , n21604 );
xor ( n21619 , n21617 , n21618 );
and ( n21620 , n21619 , n21361 );
or ( n21621 , n21616 , n21620 );
buf ( n21622 , n21621 );
not ( n21623 , n21622 );
buf ( n21624 , n21623 );
buf ( n21625 , n21624 );
not ( n21626 , n21625 );
or ( n21627 , n21613 , n21626 );
buf ( n21628 , n21627 );
buf ( n21629 , n21628 );
and ( n21630 , n21629 , n21361 );
not ( n21631 , n21630 );
and ( n21632 , n21631 , n21360 );
xor ( n21633 , n21360 , n21361 );
xor ( n21634 , n21633 , n21361 );
and ( n21635 , n21634 , n21630 );
or ( n21636 , n21632 , n21635 );
buf ( n21637 , n21636 );
and ( n21638 , n21637 , n21255 );
or ( n21639 , n21354 , n21638 );
buf ( n21640 , n21639 );
xor ( n21641 , n21343 , n21640 );
buf ( n21642 , n21641 );
buf ( n21643 , n21642 );
buf ( n21644 , n21643 );
not ( n21645 , n21644 );
buf ( n21646 , n21645 );
buf ( n21647 , n21646 );
not ( n21648 , n21647 );
buf ( n21649 , n18527 );
not ( n21650 , n14641 );
and ( n21651 , n21650 , n14647 );
buf ( n21652 , n14647 );
buf ( n21653 , n14643 );
xor ( n21654 , n21652 , n21653 );
buf ( n21655 , n14653 );
buf ( n21656 , n14944 );
and ( n21657 , n21655 , n21656 );
buf ( n21658 , n14659 );
buf ( n21659 , n14969 );
and ( n21660 , n21658 , n21659 );
buf ( n21661 , n14665 );
buf ( n21662 , n14984 );
and ( n21663 , n21661 , n21662 );
buf ( n21664 , n14671 );
buf ( n21665 , n14999 );
and ( n21666 , n21664 , n21665 );
buf ( n21667 , n14677 );
buf ( n21668 , n15014 );
and ( n21669 , n21667 , n21668 );
buf ( n21670 , n14683 );
buf ( n21671 , n15029 );
and ( n21672 , n21670 , n21671 );
buf ( n21673 , n14689 );
buf ( n21674 , n15044 );
and ( n21675 , n21673 , n21674 );
buf ( n21676 , n14695 );
buf ( n21677 , n15059 );
and ( n21678 , n21676 , n21677 );
buf ( n21679 , n14701 );
buf ( n21680 , n15074 );
and ( n21681 , n21679 , n21680 );
buf ( n21682 , n14707 );
buf ( n21683 , n15089 );
and ( n21684 , n21682 , n21683 );
buf ( n21685 , n14713 );
buf ( n21686 , n15104 );
and ( n21687 , n21685 , n21686 );
buf ( n21688 , n14719 );
buf ( n21689 , n15119 );
and ( n21690 , n21688 , n21689 );
buf ( n21691 , n14725 );
buf ( n21692 , n15456 );
and ( n21693 , n21691 , n21692 );
buf ( n21694 , n14731 );
buf ( n21695 , n15478 );
and ( n21696 , n21694 , n21695 );
buf ( n21697 , n14737 );
buf ( n21698 , n15500 );
and ( n21699 , n21697 , n21698 );
buf ( n21700 , n14743 );
buf ( n21701 , n15522 );
and ( n21702 , n21700 , n21701 );
buf ( n21703 , n14749 );
buf ( n21704 , n15544 );
and ( n21705 , n21703 , n21704 );
buf ( n21706 , n14755 );
buf ( n21707 , n15566 );
and ( n21708 , n21706 , n21707 );
buf ( n21709 , n14761 );
buf ( n21710 , n15588 );
and ( n21711 , n21709 , n21710 );
buf ( n21712 , n14767 );
buf ( n21713 , n15610 );
and ( n21714 , n21712 , n21713 );
buf ( n21715 , n14773 );
buf ( n21716 , n15632 );
and ( n21717 , n21715 , n21716 );
buf ( n21718 , n14779 );
buf ( n21719 , n15654 );
and ( n21720 , n21718 , n21719 );
buf ( n21721 , n14785 );
buf ( n21722 , n15676 );
and ( n21723 , n21721 , n21722 );
buf ( n21724 , n14791 );
buf ( n21725 , n15698 );
and ( n21726 , n21724 , n21725 );
buf ( n21727 , n14797 );
buf ( n21728 , n15720 );
and ( n21729 , n21727 , n21728 );
buf ( n21730 , n14803 );
buf ( n21731 , n15742 );
and ( n21732 , n21730 , n21731 );
buf ( n21733 , n14809 );
buf ( n21734 , n15764 );
and ( n21735 , n21733 , n21734 );
buf ( n21736 , n14815 );
buf ( n21737 , n15786 );
and ( n21738 , n21736 , n21737 );
buf ( n21739 , n14821 );
buf ( n21740 , n15808 );
and ( n21741 , n21739 , n21740 );
buf ( n21742 , n14827 );
buf ( n21743 , n15830 );
and ( n21744 , n21742 , n21743 );
and ( n21745 , n21346 , n21347 );
and ( n21746 , n21743 , n21745 );
and ( n21747 , n21742 , n21745 );
or ( n21748 , n21744 , n21746 , n21747 );
and ( n21749 , n21740 , n21748 );
and ( n21750 , n21739 , n21748 );
or ( n21751 , n21741 , n21749 , n21750 );
and ( n21752 , n21737 , n21751 );
and ( n21753 , n21736 , n21751 );
or ( n21754 , n21738 , n21752 , n21753 );
and ( n21755 , n21734 , n21754 );
and ( n21756 , n21733 , n21754 );
or ( n21757 , n21735 , n21755 , n21756 );
and ( n21758 , n21731 , n21757 );
and ( n21759 , n21730 , n21757 );
or ( n21760 , n21732 , n21758 , n21759 );
and ( n21761 , n21728 , n21760 );
and ( n21762 , n21727 , n21760 );
or ( n21763 , n21729 , n21761 , n21762 );
and ( n21764 , n21725 , n21763 );
and ( n21765 , n21724 , n21763 );
or ( n21766 , n21726 , n21764 , n21765 );
and ( n21767 , n21722 , n21766 );
and ( n21768 , n21721 , n21766 );
or ( n21769 , n21723 , n21767 , n21768 );
and ( n21770 , n21719 , n21769 );
and ( n21771 , n21718 , n21769 );
or ( n21772 , n21720 , n21770 , n21771 );
and ( n21773 , n21716 , n21772 );
and ( n21774 , n21715 , n21772 );
or ( n21775 , n21717 , n21773 , n21774 );
and ( n21776 , n21713 , n21775 );
and ( n21777 , n21712 , n21775 );
or ( n21778 , n21714 , n21776 , n21777 );
and ( n21779 , n21710 , n21778 );
and ( n21780 , n21709 , n21778 );
or ( n21781 , n21711 , n21779 , n21780 );
and ( n21782 , n21707 , n21781 );
and ( n21783 , n21706 , n21781 );
or ( n21784 , n21708 , n21782 , n21783 );
and ( n21785 , n21704 , n21784 );
and ( n21786 , n21703 , n21784 );
or ( n21787 , n21705 , n21785 , n21786 );
and ( n21788 , n21701 , n21787 );
and ( n21789 , n21700 , n21787 );
or ( n21790 , n21702 , n21788 , n21789 );
and ( n21791 , n21698 , n21790 );
and ( n21792 , n21697 , n21790 );
or ( n21793 , n21699 , n21791 , n21792 );
and ( n21794 , n21695 , n21793 );
and ( n21795 , n21694 , n21793 );
or ( n21796 , n21696 , n21794 , n21795 );
and ( n21797 , n21692 , n21796 );
and ( n21798 , n21691 , n21796 );
or ( n21799 , n21693 , n21797 , n21798 );
and ( n21800 , n21689 , n21799 );
and ( n21801 , n21688 , n21799 );
or ( n21802 , n21690 , n21800 , n21801 );
and ( n21803 , n21686 , n21802 );
and ( n21804 , n21685 , n21802 );
or ( n21805 , n21687 , n21803 , n21804 );
and ( n21806 , n21683 , n21805 );
and ( n21807 , n21682 , n21805 );
or ( n21808 , n21684 , n21806 , n21807 );
and ( n21809 , n21680 , n21808 );
and ( n21810 , n21679 , n21808 );
or ( n21811 , n21681 , n21809 , n21810 );
and ( n21812 , n21677 , n21811 );
and ( n21813 , n21676 , n21811 );
or ( n21814 , n21678 , n21812 , n21813 );
and ( n21815 , n21674 , n21814 );
and ( n21816 , n21673 , n21814 );
or ( n21817 , n21675 , n21815 , n21816 );
and ( n21818 , n21671 , n21817 );
and ( n21819 , n21670 , n21817 );
or ( n21820 , n21672 , n21818 , n21819 );
and ( n21821 , n21668 , n21820 );
and ( n21822 , n21667 , n21820 );
or ( n21823 , n21669 , n21821 , n21822 );
and ( n21824 , n21665 , n21823 );
and ( n21825 , n21664 , n21823 );
or ( n21826 , n21666 , n21824 , n21825 );
and ( n21827 , n21662 , n21826 );
and ( n21828 , n21661 , n21826 );
or ( n21829 , n21663 , n21827 , n21828 );
and ( n21830 , n21659 , n21829 );
and ( n21831 , n21658 , n21829 );
or ( n21832 , n21660 , n21830 , n21831 );
and ( n21833 , n21656 , n21832 );
and ( n21834 , n21655 , n21832 );
or ( n21835 , n21657 , n21833 , n21834 );
xor ( n21836 , n21654 , n21835 );
buf ( n21837 , n21836 );
and ( n21838 , n21837 , n14641 );
or ( n21839 , n21651 , n21838 );
and ( n21840 , n21839 , n21353 );
buf ( n21841 , n21840 );
buf ( n21842 , n21841 );
not ( n21843 , n21842 );
xor ( n21844 , n21649 , n21843 );
buf ( n21845 , n20484 );
not ( n21846 , n14641 );
and ( n21847 , n21846 , n14653 );
xor ( n21848 , n21655 , n21656 );
xor ( n21849 , n21848 , n21832 );
buf ( n21850 , n21849 );
and ( n21851 , n21850 , n14641 );
or ( n21852 , n21847 , n21851 );
and ( n21853 , n21852 , n21353 );
buf ( n21854 , n21853 );
buf ( n21855 , n21854 );
not ( n21856 , n21855 );
and ( n21857 , n21845 , n21856 );
buf ( n21858 , n20496 );
not ( n21859 , n14641 );
and ( n21860 , n21859 , n14659 );
xor ( n21861 , n21658 , n21659 );
xor ( n21862 , n21861 , n21829 );
buf ( n21863 , n21862 );
and ( n21864 , n21863 , n14641 );
or ( n21865 , n21860 , n21864 );
and ( n21866 , n21865 , n21353 );
buf ( n21867 , n21866 );
buf ( n21868 , n21867 );
not ( n21869 , n21868 );
and ( n21870 , n21858 , n21869 );
buf ( n21871 , n19458 );
not ( n21872 , n14641 );
and ( n21873 , n21872 , n14665 );
xor ( n21874 , n21661 , n21662 );
xor ( n21875 , n21874 , n21826 );
buf ( n21876 , n21875 );
and ( n21877 , n21876 , n14641 );
or ( n21878 , n21873 , n21877 );
and ( n21879 , n21878 , n21353 );
buf ( n21880 , n21879 );
buf ( n21881 , n21880 );
not ( n21882 , n21881 );
and ( n21883 , n21871 , n21882 );
buf ( n21884 , n19424 );
not ( n21885 , n14641 );
and ( n21886 , n21885 , n14671 );
xor ( n21887 , n21664 , n21665 );
xor ( n21888 , n21887 , n21823 );
buf ( n21889 , n21888 );
and ( n21890 , n21889 , n14641 );
or ( n21891 , n21886 , n21890 );
and ( n21892 , n21891 , n21353 );
buf ( n21893 , n21892 );
buf ( n21894 , n21893 );
not ( n21895 , n21894 );
and ( n21896 , n21884 , n21895 );
buf ( n21897 , n19390 );
not ( n21898 , n14641 );
and ( n21899 , n21898 , n14677 );
xor ( n21900 , n21667 , n21668 );
xor ( n21901 , n21900 , n21820 );
buf ( n21902 , n21901 );
and ( n21903 , n21902 , n14641 );
or ( n21904 , n21899 , n21903 );
and ( n21905 , n21904 , n21353 );
buf ( n21906 , n21905 );
buf ( n21907 , n21906 );
not ( n21908 , n21907 );
and ( n21909 , n21897 , n21908 );
buf ( n21910 , n19356 );
not ( n21911 , n14641 );
and ( n21912 , n21911 , n14683 );
xor ( n21913 , n21670 , n21671 );
xor ( n21914 , n21913 , n21817 );
buf ( n21915 , n21914 );
and ( n21916 , n21915 , n14641 );
or ( n21917 , n21912 , n21916 );
and ( n21918 , n21917 , n21353 );
buf ( n21919 , n21918 );
buf ( n21920 , n21919 );
not ( n21921 , n21920 );
and ( n21922 , n21910 , n21921 );
buf ( n21923 , n19323 );
not ( n21924 , n14641 );
and ( n21925 , n21924 , n14689 );
xor ( n21926 , n21673 , n21674 );
xor ( n21927 , n21926 , n21814 );
buf ( n21928 , n21927 );
and ( n21929 , n21928 , n14641 );
or ( n21930 , n21925 , n21929 );
and ( n21931 , n21930 , n21353 );
buf ( n21932 , n21931 );
buf ( n21933 , n21932 );
not ( n21934 , n21933 );
and ( n21935 , n21923 , n21934 );
buf ( n21936 , n19289 );
not ( n21937 , n14641 );
and ( n21938 , n21937 , n14695 );
xor ( n21939 , n21676 , n21677 );
xor ( n21940 , n21939 , n21811 );
buf ( n21941 , n21940 );
and ( n21942 , n21941 , n14641 );
or ( n21943 , n21938 , n21942 );
and ( n21944 , n21943 , n21353 );
buf ( n21945 , n21944 );
buf ( n21946 , n21945 );
not ( n21947 , n21946 );
and ( n21948 , n21936 , n21947 );
buf ( n21949 , n19255 );
not ( n21950 , n14641 );
and ( n21951 , n21950 , n14701 );
xor ( n21952 , n21679 , n21680 );
xor ( n21953 , n21952 , n21808 );
buf ( n21954 , n21953 );
and ( n21955 , n21954 , n14641 );
or ( n21956 , n21951 , n21955 );
and ( n21957 , n21956 , n21353 );
buf ( n21958 , n21957 );
buf ( n21959 , n21958 );
not ( n21960 , n21959 );
and ( n21961 , n21949 , n21960 );
buf ( n21962 , n19221 );
not ( n21963 , n14641 );
and ( n21964 , n21963 , n14707 );
xor ( n21965 , n21682 , n21683 );
xor ( n21966 , n21965 , n21805 );
buf ( n21967 , n21966 );
and ( n21968 , n21967 , n14641 );
or ( n21969 , n21964 , n21968 );
and ( n21970 , n21969 , n21353 );
buf ( n21971 , n21970 );
buf ( n21972 , n21971 );
not ( n21973 , n21972 );
and ( n21974 , n21962 , n21973 );
buf ( n21975 , n19187 );
not ( n21976 , n14641 );
and ( n21977 , n21976 , n14713 );
xor ( n21978 , n21685 , n21686 );
xor ( n21979 , n21978 , n21802 );
buf ( n21980 , n21979 );
and ( n21981 , n21980 , n14641 );
or ( n21982 , n21977 , n21981 );
and ( n21983 , n21982 , n21353 );
buf ( n21984 , n21983 );
buf ( n21985 , n21984 );
not ( n21986 , n21985 );
and ( n21987 , n21975 , n21986 );
buf ( n21988 , n19153 );
not ( n21989 , n14641 );
and ( n21990 , n21989 , n14719 );
xor ( n21991 , n21688 , n21689 );
xor ( n21992 , n21991 , n21799 );
buf ( n21993 , n21992 );
and ( n21994 , n21993 , n14641 );
or ( n21995 , n21990 , n21994 );
and ( n21996 , n21995 , n21353 );
not ( n21997 , n21630 );
and ( n21998 , n21997 , n21626 );
xor ( n21999 , n21626 , n21361 );
xor ( n22000 , n21612 , n21361 );
xor ( n22001 , n21598 , n21361 );
xor ( n22002 , n21584 , n21361 );
xor ( n22003 , n21570 , n21361 );
xor ( n22004 , n21556 , n21361 );
xor ( n22005 , n21542 , n21361 );
xor ( n22006 , n21528 , n21361 );
xor ( n22007 , n21514 , n21361 );
xor ( n22008 , n21500 , n21361 );
xor ( n22009 , n21486 , n21361 );
xor ( n22010 , n21472 , n21361 );
xor ( n22011 , n21458 , n21361 );
xor ( n22012 , n21444 , n21361 );
xor ( n22013 , n21430 , n21361 );
xor ( n22014 , n21416 , n21361 );
xor ( n22015 , n21402 , n21361 );
xor ( n22016 , n21388 , n21361 );
xor ( n22017 , n21374 , n21361 );
and ( n22018 , n21633 , n21361 );
and ( n22019 , n22017 , n22018 );
and ( n22020 , n22016 , n22019 );
and ( n22021 , n22015 , n22020 );
and ( n22022 , n22014 , n22021 );
and ( n22023 , n22013 , n22022 );
and ( n22024 , n22012 , n22023 );
and ( n22025 , n22011 , n22024 );
and ( n22026 , n22010 , n22025 );
and ( n22027 , n22009 , n22026 );
and ( n22028 , n22008 , n22027 );
and ( n22029 , n22007 , n22028 );
and ( n22030 , n22006 , n22029 );
and ( n22031 , n22005 , n22030 );
and ( n22032 , n22004 , n22031 );
and ( n22033 , n22003 , n22032 );
and ( n22034 , n22002 , n22033 );
and ( n22035 , n22001 , n22034 );
and ( n22036 , n22000 , n22035 );
xor ( n22037 , n21999 , n22036 );
and ( n22038 , n22037 , n21630 );
or ( n22039 , n21998 , n22038 );
buf ( n22040 , n22039 );
and ( n22041 , n22040 , n21255 );
or ( n22042 , n21996 , n22041 );
buf ( n22043 , n22042 );
not ( n22044 , n22043 );
and ( n22045 , n21988 , n22044 );
buf ( n22046 , n19119 );
not ( n22047 , n14641 );
and ( n22048 , n22047 , n14725 );
xor ( n22049 , n21691 , n21692 );
xor ( n22050 , n22049 , n21796 );
buf ( n22051 , n22050 );
and ( n22052 , n22051 , n14641 );
or ( n22053 , n22048 , n22052 );
and ( n22054 , n22053 , n21353 );
not ( n22055 , n21630 );
and ( n22056 , n22055 , n21612 );
xor ( n22057 , n22000 , n22035 );
and ( n22058 , n22057 , n21630 );
or ( n22059 , n22056 , n22058 );
buf ( n22060 , n22059 );
and ( n22061 , n22060 , n21255 );
or ( n22062 , n22054 , n22061 );
buf ( n22063 , n22062 );
not ( n22064 , n22063 );
and ( n22065 , n22046 , n22064 );
buf ( n22066 , n19085 );
not ( n22067 , n14641 );
and ( n22068 , n22067 , n14731 );
xor ( n22069 , n21694 , n21695 );
xor ( n22070 , n22069 , n21793 );
buf ( n22071 , n22070 );
and ( n22072 , n22071 , n14641 );
or ( n22073 , n22068 , n22072 );
and ( n22074 , n22073 , n21353 );
not ( n22075 , n21630 );
and ( n22076 , n22075 , n21598 );
xor ( n22077 , n22001 , n22034 );
and ( n22078 , n22077 , n21630 );
or ( n22079 , n22076 , n22078 );
buf ( n22080 , n22079 );
and ( n22081 , n22080 , n21255 );
or ( n22082 , n22074 , n22081 );
buf ( n22083 , n22082 );
not ( n22084 , n22083 );
and ( n22085 , n22066 , n22084 );
buf ( n22086 , n19051 );
not ( n22087 , n14641 );
and ( n22088 , n22087 , n14737 );
xor ( n22089 , n21697 , n21698 );
xor ( n22090 , n22089 , n21790 );
buf ( n22091 , n22090 );
and ( n22092 , n22091 , n14641 );
or ( n22093 , n22088 , n22092 );
and ( n22094 , n22093 , n21353 );
not ( n22095 , n21630 );
and ( n22096 , n22095 , n21584 );
xor ( n22097 , n22002 , n22033 );
and ( n22098 , n22097 , n21630 );
or ( n22099 , n22096 , n22098 );
buf ( n22100 , n22099 );
and ( n22101 , n22100 , n21255 );
or ( n22102 , n22094 , n22101 );
buf ( n22103 , n22102 );
not ( n22104 , n22103 );
and ( n22105 , n22086 , n22104 );
buf ( n22106 , n19017 );
not ( n22107 , n14641 );
and ( n22108 , n22107 , n14743 );
xor ( n22109 , n21700 , n21701 );
xor ( n22110 , n22109 , n21787 );
buf ( n22111 , n22110 );
and ( n22112 , n22111 , n14641 );
or ( n22113 , n22108 , n22112 );
and ( n22114 , n22113 , n21353 );
not ( n22115 , n21630 );
and ( n22116 , n22115 , n21570 );
xor ( n22117 , n22003 , n22032 );
and ( n22118 , n22117 , n21630 );
or ( n22119 , n22116 , n22118 );
buf ( n22120 , n22119 );
and ( n22121 , n22120 , n21255 );
or ( n22122 , n22114 , n22121 );
buf ( n22123 , n22122 );
not ( n22124 , n22123 );
and ( n22125 , n22106 , n22124 );
buf ( n22126 , n18983 );
not ( n22127 , n14641 );
and ( n22128 , n22127 , n14749 );
xor ( n22129 , n21703 , n21704 );
xor ( n22130 , n22129 , n21784 );
buf ( n22131 , n22130 );
and ( n22132 , n22131 , n14641 );
or ( n22133 , n22128 , n22132 );
and ( n22134 , n22133 , n21353 );
not ( n22135 , n21630 );
and ( n22136 , n22135 , n21556 );
xor ( n22137 , n22004 , n22031 );
and ( n22138 , n22137 , n21630 );
or ( n22139 , n22136 , n22138 );
buf ( n22140 , n22139 );
and ( n22141 , n22140 , n21255 );
or ( n22142 , n22134 , n22141 );
buf ( n22143 , n22142 );
not ( n22144 , n22143 );
and ( n22145 , n22126 , n22144 );
buf ( n22146 , n18949 );
not ( n22147 , n14641 );
and ( n22148 , n22147 , n14755 );
xor ( n22149 , n21706 , n21707 );
xor ( n22150 , n22149 , n21781 );
buf ( n22151 , n22150 );
and ( n22152 , n22151 , n14641 );
or ( n22153 , n22148 , n22152 );
and ( n22154 , n22153 , n21353 );
not ( n22155 , n21630 );
and ( n22156 , n22155 , n21542 );
xor ( n22157 , n22005 , n22030 );
and ( n22158 , n22157 , n21630 );
or ( n22159 , n22156 , n22158 );
buf ( n22160 , n22159 );
and ( n22161 , n22160 , n21255 );
or ( n22162 , n22154 , n22161 );
buf ( n22163 , n22162 );
not ( n22164 , n22163 );
and ( n22165 , n22146 , n22164 );
buf ( n22166 , n18915 );
not ( n22167 , n14641 );
and ( n22168 , n22167 , n14761 );
xor ( n22169 , n21709 , n21710 );
xor ( n22170 , n22169 , n21778 );
buf ( n22171 , n22170 );
and ( n22172 , n22171 , n14641 );
or ( n22173 , n22168 , n22172 );
and ( n22174 , n22173 , n21353 );
not ( n22175 , n21630 );
and ( n22176 , n22175 , n21528 );
xor ( n22177 , n22006 , n22029 );
and ( n22178 , n22177 , n21630 );
or ( n22179 , n22176 , n22178 );
buf ( n22180 , n22179 );
and ( n22181 , n22180 , n21255 );
or ( n22182 , n22174 , n22181 );
buf ( n22183 , n22182 );
not ( n22184 , n22183 );
and ( n22185 , n22166 , n22184 );
buf ( n22186 , n18881 );
not ( n22187 , n14641 );
and ( n22188 , n22187 , n14767 );
xor ( n22189 , n21712 , n21713 );
xor ( n22190 , n22189 , n21775 );
buf ( n22191 , n22190 );
and ( n22192 , n22191 , n14641 );
or ( n22193 , n22188 , n22192 );
and ( n22194 , n22193 , n21353 );
not ( n22195 , n21630 );
and ( n22196 , n22195 , n21514 );
xor ( n22197 , n22007 , n22028 );
and ( n22198 , n22197 , n21630 );
or ( n22199 , n22196 , n22198 );
buf ( n22200 , n22199 );
and ( n22201 , n22200 , n21255 );
or ( n22202 , n22194 , n22201 );
buf ( n22203 , n22202 );
not ( n22204 , n22203 );
and ( n22205 , n22186 , n22204 );
buf ( n22206 , n18847 );
not ( n22207 , n14641 );
and ( n22208 , n22207 , n14773 );
xor ( n22209 , n21715 , n21716 );
xor ( n22210 , n22209 , n21772 );
buf ( n22211 , n22210 );
and ( n22212 , n22211 , n14641 );
or ( n22213 , n22208 , n22212 );
and ( n22214 , n22213 , n21353 );
not ( n22215 , n21630 );
and ( n22216 , n22215 , n21500 );
xor ( n22217 , n22008 , n22027 );
and ( n22218 , n22217 , n21630 );
or ( n22219 , n22216 , n22218 );
buf ( n22220 , n22219 );
and ( n22221 , n22220 , n21255 );
or ( n22222 , n22214 , n22221 );
buf ( n22223 , n22222 );
not ( n22224 , n22223 );
and ( n22225 , n22206 , n22224 );
buf ( n22226 , n18813 );
not ( n22227 , n14641 );
and ( n22228 , n22227 , n14779 );
xor ( n22229 , n21718 , n21719 );
xor ( n22230 , n22229 , n21769 );
buf ( n22231 , n22230 );
and ( n22232 , n22231 , n14641 );
or ( n22233 , n22228 , n22232 );
and ( n22234 , n22233 , n21353 );
not ( n22235 , n21630 );
and ( n22236 , n22235 , n21486 );
xor ( n22237 , n22009 , n22026 );
and ( n22238 , n22237 , n21630 );
or ( n22239 , n22236 , n22238 );
buf ( n22240 , n22239 );
and ( n22241 , n22240 , n21255 );
or ( n22242 , n22234 , n22241 );
buf ( n22243 , n22242 );
not ( n22244 , n22243 );
and ( n22245 , n22226 , n22244 );
buf ( n22246 , n18779 );
not ( n22247 , n14641 );
and ( n22248 , n22247 , n14785 );
xor ( n22249 , n21721 , n21722 );
xor ( n22250 , n22249 , n21766 );
buf ( n22251 , n22250 );
and ( n22252 , n22251 , n14641 );
or ( n22253 , n22248 , n22252 );
and ( n22254 , n22253 , n21353 );
not ( n22255 , n21630 );
and ( n22256 , n22255 , n21472 );
xor ( n22257 , n22010 , n22025 );
and ( n22258 , n22257 , n21630 );
or ( n22259 , n22256 , n22258 );
buf ( n22260 , n22259 );
and ( n22261 , n22260 , n21255 );
or ( n22262 , n22254 , n22261 );
buf ( n22263 , n22262 );
not ( n22264 , n22263 );
and ( n22265 , n22246 , n22264 );
buf ( n22266 , n18745 );
not ( n22267 , n14641 );
and ( n22268 , n22267 , n14791 );
xor ( n22269 , n21724 , n21725 );
xor ( n22270 , n22269 , n21763 );
buf ( n22271 , n22270 );
and ( n22272 , n22271 , n14641 );
or ( n22273 , n22268 , n22272 );
and ( n22274 , n22273 , n21353 );
not ( n22275 , n21630 );
and ( n22276 , n22275 , n21458 );
xor ( n22277 , n22011 , n22024 );
and ( n22278 , n22277 , n21630 );
or ( n22279 , n22276 , n22278 );
buf ( n22280 , n22279 );
and ( n22281 , n22280 , n21255 );
or ( n22282 , n22274 , n22281 );
buf ( n22283 , n22282 );
not ( n22284 , n22283 );
and ( n22285 , n22266 , n22284 );
buf ( n22286 , n18711 );
not ( n22287 , n14641 );
and ( n22288 , n22287 , n14797 );
xor ( n22289 , n21727 , n21728 );
xor ( n22290 , n22289 , n21760 );
buf ( n22291 , n22290 );
and ( n22292 , n22291 , n14641 );
or ( n22293 , n22288 , n22292 );
and ( n22294 , n22293 , n21353 );
not ( n22295 , n21630 );
and ( n22296 , n22295 , n21444 );
xor ( n22297 , n22012 , n22023 );
and ( n22298 , n22297 , n21630 );
or ( n22299 , n22296 , n22298 );
buf ( n22300 , n22299 );
and ( n22301 , n22300 , n21255 );
or ( n22302 , n22294 , n22301 );
buf ( n22303 , n22302 );
not ( n22304 , n22303 );
and ( n22305 , n22286 , n22304 );
buf ( n22306 , n18677 );
not ( n22307 , n14641 );
and ( n22308 , n22307 , n14803 );
xor ( n22309 , n21730 , n21731 );
xor ( n22310 , n22309 , n21757 );
buf ( n22311 , n22310 );
and ( n22312 , n22311 , n14641 );
or ( n22313 , n22308 , n22312 );
and ( n22314 , n22313 , n21353 );
not ( n22315 , n21630 );
and ( n22316 , n22315 , n21430 );
xor ( n22317 , n22013 , n22022 );
and ( n22318 , n22317 , n21630 );
or ( n22319 , n22316 , n22318 );
buf ( n22320 , n22319 );
and ( n22321 , n22320 , n21255 );
or ( n22322 , n22314 , n22321 );
buf ( n22323 , n22322 );
not ( n22324 , n22323 );
and ( n22325 , n22306 , n22324 );
buf ( n22326 , n18643 );
not ( n22327 , n14641 );
and ( n22328 , n22327 , n14809 );
xor ( n22329 , n21733 , n21734 );
xor ( n22330 , n22329 , n21754 );
buf ( n22331 , n22330 );
and ( n22332 , n22331 , n14641 );
or ( n22333 , n22328 , n22332 );
and ( n22334 , n22333 , n21353 );
not ( n22335 , n21630 );
and ( n22336 , n22335 , n21416 );
xor ( n22337 , n22014 , n22021 );
and ( n22338 , n22337 , n21630 );
or ( n22339 , n22336 , n22338 );
buf ( n22340 , n22339 );
and ( n22341 , n22340 , n21255 );
or ( n22342 , n22334 , n22341 );
buf ( n22343 , n22342 );
not ( n22344 , n22343 );
and ( n22345 , n22326 , n22344 );
buf ( n22346 , n18610 );
not ( n22347 , n14641 );
and ( n22348 , n22347 , n14815 );
xor ( n22349 , n21736 , n21737 );
xor ( n22350 , n22349 , n21751 );
buf ( n22351 , n22350 );
and ( n22352 , n22351 , n14641 );
or ( n22353 , n22348 , n22352 );
and ( n22354 , n22353 , n21353 );
not ( n22355 , n21630 );
and ( n22356 , n22355 , n21402 );
xor ( n22357 , n22015 , n22020 );
and ( n22358 , n22357 , n21630 );
or ( n22359 , n22356 , n22358 );
buf ( n22360 , n22359 );
and ( n22361 , n22360 , n21255 );
or ( n22362 , n22354 , n22361 );
buf ( n22363 , n22362 );
not ( n22364 , n22363 );
and ( n22365 , n22346 , n22364 );
buf ( n22366 , n18577 );
not ( n22367 , n14641 );
and ( n22368 , n22367 , n14821 );
xor ( n22369 , n21739 , n21740 );
xor ( n22370 , n22369 , n21748 );
buf ( n22371 , n22370 );
and ( n22372 , n22371 , n14641 );
or ( n22373 , n22368 , n22372 );
and ( n22374 , n22373 , n21353 );
not ( n22375 , n21630 );
and ( n22376 , n22375 , n21388 );
xor ( n22377 , n22016 , n22019 );
and ( n22378 , n22377 , n21630 );
or ( n22379 , n22376 , n22378 );
buf ( n22380 , n22379 );
and ( n22381 , n22380 , n21255 );
or ( n22382 , n22374 , n22381 );
buf ( n22383 , n22382 );
not ( n22384 , n22383 );
and ( n22385 , n22366 , n22384 );
buf ( n22386 , n18546 );
not ( n22387 , n14641 );
and ( n22388 , n22387 , n14827 );
xor ( n22389 , n21742 , n21743 );
xor ( n22390 , n22389 , n21745 );
buf ( n22391 , n22390 );
and ( n22392 , n22391 , n14641 );
or ( n22393 , n22388 , n22392 );
and ( n22394 , n22393 , n21353 );
not ( n22395 , n21630 );
and ( n22396 , n22395 , n21374 );
xor ( n22397 , n22017 , n22018 );
and ( n22398 , n22397 , n21630 );
or ( n22399 , n22396 , n22398 );
buf ( n22400 , n22399 );
and ( n22401 , n22400 , n21255 );
or ( n22402 , n22394 , n22401 );
buf ( n22403 , n22402 );
not ( n22404 , n22403 );
and ( n22405 , n22386 , n22404 );
not ( n22406 , n21640 );
or ( n22407 , n21343 , n22406 );
and ( n22408 , n22404 , n22407 );
and ( n22409 , n22386 , n22407 );
or ( n22410 , n22405 , n22408 , n22409 );
and ( n22411 , n22384 , n22410 );
and ( n22412 , n22366 , n22410 );
or ( n22413 , n22385 , n22411 , n22412 );
and ( n22414 , n22364 , n22413 );
and ( n22415 , n22346 , n22413 );
or ( n22416 , n22365 , n22414 , n22415 );
and ( n22417 , n22344 , n22416 );
and ( n22418 , n22326 , n22416 );
or ( n22419 , n22345 , n22417 , n22418 );
and ( n22420 , n22324 , n22419 );
and ( n22421 , n22306 , n22419 );
or ( n22422 , n22325 , n22420 , n22421 );
and ( n22423 , n22304 , n22422 );
and ( n22424 , n22286 , n22422 );
or ( n22425 , n22305 , n22423 , n22424 );
and ( n22426 , n22284 , n22425 );
and ( n22427 , n22266 , n22425 );
or ( n22428 , n22285 , n22426 , n22427 );
and ( n22429 , n22264 , n22428 );
and ( n22430 , n22246 , n22428 );
or ( n22431 , n22265 , n22429 , n22430 );
and ( n22432 , n22244 , n22431 );
and ( n22433 , n22226 , n22431 );
or ( n22434 , n22245 , n22432 , n22433 );
and ( n22435 , n22224 , n22434 );
and ( n22436 , n22206 , n22434 );
or ( n22437 , n22225 , n22435 , n22436 );
and ( n22438 , n22204 , n22437 );
and ( n22439 , n22186 , n22437 );
or ( n22440 , n22205 , n22438 , n22439 );
and ( n22441 , n22184 , n22440 );
and ( n22442 , n22166 , n22440 );
or ( n22443 , n22185 , n22441 , n22442 );
and ( n22444 , n22164 , n22443 );
and ( n22445 , n22146 , n22443 );
or ( n22446 , n22165 , n22444 , n22445 );
and ( n22447 , n22144 , n22446 );
and ( n22448 , n22126 , n22446 );
or ( n22449 , n22145 , n22447 , n22448 );
and ( n22450 , n22124 , n22449 );
and ( n22451 , n22106 , n22449 );
or ( n22452 , n22125 , n22450 , n22451 );
and ( n22453 , n22104 , n22452 );
and ( n22454 , n22086 , n22452 );
or ( n22455 , n22105 , n22453 , n22454 );
and ( n22456 , n22084 , n22455 );
and ( n22457 , n22066 , n22455 );
or ( n22458 , n22085 , n22456 , n22457 );
and ( n22459 , n22064 , n22458 );
and ( n22460 , n22046 , n22458 );
or ( n22461 , n22065 , n22459 , n22460 );
and ( n22462 , n22044 , n22461 );
and ( n22463 , n21988 , n22461 );
or ( n22464 , n22045 , n22462 , n22463 );
and ( n22465 , n21986 , n22464 );
and ( n22466 , n21975 , n22464 );
or ( n22467 , n21987 , n22465 , n22466 );
and ( n22468 , n21973 , n22467 );
and ( n22469 , n21962 , n22467 );
or ( n22470 , n21974 , n22468 , n22469 );
and ( n22471 , n21960 , n22470 );
and ( n22472 , n21949 , n22470 );
or ( n22473 , n21961 , n22471 , n22472 );
and ( n22474 , n21947 , n22473 );
and ( n22475 , n21936 , n22473 );
or ( n22476 , n21948 , n22474 , n22475 );
and ( n22477 , n21934 , n22476 );
and ( n22478 , n21923 , n22476 );
or ( n22479 , n21935 , n22477 , n22478 );
and ( n22480 , n21921 , n22479 );
and ( n22481 , n21910 , n22479 );
or ( n22482 , n21922 , n22480 , n22481 );
and ( n22483 , n21908 , n22482 );
and ( n22484 , n21897 , n22482 );
or ( n22485 , n21909 , n22483 , n22484 );
and ( n22486 , n21895 , n22485 );
and ( n22487 , n21884 , n22485 );
or ( n22488 , n21896 , n22486 , n22487 );
and ( n22489 , n21882 , n22488 );
and ( n22490 , n21871 , n22488 );
or ( n22491 , n21883 , n22489 , n22490 );
and ( n22492 , n21869 , n22491 );
and ( n22493 , n21858 , n22491 );
or ( n22494 , n21870 , n22492 , n22493 );
and ( n22495 , n21856 , n22494 );
and ( n22496 , n21845 , n22494 );
or ( n22497 , n21857 , n22495 , n22496 );
xor ( n22498 , n21844 , n22497 );
buf ( n22499 , n22498 );
buf ( n22500 , n22499 );
not ( n22501 , n22500 );
xor ( n22502 , n22386 , n22404 );
xor ( n22503 , n22502 , n22407 );
buf ( n22504 , n22503 );
buf ( n22505 , n22504 );
and ( n22506 , n22501 , n22505 );
not ( n22507 , n22505 );
not ( n22508 , n21643 );
xor ( n22509 , n22507 , n22508 );
and ( n22510 , n22509 , n22500 );
or ( n22511 , n22506 , n22510 );
buf ( n22512 , n22511 );
not ( n22513 , n22512 );
buf ( n22514 , n22513 );
buf ( n22515 , n22514 );
not ( n22516 , n22515 );
or ( n22517 , n21648 , n22516 );
not ( n22518 , n22500 );
xor ( n22519 , n22366 , n22384 );
xor ( n22520 , n22519 , n22410 );
buf ( n22521 , n22520 );
buf ( n22522 , n22521 );
and ( n22523 , n22518 , n22522 );
not ( n22524 , n22522 );
and ( n22525 , n22507 , n22508 );
xor ( n22526 , n22524 , n22525 );
and ( n22527 , n22526 , n22500 );
or ( n22528 , n22523 , n22527 );
buf ( n22529 , n22528 );
not ( n22530 , n22529 );
buf ( n22531 , n22530 );
buf ( n22532 , n22531 );
not ( n22533 , n22532 );
or ( n22534 , n22517 , n22533 );
not ( n22535 , n22500 );
xor ( n22536 , n22346 , n22364 );
xor ( n22537 , n22536 , n22413 );
buf ( n22538 , n22537 );
buf ( n22539 , n22538 );
and ( n22540 , n22535 , n22539 );
not ( n22541 , n22539 );
and ( n22542 , n22524 , n22525 );
xor ( n22543 , n22541 , n22542 );
and ( n22544 , n22543 , n22500 );
or ( n22545 , n22540 , n22544 );
buf ( n22546 , n22545 );
not ( n22547 , n22546 );
buf ( n22548 , n22547 );
buf ( n22549 , n22548 );
not ( n22550 , n22549 );
or ( n22551 , n22534 , n22550 );
not ( n22552 , n22500 );
xor ( n22553 , n22326 , n22344 );
xor ( n22554 , n22553 , n22416 );
buf ( n22555 , n22554 );
buf ( n22556 , n22555 );
and ( n22557 , n22552 , n22556 );
not ( n22558 , n22556 );
and ( n22559 , n22541 , n22542 );
xor ( n22560 , n22558 , n22559 );
and ( n22561 , n22560 , n22500 );
or ( n22562 , n22557 , n22561 );
buf ( n22563 , n22562 );
not ( n22564 , n22563 );
buf ( n22565 , n22564 );
buf ( n22566 , n22565 );
not ( n22567 , n22566 );
or ( n22568 , n22551 , n22567 );
not ( n22569 , n22500 );
xor ( n22570 , n22306 , n22324 );
xor ( n22571 , n22570 , n22419 );
buf ( n22572 , n22571 );
buf ( n22573 , n22572 );
and ( n22574 , n22569 , n22573 );
not ( n22575 , n22573 );
and ( n22576 , n22558 , n22559 );
xor ( n22577 , n22575 , n22576 );
and ( n22578 , n22577 , n22500 );
or ( n22579 , n22574 , n22578 );
buf ( n22580 , n22579 );
not ( n22581 , n22580 );
buf ( n22582 , n22581 );
buf ( n22583 , n22582 );
not ( n22584 , n22583 );
or ( n22585 , n22568 , n22584 );
not ( n22586 , n22500 );
xor ( n22587 , n22286 , n22304 );
xor ( n22588 , n22587 , n22422 );
buf ( n22589 , n22588 );
buf ( n22590 , n22589 );
and ( n22591 , n22586 , n22590 );
not ( n22592 , n22590 );
and ( n22593 , n22575 , n22576 );
xor ( n22594 , n22592 , n22593 );
and ( n22595 , n22594 , n22500 );
or ( n22596 , n22591 , n22595 );
buf ( n22597 , n22596 );
not ( n22598 , n22597 );
buf ( n22599 , n22598 );
buf ( n22600 , n22599 );
not ( n22601 , n22600 );
or ( n22602 , n22585 , n22601 );
not ( n22603 , n22500 );
xor ( n22604 , n22266 , n22284 );
xor ( n22605 , n22604 , n22425 );
buf ( n22606 , n22605 );
buf ( n22607 , n22606 );
and ( n22608 , n22603 , n22607 );
not ( n22609 , n22607 );
and ( n22610 , n22592 , n22593 );
xor ( n22611 , n22609 , n22610 );
and ( n22612 , n22611 , n22500 );
or ( n22613 , n22608 , n22612 );
buf ( n22614 , n22613 );
not ( n22615 , n22614 );
buf ( n22616 , n22615 );
buf ( n22617 , n22616 );
not ( n22618 , n22617 );
or ( n22619 , n22602 , n22618 );
not ( n22620 , n22500 );
xor ( n22621 , n22246 , n22264 );
xor ( n22622 , n22621 , n22428 );
buf ( n22623 , n22622 );
buf ( n22624 , n22623 );
and ( n22625 , n22620 , n22624 );
not ( n22626 , n22624 );
and ( n22627 , n22609 , n22610 );
xor ( n22628 , n22626 , n22627 );
and ( n22629 , n22628 , n22500 );
or ( n22630 , n22625 , n22629 );
buf ( n22631 , n22630 );
not ( n22632 , n22631 );
buf ( n22633 , n22632 );
buf ( n22634 , n22633 );
not ( n22635 , n22634 );
or ( n22636 , n22619 , n22635 );
not ( n22637 , n22500 );
xor ( n22638 , n22226 , n22244 );
xor ( n22639 , n22638 , n22431 );
buf ( n22640 , n22639 );
buf ( n22641 , n22640 );
and ( n22642 , n22637 , n22641 );
not ( n22643 , n22641 );
and ( n22644 , n22626 , n22627 );
xor ( n22645 , n22643 , n22644 );
and ( n22646 , n22645 , n22500 );
or ( n22647 , n22642 , n22646 );
buf ( n22648 , n22647 );
not ( n22649 , n22648 );
buf ( n22650 , n22649 );
buf ( n22651 , n22650 );
not ( n22652 , n22651 );
or ( n22653 , n22636 , n22652 );
not ( n22654 , n22500 );
xor ( n22655 , n22206 , n22224 );
xor ( n22656 , n22655 , n22434 );
buf ( n22657 , n22656 );
buf ( n22658 , n22657 );
and ( n22659 , n22654 , n22658 );
not ( n22660 , n22658 );
and ( n22661 , n22643 , n22644 );
xor ( n22662 , n22660 , n22661 );
and ( n22663 , n22662 , n22500 );
or ( n22664 , n22659 , n22663 );
buf ( n22665 , n22664 );
not ( n22666 , n22665 );
buf ( n22667 , n22666 );
buf ( n22668 , n22667 );
not ( n22669 , n22668 );
or ( n22670 , n22653 , n22669 );
not ( n22671 , n22500 );
xor ( n22672 , n22186 , n22204 );
xor ( n22673 , n22672 , n22437 );
buf ( n22674 , n22673 );
buf ( n22675 , n22674 );
and ( n22676 , n22671 , n22675 );
not ( n22677 , n22675 );
and ( n22678 , n22660 , n22661 );
xor ( n22679 , n22677 , n22678 );
and ( n22680 , n22679 , n22500 );
or ( n22681 , n22676 , n22680 );
buf ( n22682 , n22681 );
not ( n22683 , n22682 );
buf ( n22684 , n22683 );
buf ( n22685 , n22684 );
not ( n22686 , n22685 );
or ( n22687 , n22670 , n22686 );
not ( n22688 , n22500 );
xor ( n22689 , n22166 , n22184 );
xor ( n22690 , n22689 , n22440 );
buf ( n22691 , n22690 );
buf ( n22692 , n22691 );
and ( n22693 , n22688 , n22692 );
not ( n22694 , n22692 );
and ( n22695 , n22677 , n22678 );
xor ( n22696 , n22694 , n22695 );
and ( n22697 , n22696 , n22500 );
or ( n22698 , n22693 , n22697 );
buf ( n22699 , n22698 );
not ( n22700 , n22699 );
buf ( n22701 , n22700 );
buf ( n22702 , n22701 );
not ( n22703 , n22702 );
or ( n22704 , n22687 , n22703 );
not ( n22705 , n22500 );
xor ( n22706 , n22146 , n22164 );
xor ( n22707 , n22706 , n22443 );
buf ( n22708 , n22707 );
buf ( n22709 , n22708 );
and ( n22710 , n22705 , n22709 );
not ( n22711 , n22709 );
and ( n22712 , n22694 , n22695 );
xor ( n22713 , n22711 , n22712 );
and ( n22714 , n22713 , n22500 );
or ( n22715 , n22710 , n22714 );
buf ( n22716 , n22715 );
not ( n22717 , n22716 );
buf ( n22718 , n22717 );
buf ( n22719 , n22718 );
not ( n22720 , n22719 );
or ( n22721 , n22704 , n22720 );
not ( n22722 , n22500 );
xor ( n22723 , n22126 , n22144 );
xor ( n22724 , n22723 , n22446 );
buf ( n22725 , n22724 );
buf ( n22726 , n22725 );
and ( n22727 , n22722 , n22726 );
not ( n22728 , n22726 );
and ( n22729 , n22711 , n22712 );
xor ( n22730 , n22728 , n22729 );
and ( n22731 , n22730 , n22500 );
or ( n22732 , n22727 , n22731 );
buf ( n22733 , n22732 );
not ( n22734 , n22733 );
buf ( n22735 , n22734 );
buf ( n22736 , n22735 );
not ( n22737 , n22736 );
or ( n22738 , n22721 , n22737 );
not ( n22739 , n22500 );
xor ( n22740 , n22106 , n22124 );
xor ( n22741 , n22740 , n22449 );
buf ( n22742 , n22741 );
buf ( n22743 , n22742 );
and ( n22744 , n22739 , n22743 );
not ( n22745 , n22743 );
and ( n22746 , n22728 , n22729 );
xor ( n22747 , n22745 , n22746 );
and ( n22748 , n22747 , n22500 );
or ( n22749 , n22744 , n22748 );
buf ( n22750 , n22749 );
not ( n22751 , n22750 );
buf ( n22752 , n22751 );
buf ( n22753 , n22752 );
not ( n22754 , n22753 );
or ( n22755 , n22738 , n22754 );
not ( n22756 , n22500 );
xor ( n22757 , n22086 , n22104 );
xor ( n22758 , n22757 , n22452 );
buf ( n22759 , n22758 );
buf ( n22760 , n22759 );
and ( n22761 , n22756 , n22760 );
not ( n22762 , n22760 );
and ( n22763 , n22745 , n22746 );
xor ( n22764 , n22762 , n22763 );
and ( n22765 , n22764 , n22500 );
or ( n22766 , n22761 , n22765 );
buf ( n22767 , n22766 );
not ( n22768 , n22767 );
buf ( n22769 , n22768 );
buf ( n22770 , n22769 );
not ( n22771 , n22770 );
or ( n22772 , n22755 , n22771 );
not ( n22773 , n22500 );
xor ( n22774 , n22066 , n22084 );
xor ( n22775 , n22774 , n22455 );
buf ( n22776 , n22775 );
buf ( n22777 , n22776 );
and ( n22778 , n22773 , n22777 );
not ( n22779 , n22777 );
and ( n22780 , n22762 , n22763 );
xor ( n22781 , n22779 , n22780 );
and ( n22782 , n22781 , n22500 );
or ( n22783 , n22778 , n22782 );
buf ( n22784 , n22783 );
not ( n22785 , n22784 );
buf ( n22786 , n22785 );
buf ( n22787 , n22786 );
not ( n22788 , n22787 );
or ( n22789 , n22772 , n22788 );
not ( n22790 , n22500 );
xor ( n22791 , n22046 , n22064 );
xor ( n22792 , n22791 , n22458 );
buf ( n22793 , n22792 );
buf ( n22794 , n22793 );
and ( n22795 , n22790 , n22794 );
not ( n22796 , n22794 );
and ( n22797 , n22779 , n22780 );
xor ( n22798 , n22796 , n22797 );
and ( n22799 , n22798 , n22500 );
or ( n22800 , n22795 , n22799 );
buf ( n22801 , n22800 );
not ( n22802 , n22801 );
buf ( n22803 , n22802 );
buf ( n22804 , n22803 );
not ( n22805 , n22804 );
or ( n22806 , n22789 , n22805 );
not ( n22807 , n22500 );
xor ( n22808 , n21988 , n22044 );
xor ( n22809 , n22808 , n22461 );
buf ( n22810 , n22809 );
buf ( n22811 , n22810 );
and ( n22812 , n22807 , n22811 );
not ( n22813 , n22811 );
and ( n22814 , n22796 , n22797 );
xor ( n22815 , n22813 , n22814 );
and ( n22816 , n22815 , n22500 );
or ( n22817 , n22812 , n22816 );
buf ( n22818 , n22817 );
not ( n22819 , n22818 );
buf ( n22820 , n22819 );
buf ( n22821 , n22820 );
not ( n22822 , n22821 );
or ( n22823 , n22806 , n22822 );
not ( n22824 , n22500 );
xor ( n22825 , n21975 , n21986 );
xor ( n22826 , n22825 , n22464 );
buf ( n22827 , n22826 );
buf ( n22828 , n22827 );
and ( n22829 , n22824 , n22828 );
not ( n22830 , n22828 );
and ( n22831 , n22813 , n22814 );
xor ( n22832 , n22830 , n22831 );
and ( n22833 , n22832 , n22500 );
or ( n22834 , n22829 , n22833 );
buf ( n22835 , n22834 );
not ( n22836 , n22835 );
buf ( n22837 , n22836 );
buf ( n22838 , n22837 );
not ( n22839 , n22838 );
or ( n22840 , n22823 , n22839 );
not ( n22841 , n22500 );
xor ( n22842 , n21962 , n21973 );
xor ( n22843 , n22842 , n22467 );
buf ( n22844 , n22843 );
buf ( n22845 , n22844 );
and ( n22846 , n22841 , n22845 );
not ( n22847 , n22845 );
and ( n22848 , n22830 , n22831 );
xor ( n22849 , n22847 , n22848 );
and ( n22850 , n22849 , n22500 );
or ( n22851 , n22846 , n22850 );
buf ( n22852 , n22851 );
not ( n22853 , n22852 );
buf ( n22854 , n22853 );
buf ( n22855 , n22854 );
not ( n22856 , n22855 );
or ( n22857 , n22840 , n22856 );
not ( n22858 , n22500 );
xor ( n22859 , n21949 , n21960 );
xor ( n22860 , n22859 , n22470 );
buf ( n22861 , n22860 );
buf ( n22862 , n22861 );
and ( n22863 , n22858 , n22862 );
not ( n22864 , n22862 );
and ( n22865 , n22847 , n22848 );
xor ( n22866 , n22864 , n22865 );
and ( n22867 , n22866 , n22500 );
or ( n22868 , n22863 , n22867 );
buf ( n22869 , n22868 );
not ( n22870 , n22869 );
buf ( n22871 , n22870 );
buf ( n22872 , n22871 );
not ( n22873 , n22872 );
or ( n22874 , n22857 , n22873 );
not ( n22875 , n22500 );
xor ( n22876 , n21936 , n21947 );
xor ( n22877 , n22876 , n22473 );
buf ( n22878 , n22877 );
buf ( n22879 , n22878 );
and ( n22880 , n22875 , n22879 );
not ( n22881 , n22879 );
and ( n22882 , n22864 , n22865 );
xor ( n22883 , n22881 , n22882 );
and ( n22884 , n22883 , n22500 );
or ( n22885 , n22880 , n22884 );
buf ( n22886 , n22885 );
not ( n22887 , n22886 );
buf ( n22888 , n22887 );
buf ( n22889 , n22888 );
not ( n22890 , n22889 );
or ( n22891 , n22874 , n22890 );
not ( n22892 , n22500 );
xor ( n22893 , n21923 , n21934 );
xor ( n22894 , n22893 , n22476 );
buf ( n22895 , n22894 );
buf ( n22896 , n22895 );
and ( n22897 , n22892 , n22896 );
not ( n22898 , n22896 );
and ( n22899 , n22881 , n22882 );
xor ( n22900 , n22898 , n22899 );
and ( n22901 , n22900 , n22500 );
or ( n22902 , n22897 , n22901 );
buf ( n22903 , n22902 );
not ( n22904 , n22903 );
buf ( n22905 , n22904 );
buf ( n22906 , n22905 );
not ( n22907 , n22906 );
or ( n22908 , n22891 , n22907 );
not ( n22909 , n22500 );
xor ( n22910 , n21910 , n21921 );
xor ( n22911 , n22910 , n22479 );
buf ( n22912 , n22911 );
buf ( n22913 , n22912 );
and ( n22914 , n22909 , n22913 );
not ( n22915 , n22913 );
and ( n22916 , n22898 , n22899 );
xor ( n22917 , n22915 , n22916 );
and ( n22918 , n22917 , n22500 );
or ( n22919 , n22914 , n22918 );
buf ( n22920 , n22919 );
not ( n22921 , n22920 );
buf ( n22922 , n22921 );
buf ( n22923 , n22922 );
not ( n22924 , n22923 );
or ( n22925 , n22908 , n22924 );
not ( n22926 , n22500 );
xor ( n22927 , n21897 , n21908 );
xor ( n22928 , n22927 , n22482 );
buf ( n22929 , n22928 );
buf ( n22930 , n22929 );
and ( n22931 , n22926 , n22930 );
not ( n22932 , n22930 );
and ( n22933 , n22915 , n22916 );
xor ( n22934 , n22932 , n22933 );
and ( n22935 , n22934 , n22500 );
or ( n22936 , n22931 , n22935 );
buf ( n22937 , n22936 );
not ( n22938 , n22937 );
buf ( n22939 , n22938 );
buf ( n22940 , n22939 );
not ( n22941 , n22940 );
or ( n22942 , n22925 , n22941 );
not ( n22943 , n22500 );
xor ( n22944 , n21884 , n21895 );
xor ( n22945 , n22944 , n22485 );
buf ( n22946 , n22945 );
buf ( n22947 , n22946 );
and ( n22948 , n22943 , n22947 );
not ( n22949 , n22947 );
and ( n22950 , n22932 , n22933 );
xor ( n22951 , n22949 , n22950 );
and ( n22952 , n22951 , n22500 );
or ( n22953 , n22948 , n22952 );
buf ( n22954 , n22953 );
not ( n22955 , n22954 );
buf ( n22956 , n22955 );
buf ( n22957 , n22956 );
not ( n22958 , n22957 );
or ( n22959 , n22942 , n22958 );
not ( n22960 , n22500 );
xor ( n22961 , n21871 , n21882 );
xor ( n22962 , n22961 , n22488 );
buf ( n22963 , n22962 );
buf ( n22964 , n22963 );
and ( n22965 , n22960 , n22964 );
not ( n22966 , n22964 );
and ( n22967 , n22949 , n22950 );
xor ( n22968 , n22966 , n22967 );
and ( n22969 , n22968 , n22500 );
or ( n22970 , n22965 , n22969 );
buf ( n22971 , n22970 );
not ( n22972 , n22971 );
buf ( n22973 , n22972 );
buf ( n22974 , n22973 );
not ( n22975 , n22974 );
or ( n22976 , n22959 , n22975 );
not ( n22977 , n22500 );
xor ( n22978 , n21858 , n21869 );
xor ( n22979 , n22978 , n22491 );
buf ( n22980 , n22979 );
buf ( n22981 , n22980 );
and ( n22982 , n22977 , n22981 );
not ( n22983 , n22981 );
and ( n22984 , n22966 , n22967 );
xor ( n22985 , n22983 , n22984 );
and ( n22986 , n22985 , n22500 );
or ( n22987 , n22982 , n22986 );
buf ( n22988 , n22987 );
not ( n22989 , n22988 );
buf ( n22990 , n22989 );
buf ( n22991 , n22990 );
not ( n22992 , n22991 );
or ( n22993 , n22976 , n22992 );
buf ( n22994 , n22993 );
buf ( n22995 , n22994 );
and ( n22996 , n22995 , n22500 );
not ( n22997 , n22996 );
and ( n22998 , n22997 , n22924 );
xor ( n22999 , n22924 , n22500 );
xor ( n23000 , n22907 , n22500 );
xor ( n23001 , n22890 , n22500 );
xor ( n23002 , n22873 , n22500 );
xor ( n23003 , n22856 , n22500 );
xor ( n23004 , n22839 , n22500 );
xor ( n23005 , n22822 , n22500 );
xor ( n23006 , n22805 , n22500 );
xor ( n23007 , n22788 , n22500 );
xor ( n23008 , n22771 , n22500 );
xor ( n23009 , n22754 , n22500 );
xor ( n23010 , n22737 , n22500 );
xor ( n23011 , n22720 , n22500 );
xor ( n23012 , n22703 , n22500 );
xor ( n23013 , n22686 , n22500 );
xor ( n23014 , n22669 , n22500 );
xor ( n23015 , n22652 , n22500 );
xor ( n23016 , n22635 , n22500 );
xor ( n23017 , n22618 , n22500 );
xor ( n23018 , n22601 , n22500 );
xor ( n23019 , n22584 , n22500 );
xor ( n23020 , n22567 , n22500 );
xor ( n23021 , n22550 , n22500 );
xor ( n23022 , n22533 , n22500 );
xor ( n23023 , n22516 , n22500 );
xor ( n23024 , n21648 , n22500 );
and ( n23025 , n23024 , n22500 );
and ( n23026 , n23023 , n23025 );
and ( n23027 , n23022 , n23026 );
and ( n23028 , n23021 , n23027 );
and ( n23029 , n23020 , n23028 );
and ( n23030 , n23019 , n23029 );
and ( n23031 , n23018 , n23030 );
and ( n23032 , n23017 , n23031 );
and ( n23033 , n23016 , n23032 );
and ( n23034 , n23015 , n23033 );
and ( n23035 , n23014 , n23034 );
and ( n23036 , n23013 , n23035 );
and ( n23037 , n23012 , n23036 );
and ( n23038 , n23011 , n23037 );
and ( n23039 , n23010 , n23038 );
and ( n23040 , n23009 , n23039 );
and ( n23041 , n23008 , n23040 );
and ( n23042 , n23007 , n23041 );
and ( n23043 , n23006 , n23042 );
and ( n23044 , n23005 , n23043 );
and ( n23045 , n23004 , n23044 );
and ( n23046 , n23003 , n23045 );
and ( n23047 , n23002 , n23046 );
and ( n23048 , n23001 , n23047 );
and ( n23049 , n23000 , n23048 );
xor ( n23050 , n22999 , n23049 );
and ( n23051 , n23050 , n22996 );
or ( n23052 , n22998 , n23051 );
buf ( n23053 , n23052 );
and ( n23054 , n23053 , n21330 );
and ( n23055 , n17453 , n21338 );
or ( n23056 , n23054 , n23055 );
not ( n23057 , n17867 );
and ( n23058 , n17869 , n17850 , n17859 , n23057 );
and ( n23059 , n17842 , n17850 , n17859 , n23057 );
or ( n23060 , n23058 , n23059 );
nor ( n23061 , n17869 , n17850 , n17859 , n23057 );
or ( n23062 , n23060 , n23061 );
nor ( n23063 , n17869 , n17851 , n17859 , n23057 );
or ( n23064 , n23062 , n23063 );
and ( n23065 , n23056 , n23064 );
buf ( n23066 , n18514 );
buf ( n23067 , n21639 );
xor ( n23068 , n23066 , n23067 );
buf ( n23069 , n23068 );
buf ( n23070 , n23069 );
buf ( n23071 , n23070 );
not ( n23072 , n23071 );
buf ( n23073 , n23072 );
buf ( n23074 , n23073 );
not ( n23075 , n23074 );
buf ( n23076 , n18527 );
buf ( n23077 , n21841 );
xor ( n23078 , n23076 , n23077 );
buf ( n23079 , n20484 );
buf ( n23080 , n21854 );
and ( n23081 , n23079 , n23080 );
buf ( n23082 , n20496 );
buf ( n23083 , n21867 );
and ( n23084 , n23082 , n23083 );
buf ( n23085 , n19458 );
buf ( n23086 , n21880 );
and ( n23087 , n23085 , n23086 );
buf ( n23088 , n19424 );
buf ( n23089 , n21893 );
and ( n23090 , n23088 , n23089 );
buf ( n23091 , n19390 );
buf ( n23092 , n21906 );
and ( n23093 , n23091 , n23092 );
buf ( n23094 , n19356 );
buf ( n23095 , n21919 );
and ( n23096 , n23094 , n23095 );
buf ( n23097 , n19323 );
buf ( n23098 , n21932 );
and ( n23099 , n23097 , n23098 );
buf ( n23100 , n19289 );
buf ( n23101 , n21945 );
and ( n23102 , n23100 , n23101 );
buf ( n23103 , n19255 );
buf ( n23104 , n21958 );
and ( n23105 , n23103 , n23104 );
buf ( n23106 , n19221 );
buf ( n23107 , n21971 );
and ( n23108 , n23106 , n23107 );
buf ( n23109 , n19187 );
buf ( n23110 , n21984 );
and ( n23111 , n23109 , n23110 );
buf ( n23112 , n19153 );
buf ( n23113 , n22042 );
and ( n23114 , n23112 , n23113 );
buf ( n23115 , n19119 );
buf ( n23116 , n22062 );
and ( n23117 , n23115 , n23116 );
buf ( n23118 , n19085 );
buf ( n23119 , n22082 );
and ( n23120 , n23118 , n23119 );
buf ( n23121 , n19051 );
buf ( n23122 , n22102 );
and ( n23123 , n23121 , n23122 );
buf ( n23124 , n19017 );
buf ( n23125 , n22122 );
and ( n23126 , n23124 , n23125 );
buf ( n23127 , n18983 );
buf ( n23128 , n22142 );
and ( n23129 , n23127 , n23128 );
buf ( n23130 , n18949 );
buf ( n23131 , n22162 );
and ( n23132 , n23130 , n23131 );
buf ( n23133 , n18915 );
buf ( n23134 , n22182 );
and ( n23135 , n23133 , n23134 );
buf ( n23136 , n18881 );
buf ( n23137 , n22202 );
and ( n23138 , n23136 , n23137 );
buf ( n23139 , n18847 );
buf ( n23140 , n22222 );
and ( n23141 , n23139 , n23140 );
buf ( n23142 , n18813 );
buf ( n23143 , n22242 );
and ( n23144 , n23142 , n23143 );
buf ( n23145 , n18779 );
buf ( n23146 , n22262 );
and ( n23147 , n23145 , n23146 );
buf ( n23148 , n18745 );
buf ( n23149 , n22282 );
and ( n23150 , n23148 , n23149 );
buf ( n23151 , n18711 );
buf ( n23152 , n22302 );
and ( n23153 , n23151 , n23152 );
buf ( n23154 , n18677 );
buf ( n23155 , n22322 );
and ( n23156 , n23154 , n23155 );
buf ( n23157 , n18643 );
buf ( n23158 , n22342 );
and ( n23159 , n23157 , n23158 );
buf ( n23160 , n18610 );
buf ( n23161 , n22362 );
and ( n23162 , n23160 , n23161 );
buf ( n23163 , n18577 );
buf ( n23164 , n22382 );
and ( n23165 , n23163 , n23164 );
buf ( n23166 , n18546 );
buf ( n23167 , n22402 );
and ( n23168 , n23166 , n23167 );
and ( n23169 , n23066 , n23067 );
and ( n23170 , n23167 , n23169 );
and ( n23171 , n23166 , n23169 );
or ( n23172 , n23168 , n23170 , n23171 );
and ( n23173 , n23164 , n23172 );
and ( n23174 , n23163 , n23172 );
or ( n23175 , n23165 , n23173 , n23174 );
and ( n23176 , n23161 , n23175 );
and ( n23177 , n23160 , n23175 );
or ( n23178 , n23162 , n23176 , n23177 );
and ( n23179 , n23158 , n23178 );
and ( n23180 , n23157 , n23178 );
or ( n23181 , n23159 , n23179 , n23180 );
and ( n23182 , n23155 , n23181 );
and ( n23183 , n23154 , n23181 );
or ( n23184 , n23156 , n23182 , n23183 );
and ( n23185 , n23152 , n23184 );
and ( n23186 , n23151 , n23184 );
or ( n23187 , n23153 , n23185 , n23186 );
and ( n23188 , n23149 , n23187 );
and ( n23189 , n23148 , n23187 );
or ( n23190 , n23150 , n23188 , n23189 );
and ( n23191 , n23146 , n23190 );
and ( n23192 , n23145 , n23190 );
or ( n23193 , n23147 , n23191 , n23192 );
and ( n23194 , n23143 , n23193 );
and ( n23195 , n23142 , n23193 );
or ( n23196 , n23144 , n23194 , n23195 );
and ( n23197 , n23140 , n23196 );
and ( n23198 , n23139 , n23196 );
or ( n23199 , n23141 , n23197 , n23198 );
and ( n23200 , n23137 , n23199 );
and ( n23201 , n23136 , n23199 );
or ( n23202 , n23138 , n23200 , n23201 );
and ( n23203 , n23134 , n23202 );
and ( n23204 , n23133 , n23202 );
or ( n23205 , n23135 , n23203 , n23204 );
and ( n23206 , n23131 , n23205 );
and ( n23207 , n23130 , n23205 );
or ( n23208 , n23132 , n23206 , n23207 );
and ( n23209 , n23128 , n23208 );
and ( n23210 , n23127 , n23208 );
or ( n23211 , n23129 , n23209 , n23210 );
and ( n23212 , n23125 , n23211 );
and ( n23213 , n23124 , n23211 );
or ( n23214 , n23126 , n23212 , n23213 );
and ( n23215 , n23122 , n23214 );
and ( n23216 , n23121 , n23214 );
or ( n23217 , n23123 , n23215 , n23216 );
and ( n23218 , n23119 , n23217 );
and ( n23219 , n23118 , n23217 );
or ( n23220 , n23120 , n23218 , n23219 );
and ( n23221 , n23116 , n23220 );
and ( n23222 , n23115 , n23220 );
or ( n23223 , n23117 , n23221 , n23222 );
and ( n23224 , n23113 , n23223 );
and ( n23225 , n23112 , n23223 );
or ( n23226 , n23114 , n23224 , n23225 );
and ( n23227 , n23110 , n23226 );
and ( n23228 , n23109 , n23226 );
or ( n23229 , n23111 , n23227 , n23228 );
and ( n23230 , n23107 , n23229 );
and ( n23231 , n23106 , n23229 );
or ( n23232 , n23108 , n23230 , n23231 );
and ( n23233 , n23104 , n23232 );
and ( n23234 , n23103 , n23232 );
or ( n23235 , n23105 , n23233 , n23234 );
and ( n23236 , n23101 , n23235 );
and ( n23237 , n23100 , n23235 );
or ( n23238 , n23102 , n23236 , n23237 );
and ( n23239 , n23098 , n23238 );
and ( n23240 , n23097 , n23238 );
or ( n23241 , n23099 , n23239 , n23240 );
and ( n23242 , n23095 , n23241 );
and ( n23243 , n23094 , n23241 );
or ( n23244 , n23096 , n23242 , n23243 );
and ( n23245 , n23092 , n23244 );
and ( n23246 , n23091 , n23244 );
or ( n23247 , n23093 , n23245 , n23246 );
and ( n23248 , n23089 , n23247 );
and ( n23249 , n23088 , n23247 );
or ( n23250 , n23090 , n23248 , n23249 );
and ( n23251 , n23086 , n23250 );
and ( n23252 , n23085 , n23250 );
or ( n23253 , n23087 , n23251 , n23252 );
and ( n23254 , n23083 , n23253 );
and ( n23255 , n23082 , n23253 );
or ( n23256 , n23084 , n23254 , n23255 );
and ( n23257 , n23080 , n23256 );
and ( n23258 , n23079 , n23256 );
or ( n23259 , n23081 , n23257 , n23258 );
xor ( n23260 , n23078 , n23259 );
buf ( n23261 , n23260 );
buf ( n23262 , n23261 );
not ( n23263 , n23262 );
xor ( n23264 , n23166 , n23167 );
xor ( n23265 , n23264 , n23169 );
buf ( n23266 , n23265 );
buf ( n23267 , n23266 );
and ( n23268 , n23263 , n23267 );
not ( n23269 , n23267 );
not ( n23270 , n23070 );
xor ( n23271 , n23269 , n23270 );
and ( n23272 , n23271 , n23262 );
or ( n23273 , n23268 , n23272 );
buf ( n23274 , n23273 );
not ( n23275 , n23274 );
buf ( n23276 , n23275 );
buf ( n23277 , n23276 );
not ( n23278 , n23277 );
or ( n23279 , n23075 , n23278 );
not ( n23280 , n23262 );
xor ( n23281 , n23163 , n23164 );
xor ( n23282 , n23281 , n23172 );
buf ( n23283 , n23282 );
buf ( n23284 , n23283 );
and ( n23285 , n23280 , n23284 );
not ( n23286 , n23284 );
and ( n23287 , n23269 , n23270 );
xor ( n23288 , n23286 , n23287 );
and ( n23289 , n23288 , n23262 );
or ( n23290 , n23285 , n23289 );
buf ( n23291 , n23290 );
not ( n23292 , n23291 );
buf ( n23293 , n23292 );
buf ( n23294 , n23293 );
not ( n23295 , n23294 );
or ( n23296 , n23279 , n23295 );
not ( n23297 , n23262 );
xor ( n23298 , n23160 , n23161 );
xor ( n23299 , n23298 , n23175 );
buf ( n23300 , n23299 );
buf ( n23301 , n23300 );
and ( n23302 , n23297 , n23301 );
not ( n23303 , n23301 );
and ( n23304 , n23286 , n23287 );
xor ( n23305 , n23303 , n23304 );
and ( n23306 , n23305 , n23262 );
or ( n23307 , n23302 , n23306 );
buf ( n23308 , n23307 );
not ( n23309 , n23308 );
buf ( n23310 , n23309 );
buf ( n23311 , n23310 );
not ( n23312 , n23311 );
or ( n23313 , n23296 , n23312 );
not ( n23314 , n23262 );
xor ( n23315 , n23157 , n23158 );
xor ( n23316 , n23315 , n23178 );
buf ( n23317 , n23316 );
buf ( n23318 , n23317 );
and ( n23319 , n23314 , n23318 );
not ( n23320 , n23318 );
and ( n23321 , n23303 , n23304 );
xor ( n23322 , n23320 , n23321 );
and ( n23323 , n23322 , n23262 );
or ( n23324 , n23319 , n23323 );
buf ( n23325 , n23324 );
not ( n23326 , n23325 );
buf ( n23327 , n23326 );
buf ( n23328 , n23327 );
not ( n23329 , n23328 );
or ( n23330 , n23313 , n23329 );
not ( n23331 , n23262 );
xor ( n23332 , n23154 , n23155 );
xor ( n23333 , n23332 , n23181 );
buf ( n23334 , n23333 );
buf ( n23335 , n23334 );
and ( n23336 , n23331 , n23335 );
not ( n23337 , n23335 );
and ( n23338 , n23320 , n23321 );
xor ( n23339 , n23337 , n23338 );
and ( n23340 , n23339 , n23262 );
or ( n23341 , n23336 , n23340 );
buf ( n23342 , n23341 );
not ( n23343 , n23342 );
buf ( n23344 , n23343 );
buf ( n23345 , n23344 );
not ( n23346 , n23345 );
or ( n23347 , n23330 , n23346 );
not ( n23348 , n23262 );
xor ( n23349 , n23151 , n23152 );
xor ( n23350 , n23349 , n23184 );
buf ( n23351 , n23350 );
buf ( n23352 , n23351 );
and ( n23353 , n23348 , n23352 );
not ( n23354 , n23352 );
and ( n23355 , n23337 , n23338 );
xor ( n23356 , n23354 , n23355 );
and ( n23357 , n23356 , n23262 );
or ( n23358 , n23353 , n23357 );
buf ( n23359 , n23358 );
not ( n23360 , n23359 );
buf ( n23361 , n23360 );
buf ( n23362 , n23361 );
not ( n23363 , n23362 );
or ( n23364 , n23347 , n23363 );
not ( n23365 , n23262 );
xor ( n23366 , n23148 , n23149 );
xor ( n23367 , n23366 , n23187 );
buf ( n23368 , n23367 );
buf ( n23369 , n23368 );
and ( n23370 , n23365 , n23369 );
not ( n23371 , n23369 );
and ( n23372 , n23354 , n23355 );
xor ( n23373 , n23371 , n23372 );
and ( n23374 , n23373 , n23262 );
or ( n23375 , n23370 , n23374 );
buf ( n23376 , n23375 );
not ( n23377 , n23376 );
buf ( n23378 , n23377 );
buf ( n23379 , n23378 );
not ( n23380 , n23379 );
or ( n23381 , n23364 , n23380 );
not ( n23382 , n23262 );
xor ( n23383 , n23145 , n23146 );
xor ( n23384 , n23383 , n23190 );
buf ( n23385 , n23384 );
buf ( n23386 , n23385 );
and ( n23387 , n23382 , n23386 );
not ( n23388 , n23386 );
and ( n23389 , n23371 , n23372 );
xor ( n23390 , n23388 , n23389 );
and ( n23391 , n23390 , n23262 );
or ( n23392 , n23387 , n23391 );
buf ( n23393 , n23392 );
not ( n23394 , n23393 );
buf ( n23395 , n23394 );
buf ( n23396 , n23395 );
not ( n23397 , n23396 );
or ( n23398 , n23381 , n23397 );
not ( n23399 , n23262 );
xor ( n23400 , n23142 , n23143 );
xor ( n23401 , n23400 , n23193 );
buf ( n23402 , n23401 );
buf ( n23403 , n23402 );
and ( n23404 , n23399 , n23403 );
not ( n23405 , n23403 );
and ( n23406 , n23388 , n23389 );
xor ( n23407 , n23405 , n23406 );
and ( n23408 , n23407 , n23262 );
or ( n23409 , n23404 , n23408 );
buf ( n23410 , n23409 );
not ( n23411 , n23410 );
buf ( n23412 , n23411 );
buf ( n23413 , n23412 );
not ( n23414 , n23413 );
or ( n23415 , n23398 , n23414 );
not ( n23416 , n23262 );
xor ( n23417 , n23139 , n23140 );
xor ( n23418 , n23417 , n23196 );
buf ( n23419 , n23418 );
buf ( n23420 , n23419 );
and ( n23421 , n23416 , n23420 );
not ( n23422 , n23420 );
and ( n23423 , n23405 , n23406 );
xor ( n23424 , n23422 , n23423 );
and ( n23425 , n23424 , n23262 );
or ( n23426 , n23421 , n23425 );
buf ( n23427 , n23426 );
not ( n23428 , n23427 );
buf ( n23429 , n23428 );
buf ( n23430 , n23429 );
not ( n23431 , n23430 );
or ( n23432 , n23415 , n23431 );
not ( n23433 , n23262 );
xor ( n23434 , n23136 , n23137 );
xor ( n23435 , n23434 , n23199 );
buf ( n23436 , n23435 );
buf ( n23437 , n23436 );
and ( n23438 , n23433 , n23437 );
not ( n23439 , n23437 );
and ( n23440 , n23422 , n23423 );
xor ( n23441 , n23439 , n23440 );
and ( n23442 , n23441 , n23262 );
or ( n23443 , n23438 , n23442 );
buf ( n23444 , n23443 );
not ( n23445 , n23444 );
buf ( n23446 , n23445 );
buf ( n23447 , n23446 );
not ( n23448 , n23447 );
or ( n23449 , n23432 , n23448 );
not ( n23450 , n23262 );
xor ( n23451 , n23133 , n23134 );
xor ( n23452 , n23451 , n23202 );
buf ( n23453 , n23452 );
buf ( n23454 , n23453 );
and ( n23455 , n23450 , n23454 );
not ( n23456 , n23454 );
and ( n23457 , n23439 , n23440 );
xor ( n23458 , n23456 , n23457 );
and ( n23459 , n23458 , n23262 );
or ( n23460 , n23455 , n23459 );
buf ( n23461 , n23460 );
not ( n23462 , n23461 );
buf ( n23463 , n23462 );
buf ( n23464 , n23463 );
not ( n23465 , n23464 );
or ( n23466 , n23449 , n23465 );
not ( n23467 , n23262 );
xor ( n23468 , n23130 , n23131 );
xor ( n23469 , n23468 , n23205 );
buf ( n23470 , n23469 );
buf ( n23471 , n23470 );
and ( n23472 , n23467 , n23471 );
not ( n23473 , n23471 );
and ( n23474 , n23456 , n23457 );
xor ( n23475 , n23473 , n23474 );
and ( n23476 , n23475 , n23262 );
or ( n23477 , n23472 , n23476 );
buf ( n23478 , n23477 );
not ( n23479 , n23478 );
buf ( n23480 , n23479 );
buf ( n23481 , n23480 );
not ( n23482 , n23481 );
or ( n23483 , n23466 , n23482 );
not ( n23484 , n23262 );
xor ( n23485 , n23127 , n23128 );
xor ( n23486 , n23485 , n23208 );
buf ( n23487 , n23486 );
buf ( n23488 , n23487 );
and ( n23489 , n23484 , n23488 );
not ( n23490 , n23488 );
and ( n23491 , n23473 , n23474 );
xor ( n23492 , n23490 , n23491 );
and ( n23493 , n23492 , n23262 );
or ( n23494 , n23489 , n23493 );
buf ( n23495 , n23494 );
not ( n23496 , n23495 );
buf ( n23497 , n23496 );
buf ( n23498 , n23497 );
not ( n23499 , n23498 );
or ( n23500 , n23483 , n23499 );
not ( n23501 , n23262 );
xor ( n23502 , n23124 , n23125 );
xor ( n23503 , n23502 , n23211 );
buf ( n23504 , n23503 );
buf ( n23505 , n23504 );
and ( n23506 , n23501 , n23505 );
not ( n23507 , n23505 );
and ( n23508 , n23490 , n23491 );
xor ( n23509 , n23507 , n23508 );
and ( n23510 , n23509 , n23262 );
or ( n23511 , n23506 , n23510 );
buf ( n23512 , n23511 );
not ( n23513 , n23512 );
buf ( n23514 , n23513 );
buf ( n23515 , n23514 );
not ( n23516 , n23515 );
or ( n23517 , n23500 , n23516 );
not ( n23518 , n23262 );
xor ( n23519 , n23121 , n23122 );
xor ( n23520 , n23519 , n23214 );
buf ( n23521 , n23520 );
buf ( n23522 , n23521 );
and ( n23523 , n23518 , n23522 );
not ( n23524 , n23522 );
and ( n23525 , n23507 , n23508 );
xor ( n23526 , n23524 , n23525 );
and ( n23527 , n23526 , n23262 );
or ( n23528 , n23523 , n23527 );
buf ( n23529 , n23528 );
not ( n23530 , n23529 );
buf ( n23531 , n23530 );
buf ( n23532 , n23531 );
not ( n23533 , n23532 );
or ( n23534 , n23517 , n23533 );
not ( n23535 , n23262 );
xor ( n23536 , n23118 , n23119 );
xor ( n23537 , n23536 , n23217 );
buf ( n23538 , n23537 );
buf ( n23539 , n23538 );
and ( n23540 , n23535 , n23539 );
not ( n23541 , n23539 );
and ( n23542 , n23524 , n23525 );
xor ( n23543 , n23541 , n23542 );
and ( n23544 , n23543 , n23262 );
or ( n23545 , n23540 , n23544 );
buf ( n23546 , n23545 );
not ( n23547 , n23546 );
buf ( n23548 , n23547 );
buf ( n23549 , n23548 );
not ( n23550 , n23549 );
or ( n23551 , n23534 , n23550 );
not ( n23552 , n23262 );
xor ( n23553 , n23115 , n23116 );
xor ( n23554 , n23553 , n23220 );
buf ( n23555 , n23554 );
buf ( n23556 , n23555 );
and ( n23557 , n23552 , n23556 );
not ( n23558 , n23556 );
and ( n23559 , n23541 , n23542 );
xor ( n23560 , n23558 , n23559 );
and ( n23561 , n23560 , n23262 );
or ( n23562 , n23557 , n23561 );
buf ( n23563 , n23562 );
not ( n23564 , n23563 );
buf ( n23565 , n23564 );
buf ( n23566 , n23565 );
not ( n23567 , n23566 );
or ( n23568 , n23551 , n23567 );
not ( n23569 , n23262 );
xor ( n23570 , n23112 , n23113 );
xor ( n23571 , n23570 , n23223 );
buf ( n23572 , n23571 );
buf ( n23573 , n23572 );
and ( n23574 , n23569 , n23573 );
not ( n23575 , n23573 );
and ( n23576 , n23558 , n23559 );
xor ( n23577 , n23575 , n23576 );
and ( n23578 , n23577 , n23262 );
or ( n23579 , n23574 , n23578 );
buf ( n23580 , n23579 );
not ( n23581 , n23580 );
buf ( n23582 , n23581 );
buf ( n23583 , n23582 );
not ( n23584 , n23583 );
or ( n23585 , n23568 , n23584 );
not ( n23586 , n23262 );
xor ( n23587 , n23109 , n23110 );
xor ( n23588 , n23587 , n23226 );
buf ( n23589 , n23588 );
buf ( n23590 , n23589 );
and ( n23591 , n23586 , n23590 );
not ( n23592 , n23590 );
and ( n23593 , n23575 , n23576 );
xor ( n23594 , n23592 , n23593 );
and ( n23595 , n23594 , n23262 );
or ( n23596 , n23591 , n23595 );
buf ( n23597 , n23596 );
not ( n23598 , n23597 );
buf ( n23599 , n23598 );
buf ( n23600 , n23599 );
not ( n23601 , n23600 );
or ( n23602 , n23585 , n23601 );
not ( n23603 , n23262 );
xor ( n23604 , n23106 , n23107 );
xor ( n23605 , n23604 , n23229 );
buf ( n23606 , n23605 );
buf ( n23607 , n23606 );
and ( n23608 , n23603 , n23607 );
not ( n23609 , n23607 );
and ( n23610 , n23592 , n23593 );
xor ( n23611 , n23609 , n23610 );
and ( n23612 , n23611 , n23262 );
or ( n23613 , n23608 , n23612 );
buf ( n23614 , n23613 );
not ( n23615 , n23614 );
buf ( n23616 , n23615 );
buf ( n23617 , n23616 );
not ( n23618 , n23617 );
or ( n23619 , n23602 , n23618 );
not ( n23620 , n23262 );
xor ( n23621 , n23103 , n23104 );
xor ( n23622 , n23621 , n23232 );
buf ( n23623 , n23622 );
buf ( n23624 , n23623 );
and ( n23625 , n23620 , n23624 );
not ( n23626 , n23624 );
and ( n23627 , n23609 , n23610 );
xor ( n23628 , n23626 , n23627 );
and ( n23629 , n23628 , n23262 );
or ( n23630 , n23625 , n23629 );
buf ( n23631 , n23630 );
not ( n23632 , n23631 );
buf ( n23633 , n23632 );
buf ( n23634 , n23633 );
not ( n23635 , n23634 );
or ( n23636 , n23619 , n23635 );
not ( n23637 , n23262 );
xor ( n23638 , n23100 , n23101 );
xor ( n23639 , n23638 , n23235 );
buf ( n23640 , n23639 );
buf ( n23641 , n23640 );
and ( n23642 , n23637 , n23641 );
not ( n23643 , n23641 );
and ( n23644 , n23626 , n23627 );
xor ( n23645 , n23643 , n23644 );
and ( n23646 , n23645 , n23262 );
or ( n23647 , n23642 , n23646 );
buf ( n23648 , n23647 );
not ( n23649 , n23648 );
buf ( n23650 , n23649 );
buf ( n23651 , n23650 );
not ( n23652 , n23651 );
or ( n23653 , n23636 , n23652 );
not ( n23654 , n23262 );
xor ( n23655 , n23097 , n23098 );
xor ( n23656 , n23655 , n23238 );
buf ( n23657 , n23656 );
buf ( n23658 , n23657 );
and ( n23659 , n23654 , n23658 );
not ( n23660 , n23658 );
and ( n23661 , n23643 , n23644 );
xor ( n23662 , n23660 , n23661 );
and ( n23663 , n23662 , n23262 );
or ( n23664 , n23659 , n23663 );
buf ( n23665 , n23664 );
not ( n23666 , n23665 );
buf ( n23667 , n23666 );
buf ( n23668 , n23667 );
not ( n23669 , n23668 );
or ( n23670 , n23653 , n23669 );
not ( n23671 , n23262 );
xor ( n23672 , n23094 , n23095 );
xor ( n23673 , n23672 , n23241 );
buf ( n23674 , n23673 );
buf ( n23675 , n23674 );
and ( n23676 , n23671 , n23675 );
not ( n23677 , n23675 );
and ( n23678 , n23660 , n23661 );
xor ( n23679 , n23677 , n23678 );
and ( n23680 , n23679 , n23262 );
or ( n23681 , n23676 , n23680 );
buf ( n23682 , n23681 );
not ( n23683 , n23682 );
buf ( n23684 , n23683 );
buf ( n23685 , n23684 );
not ( n23686 , n23685 );
or ( n23687 , n23670 , n23686 );
not ( n23688 , n23262 );
xor ( n23689 , n23091 , n23092 );
xor ( n23690 , n23689 , n23244 );
buf ( n23691 , n23690 );
buf ( n23692 , n23691 );
and ( n23693 , n23688 , n23692 );
not ( n23694 , n23692 );
and ( n23695 , n23677 , n23678 );
xor ( n23696 , n23694 , n23695 );
and ( n23697 , n23696 , n23262 );
or ( n23698 , n23693 , n23697 );
buf ( n23699 , n23698 );
not ( n23700 , n23699 );
buf ( n23701 , n23700 );
buf ( n23702 , n23701 );
not ( n23703 , n23702 );
or ( n23704 , n23687 , n23703 );
not ( n23705 , n23262 );
xor ( n23706 , n23088 , n23089 );
xor ( n23707 , n23706 , n23247 );
buf ( n23708 , n23707 );
buf ( n23709 , n23708 );
and ( n23710 , n23705 , n23709 );
not ( n23711 , n23709 );
and ( n23712 , n23694 , n23695 );
xor ( n23713 , n23711 , n23712 );
and ( n23714 , n23713 , n23262 );
or ( n23715 , n23710 , n23714 );
buf ( n23716 , n23715 );
not ( n23717 , n23716 );
buf ( n23718 , n23717 );
buf ( n23719 , n23718 );
not ( n23720 , n23719 );
or ( n23721 , n23704 , n23720 );
not ( n23722 , n23262 );
xor ( n23723 , n23085 , n23086 );
xor ( n23724 , n23723 , n23250 );
buf ( n23725 , n23724 );
buf ( n23726 , n23725 );
and ( n23727 , n23722 , n23726 );
not ( n23728 , n23726 );
and ( n23729 , n23711 , n23712 );
xor ( n23730 , n23728 , n23729 );
and ( n23731 , n23730 , n23262 );
or ( n23732 , n23727 , n23731 );
buf ( n23733 , n23732 );
not ( n23734 , n23733 );
buf ( n23735 , n23734 );
buf ( n23736 , n23735 );
not ( n23737 , n23736 );
or ( n23738 , n23721 , n23737 );
not ( n23739 , n23262 );
xor ( n23740 , n23082 , n23083 );
xor ( n23741 , n23740 , n23253 );
buf ( n23742 , n23741 );
buf ( n23743 , n23742 );
and ( n23744 , n23739 , n23743 );
not ( n23745 , n23743 );
and ( n23746 , n23728 , n23729 );
xor ( n23747 , n23745 , n23746 );
and ( n23748 , n23747 , n23262 );
or ( n23749 , n23744 , n23748 );
buf ( n23750 , n23749 );
not ( n23751 , n23750 );
buf ( n23752 , n23751 );
buf ( n23753 , n23752 );
not ( n23754 , n23753 );
or ( n23755 , n23738 , n23754 );
buf ( n23756 , n23755 );
buf ( n23757 , n23756 );
and ( n23758 , n23757 , n23262 );
not ( n23759 , n23758 );
and ( n23760 , n23759 , n23686 );
xor ( n23761 , n23686 , n23262 );
xor ( n23762 , n23669 , n23262 );
xor ( n23763 , n23652 , n23262 );
xor ( n23764 , n23635 , n23262 );
xor ( n23765 , n23618 , n23262 );
xor ( n23766 , n23601 , n23262 );
xor ( n23767 , n23584 , n23262 );
xor ( n23768 , n23567 , n23262 );
xor ( n23769 , n23550 , n23262 );
xor ( n23770 , n23533 , n23262 );
xor ( n23771 , n23516 , n23262 );
xor ( n23772 , n23499 , n23262 );
xor ( n23773 , n23482 , n23262 );
xor ( n23774 , n23465 , n23262 );
xor ( n23775 , n23448 , n23262 );
xor ( n23776 , n23431 , n23262 );
xor ( n23777 , n23414 , n23262 );
xor ( n23778 , n23397 , n23262 );
xor ( n23779 , n23380 , n23262 );
xor ( n23780 , n23363 , n23262 );
xor ( n23781 , n23346 , n23262 );
xor ( n23782 , n23329 , n23262 );
xor ( n23783 , n23312 , n23262 );
xor ( n23784 , n23295 , n23262 );
xor ( n23785 , n23278 , n23262 );
xor ( n23786 , n23075 , n23262 );
and ( n23787 , n23786 , n23262 );
and ( n23788 , n23785 , n23787 );
and ( n23789 , n23784 , n23788 );
and ( n23790 , n23783 , n23789 );
and ( n23791 , n23782 , n23790 );
and ( n23792 , n23781 , n23791 );
and ( n23793 , n23780 , n23792 );
and ( n23794 , n23779 , n23793 );
and ( n23795 , n23778 , n23794 );
and ( n23796 , n23777 , n23795 );
and ( n23797 , n23776 , n23796 );
and ( n23798 , n23775 , n23797 );
and ( n23799 , n23774 , n23798 );
and ( n23800 , n23773 , n23799 );
and ( n23801 , n23772 , n23800 );
and ( n23802 , n23771 , n23801 );
and ( n23803 , n23770 , n23802 );
and ( n23804 , n23769 , n23803 );
and ( n23805 , n23768 , n23804 );
and ( n23806 , n23767 , n23805 );
and ( n23807 , n23766 , n23806 );
and ( n23808 , n23765 , n23807 );
and ( n23809 , n23764 , n23808 );
and ( n23810 , n23763 , n23809 );
and ( n23811 , n23762 , n23810 );
xor ( n23812 , n23761 , n23811 );
and ( n23813 , n23812 , n23758 );
or ( n23814 , n23760 , n23813 );
buf ( n23815 , n23814 );
and ( n23816 , n23815 , n21330 );
and ( n23817 , n17453 , n21338 );
or ( n23818 , n23816 , n23817 );
and ( n23819 , n17869 , n17851 , n17859 , n23057 );
and ( n23820 , n17842 , n17851 , n17859 , n23057 );
or ( n23821 , n23819 , n23820 );
nor ( n23822 , n17842 , n17850 , n17859 , n23057 );
or ( n23823 , n23821 , n23822 );
nor ( n23824 , n17842 , n17851 , n17859 , n23057 );
or ( n23825 , n23823 , n23824 );
and ( n23826 , n23818 , n23825 );
and ( n23827 , n21919 , n21330 );
and ( n23828 , n17453 , n21338 );
or ( n23829 , n23827 , n23828 );
nor ( n23830 , n17842 , n17851 , n17859 , n17867 );
nor ( n23831 , n17869 , n17851 , n17859 , n17867 );
or ( n23832 , n23830 , n23831 );
and ( n23833 , n23829 , n23832 );
nor ( n23834 , n17869 , n17850 , n17859 , n17867 );
and ( n23835 , n19349 , n23834 );
buf ( n23836 , n21919 );
not ( n23837 , n23836 );
buf ( n23838 , n21932 );
not ( n23839 , n23838 );
buf ( n23840 , n21945 );
not ( n23841 , n23840 );
buf ( n23842 , n21958 );
not ( n23843 , n23842 );
buf ( n23844 , n21971 );
not ( n23845 , n23844 );
buf ( n23846 , n21984 );
not ( n23847 , n23846 );
buf ( n23848 , n22042 );
not ( n23849 , n23848 );
buf ( n23850 , n22062 );
not ( n23851 , n23850 );
buf ( n23852 , n22082 );
not ( n23853 , n23852 );
buf ( n23854 , n22102 );
not ( n23855 , n23854 );
buf ( n23856 , n22122 );
not ( n23857 , n23856 );
buf ( n23858 , n22142 );
not ( n23859 , n23858 );
buf ( n23860 , n22162 );
not ( n23861 , n23860 );
buf ( n23862 , n22182 );
not ( n23863 , n23862 );
buf ( n23864 , n22202 );
not ( n23865 , n23864 );
buf ( n23866 , n22222 );
not ( n23867 , n23866 );
buf ( n23868 , n22242 );
not ( n23869 , n23868 );
buf ( n23870 , n22262 );
not ( n23871 , n23870 );
buf ( n23872 , n22282 );
not ( n23873 , n23872 );
buf ( n23874 , n22302 );
not ( n23875 , n23874 );
buf ( n23876 , n22322 );
not ( n23877 , n23876 );
buf ( n23878 , n22342 );
not ( n23879 , n23878 );
buf ( n23880 , n22362 );
not ( n23881 , n23880 );
buf ( n23882 , n22382 );
not ( n23883 , n23882 );
buf ( n23884 , n22402 );
not ( n23885 , n23884 );
buf ( n23886 , n21639 );
not ( n23887 , n23886 );
and ( n23888 , n23885 , n23887 );
and ( n23889 , n23883 , n23888 );
and ( n23890 , n23881 , n23889 );
and ( n23891 , n23879 , n23890 );
and ( n23892 , n23877 , n23891 );
and ( n23893 , n23875 , n23892 );
and ( n23894 , n23873 , n23893 );
and ( n23895 , n23871 , n23894 );
and ( n23896 , n23869 , n23895 );
and ( n23897 , n23867 , n23896 );
and ( n23898 , n23865 , n23897 );
and ( n23899 , n23863 , n23898 );
and ( n23900 , n23861 , n23899 );
and ( n23901 , n23859 , n23900 );
and ( n23902 , n23857 , n23901 );
and ( n23903 , n23855 , n23902 );
and ( n23904 , n23853 , n23903 );
and ( n23905 , n23851 , n23904 );
and ( n23906 , n23849 , n23905 );
and ( n23907 , n23847 , n23906 );
and ( n23908 , n23845 , n23907 );
and ( n23909 , n23843 , n23908 );
and ( n23910 , n23841 , n23909 );
and ( n23911 , n23839 , n23910 );
xor ( n23912 , n23837 , n23911 );
buf ( n23913 , n23912 );
and ( n23914 , n23913 , n21330 );
and ( n23915 , n17453 , n21338 );
or ( n23916 , n23914 , n23915 );
nor ( n23917 , n17842 , n17850 , n17859 , n17867 );
and ( n23918 , n23916 , n23917 );
or ( n23919 , n17874 , n21342 , n23065 , n23826 , n23833 , n23835 , n23918 );
and ( n23920 , n17452 , n23919 );
and ( n23921 , n17453 , n17451 );
or ( n23922 , n23920 , n23921 );
buf ( n23923 , RI210cfd40_236);
buf ( n23924 , n23923 );
and ( n23925 , n23922 , n23924 );
not ( n23926 , n23923 );
and ( n23927 , n17453 , n23926 );
or ( n23928 , n23925 , n23927 );
buf ( n23929 , n23928 );
buf ( n23930 , n23929 );
buf ( n23931 , RI210c9b48_275);
buf ( n23932 , n23931 );
not ( n23933 , n23932 );
buf ( n23934 , RI210ca3b8_274);
buf ( n23935 , n23934 );
not ( n23936 , n23935 );
buf ( n23937 , RI210ca4a8_272);
buf ( n23938 , n23937 );
not ( n23939 , n23938 );
buf ( n23940 , RI210ca520_271);
buf ( n23941 , n23940 );
not ( n23942 , n23941 );
buf ( n23943 , RI210cad90_270);
buf ( n23944 , n23943 );
not ( n23945 , n23944 );
buf ( n23946 , RI210cae08_269);
buf ( n23947 , n23946 );
not ( n23948 , n23947 );
buf ( n23949 , RI210cae80_268);
buf ( n23950 , n23949 );
not ( n23951 , n23950 );
buf ( n23952 , RI210caef8_267);
buf ( n23953 , n23952 );
not ( n23954 , n23953 );
buf ( n23955 , RI210cb768_266);
buf ( n23956 , n23955 );
not ( n23957 , n23956 );
buf ( n23958 , RI210cb7e0_265);
buf ( n23959 , n23958 );
not ( n23960 , n23959 );
buf ( n23961 , RI210cb858_264);
buf ( n23962 , n23961 );
not ( n23963 , n23962 );
buf ( n23964 , RI210cb8d0_263);
buf ( n23965 , n23964 );
not ( n23966 , n23965 );
buf ( n23967 , RI210cc1b8_261);
buf ( n23968 , n23967 );
not ( n23969 , n23968 );
buf ( n23970 , RI210cc230_260);
buf ( n23971 , n23970 );
not ( n23972 , n23971 );
buf ( n23973 , RI210cc2a8_259);
buf ( n23974 , n23973 );
not ( n23975 , n23974 );
buf ( n23976 , RI210ccb18_258);
buf ( n23977 , n23976 );
not ( n23978 , n23977 );
buf ( n23979 , RI210ccb90_257);
buf ( n23980 , n23979 );
not ( n23981 , n23980 );
buf ( n23982 , RI210ccc08_256);
buf ( n23983 , n23982 );
not ( n23984 , n23983 );
buf ( n23985 , RI210ccc80_255);
buf ( n23986 , n23985 );
not ( n23987 , n23986 );
buf ( n23988 , RI210cd4f0_254);
buf ( n23989 , n23988 );
not ( n23990 , n23989 );
buf ( n23991 , RI210cd568_253);
buf ( n23992 , n23991 );
not ( n23993 , n23992 );
buf ( n23994 , RI210cd5e0_252);
buf ( n23995 , n23994 );
not ( n23996 , n23995 );
buf ( n23997 , RI210c07a0_282);
buf ( n23998 , n23997 );
not ( n23999 , n23998 );
buf ( n24000 , RI210c0818_281);
buf ( n24001 , n24000 );
not ( n24002 , n24001 );
buf ( n24003 , RI210c2078_280);
buf ( n24004 , n24003 );
not ( n24005 , n24004 );
buf ( n24006 , RI210c9170_279);
buf ( n24007 , n24006 );
not ( n24008 , n24007 );
buf ( n24009 , RI210c91e8_278);
buf ( n24010 , n24009 );
not ( n24011 , n24010 );
buf ( n24012 , RI210c9a58_277);
buf ( n24013 , n24012 );
not ( n24014 , n24013 );
buf ( n24015 , RI210c9ad0_276);
buf ( n24016 , n24015 );
not ( n24017 , n24016 );
buf ( n24018 , RI210ca430_273);
buf ( n24019 , n24018 );
not ( n24020 , n24019 );
buf ( n24021 , RI210cc140_262);
buf ( n24022 , n24021 );
not ( n24023 , n24022 );
buf ( n24024 , RI210cd658_251);
buf ( n24025 , n24024 );
not ( n24026 , n24025 );
and ( n24027 , n24023 , n24026 );
and ( n24028 , n24020 , n24027 );
and ( n24029 , n24017 , n24028 );
and ( n24030 , n24014 , n24029 );
and ( n24031 , n24011 , n24030 );
and ( n24032 , n24008 , n24031 );
and ( n24033 , n24005 , n24032 );
and ( n24034 , n24002 , n24033 );
and ( n24035 , n23999 , n24034 );
and ( n24036 , n23996 , n24035 );
and ( n24037 , n23993 , n24036 );
and ( n24038 , n23990 , n24037 );
and ( n24039 , n23987 , n24038 );
and ( n24040 , n23984 , n24039 );
and ( n24041 , n23981 , n24040 );
and ( n24042 , n23978 , n24041 );
and ( n24043 , n23975 , n24042 );
and ( n24044 , n23972 , n24043 );
and ( n24045 , n23969 , n24044 );
and ( n24046 , n23966 , n24045 );
and ( n24047 , n23963 , n24046 );
and ( n24048 , n23960 , n24047 );
and ( n24049 , n23957 , n24048 );
and ( n24050 , n23954 , n24049 );
and ( n24051 , n23951 , n24050 );
and ( n24052 , n23948 , n24051 );
and ( n24053 , n23945 , n24052 );
and ( n24054 , n23942 , n24053 );
and ( n24055 , n23939 , n24054 );
and ( n24056 , n23936 , n24055 );
xor ( n24057 , n23933 , n24056 );
buf ( n24058 , n24057 );
buf ( n24059 , n23931 );
and ( n24060 , n24058 , n24059 );
or ( n24061 , C0 , n24060 );
buf ( n24062 , n24061 );
not ( n24063 , n24062 );
not ( n24064 , n24059 );
and ( n24065 , n24064 , n23955 );
xor ( n24066 , n23957 , n24048 );
buf ( n24067 , n24066 );
and ( n24068 , n24067 , n24059 );
or ( n24069 , n24065 , n24068 );
buf ( n24070 , n24069 );
and ( n24071 , n24063 , n24070 );
not ( n24072 , n24070 );
not ( n24073 , n24059 );
and ( n24074 , n24073 , n23958 );
xor ( n24075 , n23960 , n24047 );
buf ( n24076 , n24075 );
and ( n24077 , n24076 , n24059 );
or ( n24078 , n24074 , n24077 );
buf ( n24079 , n24078 );
not ( n24080 , n24079 );
not ( n24081 , n24059 );
and ( n24082 , n24081 , n23961 );
xor ( n24083 , n23963 , n24046 );
buf ( n24084 , n24083 );
and ( n24085 , n24084 , n24059 );
or ( n24086 , n24082 , n24085 );
buf ( n24087 , n24086 );
not ( n24088 , n24087 );
not ( n24089 , n24059 );
and ( n24090 , n24089 , n23964 );
xor ( n24091 , n23966 , n24045 );
buf ( n24092 , n24091 );
and ( n24093 , n24092 , n24059 );
or ( n24094 , n24090 , n24093 );
buf ( n24095 , n24094 );
not ( n24096 , n24095 );
not ( n24097 , n24059 );
and ( n24098 , n24097 , n23967 );
xor ( n24099 , n23969 , n24044 );
buf ( n24100 , n24099 );
and ( n24101 , n24100 , n24059 );
or ( n24102 , n24098 , n24101 );
buf ( n24103 , n24102 );
not ( n24104 , n24103 );
not ( n24105 , n24059 );
and ( n24106 , n24105 , n23970 );
xor ( n24107 , n23972 , n24043 );
buf ( n24108 , n24107 );
and ( n24109 , n24108 , n24059 );
or ( n24110 , n24106 , n24109 );
buf ( n24111 , n24110 );
not ( n24112 , n24111 );
not ( n24113 , n24059 );
and ( n24114 , n24113 , n23973 );
xor ( n24115 , n23975 , n24042 );
buf ( n24116 , n24115 );
and ( n24117 , n24116 , n24059 );
or ( n24118 , n24114 , n24117 );
buf ( n24119 , n24118 );
not ( n24120 , n24119 );
not ( n24121 , n24059 );
and ( n24122 , n24121 , n23976 );
xor ( n24123 , n23978 , n24041 );
buf ( n24124 , n24123 );
and ( n24125 , n24124 , n24059 );
or ( n24126 , n24122 , n24125 );
buf ( n24127 , n24126 );
not ( n24128 , n24127 );
not ( n24129 , n24059 );
and ( n24130 , n24129 , n23979 );
xor ( n24131 , n23981 , n24040 );
buf ( n24132 , n24131 );
and ( n24133 , n24132 , n24059 );
or ( n24134 , n24130 , n24133 );
buf ( n24135 , n24134 );
not ( n24136 , n24135 );
not ( n24137 , n24059 );
and ( n24138 , n24137 , n23982 );
xor ( n24139 , n23984 , n24039 );
buf ( n24140 , n24139 );
and ( n24141 , n24140 , n24059 );
or ( n24142 , n24138 , n24141 );
buf ( n24143 , n24142 );
not ( n24144 , n24143 );
not ( n24145 , n24059 );
and ( n24146 , n24145 , n23985 );
xor ( n24147 , n23987 , n24038 );
buf ( n24148 , n24147 );
and ( n24149 , n24148 , n24059 );
or ( n24150 , n24146 , n24149 );
buf ( n24151 , n24150 );
not ( n24152 , n24151 );
not ( n24153 , n24059 );
and ( n24154 , n24153 , n23988 );
xor ( n24155 , n23990 , n24037 );
buf ( n24156 , n24155 );
and ( n24157 , n24156 , n24059 );
or ( n24158 , n24154 , n24157 );
buf ( n24159 , n24158 );
not ( n24160 , n24159 );
not ( n24161 , n24059 );
and ( n24162 , n24161 , n23991 );
xor ( n24163 , n23993 , n24036 );
buf ( n24164 , n24163 );
and ( n24165 , n24164 , n24059 );
or ( n24166 , n24162 , n24165 );
buf ( n24167 , n24166 );
not ( n24168 , n24167 );
not ( n24169 , n24059 );
and ( n24170 , n24169 , n23994 );
xor ( n24171 , n23996 , n24035 );
buf ( n24172 , n24171 );
and ( n24173 , n24172 , n24059 );
or ( n24174 , n24170 , n24173 );
buf ( n24175 , n24174 );
not ( n24176 , n24175 );
not ( n24177 , n24059 );
and ( n24178 , n24177 , n23997 );
xor ( n24179 , n23999 , n24034 );
buf ( n24180 , n24179 );
and ( n24181 , n24180 , n24059 );
or ( n24182 , n24178 , n24181 );
buf ( n24183 , n24182 );
not ( n24184 , n24183 );
not ( n24185 , n24059 );
and ( n24186 , n24185 , n24000 );
xor ( n24187 , n24002 , n24033 );
buf ( n24188 , n24187 );
and ( n24189 , n24188 , n24059 );
or ( n24190 , n24186 , n24189 );
buf ( n24191 , n24190 );
not ( n24192 , n24191 );
not ( n24193 , n24059 );
and ( n24194 , n24193 , n24003 );
xor ( n24195 , n24005 , n24032 );
buf ( n24196 , n24195 );
and ( n24197 , n24196 , n24059 );
or ( n24198 , n24194 , n24197 );
buf ( n24199 , n24198 );
not ( n24200 , n24199 );
not ( n24201 , n24059 );
and ( n24202 , n24201 , n24006 );
xor ( n24203 , n24008 , n24031 );
buf ( n24204 , n24203 );
and ( n24205 , n24204 , n24059 );
or ( n24206 , n24202 , n24205 );
buf ( n24207 , n24206 );
not ( n24208 , n24207 );
not ( n24209 , n24059 );
and ( n24210 , n24209 , n24009 );
xor ( n24211 , n24011 , n24030 );
buf ( n24212 , n24211 );
and ( n24213 , n24212 , n24059 );
or ( n24214 , n24210 , n24213 );
buf ( n24215 , n24214 );
not ( n24216 , n24215 );
not ( n24217 , n24059 );
and ( n24218 , n24217 , n24012 );
xor ( n24219 , n24014 , n24029 );
buf ( n24220 , n24219 );
and ( n24221 , n24220 , n24059 );
or ( n24222 , n24218 , n24221 );
buf ( n24223 , n24222 );
not ( n24224 , n24223 );
not ( n24225 , n24059 );
and ( n24226 , n24225 , n24015 );
xor ( n24227 , n24017 , n24028 );
buf ( n24228 , n24227 );
and ( n24229 , n24228 , n24059 );
or ( n24230 , n24226 , n24229 );
buf ( n24231 , n24230 );
not ( n24232 , n24231 );
not ( n24233 , n24059 );
and ( n24234 , n24233 , n24018 );
xor ( n24235 , n24020 , n24027 );
buf ( n24236 , n24235 );
and ( n24237 , n24236 , n24059 );
or ( n24238 , n24234 , n24237 );
buf ( n24239 , n24238 );
not ( n24240 , n24239 );
not ( n24241 , n24059 );
and ( n24242 , n24241 , n24021 );
xor ( n24243 , n24023 , n24026 );
buf ( n24244 , n24243 );
and ( n24245 , n24244 , n24059 );
or ( n24246 , n24242 , n24245 );
buf ( n24247 , n24246 );
not ( n24248 , n24247 );
buf ( n24249 , n24024 );
buf ( n24250 , n24249 );
not ( n24251 , n24250 );
and ( n24252 , n24248 , n24251 );
and ( n24253 , n24240 , n24252 );
and ( n24254 , n24232 , n24253 );
and ( n24255 , n24224 , n24254 );
and ( n24256 , n24216 , n24255 );
and ( n24257 , n24208 , n24256 );
and ( n24258 , n24200 , n24257 );
and ( n24259 , n24192 , n24258 );
and ( n24260 , n24184 , n24259 );
and ( n24261 , n24176 , n24260 );
and ( n24262 , n24168 , n24261 );
and ( n24263 , n24160 , n24262 );
and ( n24264 , n24152 , n24263 );
and ( n24265 , n24144 , n24264 );
and ( n24266 , n24136 , n24265 );
and ( n24267 , n24128 , n24266 );
and ( n24268 , n24120 , n24267 );
and ( n24269 , n24112 , n24268 );
and ( n24270 , n24104 , n24269 );
and ( n24271 , n24096 , n24270 );
and ( n24272 , n24088 , n24271 );
and ( n24273 , n24080 , n24272 );
xor ( n24274 , n24072 , n24273 );
and ( n24275 , n24274 , n24062 );
or ( n24276 , n24071 , n24275 );
buf ( n24277 , n24276 );
not ( n24278 , n24277 );
buf ( n24279 , n24278 );
buf ( n24280 , n24279 );
not ( n24281 , n24280 );
buf ( n24282 , n24281 );
buf ( n24283 , n24282 );
not ( n24284 , n24283 );
buf ( n24285 , n24284 );
buf ( n24286 , n24285 );
not ( n24287 , n24286 );
or ( n24288 , n24287 , C0 );
or ( n24289 , n24288 , C0 );
or ( n24290 , n24289 , C0 );
or ( n24291 , n24290 , C0 );
or ( n24292 , n24291 , C0 );
or ( n24293 , n24292 , C0 );
or ( n24294 , n24293 , C0 );
or ( n24295 , n24294 , C0 );
or ( n24296 , n24295 , C0 );
or ( n24297 , n24296 , C0 );
or ( n24298 , n24297 , C0 );
or ( n24299 , n24298 , C0 );
or ( n24300 , n24299 , C0 );
or ( n24301 , n24300 , C0 );
or ( n24302 , n24301 , C0 );
or ( n24303 , n24302 , C0 );
or ( n24304 , n24303 , C0 );
or ( n24305 , n24304 , C0 );
or ( n24306 , n24305 , C0 );
or ( n24307 , n24306 , C0 );
or ( n24308 , n24307 , C0 );
or ( n24309 , n24308 , C0 );
or ( n24310 , n24309 , C0 );
or ( n24311 , n24310 , C0 );
or ( n24312 , n24311 , C0 );
or ( n24313 , n24312 , C0 );
or ( n24314 , n24313 , C0 );
or ( n24315 , n24314 , C0 );
or ( n24316 , n24315 , C0 );
or ( n24317 , n24316 , C0 );
buf ( n24318 , n24317 );
not ( n24319 , n24062 );
not ( n24320 , n24059 );
and ( n24321 , n24320 , n23934 );
xor ( n24322 , n23936 , n24055 );
buf ( n24323 , n24322 );
and ( n24324 , n24323 , n24059 );
or ( n24325 , n24321 , n24324 );
buf ( n24326 , n24325 );
not ( n24327 , n24326 );
not ( n24328 , n24059 );
and ( n24329 , n24328 , n23937 );
xor ( n24330 , n23939 , n24054 );
buf ( n24331 , n24330 );
and ( n24332 , n24331 , n24059 );
or ( n24333 , n24329 , n24332 );
buf ( n24334 , n24333 );
not ( n24335 , n24334 );
not ( n24336 , n24059 );
and ( n24337 , n24336 , n23940 );
xor ( n24338 , n23942 , n24053 );
buf ( n24339 , n24338 );
and ( n24340 , n24339 , n24059 );
or ( n24341 , n24337 , n24340 );
buf ( n24342 , n24341 );
not ( n24343 , n24342 );
not ( n24344 , n24059 );
and ( n24345 , n24344 , n23943 );
xor ( n24346 , n23945 , n24052 );
buf ( n24347 , n24346 );
and ( n24348 , n24347 , n24059 );
or ( n24349 , n24345 , n24348 );
buf ( n24350 , n24349 );
not ( n24351 , n24350 );
not ( n24352 , n24059 );
and ( n24353 , n24352 , n23946 );
xor ( n24354 , n23948 , n24051 );
buf ( n24355 , n24354 );
and ( n24356 , n24355 , n24059 );
or ( n24357 , n24353 , n24356 );
buf ( n24358 , n24357 );
not ( n24359 , n24358 );
not ( n24360 , n24059 );
and ( n24361 , n24360 , n23949 );
xor ( n24362 , n23951 , n24050 );
buf ( n24363 , n24362 );
and ( n24364 , n24363 , n24059 );
or ( n24365 , n24361 , n24364 );
buf ( n24366 , n24365 );
not ( n24367 , n24366 );
not ( n24368 , n24059 );
and ( n24369 , n24368 , n23952 );
xor ( n24370 , n23954 , n24049 );
buf ( n24371 , n24370 );
and ( n24372 , n24371 , n24059 );
or ( n24373 , n24369 , n24372 );
buf ( n24374 , n24373 );
not ( n24375 , n24374 );
and ( n24376 , n24072 , n24273 );
and ( n24377 , n24375 , n24376 );
and ( n24378 , n24367 , n24377 );
and ( n24379 , n24359 , n24378 );
and ( n24380 , n24351 , n24379 );
and ( n24381 , n24343 , n24380 );
and ( n24382 , n24335 , n24381 );
and ( n24383 , n24327 , n24382 );
xor ( n24384 , n24319 , n24383 );
buf ( n24385 , n24062 );
and ( n24386 , n24384 , n24385 );
or ( n24387 , C0 , n24386 );
buf ( n24388 , n24387 );
not ( n24389 , n24388 );
buf ( n24390 , n24389 );
buf ( n24391 , n24390 );
not ( n24392 , n24391 );
buf ( n24393 , n24392 );
not ( n24394 , n24393 );
buf ( n24395 , n24394 );
not ( n24396 , n24062 );
and ( n24397 , n24396 , n24326 );
xor ( n24398 , n24327 , n24382 );
and ( n24399 , n24398 , n24062 );
or ( n24400 , n24397 , n24399 );
buf ( n24401 , n24400 );
not ( n24402 , n24401 );
buf ( n24403 , n24402 );
buf ( n24404 , n24403 );
not ( n24405 , n24404 );
buf ( n24406 , n24405 );
not ( n24407 , n24406 );
buf ( n24408 , n24407 );
not ( n24409 , n24062 );
and ( n24410 , n24409 , n24334 );
xor ( n24411 , n24335 , n24381 );
and ( n24412 , n24411 , n24062 );
or ( n24413 , n24410 , n24412 );
buf ( n24414 , n24413 );
not ( n24415 , n24414 );
buf ( n24416 , n24415 );
buf ( n24417 , n24416 );
not ( n24418 , n24417 );
buf ( n24419 , n24418 );
not ( n24420 , n24419 );
buf ( n24421 , n24420 );
not ( n24422 , n24062 );
and ( n24423 , n24422 , n24342 );
xor ( n24424 , n24343 , n24380 );
and ( n24425 , n24424 , n24062 );
or ( n24426 , n24423 , n24425 );
buf ( n24427 , n24426 );
not ( n24428 , n24427 );
buf ( n24429 , n24428 );
buf ( n24430 , n24429 );
not ( n24431 , n24430 );
buf ( n24432 , n24431 );
not ( n24433 , n24432 );
buf ( n24434 , n24433 );
not ( n24435 , n24062 );
and ( n24436 , n24435 , n24350 );
xor ( n24437 , n24351 , n24379 );
and ( n24438 , n24437 , n24062 );
or ( n24439 , n24436 , n24438 );
buf ( n24440 , n24439 );
not ( n24441 , n24440 );
buf ( n24442 , n24441 );
buf ( n24443 , n24442 );
not ( n24444 , n24443 );
buf ( n24445 , n24444 );
not ( n24446 , n24445 );
buf ( n24447 , n24446 );
not ( n24448 , n24062 );
and ( n24449 , n24448 , n24358 );
xor ( n24450 , n24359 , n24378 );
and ( n24451 , n24450 , n24062 );
or ( n24452 , n24449 , n24451 );
buf ( n24453 , n24452 );
not ( n24454 , n24453 );
buf ( n24455 , n24454 );
buf ( n24456 , n24455 );
not ( n24457 , n24456 );
buf ( n24458 , n24457 );
not ( n24459 , n24458 );
buf ( n24460 , n24459 );
not ( n24461 , n24062 );
and ( n24462 , n24461 , n24366 );
xor ( n24463 , n24367 , n24377 );
and ( n24464 , n24463 , n24062 );
or ( n24465 , n24462 , n24464 );
buf ( n24466 , n24465 );
not ( n24467 , n24466 );
buf ( n24468 , n24467 );
buf ( n24469 , n24468 );
not ( n24470 , n24469 );
buf ( n24471 , n24470 );
not ( n24472 , n24471 );
buf ( n24473 , n24472 );
not ( n24474 , n24062 );
and ( n24475 , n24474 , n24374 );
xor ( n24476 , n24375 , n24376 );
and ( n24477 , n24476 , n24062 );
or ( n24478 , n24475 , n24477 );
buf ( n24479 , n24478 );
not ( n24480 , n24479 );
buf ( n24481 , n24480 );
buf ( n24482 , n24481 );
not ( n24483 , n24482 );
buf ( n24484 , n24483 );
not ( n24485 , n24484 );
buf ( n24486 , n24485 );
not ( n24487 , n24282 );
buf ( n24488 , n24487 );
and ( n24489 , n24486 , n24488 );
and ( n24490 , n24473 , n24489 );
and ( n24491 , n24460 , n24490 );
and ( n24492 , n24447 , n24491 );
and ( n24493 , n24434 , n24492 );
and ( n24494 , n24421 , n24493 );
and ( n24495 , n24408 , n24494 );
and ( n24496 , n24395 , n24495 );
not ( n24497 , n24496 );
buf ( n24498 , n24497 );
buf ( n24499 , n24062 );
and ( n24500 , n24498 , n24499 );
or ( n24501 , C0 , n24500 );
buf ( n24502 , n24501 );
buf ( n24503 , n24502 );
and ( n24504 , n24318 , n24503 );
not ( n24505 , n24504 );
and ( n24506 , n24505 , n24287 );
xor ( n24507 , n24287 , n24503 );
xor ( n24508 , n24507 , n24503 );
and ( n24509 , n24508 , n24504 );
or ( n24510 , n24506 , n24509 );
buf ( n24511 , n24510 );
buf ( n24512 , n24061 );
not ( n24513 , n24512 );
buf ( n24514 , n24373 );
and ( n24515 , n24513 , n24514 );
not ( n24516 , n24514 );
buf ( n24517 , n24069 );
not ( n24518 , n24517 );
buf ( n24519 , n24078 );
not ( n24520 , n24519 );
buf ( n24521 , n24086 );
not ( n24522 , n24521 );
buf ( n24523 , n24094 );
not ( n24524 , n24523 );
buf ( n24525 , n24102 );
not ( n24526 , n24525 );
buf ( n24527 , n24110 );
not ( n24528 , n24527 );
buf ( n24529 , n24118 );
not ( n24530 , n24529 );
buf ( n24531 , n24126 );
not ( n24532 , n24531 );
buf ( n24533 , n24134 );
not ( n24534 , n24533 );
buf ( n24535 , n24142 );
not ( n24536 , n24535 );
buf ( n24537 , n24150 );
not ( n24538 , n24537 );
buf ( n24539 , n24158 );
not ( n24540 , n24539 );
buf ( n24541 , n24166 );
not ( n24542 , n24541 );
buf ( n24543 , n24174 );
not ( n24544 , n24543 );
buf ( n24545 , n24182 );
not ( n24546 , n24545 );
buf ( n24547 , n24190 );
not ( n24548 , n24547 );
buf ( n24549 , n24198 );
not ( n24550 , n24549 );
buf ( n24551 , n24206 );
not ( n24552 , n24551 );
buf ( n24553 , n24214 );
not ( n24554 , n24553 );
buf ( n24555 , n24222 );
not ( n24556 , n24555 );
buf ( n24557 , n24230 );
not ( n24558 , n24557 );
buf ( n24559 , n24238 );
not ( n24560 , n24559 );
buf ( n24561 , n24246 );
not ( n24562 , n24561 );
buf ( n24563 , n24249 );
not ( n24564 , n24563 );
and ( n24565 , n24562 , n24564 );
and ( n24566 , n24560 , n24565 );
and ( n24567 , n24558 , n24566 );
and ( n24568 , n24556 , n24567 );
and ( n24569 , n24554 , n24568 );
and ( n24570 , n24552 , n24569 );
and ( n24571 , n24550 , n24570 );
and ( n24572 , n24548 , n24571 );
and ( n24573 , n24546 , n24572 );
and ( n24574 , n24544 , n24573 );
and ( n24575 , n24542 , n24574 );
and ( n24576 , n24540 , n24575 );
and ( n24577 , n24538 , n24576 );
and ( n24578 , n24536 , n24577 );
and ( n24579 , n24534 , n24578 );
and ( n24580 , n24532 , n24579 );
and ( n24581 , n24530 , n24580 );
and ( n24582 , n24528 , n24581 );
and ( n24583 , n24526 , n24582 );
and ( n24584 , n24524 , n24583 );
and ( n24585 , n24522 , n24584 );
and ( n24586 , n24520 , n24585 );
and ( n24587 , n24518 , n24586 );
xor ( n24588 , n24516 , n24587 );
and ( n24589 , n24588 , n24512 );
or ( n24590 , n24515 , n24589 );
buf ( n24591 , n24590 );
not ( n24592 , n24591 );
buf ( n24593 , n24592 );
buf ( n24594 , n24593 );
not ( n24595 , n24594 );
buf ( n24596 , n24595 );
buf ( n24597 , n24596 );
buf ( n24598 , n24597 );
not ( n24599 , n24598 );
buf ( n24600 , n24599 );
buf ( n24601 , n24600 );
not ( n24602 , n24601 );
not ( n24603 , n24512 );
buf ( n24604 , n24325 );
not ( n24605 , n24604 );
buf ( n24606 , n24333 );
not ( n24607 , n24606 );
buf ( n24608 , n24341 );
not ( n24609 , n24608 );
buf ( n24610 , n24349 );
not ( n24611 , n24610 );
buf ( n24612 , n24357 );
not ( n24613 , n24612 );
buf ( n24614 , n24365 );
not ( n24615 , n24614 );
and ( n24616 , n24516 , n24587 );
and ( n24617 , n24615 , n24616 );
and ( n24618 , n24613 , n24617 );
and ( n24619 , n24611 , n24618 );
and ( n24620 , n24609 , n24619 );
and ( n24621 , n24607 , n24620 );
and ( n24622 , n24605 , n24621 );
xor ( n24623 , n24603 , n24622 );
buf ( n24624 , n24512 );
and ( n24625 , n24623 , n24624 );
or ( n24626 , C0 , n24625 );
buf ( n24627 , n24626 );
not ( n24628 , n24627 );
buf ( n24629 , n24628 );
buf ( n24630 , n24629 );
not ( n24631 , n24630 );
buf ( n24632 , n24631 );
not ( n24633 , n24632 );
buf ( n24634 , n24633 );
not ( n24635 , n24512 );
and ( n24636 , n24635 , n24604 );
xor ( n24637 , n24605 , n24621 );
and ( n24638 , n24637 , n24512 );
or ( n24639 , n24636 , n24638 );
buf ( n24640 , n24639 );
not ( n24641 , n24640 );
buf ( n24642 , n24641 );
buf ( n24643 , n24642 );
not ( n24644 , n24643 );
buf ( n24645 , n24644 );
not ( n24646 , n24645 );
buf ( n24647 , n24646 );
not ( n24648 , n24512 );
and ( n24649 , n24648 , n24606 );
xor ( n24650 , n24607 , n24620 );
and ( n24651 , n24650 , n24512 );
or ( n24652 , n24649 , n24651 );
buf ( n24653 , n24652 );
not ( n24654 , n24653 );
buf ( n24655 , n24654 );
buf ( n24656 , n24655 );
not ( n24657 , n24656 );
buf ( n24658 , n24657 );
not ( n24659 , n24658 );
buf ( n24660 , n24659 );
not ( n24661 , n24512 );
and ( n24662 , n24661 , n24608 );
xor ( n24663 , n24609 , n24619 );
and ( n24664 , n24663 , n24512 );
or ( n24665 , n24662 , n24664 );
buf ( n24666 , n24665 );
not ( n24667 , n24666 );
buf ( n24668 , n24667 );
buf ( n24669 , n24668 );
not ( n24670 , n24669 );
buf ( n24671 , n24670 );
not ( n24672 , n24671 );
buf ( n24673 , n24672 );
not ( n24674 , n24512 );
and ( n24675 , n24674 , n24610 );
xor ( n24676 , n24611 , n24618 );
and ( n24677 , n24676 , n24512 );
or ( n24678 , n24675 , n24677 );
buf ( n24679 , n24678 );
not ( n24680 , n24679 );
buf ( n24681 , n24680 );
buf ( n24682 , n24681 );
not ( n24683 , n24682 );
buf ( n24684 , n24683 );
not ( n24685 , n24684 );
buf ( n24686 , n24685 );
not ( n24687 , n24512 );
and ( n24688 , n24687 , n24612 );
xor ( n24689 , n24613 , n24617 );
and ( n24690 , n24689 , n24512 );
or ( n24691 , n24688 , n24690 );
buf ( n24692 , n24691 );
not ( n24693 , n24692 );
buf ( n24694 , n24693 );
buf ( n24695 , n24694 );
not ( n24696 , n24695 );
buf ( n24697 , n24696 );
not ( n24698 , n24697 );
buf ( n24699 , n24698 );
not ( n24700 , n24512 );
and ( n24701 , n24700 , n24614 );
xor ( n24702 , n24615 , n24616 );
and ( n24703 , n24702 , n24512 );
or ( n24704 , n24701 , n24703 );
buf ( n24705 , n24704 );
not ( n24706 , n24705 );
buf ( n24707 , n24706 );
buf ( n24708 , n24707 );
not ( n24709 , n24708 );
buf ( n24710 , n24709 );
not ( n24711 , n24710 );
buf ( n24712 , n24711 );
not ( n24713 , n24596 );
buf ( n24714 , n24713 );
and ( n24715 , n24712 , n24714 );
and ( n24716 , n24699 , n24715 );
and ( n24717 , n24686 , n24716 );
and ( n24718 , n24673 , n24717 );
and ( n24719 , n24660 , n24718 );
and ( n24720 , n24647 , n24719 );
and ( n24721 , n24634 , n24720 );
not ( n24722 , n24721 );
buf ( n24723 , n24722 );
buf ( n24724 , n24512 );
and ( n24725 , n24723 , n24724 );
or ( n24726 , C0 , n24725 );
buf ( n24727 , n24726 );
buf ( n24728 , n24727 );
not ( n24729 , n24728 );
not ( n24730 , n24724 );
buf ( n24731 , n24710 );
and ( n24732 , n24730 , n24731 );
xor ( n24733 , n24712 , n24714 );
buf ( n24734 , n24733 );
and ( n24735 , n24734 , n24724 );
or ( n24736 , n24732 , n24735 );
buf ( n24737 , n24736 );
buf ( n24738 , n24737 );
and ( n24739 , n24729 , n24738 );
not ( n24740 , n24738 );
not ( n24741 , n24597 );
xor ( n24742 , n24740 , n24741 );
and ( n24743 , n24742 , n24728 );
or ( n24744 , n24739 , n24743 );
buf ( n24745 , n24744 );
not ( n24746 , n24745 );
buf ( n24747 , n24746 );
buf ( n24748 , n24747 );
not ( n24749 , n24748 );
or ( n24750 , n24602 , n24749 );
not ( n24751 , n24728 );
not ( n24752 , n24724 );
buf ( n24753 , n24697 );
and ( n24754 , n24752 , n24753 );
xor ( n24755 , n24699 , n24715 );
buf ( n24756 , n24755 );
and ( n24757 , n24756 , n24724 );
or ( n24758 , n24754 , n24757 );
buf ( n24759 , n24758 );
buf ( n24760 , n24759 );
and ( n24761 , n24751 , n24760 );
not ( n24762 , n24760 );
and ( n24763 , n24740 , n24741 );
xor ( n24764 , n24762 , n24763 );
and ( n24765 , n24764 , n24728 );
or ( n24766 , n24761 , n24765 );
buf ( n24767 , n24766 );
not ( n24768 , n24767 );
buf ( n24769 , n24768 );
buf ( n24770 , n24769 );
not ( n24771 , n24770 );
or ( n24772 , n24750 , n24771 );
buf ( n24773 , n24772 );
buf ( n24774 , n24773 );
and ( n24775 , n24774 , n24728 );
not ( n24776 , n24775 );
and ( n24777 , n24776 , n24602 );
xor ( n24778 , n24602 , n24728 );
xor ( n24779 , n24778 , n24728 );
and ( n24780 , n24779 , n24775 );
or ( n24781 , n24777 , n24780 );
buf ( n24782 , n24781 );
not ( n24783 , n24775 );
and ( n24784 , n24783 , n24749 );
xor ( n24785 , n24749 , n24728 );
and ( n24786 , n24778 , n24728 );
xor ( n24787 , n24785 , n24786 );
and ( n24788 , n24787 , n24775 );
or ( n24789 , n24784 , n24788 );
buf ( n24790 , n24789 );
not ( n24791 , n24775 );
and ( n24792 , n24791 , n24771 );
xor ( n24793 , n24771 , n24728 );
and ( n24794 , n24785 , n24786 );
xor ( n24795 , n24793 , n24794 );
and ( n24796 , n24795 , n24775 );
or ( n24797 , n24792 , n24796 );
buf ( n24798 , n24797 );
and ( n24799 , n24782 , n24790 , n24798 );
or ( n24800 , n24511 , n24799 );
not ( n24801 , n24800 );
buf ( n24802 , RI2107f4a8_454);
buf ( n24803 , n24061 );
not ( n24804 , n24803 );
buf ( n24805 , n24102 );
and ( n24806 , n24804 , n24805 );
not ( n24807 , n24805 );
buf ( n24808 , n24110 );
not ( n24809 , n24808 );
buf ( n24810 , n24118 );
not ( n24811 , n24810 );
buf ( n24812 , n24126 );
not ( n24813 , n24812 );
buf ( n24814 , n24134 );
not ( n24815 , n24814 );
buf ( n24816 , n24142 );
not ( n24817 , n24816 );
buf ( n24818 , n24150 );
not ( n24819 , n24818 );
buf ( n24820 , n24158 );
not ( n24821 , n24820 );
buf ( n24822 , n24166 );
not ( n24823 , n24822 );
buf ( n24824 , n24174 );
not ( n24825 , n24824 );
buf ( n24826 , n24182 );
not ( n24827 , n24826 );
buf ( n24828 , n24190 );
not ( n24829 , n24828 );
buf ( n24830 , n24198 );
not ( n24831 , n24830 );
buf ( n24832 , n24206 );
not ( n24833 , n24832 );
buf ( n24834 , n24214 );
not ( n24835 , n24834 );
buf ( n24836 , n24222 );
not ( n24837 , n24836 );
buf ( n24838 , n24230 );
not ( n24839 , n24838 );
buf ( n24840 , n24238 );
not ( n24841 , n24840 );
buf ( n24842 , n24246 );
not ( n24843 , n24842 );
buf ( n24844 , n24249 );
not ( n24845 , n24844 );
and ( n24846 , n24843 , n24845 );
and ( n24847 , n24841 , n24846 );
and ( n24848 , n24839 , n24847 );
and ( n24849 , n24837 , n24848 );
and ( n24850 , n24835 , n24849 );
and ( n24851 , n24833 , n24850 );
and ( n24852 , n24831 , n24851 );
and ( n24853 , n24829 , n24852 );
and ( n24854 , n24827 , n24853 );
and ( n24855 , n24825 , n24854 );
and ( n24856 , n24823 , n24855 );
and ( n24857 , n24821 , n24856 );
and ( n24858 , n24819 , n24857 );
and ( n24859 , n24817 , n24858 );
and ( n24860 , n24815 , n24859 );
and ( n24861 , n24813 , n24860 );
and ( n24862 , n24811 , n24861 );
and ( n24863 , n24809 , n24862 );
xor ( n24864 , n24807 , n24863 );
and ( n24865 , n24864 , n24803 );
or ( n24866 , n24806 , n24865 );
buf ( n24867 , n24866 );
not ( n24868 , n24867 );
buf ( n24869 , n24868 );
buf ( n24870 , n24869 );
not ( n24871 , n24870 );
buf ( n24872 , n24871 );
buf ( n24873 , n24872 );
buf ( n24874 , n24873 );
not ( n24875 , n24874 );
buf ( n24876 , n24875 );
buf ( n24877 , n24876 );
not ( n24878 , n24877 );
not ( n24879 , n24803 );
buf ( n24880 , n24325 );
not ( n24881 , n24880 );
buf ( n24882 , n24333 );
not ( n24883 , n24882 );
buf ( n24884 , n24341 );
not ( n24885 , n24884 );
buf ( n24886 , n24349 );
not ( n24887 , n24886 );
buf ( n24888 , n24357 );
not ( n24889 , n24888 );
buf ( n24890 , n24365 );
not ( n24891 , n24890 );
buf ( n24892 , n24373 );
not ( n24893 , n24892 );
buf ( n24894 , n24069 );
not ( n24895 , n24894 );
buf ( n24896 , n24078 );
not ( n24897 , n24896 );
buf ( n24898 , n24086 );
not ( n24899 , n24898 );
buf ( n24900 , n24094 );
not ( n24901 , n24900 );
and ( n24902 , n24807 , n24863 );
and ( n24903 , n24901 , n24902 );
and ( n24904 , n24899 , n24903 );
and ( n24905 , n24897 , n24904 );
and ( n24906 , n24895 , n24905 );
and ( n24907 , n24893 , n24906 );
and ( n24908 , n24891 , n24907 );
and ( n24909 , n24889 , n24908 );
and ( n24910 , n24887 , n24909 );
and ( n24911 , n24885 , n24910 );
and ( n24912 , n24883 , n24911 );
and ( n24913 , n24881 , n24912 );
xor ( n24914 , n24879 , n24913 );
buf ( n24915 , n24803 );
and ( n24916 , n24914 , n24915 );
or ( n24917 , C0 , n24916 );
buf ( n24918 , n24917 );
not ( n24919 , n24918 );
buf ( n24920 , n24919 );
buf ( n24921 , n24920 );
not ( n24922 , n24921 );
buf ( n24923 , n24922 );
not ( n24924 , n24923 );
buf ( n24925 , n24924 );
not ( n24926 , n24803 );
and ( n24927 , n24926 , n24880 );
xor ( n24928 , n24881 , n24912 );
and ( n24929 , n24928 , n24803 );
or ( n24930 , n24927 , n24929 );
buf ( n24931 , n24930 );
not ( n24932 , n24931 );
buf ( n24933 , n24932 );
buf ( n24934 , n24933 );
not ( n24935 , n24934 );
buf ( n24936 , n24935 );
not ( n24937 , n24936 );
buf ( n24938 , n24937 );
not ( n24939 , n24803 );
and ( n24940 , n24939 , n24882 );
xor ( n24941 , n24883 , n24911 );
and ( n24942 , n24941 , n24803 );
or ( n24943 , n24940 , n24942 );
buf ( n24944 , n24943 );
not ( n24945 , n24944 );
buf ( n24946 , n24945 );
buf ( n24947 , n24946 );
not ( n24948 , n24947 );
buf ( n24949 , n24948 );
not ( n24950 , n24949 );
buf ( n24951 , n24950 );
not ( n24952 , n24803 );
and ( n24953 , n24952 , n24884 );
xor ( n24954 , n24885 , n24910 );
and ( n24955 , n24954 , n24803 );
or ( n24956 , n24953 , n24955 );
buf ( n24957 , n24956 );
not ( n24958 , n24957 );
buf ( n24959 , n24958 );
buf ( n24960 , n24959 );
not ( n24961 , n24960 );
buf ( n24962 , n24961 );
not ( n24963 , n24962 );
buf ( n24964 , n24963 );
not ( n24965 , n24803 );
and ( n24966 , n24965 , n24886 );
xor ( n24967 , n24887 , n24909 );
and ( n24968 , n24967 , n24803 );
or ( n24969 , n24966 , n24968 );
buf ( n24970 , n24969 );
not ( n24971 , n24970 );
buf ( n24972 , n24971 );
buf ( n24973 , n24972 );
not ( n24974 , n24973 );
buf ( n24975 , n24974 );
not ( n24976 , n24975 );
buf ( n24977 , n24976 );
not ( n24978 , n24803 );
and ( n24979 , n24978 , n24888 );
xor ( n24980 , n24889 , n24908 );
and ( n24981 , n24980 , n24803 );
or ( n24982 , n24979 , n24981 );
buf ( n24983 , n24982 );
not ( n24984 , n24983 );
buf ( n24985 , n24984 );
buf ( n24986 , n24985 );
not ( n24987 , n24986 );
buf ( n24988 , n24987 );
not ( n24989 , n24988 );
buf ( n24990 , n24989 );
not ( n24991 , n24803 );
and ( n24992 , n24991 , n24890 );
xor ( n24993 , n24891 , n24907 );
and ( n24994 , n24993 , n24803 );
or ( n24995 , n24992 , n24994 );
buf ( n24996 , n24995 );
not ( n24997 , n24996 );
buf ( n24998 , n24997 );
buf ( n24999 , n24998 );
not ( n25000 , n24999 );
buf ( n25001 , n25000 );
not ( n25002 , n25001 );
buf ( n25003 , n25002 );
not ( n25004 , n24803 );
and ( n25005 , n25004 , n24892 );
xor ( n25006 , n24893 , n24906 );
and ( n25007 , n25006 , n24803 );
or ( n25008 , n25005 , n25007 );
buf ( n25009 , n25008 );
not ( n25010 , n25009 );
buf ( n25011 , n25010 );
buf ( n25012 , n25011 );
not ( n25013 , n25012 );
buf ( n25014 , n25013 );
not ( n25015 , n25014 );
buf ( n25016 , n25015 );
not ( n25017 , n24803 );
and ( n25018 , n25017 , n24894 );
xor ( n25019 , n24895 , n24905 );
and ( n25020 , n25019 , n24803 );
or ( n25021 , n25018 , n25020 );
buf ( n25022 , n25021 );
not ( n25023 , n25022 );
buf ( n25024 , n25023 );
buf ( n25025 , n25024 );
not ( n25026 , n25025 );
buf ( n25027 , n25026 );
not ( n25028 , n25027 );
buf ( n25029 , n25028 );
not ( n25030 , n24803 );
and ( n25031 , n25030 , n24896 );
xor ( n25032 , n24897 , n24904 );
and ( n25033 , n25032 , n24803 );
or ( n25034 , n25031 , n25033 );
buf ( n25035 , n25034 );
not ( n25036 , n25035 );
buf ( n25037 , n25036 );
buf ( n25038 , n25037 );
not ( n25039 , n25038 );
buf ( n25040 , n25039 );
not ( n25041 , n25040 );
buf ( n25042 , n25041 );
not ( n25043 , n24803 );
and ( n25044 , n25043 , n24898 );
xor ( n25045 , n24899 , n24903 );
and ( n25046 , n25045 , n24803 );
or ( n25047 , n25044 , n25046 );
buf ( n25048 , n25047 );
not ( n25049 , n25048 );
buf ( n25050 , n25049 );
buf ( n25051 , n25050 );
not ( n25052 , n25051 );
buf ( n25053 , n25052 );
not ( n25054 , n25053 );
buf ( n25055 , n25054 );
not ( n25056 , n24803 );
and ( n25057 , n25056 , n24900 );
xor ( n25058 , n24901 , n24902 );
and ( n25059 , n25058 , n24803 );
or ( n25060 , n25057 , n25059 );
buf ( n25061 , n25060 );
not ( n25062 , n25061 );
buf ( n25063 , n25062 );
buf ( n25064 , n25063 );
not ( n25065 , n25064 );
buf ( n25066 , n25065 );
not ( n25067 , n25066 );
buf ( n25068 , n25067 );
not ( n25069 , n24872 );
buf ( n25070 , n25069 );
and ( n25071 , n25068 , n25070 );
and ( n25072 , n25055 , n25071 );
and ( n25073 , n25042 , n25072 );
and ( n25074 , n25029 , n25073 );
and ( n25075 , n25016 , n25074 );
and ( n25076 , n25003 , n25075 );
and ( n25077 , n24990 , n25076 );
and ( n25078 , n24977 , n25077 );
and ( n25079 , n24964 , n25078 );
and ( n25080 , n24951 , n25079 );
and ( n25081 , n24938 , n25080 );
and ( n25082 , n24925 , n25081 );
not ( n25083 , n25082 );
buf ( n25084 , n25083 );
buf ( n25085 , n24803 );
and ( n25086 , n25084 , n25085 );
or ( n25087 , C0 , n25086 );
buf ( n25088 , n25087 );
buf ( n25089 , n25088 );
not ( n25090 , n25089 );
not ( n25091 , n25085 );
buf ( n25092 , n25066 );
and ( n25093 , n25091 , n25092 );
xor ( n25094 , n25068 , n25070 );
buf ( n25095 , n25094 );
and ( n25096 , n25095 , n25085 );
or ( n25097 , n25093 , n25096 );
buf ( n25098 , n25097 );
buf ( n25099 , n25098 );
and ( n25100 , n25090 , n25099 );
not ( n25101 , n25099 );
not ( n25102 , n24873 );
xor ( n25103 , n25101 , n25102 );
and ( n25104 , n25103 , n25089 );
or ( n25105 , n25100 , n25104 );
buf ( n25106 , n25105 );
not ( n25107 , n25106 );
buf ( n25108 , n25107 );
buf ( n25109 , n25108 );
not ( n25110 , n25109 );
or ( n25111 , n24878 , n25110 );
not ( n25112 , n25089 );
not ( n25113 , n25085 );
buf ( n25114 , n25053 );
and ( n25115 , n25113 , n25114 );
xor ( n25116 , n25055 , n25071 );
buf ( n25117 , n25116 );
and ( n25118 , n25117 , n25085 );
or ( n25119 , n25115 , n25118 );
buf ( n25120 , n25119 );
buf ( n25121 , n25120 );
and ( n25122 , n25112 , n25121 );
not ( n25123 , n25121 );
and ( n25124 , n25101 , n25102 );
xor ( n25125 , n25123 , n25124 );
and ( n25126 , n25125 , n25089 );
or ( n25127 , n25122 , n25126 );
buf ( n25128 , n25127 );
not ( n25129 , n25128 );
buf ( n25130 , n25129 );
buf ( n25131 , n25130 );
not ( n25132 , n25131 );
or ( n25133 , n25111 , n25132 );
not ( n25134 , n25089 );
not ( n25135 , n25085 );
buf ( n25136 , n25040 );
and ( n25137 , n25135 , n25136 );
xor ( n25138 , n25042 , n25072 );
buf ( n25139 , n25138 );
and ( n25140 , n25139 , n25085 );
or ( n25141 , n25137 , n25140 );
buf ( n25142 , n25141 );
buf ( n25143 , n25142 );
and ( n25144 , n25134 , n25143 );
not ( n25145 , n25143 );
and ( n25146 , n25123 , n25124 );
xor ( n25147 , n25145 , n25146 );
and ( n25148 , n25147 , n25089 );
or ( n25149 , n25144 , n25148 );
buf ( n25150 , n25149 );
not ( n25151 , n25150 );
buf ( n25152 , n25151 );
buf ( n25153 , n25152 );
not ( n25154 , n25153 );
or ( n25155 , n25133 , n25154 );
or ( n25156 , n25155 , C0 );
or ( n25157 , n25156 , C0 );
or ( n25158 , n25157 , C0 );
or ( n25159 , n25158 , C0 );
or ( n25160 , n25159 , C0 );
or ( n25161 , n25160 , C0 );
or ( n25162 , n25161 , C0 );
or ( n25163 , n25162 , C0 );
or ( n25164 , n25163 , C0 );
or ( n25165 , n25164 , C0 );
or ( n25166 , n25165 , C0 );
or ( n25167 , n25166 , C0 );
or ( n25168 , n25167 , C0 );
or ( n25169 , n25168 , C0 );
or ( n25170 , n25169 , C0 );
or ( n25171 , n25170 , C0 );
or ( n25172 , n25171 , C0 );
or ( n25173 , n25172 , C0 );
or ( n25174 , n25173 , C0 );
or ( n25175 , n25174 , C0 );
or ( n25176 , n25175 , C0 );
or ( n25177 , n25176 , C0 );
or ( n25178 , n25177 , C0 );
or ( n25179 , n25178 , C0 );
or ( n25180 , n25179 , C0 );
or ( n25181 , n25180 , C0 );
or ( n25182 , n25181 , C0 );
buf ( n25183 , n25182 );
and ( n25184 , n25183 , n25089 );
not ( n25185 , n25184 );
and ( n25186 , n25185 , n24878 );
xor ( n25187 , n24878 , n25089 );
xor ( n25188 , n25187 , n25089 );
and ( n25189 , n25188 , n25184 );
or ( n25190 , n25186 , n25189 );
buf ( n25191 , n25190 );
not ( n25192 , n25184 );
and ( n25193 , n25192 , n25110 );
xor ( n25194 , n25110 , n25089 );
and ( n25195 , n25187 , n25089 );
xor ( n25196 , n25194 , n25195 );
and ( n25197 , n25196 , n25184 );
or ( n25198 , n25193 , n25197 );
buf ( n25199 , n25198 );
not ( n25200 , n25199 );
not ( n25201 , n25184 );
and ( n25202 , n25201 , n25132 );
xor ( n25203 , n25132 , n25089 );
and ( n25204 , n25194 , n25195 );
xor ( n25205 , n25203 , n25204 );
and ( n25206 , n25205 , n25184 );
or ( n25207 , n25202 , n25206 );
buf ( n25208 , n25207 );
not ( n25209 , n25184 );
and ( n25210 , n25209 , n25154 );
xor ( n25211 , n25154 , n25089 );
and ( n25212 , n25203 , n25204 );
xor ( n25213 , n25211 , n25212 );
and ( n25214 , n25213 , n25184 );
or ( n25215 , n25210 , n25214 );
buf ( n25216 , n25215 );
and ( n25217 , n25191 , n25200 , n25208 , n25216 );
not ( n25218 , n25191 );
and ( n25219 , n25218 , n25199 , n25208 , n25216 );
or ( n25220 , n25217 , n25219 );
and ( n25221 , n25191 , n25199 , n25208 , n25216 );
or ( n25222 , n25220 , n25221 );
and ( n25223 , n24802 , n25222 );
buf ( n25224 , RI210aeb90_395);
buf ( n25225 , n25224 );
buf ( n25226 , n25225 );
not ( n25227 , n25226 );
buf ( n25228 , n25227 );
buf ( n25229 , n25228 );
not ( n25230 , n25229 );
buf ( n25231 , GI20471ac0_434);
buf ( n25232 , n25231 );
not ( n25233 , n25232 );
buf ( n25234 , RI2107f340_457);
buf ( n25235 , n25234 );
and ( n25236 , n25233 , n25235 );
not ( n25237 , n25235 );
not ( n25238 , n25225 );
xor ( n25239 , n25237 , n25238 );
and ( n25240 , n25239 , n25232 );
or ( n25241 , n25236 , n25240 );
buf ( n25242 , n25241 );
not ( n25243 , n25242 );
buf ( n25244 , n25243 );
buf ( n25245 , n25244 );
not ( n25246 , n25245 );
or ( n25247 , n25230 , n25246 );
not ( n25248 , n25232 );
buf ( n25249 , RI2107e878_458);
buf ( n25250 , n25249 );
and ( n25251 , n25248 , n25250 );
not ( n25252 , n25250 );
and ( n25253 , n25237 , n25238 );
xor ( n25254 , n25252 , n25253 );
and ( n25255 , n25254 , n25232 );
or ( n25256 , n25251 , n25255 );
buf ( n25257 , n25256 );
not ( n25258 , n25257 );
buf ( n25259 , n25258 );
buf ( n25260 , n25259 );
not ( n25261 , n25260 );
or ( n25262 , n25247 , n25261 );
not ( n25263 , n25232 );
buf ( n25264 , RI21084f20_415);
buf ( n25265 , n25264 );
and ( n25266 , n25263 , n25265 );
not ( n25267 , n25265 );
and ( n25268 , n25252 , n25253 );
xor ( n25269 , n25267 , n25268 );
and ( n25270 , n25269 , n25232 );
or ( n25271 , n25266 , n25270 );
buf ( n25272 , n25271 );
not ( n25273 , n25272 );
buf ( n25274 , n25273 );
buf ( n25275 , n25274 );
not ( n25276 , n25275 );
or ( n25277 , n25262 , n25276 );
not ( n25278 , n25232 );
buf ( n25279 , RI21084458_416);
buf ( n25280 , n25279 );
and ( n25281 , n25278 , n25280 );
not ( n25282 , n25280 );
and ( n25283 , n25267 , n25268 );
xor ( n25284 , n25282 , n25283 );
and ( n25285 , n25284 , n25232 );
or ( n25286 , n25281 , n25285 );
buf ( n25287 , n25286 );
not ( n25288 , n25287 );
buf ( n25289 , n25288 );
buf ( n25290 , n25289 );
not ( n25291 , n25290 );
or ( n25292 , n25277 , n25291 );
not ( n25293 , n25232 );
buf ( n25294 , RI2107e800_459);
buf ( n25295 , n25294 );
and ( n25296 , n25293 , n25295 );
not ( n25297 , n25295 );
and ( n25298 , n25282 , n25283 );
xor ( n25299 , n25297 , n25298 );
and ( n25300 , n25299 , n25232 );
or ( n25301 , n25296 , n25300 );
buf ( n25302 , n25301 );
not ( n25303 , n25302 );
buf ( n25304 , n25303 );
buf ( n25305 , n25304 );
not ( n25306 , n25305 );
or ( n25307 , n25292 , n25306 );
not ( n25308 , n25232 );
buf ( n25309 , RI2107e788_460);
buf ( n25310 , n25309 );
and ( n25311 , n25308 , n25310 );
not ( n25312 , n25310 );
and ( n25313 , n25297 , n25298 );
xor ( n25314 , n25312 , n25313 );
and ( n25315 , n25314 , n25232 );
or ( n25316 , n25311 , n25315 );
buf ( n25317 , n25316 );
not ( n25318 , n25317 );
buf ( n25319 , n25318 );
buf ( n25320 , n25319 );
not ( n25321 , n25320 );
or ( n25322 , n25307 , n25321 );
not ( n25323 , n25232 );
buf ( n25324 , RI2107e710_461);
buf ( n25325 , n25324 );
and ( n25326 , n25323 , n25325 );
not ( n25327 , n25325 );
and ( n25328 , n25312 , n25313 );
xor ( n25329 , n25327 , n25328 );
and ( n25330 , n25329 , n25232 );
or ( n25331 , n25326 , n25330 );
buf ( n25332 , n25331 );
not ( n25333 , n25332 );
buf ( n25334 , n25333 );
buf ( n25335 , n25334 );
not ( n25336 , n25335 );
or ( n25337 , n25322 , n25336 );
not ( n25338 , n25232 );
buf ( n25339 , RI2107e698_462);
buf ( n25340 , n25339 );
and ( n25341 , n25338 , n25340 );
not ( n25342 , n25340 );
and ( n25343 , n25327 , n25328 );
xor ( n25344 , n25342 , n25343 );
and ( n25345 , n25344 , n25232 );
or ( n25346 , n25341 , n25345 );
buf ( n25347 , n25346 );
not ( n25348 , n25347 );
buf ( n25349 , n25348 );
buf ( n25350 , n25349 );
not ( n25351 , n25350 );
or ( n25352 , n25337 , n25351 );
not ( n25353 , n25232 );
buf ( n25354 , RI210843e0_417);
buf ( n25355 , n25354 );
and ( n25356 , n25353 , n25355 );
not ( n25357 , n25355 );
and ( n25358 , n25342 , n25343 );
xor ( n25359 , n25357 , n25358 );
and ( n25360 , n25359 , n25232 );
or ( n25361 , n25356 , n25360 );
buf ( n25362 , n25361 );
not ( n25363 , n25362 );
buf ( n25364 , n25363 );
buf ( n25365 , n25364 );
not ( n25366 , n25365 );
or ( n25367 , n25352 , n25366 );
not ( n25368 , n25232 );
buf ( n25369 , RI210a63a0_396);
buf ( n25370 , n25369 );
and ( n25371 , n25368 , n25370 );
not ( n25372 , n25370 );
and ( n25373 , n25357 , n25358 );
xor ( n25374 , n25372 , n25373 );
and ( n25375 , n25374 , n25232 );
or ( n25376 , n25371 , n25375 );
buf ( n25377 , n25376 );
not ( n25378 , n25377 );
buf ( n25379 , n25378 );
buf ( n25380 , n25379 );
not ( n25381 , n25380 );
or ( n25382 , n25367 , n25381 );
not ( n25383 , n25232 );
buf ( n25384 , RI21086e10_397);
buf ( n25385 , n25384 );
and ( n25386 , n25383 , n25385 );
not ( n25387 , n25385 );
and ( n25388 , n25372 , n25373 );
xor ( n25389 , n25387 , n25388 );
and ( n25390 , n25389 , n25232 );
or ( n25391 , n25386 , n25390 );
buf ( n25392 , n25391 );
not ( n25393 , n25392 );
buf ( n25394 , n25393 );
buf ( n25395 , n25394 );
not ( n25396 , n25395 );
or ( n25397 , n25382 , n25396 );
not ( n25398 , n25232 );
buf ( n25399 , RI21086bb8_398);
buf ( n25400 , n25399 );
and ( n25401 , n25398 , n25400 );
not ( n25402 , n25400 );
and ( n25403 , n25387 , n25388 );
xor ( n25404 , n25402 , n25403 );
and ( n25405 , n25404 , n25232 );
or ( n25406 , n25401 , n25405 );
buf ( n25407 , n25406 );
not ( n25408 , n25407 );
buf ( n25409 , n25408 );
buf ( n25410 , n25409 );
not ( n25411 , n25410 );
or ( n25412 , n25397 , n25411 );
not ( n25413 , n25232 );
buf ( n25414 , RI21086b40_399);
buf ( n25415 , n25414 );
and ( n25416 , n25413 , n25415 );
not ( n25417 , n25415 );
and ( n25418 , n25402 , n25403 );
xor ( n25419 , n25417 , n25418 );
and ( n25420 , n25419 , n25232 );
or ( n25421 , n25416 , n25420 );
buf ( n25422 , n25421 );
not ( n25423 , n25422 );
buf ( n25424 , n25423 );
buf ( n25425 , n25424 );
not ( n25426 , n25425 );
or ( n25427 , n25412 , n25426 );
not ( n25428 , n25232 );
buf ( n25429 , RI21086ac8_400);
buf ( n25430 , n25429 );
and ( n25431 , n25428 , n25430 );
not ( n25432 , n25430 );
and ( n25433 , n25417 , n25418 );
xor ( n25434 , n25432 , n25433 );
and ( n25435 , n25434 , n25232 );
or ( n25436 , n25431 , n25435 );
buf ( n25437 , n25436 );
not ( n25438 , n25437 );
buf ( n25439 , n25438 );
buf ( n25440 , n25439 );
not ( n25441 , n25440 );
or ( n25442 , n25427 , n25441 );
not ( n25443 , n25232 );
buf ( n25444 , RI21086a50_401);
buf ( n25445 , n25444 );
and ( n25446 , n25443 , n25445 );
not ( n25447 , n25445 );
and ( n25448 , n25432 , n25433 );
xor ( n25449 , n25447 , n25448 );
and ( n25450 , n25449 , n25232 );
or ( n25451 , n25446 , n25450 );
buf ( n25452 , n25451 );
not ( n25453 , n25452 );
buf ( n25454 , n25453 );
buf ( n25455 , n25454 );
not ( n25456 , n25455 );
or ( n25457 , n25442 , n25456 );
not ( n25458 , n25232 );
buf ( n25459 , RI210869d8_402);
buf ( n25460 , n25459 );
and ( n25461 , n25458 , n25460 );
not ( n25462 , n25460 );
and ( n25463 , n25447 , n25448 );
xor ( n25464 , n25462 , n25463 );
and ( n25465 , n25464 , n25232 );
or ( n25466 , n25461 , n25465 );
buf ( n25467 , n25466 );
not ( n25468 , n25467 );
buf ( n25469 , n25468 );
buf ( n25470 , n25469 );
not ( n25471 , n25470 );
or ( n25472 , n25457 , n25471 );
not ( n25473 , n25232 );
buf ( n25474 , RI21086960_403);
buf ( n25475 , n25474 );
and ( n25476 , n25473 , n25475 );
not ( n25477 , n25475 );
and ( n25478 , n25462 , n25463 );
xor ( n25479 , n25477 , n25478 );
and ( n25480 , n25479 , n25232 );
or ( n25481 , n25476 , n25480 );
buf ( n25482 , n25481 );
not ( n25483 , n25482 );
buf ( n25484 , n25483 );
buf ( n25485 , n25484 );
not ( n25486 , n25485 );
or ( n25487 , n25472 , n25486 );
not ( n25488 , n25232 );
buf ( n25489 , RI21085e98_404);
buf ( n25490 , n25489 );
and ( n25491 , n25488 , n25490 );
not ( n25492 , n25490 );
and ( n25493 , n25477 , n25478 );
xor ( n25494 , n25492 , n25493 );
and ( n25495 , n25494 , n25232 );
or ( n25496 , n25491 , n25495 );
buf ( n25497 , n25496 );
not ( n25498 , n25497 );
buf ( n25499 , n25498 );
buf ( n25500 , n25499 );
not ( n25501 , n25500 );
or ( n25502 , n25487 , n25501 );
not ( n25503 , n25232 );
buf ( n25504 , RI21085e20_405);
buf ( n25505 , n25504 );
and ( n25506 , n25503 , n25505 );
not ( n25507 , n25505 );
and ( n25508 , n25492 , n25493 );
xor ( n25509 , n25507 , n25508 );
and ( n25510 , n25509 , n25232 );
or ( n25511 , n25506 , n25510 );
buf ( n25512 , n25511 );
not ( n25513 , n25512 );
buf ( n25514 , n25513 );
buf ( n25515 , n25514 );
not ( n25516 , n25515 );
or ( n25517 , n25502 , n25516 );
not ( n25518 , n25232 );
buf ( n25519 , RI21085da8_406);
buf ( n25520 , n25519 );
and ( n25521 , n25518 , n25520 );
not ( n25522 , n25520 );
and ( n25523 , n25507 , n25508 );
xor ( n25524 , n25522 , n25523 );
and ( n25525 , n25524 , n25232 );
or ( n25526 , n25521 , n25525 );
buf ( n25527 , n25526 );
not ( n25528 , n25527 );
buf ( n25529 , n25528 );
buf ( n25530 , n25529 );
not ( n25531 , n25530 );
or ( n25532 , n25517 , n25531 );
not ( n25533 , n25232 );
buf ( n25534 , RI21085d30_407);
buf ( n25535 , n25534 );
and ( n25536 , n25533 , n25535 );
not ( n25537 , n25535 );
and ( n25538 , n25522 , n25523 );
xor ( n25539 , n25537 , n25538 );
and ( n25540 , n25539 , n25232 );
or ( n25541 , n25536 , n25540 );
buf ( n25542 , n25541 );
not ( n25543 , n25542 );
buf ( n25544 , n25543 );
buf ( n25545 , n25544 );
not ( n25546 , n25545 );
or ( n25547 , n25532 , n25546 );
not ( n25548 , n25232 );
buf ( n25549 , RI21085cb8_408);
buf ( n25550 , n25549 );
and ( n25551 , n25548 , n25550 );
not ( n25552 , n25550 );
and ( n25553 , n25537 , n25538 );
xor ( n25554 , n25552 , n25553 );
and ( n25555 , n25554 , n25232 );
or ( n25556 , n25551 , n25555 );
buf ( n25557 , n25556 );
not ( n25558 , n25557 );
buf ( n25559 , n25558 );
buf ( n25560 , n25559 );
not ( n25561 , n25560 );
or ( n25562 , n25547 , n25561 );
not ( n25563 , n25232 );
buf ( n25564 , RI21085c40_409);
buf ( n25565 , n25564 );
and ( n25566 , n25563 , n25565 );
not ( n25567 , n25565 );
and ( n25568 , n25552 , n25553 );
xor ( n25569 , n25567 , n25568 );
and ( n25570 , n25569 , n25232 );
or ( n25571 , n25566 , n25570 );
buf ( n25572 , n25571 );
not ( n25573 , n25572 );
buf ( n25574 , n25573 );
buf ( n25575 , n25574 );
not ( n25576 , n25575 );
or ( n25577 , n25562 , n25576 );
not ( n25578 , n25232 );
buf ( n25579 , RI21085178_410);
buf ( n25580 , n25579 );
and ( n25581 , n25578 , n25580 );
not ( n25582 , n25580 );
and ( n25583 , n25567 , n25568 );
xor ( n25584 , n25582 , n25583 );
and ( n25585 , n25584 , n25232 );
or ( n25586 , n25581 , n25585 );
buf ( n25587 , n25586 );
not ( n25588 , n25587 );
buf ( n25589 , n25588 );
buf ( n25590 , n25589 );
not ( n25591 , n25590 );
or ( n25592 , n25577 , n25591 );
not ( n25593 , n25232 );
buf ( n25594 , RI21085100_411);
buf ( n25595 , n25594 );
and ( n25596 , n25593 , n25595 );
not ( n25597 , n25595 );
and ( n25598 , n25582 , n25583 );
xor ( n25599 , n25597 , n25598 );
and ( n25600 , n25599 , n25232 );
or ( n25601 , n25596 , n25600 );
buf ( n25602 , n25601 );
not ( n25603 , n25602 );
buf ( n25604 , n25603 );
buf ( n25605 , n25604 );
not ( n25606 , n25605 );
or ( n25607 , n25592 , n25606 );
not ( n25608 , n25232 );
buf ( n25609 , RI21085088_412);
buf ( n25610 , n25609 );
and ( n25611 , n25608 , n25610 );
not ( n25612 , n25610 );
and ( n25613 , n25597 , n25598 );
xor ( n25614 , n25612 , n25613 );
and ( n25615 , n25614 , n25232 );
or ( n25616 , n25611 , n25615 );
buf ( n25617 , n25616 );
not ( n25618 , n25617 );
buf ( n25619 , n25618 );
buf ( n25620 , n25619 );
not ( n25621 , n25620 );
or ( n25622 , n25607 , n25621 );
not ( n25623 , n25232 );
buf ( n25624 , RI21085010_413);
buf ( n25625 , n25624 );
and ( n25626 , n25623 , n25625 );
not ( n25627 , n25625 );
and ( n25628 , n25612 , n25613 );
xor ( n25629 , n25627 , n25628 );
and ( n25630 , n25629 , n25232 );
or ( n25631 , n25626 , n25630 );
buf ( n25632 , n25631 );
not ( n25633 , n25632 );
buf ( n25634 , n25633 );
buf ( n25635 , n25634 );
not ( n25636 , n25635 );
or ( n25637 , n25622 , n25636 );
not ( n25638 , n25232 );
buf ( n25639 , RI21084f98_414);
buf ( n25640 , n25639 );
and ( n25641 , n25638 , n25640 );
not ( n25642 , n25640 );
and ( n25643 , n25627 , n25628 );
xor ( n25644 , n25642 , n25643 );
and ( n25645 , n25644 , n25232 );
or ( n25646 , n25641 , n25645 );
buf ( n25647 , n25646 );
not ( n25648 , n25647 );
buf ( n25649 , n25648 );
buf ( n25650 , n25649 );
not ( n25651 , n25650 );
or ( n25652 , n25637 , n25651 );
buf ( n25653 , n25652 );
buf ( n25654 , n25653 );
and ( n25655 , n25654 , n25232 );
not ( n25656 , n25655 );
and ( n25657 , n25656 , n25230 );
xor ( n25658 , n25230 , n25232 );
xor ( n25659 , n25658 , n25232 );
and ( n25660 , n25659 , n25655 );
or ( n25661 , n25657 , n25660 );
buf ( n25662 , n25661 );
buf ( n25663 , n25662 );
buf ( n25664 , n24061 );
not ( n25665 , n25664 );
buf ( n25666 , n24333 );
and ( n25667 , n25665 , n25666 );
not ( n25668 , n25666 );
buf ( n25669 , n24341 );
not ( n25670 , n25669 );
buf ( n25671 , n24349 );
not ( n25672 , n25671 );
buf ( n25673 , n24357 );
not ( n25674 , n25673 );
buf ( n25675 , n24365 );
not ( n25676 , n25675 );
buf ( n25677 , n24373 );
not ( n25678 , n25677 );
buf ( n25679 , n24069 );
not ( n25680 , n25679 );
buf ( n25681 , n24078 );
not ( n25682 , n25681 );
buf ( n25683 , n24086 );
not ( n25684 , n25683 );
buf ( n25685 , n24094 );
not ( n25686 , n25685 );
buf ( n25687 , n24102 );
not ( n25688 , n25687 );
buf ( n25689 , n24110 );
not ( n25690 , n25689 );
buf ( n25691 , n24118 );
not ( n25692 , n25691 );
buf ( n25693 , n24126 );
not ( n25694 , n25693 );
buf ( n25695 , n24134 );
not ( n25696 , n25695 );
buf ( n25697 , n24142 );
not ( n25698 , n25697 );
buf ( n25699 , n24150 );
not ( n25700 , n25699 );
buf ( n25701 , n24158 );
not ( n25702 , n25701 );
buf ( n25703 , n24166 );
not ( n25704 , n25703 );
buf ( n25705 , n24174 );
not ( n25706 , n25705 );
buf ( n25707 , n24182 );
not ( n25708 , n25707 );
buf ( n25709 , n24190 );
not ( n25710 , n25709 );
buf ( n25711 , n24198 );
not ( n25712 , n25711 );
buf ( n25713 , n24206 );
not ( n25714 , n25713 );
buf ( n25715 , n24214 );
not ( n25716 , n25715 );
buf ( n25717 , n24222 );
not ( n25718 , n25717 );
buf ( n25719 , n24230 );
not ( n25720 , n25719 );
buf ( n25721 , n24238 );
not ( n25722 , n25721 );
buf ( n25723 , n24246 );
not ( n25724 , n25723 );
buf ( n25725 , n24249 );
not ( n25726 , n25725 );
and ( n25727 , n25724 , n25726 );
and ( n25728 , n25722 , n25727 );
and ( n25729 , n25720 , n25728 );
and ( n25730 , n25718 , n25729 );
and ( n25731 , n25716 , n25730 );
and ( n25732 , n25714 , n25731 );
and ( n25733 , n25712 , n25732 );
and ( n25734 , n25710 , n25733 );
and ( n25735 , n25708 , n25734 );
and ( n25736 , n25706 , n25735 );
and ( n25737 , n25704 , n25736 );
and ( n25738 , n25702 , n25737 );
and ( n25739 , n25700 , n25738 );
and ( n25740 , n25698 , n25739 );
and ( n25741 , n25696 , n25740 );
and ( n25742 , n25694 , n25741 );
and ( n25743 , n25692 , n25742 );
and ( n25744 , n25690 , n25743 );
and ( n25745 , n25688 , n25744 );
and ( n25746 , n25686 , n25745 );
and ( n25747 , n25684 , n25746 );
and ( n25748 , n25682 , n25747 );
and ( n25749 , n25680 , n25748 );
and ( n25750 , n25678 , n25749 );
and ( n25751 , n25676 , n25750 );
and ( n25752 , n25674 , n25751 );
and ( n25753 , n25672 , n25752 );
and ( n25754 , n25670 , n25753 );
xor ( n25755 , n25668 , n25754 );
and ( n25756 , n25755 , n25664 );
or ( n25757 , n25667 , n25756 );
buf ( n25758 , n25757 );
not ( n25759 , n25758 );
buf ( n25760 , n25759 );
buf ( n25761 , n25760 );
not ( n25762 , n25761 );
buf ( n25763 , n25762 );
buf ( n25764 , n25763 );
buf ( n25765 , n25764 );
not ( n25766 , n25765 );
buf ( n25767 , n25766 );
buf ( n25768 , n25767 );
not ( n25769 , n25768 );
not ( n25770 , n25664 );
buf ( n25771 , n24325 );
not ( n25772 , n25771 );
and ( n25773 , n25668 , n25754 );
and ( n25774 , n25772 , n25773 );
xor ( n25775 , n25770 , n25774 );
buf ( n25776 , n25664 );
and ( n25777 , n25775 , n25776 );
or ( n25778 , C0 , n25777 );
buf ( n25779 , n25778 );
not ( n25780 , n25779 );
buf ( n25781 , n25780 );
buf ( n25782 , n25781 );
not ( n25783 , n25782 );
buf ( n25784 , n25783 );
not ( n25785 , n25784 );
buf ( n25786 , n25785 );
not ( n25787 , n25664 );
and ( n25788 , n25787 , n25771 );
xor ( n25789 , n25772 , n25773 );
and ( n25790 , n25789 , n25664 );
or ( n25791 , n25788 , n25790 );
buf ( n25792 , n25791 );
not ( n25793 , n25792 );
buf ( n25794 , n25793 );
buf ( n25795 , n25794 );
not ( n25796 , n25795 );
buf ( n25797 , n25796 );
not ( n25798 , n25797 );
buf ( n25799 , n25798 );
not ( n25800 , n25763 );
buf ( n25801 , n25800 );
and ( n25802 , n25799 , n25801 );
and ( n25803 , n25786 , n25802 );
not ( n25804 , n25803 );
buf ( n25805 , n25804 );
buf ( n25806 , n25664 );
and ( n25807 , n25805 , n25806 );
or ( n25808 , C0 , n25807 );
buf ( n25809 , n25808 );
buf ( n25810 , n25809 );
not ( n25811 , n25810 );
not ( n25812 , n25806 );
buf ( n25813 , n25797 );
and ( n25814 , n25812 , n25813 );
xor ( n25815 , n25799 , n25801 );
buf ( n25816 , n25815 );
and ( n25817 , n25816 , n25806 );
or ( n25818 , n25814 , n25817 );
buf ( n25819 , n25818 );
buf ( n25820 , n25819 );
and ( n25821 , n25811 , n25820 );
not ( n25822 , n25820 );
not ( n25823 , n25764 );
xor ( n25824 , n25822 , n25823 );
and ( n25825 , n25824 , n25810 );
or ( n25826 , n25821 , n25825 );
buf ( n25827 , n25826 );
not ( n25828 , n25827 );
buf ( n25829 , n25828 );
buf ( n25830 , n25829 );
not ( n25831 , n25830 );
or ( n25832 , n25769 , n25831 );
buf ( n25833 , n25832 );
buf ( n25834 , n25833 );
and ( n25835 , n25834 , n25810 );
not ( n25836 , n25835 );
and ( n25837 , n25836 , n25769 );
xor ( n25838 , n25769 , n25810 );
xor ( n25839 , n25838 , n25810 );
and ( n25840 , n25839 , n25835 );
or ( n25841 , n25837 , n25840 );
buf ( n25842 , n25841 );
not ( n25843 , n25835 );
and ( n25844 , n25843 , n25831 );
xor ( n25845 , n25831 , n25810 );
and ( n25846 , n25838 , n25810 );
xor ( n25847 , n25845 , n25846 );
and ( n25848 , n25847 , n25835 );
or ( n25849 , n25844 , n25848 );
buf ( n25850 , n25849 );
and ( n25851 , n25842 , n25850 );
and ( n25852 , n25663 , n25851 );
buf ( n25853 , RI210b2538_374);
not ( n25854 , n25842 );
and ( n25855 , n25854 , n25850 );
and ( n25856 , n25853 , n25855 );
buf ( n25857 , RI210b43b0_360);
nor ( n25858 , n25854 , n25850 );
and ( n25859 , n25857 , n25858 );
buf ( n25860 , RI210b7f38_335);
nor ( n25861 , n25842 , n25850 );
and ( n25862 , n25860 , n25861 );
or ( n25863 , n25852 , n25856 , n25859 , n25862 );
buf ( n25864 , n25863 );
buf ( n25865 , n25864 );
not ( n25866 , n25865 );
buf ( n25867 , n25866 );
buf ( n25868 , n25867 );
not ( n25869 , n25868 );
buf ( n25870 , RI210afec8_388);
and ( n25871 , n25870 , n25855 );
buf ( n25872 , RI210b2628_372);
and ( n25873 , n25872 , n25858 );
buf ( n25874 , RI210b4d88_356);
and ( n25875 , n25874 , n25861 );
or ( n25876 , C0 , n25871 , n25873 , n25875 );
buf ( n25877 , n25876 );
not ( n25878 , n25877 );
not ( n25879 , n25655 );
and ( n25880 , n25879 , n25246 );
xor ( n25881 , n25246 , n25232 );
and ( n25882 , n25658 , n25232 );
xor ( n25883 , n25881 , n25882 );
and ( n25884 , n25883 , n25655 );
or ( n25885 , n25880 , n25884 );
buf ( n25886 , n25885 );
buf ( n25887 , n25886 );
and ( n25888 , n25887 , n25851 );
and ( n25889 , n24802 , n25855 );
buf ( n25890 , RI21081b18_438);
and ( n25891 , n25890 , n25858 );
buf ( n25892 , RI210b6b88_343);
and ( n25893 , n25892 , n25861 );
or ( n25894 , n25888 , n25889 , n25891 , n25893 );
buf ( n25895 , n25894 );
and ( n25896 , n25878 , n25895 );
not ( n25897 , n25895 );
not ( n25898 , n25864 );
xor ( n25899 , n25897 , n25898 );
and ( n25900 , n25899 , n25877 );
or ( n25901 , n25896 , n25900 );
buf ( n25902 , n25901 );
not ( n25903 , n25902 );
buf ( n25904 , n25903 );
buf ( n25905 , n25904 );
not ( n25906 , n25905 );
or ( n25907 , n25869 , n25906 );
not ( n25908 , n25877 );
not ( n25909 , n25655 );
and ( n25910 , n25909 , n25261 );
xor ( n25911 , n25261 , n25232 );
and ( n25912 , n25881 , n25882 );
xor ( n25913 , n25911 , n25912 );
and ( n25914 , n25913 , n25655 );
or ( n25915 , n25910 , n25914 );
buf ( n25916 , n25915 );
buf ( n25917 , n25916 );
and ( n25918 , n25917 , n25851 );
buf ( n25919 , RI210b07b0_386);
and ( n25920 , n25919 , n25855 );
buf ( n25921 , RI21081aa0_439);
and ( n25922 , n25921 , n25858 );
buf ( n25923 , RI210b5670_354);
and ( n25924 , n25923 , n25861 );
or ( n25925 , n25918 , n25920 , n25922 , n25924 );
buf ( n25926 , n25925 );
and ( n25927 , n25908 , n25926 );
not ( n25928 , n25926 );
and ( n25929 , n25897 , n25898 );
xor ( n25930 , n25928 , n25929 );
and ( n25931 , n25930 , n25877 );
or ( n25932 , n25927 , n25931 );
buf ( n25933 , n25932 );
not ( n25934 , n25933 );
buf ( n25935 , n25934 );
buf ( n25936 , n25935 );
not ( n25937 , n25936 );
or ( n25938 , n25907 , n25937 );
not ( n25939 , n25877 );
not ( n25940 , n25655 );
and ( n25941 , n25940 , n25276 );
xor ( n25942 , n25276 , n25232 );
and ( n25943 , n25911 , n25912 );
xor ( n25944 , n25942 , n25943 );
and ( n25945 , n25944 , n25655 );
or ( n25946 , n25941 , n25945 );
buf ( n25947 , n25946 );
buf ( n25948 , n25947 );
not ( n25949 , n25948 );
buf ( n25950 , n25949 );
and ( n25951 , n25950 , n25851 );
buf ( n25952 , RI210afe50_389);
and ( n25953 , n25952 , n25855 );
buf ( n25954 , RI21080fd8_440);
and ( n25955 , n25954 , n25858 );
buf ( n25956 , RI21083648_424);
and ( n25957 , n25956 , n25861 );
or ( n25958 , n25951 , n25953 , n25955 , n25957 );
buf ( n25959 , n25958 );
and ( n25960 , n25939 , n25959 );
not ( n25961 , n25959 );
and ( n25962 , n25928 , n25929 );
xor ( n25963 , n25961 , n25962 );
and ( n25964 , n25963 , n25877 );
or ( n25965 , n25960 , n25964 );
buf ( n25966 , n25965 );
not ( n25967 , n25966 );
buf ( n25968 , n25967 );
buf ( n25969 , n25968 );
not ( n25970 , n25969 );
or ( n25971 , n25938 , n25970 );
not ( n25972 , n25877 );
not ( n25973 , n25655 );
and ( n25974 , n25973 , n25291 );
xor ( n25975 , n25291 , n25232 );
and ( n25976 , n25942 , n25943 );
xor ( n25977 , n25975 , n25976 );
and ( n25978 , n25977 , n25655 );
or ( n25979 , n25974 , n25978 );
buf ( n25980 , n25979 );
buf ( n25981 , n25980 );
xor ( n25982 , n25981 , n25948 );
buf ( n25983 , n25982 );
and ( n25984 , n25983 , n25851 );
buf ( n25985 , RI2107f3b8_456);
and ( n25986 , n25985 , n25855 );
buf ( n25987 , RI21080f60_441);
and ( n25988 , n25987 , n25858 );
buf ( n25989 , RI210835d0_425);
and ( n25990 , n25989 , n25861 );
or ( n25991 , n25984 , n25986 , n25988 , n25990 );
buf ( n25992 , n25991 );
and ( n25993 , n25972 , n25992 );
not ( n25994 , n25992 );
and ( n25995 , n25961 , n25962 );
xor ( n25996 , n25994 , n25995 );
and ( n25997 , n25996 , n25877 );
or ( n25998 , n25993 , n25997 );
buf ( n25999 , n25998 );
not ( n26000 , n25999 );
buf ( n26001 , n26000 );
buf ( n26002 , n26001 );
not ( n26003 , n26002 );
or ( n26004 , n25971 , n26003 );
not ( n26005 , n25877 );
not ( n26006 , n25655 );
and ( n26007 , n26006 , n25306 );
xor ( n26008 , n25306 , n25232 );
and ( n26009 , n25975 , n25976 );
xor ( n26010 , n26008 , n26009 );
and ( n26011 , n26010 , n25655 );
or ( n26012 , n26007 , n26011 );
buf ( n26013 , n26012 );
buf ( n26014 , n26013 );
and ( n26015 , n25981 , n25948 );
xor ( n26016 , n26014 , n26015 );
buf ( n26017 , n26016 );
and ( n26018 , n26017 , n25851 );
buf ( n26019 , RI210afdd8_390);
and ( n26020 , n26019 , n25855 );
buf ( n26021 , RI21080ee8_442);
and ( n26022 , n26021 , n25858 );
buf ( n26023 , RI210b4d10_357);
and ( n26024 , n26023 , n25861 );
or ( n26025 , n26018 , n26020 , n26022 , n26024 );
buf ( n26026 , n26025 );
and ( n26027 , n26005 , n26026 );
not ( n26028 , n26026 );
and ( n26029 , n25994 , n25995 );
xor ( n26030 , n26028 , n26029 );
and ( n26031 , n26030 , n25877 );
or ( n26032 , n26027 , n26031 );
buf ( n26033 , n26032 );
not ( n26034 , n26033 );
buf ( n26035 , n26034 );
buf ( n26036 , n26035 );
not ( n26037 , n26036 );
or ( n26038 , n26004 , n26037 );
not ( n26039 , n25877 );
not ( n26040 , n25655 );
and ( n26041 , n26040 , n25321 );
xor ( n26042 , n25321 , n25232 );
and ( n26043 , n26008 , n26009 );
xor ( n26044 , n26042 , n26043 );
and ( n26045 , n26044 , n25655 );
or ( n26046 , n26041 , n26045 );
buf ( n26047 , n26046 );
buf ( n26048 , n26047 );
and ( n26049 , n26014 , n26015 );
xor ( n26050 , n26048 , n26049 );
buf ( n26051 , n26050 );
and ( n26052 , n26051 , n25851 );
buf ( n26053 , RI210af568_391);
and ( n26054 , n26053 , n25855 );
buf ( n26055 , RI21080e70_443);
and ( n26056 , n26055 , n25858 );
buf ( n26057 , RI210b4c98_358);
and ( n26058 , n26057 , n25861 );
or ( n26059 , n26052 , n26054 , n26056 , n26058 );
buf ( n26060 , n26059 );
and ( n26061 , n26039 , n26060 );
not ( n26062 , n26060 );
and ( n26063 , n26028 , n26029 );
xor ( n26064 , n26062 , n26063 );
and ( n26065 , n26064 , n25877 );
or ( n26066 , n26061 , n26065 );
buf ( n26067 , n26066 );
not ( n26068 , n26067 );
buf ( n26069 , n26068 );
buf ( n26070 , n26069 );
not ( n26071 , n26070 );
or ( n26072 , n26038 , n26071 );
not ( n26073 , n25877 );
not ( n26074 , n25655 );
and ( n26075 , n26074 , n25336 );
xor ( n26076 , n25336 , n25232 );
and ( n26077 , n26042 , n26043 );
xor ( n26078 , n26076 , n26077 );
and ( n26079 , n26078 , n25655 );
or ( n26080 , n26075 , n26079 );
buf ( n26081 , n26080 );
buf ( n26082 , n26081 );
and ( n26083 , n26048 , n26049 );
xor ( n26084 , n26082 , n26083 );
buf ( n26085 , n26084 );
and ( n26086 , n26085 , n25851 );
buf ( n26087 , RI210af4f0_392);
and ( n26088 , n26087 , n25855 );
buf ( n26089 , RI21080df8_444);
and ( n26090 , n26089 , n25858 );
buf ( n26091 , RI21083558_426);
and ( n26092 , n26091 , n25861 );
or ( n26093 , n26086 , n26088 , n26090 , n26092 );
buf ( n26094 , n26093 );
and ( n26095 , n26073 , n26094 );
not ( n26096 , n26094 );
and ( n26097 , n26062 , n26063 );
xor ( n26098 , n26096 , n26097 );
and ( n26099 , n26098 , n25877 );
or ( n26100 , n26095 , n26099 );
buf ( n26101 , n26100 );
not ( n26102 , n26101 );
buf ( n26103 , n26102 );
buf ( n26104 , n26103 );
not ( n26105 , n26104 );
or ( n26106 , n26072 , n26105 );
not ( n26107 , n25877 );
not ( n26108 , n25655 );
and ( n26109 , n26108 , n25351 );
xor ( n26110 , n25351 , n25232 );
and ( n26111 , n26076 , n26077 );
xor ( n26112 , n26110 , n26111 );
and ( n26113 , n26112 , n25655 );
or ( n26114 , n26109 , n26113 );
buf ( n26115 , n26114 );
buf ( n26116 , n26115 );
and ( n26117 , n26082 , n26083 );
xor ( n26118 , n26116 , n26117 );
buf ( n26119 , n26118 );
and ( n26120 , n26119 , n25851 );
buf ( n26121 , RI210af478_393);
and ( n26122 , n26121 , n25855 );
buf ( n26123 , RI21080d80_445);
and ( n26124 , n26123 , n25858 );
buf ( n26125 , RI210834e0_427);
and ( n26126 , n26125 , n25861 );
or ( n26127 , n26120 , n26122 , n26124 , n26126 );
buf ( n26128 , n26127 );
and ( n26129 , n26107 , n26128 );
not ( n26130 , n26128 );
and ( n26131 , n26096 , n26097 );
xor ( n26132 , n26130 , n26131 );
and ( n26133 , n26132 , n25877 );
or ( n26134 , n26129 , n26133 );
buf ( n26135 , n26134 );
not ( n26136 , n26135 );
buf ( n26137 , n26136 );
buf ( n26138 , n26137 );
not ( n26139 , n26138 );
or ( n26140 , n26106 , n26139 );
not ( n26141 , n25877 );
not ( n26142 , n25655 );
and ( n26143 , n26142 , n25366 );
xor ( n26144 , n25366 , n25232 );
and ( n26145 , n26110 , n26111 );
xor ( n26146 , n26144 , n26145 );
and ( n26147 , n26146 , n25655 );
or ( n26148 , n26143 , n26147 );
buf ( n26149 , n26148 );
buf ( n26150 , n26149 );
and ( n26151 , n26116 , n26117 );
xor ( n26152 , n26150 , n26151 );
buf ( n26153 , n26152 );
and ( n26154 , n26153 , n25851 );
buf ( n26155 , RI210aec08_394);
and ( n26156 , n26155 , n25855 );
buf ( n26157 , RI210b25b0_373);
and ( n26158 , n26157 , n25858 );
buf ( n26159 , RI210b4428_359);
and ( n26160 , n26159 , n25861 );
or ( n26161 , n26154 , n26156 , n26158 , n26160 );
buf ( n26162 , n26161 );
and ( n26163 , n26141 , n26162 );
not ( n26164 , n26162 );
and ( n26165 , n26130 , n26131 );
xor ( n26166 , n26164 , n26165 );
and ( n26167 , n26166 , n25877 );
or ( n26168 , n26163 , n26167 );
buf ( n26169 , n26168 );
not ( n26170 , n26169 );
buf ( n26171 , n26170 );
buf ( n26172 , n26171 );
not ( n26173 , n26172 );
or ( n26174 , n26140 , n26173 );
not ( n26175 , n25877 );
not ( n26176 , n25655 );
and ( n26177 , n26176 , n25381 );
xor ( n26178 , n25381 , n25232 );
and ( n26179 , n26144 , n26145 );
xor ( n26180 , n26178 , n26179 );
and ( n26181 , n26180 , n25655 );
or ( n26182 , n26177 , n26181 );
buf ( n26183 , n26182 );
buf ( n26184 , n26183 );
and ( n26185 , n26150 , n26151 );
xor ( n26186 , n26184 , n26185 );
buf ( n26187 , n26186 );
and ( n26188 , n26187 , n25851 );
buf ( n26189 , RI210b1cc8_375);
and ( n26190 , n26189 , n25855 );
buf ( n26191 , RI21082a18_428);
and ( n26192 , n26191 , n25858 );
buf ( n26193 , RI210b7ec0_336);
and ( n26194 , n26193 , n25861 );
or ( n26195 , n26188 , n26190 , n26192 , n26194 );
buf ( n26196 , n26195 );
and ( n26197 , n26175 , n26196 );
not ( n26198 , n26196 );
and ( n26199 , n26164 , n26165 );
xor ( n26200 , n26198 , n26199 );
and ( n26201 , n26200 , n25877 );
or ( n26202 , n26197 , n26201 );
buf ( n26203 , n26202 );
not ( n26204 , n26203 );
buf ( n26205 , n26204 );
buf ( n26206 , n26205 );
not ( n26207 , n26206 );
or ( n26208 , n26174 , n26207 );
not ( n26209 , n25877 );
not ( n26210 , n25655 );
and ( n26211 , n26210 , n25396 );
xor ( n26212 , n25396 , n25232 );
and ( n26213 , n26178 , n26179 );
xor ( n26214 , n26212 , n26213 );
and ( n26215 , n26214 , n25655 );
or ( n26216 , n26211 , n26215 );
buf ( n26217 , n26216 );
buf ( n26218 , n26217 );
and ( n26219 , n26184 , n26185 );
xor ( n26220 , n26218 , n26219 );
buf ( n26221 , n26220 );
and ( n26222 , n26221 , n25851 );
buf ( n26223 , RI210802b8_446);
and ( n26224 , n26223 , n25855 );
buf ( n26225 , RI210829a0_429);
and ( n26226 , n26225 , n25858 );
buf ( n26227 , RI210b7e48_337);
and ( n26228 , n26227 , n25861 );
or ( n26229 , n26222 , n26224 , n26226 , n26228 );
buf ( n26230 , n26229 );
and ( n26231 , n26209 , n26230 );
not ( n26232 , n26230 );
and ( n26233 , n26198 , n26199 );
xor ( n26234 , n26232 , n26233 );
and ( n26235 , n26234 , n25877 );
or ( n26236 , n26231 , n26235 );
buf ( n26237 , n26236 );
not ( n26238 , n26237 );
buf ( n26239 , n26238 );
buf ( n26240 , n26239 );
not ( n26241 , n26240 );
or ( n26242 , n26208 , n26241 );
not ( n26243 , n25877 );
not ( n26244 , n25655 );
and ( n26245 , n26244 , n25411 );
xor ( n26246 , n25411 , n25232 );
and ( n26247 , n26212 , n26213 );
xor ( n26248 , n26246 , n26247 );
and ( n26249 , n26248 , n25655 );
or ( n26250 , n26245 , n26249 );
buf ( n26251 , n26250 );
buf ( n26252 , n26251 );
and ( n26253 , n26218 , n26219 );
xor ( n26254 , n26252 , n26253 );
buf ( n26255 , n26254 );
and ( n26256 , n26255 , n25851 );
buf ( n26257 , RI21080240_447);
and ( n26258 , n26257 , n25855 );
buf ( n26259 , RI21082928_430);
and ( n26260 , n26259 , n25858 );
buf ( n26261 , RI210b7dd0_338);
and ( n26262 , n26261 , n25861 );
or ( n26263 , n26256 , n26258 , n26260 , n26262 );
buf ( n26264 , n26263 );
and ( n26265 , n26243 , n26264 );
not ( n26266 , n26264 );
and ( n26267 , n26232 , n26233 );
xor ( n26268 , n26266 , n26267 );
and ( n26269 , n26268 , n25877 );
or ( n26270 , n26265 , n26269 );
buf ( n26271 , n26270 );
not ( n26272 , n26271 );
buf ( n26273 , n26272 );
buf ( n26274 , n26273 );
not ( n26275 , n26274 );
or ( n26276 , n26242 , n26275 );
not ( n26277 , n25877 );
not ( n26278 , n25655 );
and ( n26279 , n26278 , n25426 );
xor ( n26280 , n25426 , n25232 );
and ( n26281 , n26246 , n26247 );
xor ( n26282 , n26280 , n26281 );
and ( n26283 , n26282 , n25655 );
or ( n26284 , n26279 , n26283 );
buf ( n26285 , n26284 );
buf ( n26286 , n26285 );
and ( n26287 , n26252 , n26253 );
xor ( n26288 , n26286 , n26287 );
buf ( n26289 , n26288 );
and ( n26290 , n26289 , n25851 );
buf ( n26291 , RI210801c8_448);
and ( n26292 , n26291 , n25855 );
buf ( n26293 , RI210828b0_431);
and ( n26294 , n26293 , n25858 );
buf ( n26295 , RI210b7560_339);
and ( n26296 , n26295 , n25861 );
or ( n26297 , n26290 , n26292 , n26294 , n26296 );
buf ( n26298 , n26297 );
and ( n26299 , n26277 , n26298 );
not ( n26300 , n26298 );
and ( n26301 , n26266 , n26267 );
xor ( n26302 , n26300 , n26301 );
and ( n26303 , n26302 , n25877 );
or ( n26304 , n26299 , n26303 );
buf ( n26305 , n26304 );
not ( n26306 , n26305 );
buf ( n26307 , n26306 );
buf ( n26308 , n26307 );
not ( n26309 , n26308 );
or ( n26310 , n26276 , n26309 );
not ( n26311 , n25877 );
not ( n26312 , n25655 );
and ( n26313 , n26312 , n25441 );
xor ( n26314 , n25441 , n25232 );
and ( n26315 , n26280 , n26281 );
xor ( n26316 , n26314 , n26315 );
and ( n26317 , n26316 , n25655 );
or ( n26318 , n26313 , n26317 );
buf ( n26319 , n26318 );
buf ( n26320 , n26319 );
and ( n26321 , n26286 , n26287 );
xor ( n26322 , n26320 , n26321 );
buf ( n26323 , n26322 );
and ( n26324 , n26323 , n25851 );
buf ( n26325 , RI21080150_449);
and ( n26326 , n26325 , n25855 );
buf ( n26327 , RI21082838_432);
and ( n26328 , n26327 , n25858 );
buf ( n26329 , RI210b74e8_340);
and ( n26330 , n26329 , n25861 );
or ( n26331 , n26324 , n26326 , n26328 , n26330 );
buf ( n26332 , n26331 );
and ( n26333 , n26311 , n26332 );
not ( n26334 , n26332 );
and ( n26335 , n26300 , n26301 );
xor ( n26336 , n26334 , n26335 );
and ( n26337 , n26336 , n25877 );
or ( n26338 , n26333 , n26337 );
buf ( n26339 , n26338 );
not ( n26340 , n26339 );
buf ( n26341 , n26340 );
buf ( n26342 , n26341 );
not ( n26343 , n26342 );
or ( n26344 , n26310 , n26343 );
not ( n26345 , n25877 );
not ( n26346 , n25655 );
and ( n26347 , n26346 , n25456 );
xor ( n26348 , n25456 , n25232 );
and ( n26349 , n26314 , n26315 );
xor ( n26350 , n26348 , n26349 );
and ( n26351 , n26350 , n25655 );
or ( n26352 , n26347 , n26351 );
buf ( n26353 , n26352 );
buf ( n26354 , n26353 );
and ( n26355 , n26320 , n26321 );
xor ( n26356 , n26354 , n26355 );
buf ( n26357 , n26356 );
and ( n26358 , n26357 , n25851 );
buf ( n26359 , RI210800d8_450);
and ( n26360 , n26359 , n25855 );
buf ( n26361 , RI210827c0_433);
and ( n26362 , n26361 , n25858 );
buf ( n26363 , RI210b7470_341);
and ( n26364 , n26363 , n25861 );
or ( n26365 , n26358 , n26360 , n26362 , n26364 );
buf ( n26366 , n26365 );
and ( n26367 , n26345 , n26366 );
not ( n26368 , n26366 );
and ( n26369 , n26334 , n26335 );
xor ( n26370 , n26368 , n26369 );
and ( n26371 , n26370 , n25877 );
or ( n26372 , n26367 , n26371 );
buf ( n26373 , n26372 );
not ( n26374 , n26373 );
buf ( n26375 , n26374 );
buf ( n26376 , n26375 );
not ( n26377 , n26376 );
or ( n26378 , n26344 , n26377 );
not ( n26379 , n25877 );
not ( n26380 , n25655 );
and ( n26381 , n26380 , n25471 );
xor ( n26382 , n25471 , n25232 );
and ( n26383 , n26348 , n26349 );
xor ( n26384 , n26382 , n26383 );
and ( n26385 , n26384 , n25655 );
or ( n26386 , n26381 , n26385 );
buf ( n26387 , n26386 );
buf ( n26388 , n26387 );
and ( n26389 , n26354 , n26355 );
xor ( n26390 , n26388 , n26389 );
buf ( n26391 , n26390 );
and ( n26392 , n26391 , n25851 );
buf ( n26393 , RI21080060_451);
and ( n26394 , n26393 , n25855 );
buf ( n26395 , RI21081cf8_434);
and ( n26396 , n26395 , n25858 );
buf ( n26397 , RI21084200_421);
and ( n26398 , n26397 , n25861 );
or ( n26399 , n26392 , n26394 , n26396 , n26398 );
buf ( n26400 , n26399 );
and ( n26401 , n26379 , n26400 );
not ( n26402 , n26400 );
and ( n26403 , n26368 , n26369 );
xor ( n26404 , n26402 , n26403 );
and ( n26405 , n26404 , n25877 );
or ( n26406 , n26401 , n26405 );
buf ( n26407 , n26406 );
not ( n26408 , n26407 );
buf ( n26409 , n26408 );
buf ( n26410 , n26409 );
not ( n26411 , n26410 );
or ( n26412 , n26378 , n26411 );
not ( n26413 , n25877 );
not ( n26414 , n25655 );
and ( n26415 , n26414 , n25486 );
xor ( n26416 , n25486 , n25232 );
and ( n26417 , n26382 , n26383 );
xor ( n26418 , n26416 , n26417 );
and ( n26419 , n26418 , n25655 );
or ( n26420 , n26415 , n26419 );
buf ( n26421 , n26420 );
buf ( n26422 , n26421 );
and ( n26423 , n26388 , n26389 );
xor ( n26424 , n26422 , n26423 );
buf ( n26425 , n26424 );
and ( n26426 , n26425 , n25851 );
buf ( n26427 , RI2107f598_452);
and ( n26428 , n26427 , n25855 );
buf ( n26429 , RI21081c80_435);
and ( n26430 , n26429 , n25858 );
buf ( n26431 , RI21083738_422);
and ( n26432 , n26431 , n25861 );
or ( n26433 , n26426 , n26428 , n26430 , n26432 );
buf ( n26434 , n26433 );
and ( n26435 , n26413 , n26434 );
not ( n26436 , n26434 );
and ( n26437 , n26402 , n26403 );
xor ( n26438 , n26436 , n26437 );
and ( n26439 , n26438 , n25877 );
or ( n26440 , n26435 , n26439 );
buf ( n26441 , n26440 );
not ( n26442 , n26441 );
buf ( n26443 , n26442 );
buf ( n26444 , n26443 );
not ( n26445 , n26444 );
or ( n26446 , n26412 , n26445 );
not ( n26447 , n25877 );
not ( n26448 , n25655 );
and ( n26449 , n26448 , n25501 );
xor ( n26450 , n25501 , n25232 );
and ( n26451 , n26416 , n26417 );
xor ( n26452 , n26450 , n26451 );
and ( n26453 , n26452 , n25655 );
or ( n26454 , n26449 , n26453 );
buf ( n26455 , n26454 );
buf ( n26456 , n26455 );
and ( n26457 , n26422 , n26423 );
xor ( n26458 , n26456 , n26457 );
buf ( n26459 , n26458 );
and ( n26460 , n26459 , n25851 );
buf ( n26461 , RI210b1c50_376);
and ( n26462 , n26461 , n25855 );
buf ( n26463 , RI21081c08_436);
and ( n26464 , n26463 , n25858 );
buf ( n26465 , RI210836c0_423);
and ( n26466 , n26465 , n25861 );
or ( n26467 , n26460 , n26462 , n26464 , n26466 );
buf ( n26468 , n26467 );
and ( n26469 , n26447 , n26468 );
not ( n26470 , n26468 );
and ( n26471 , n26436 , n26437 );
xor ( n26472 , n26470 , n26471 );
and ( n26473 , n26472 , n25877 );
or ( n26474 , n26469 , n26473 );
buf ( n26475 , n26474 );
not ( n26476 , n26475 );
buf ( n26477 , n26476 );
buf ( n26478 , n26477 );
not ( n26479 , n26478 );
or ( n26480 , n26446 , n26479 );
not ( n26481 , n25877 );
not ( n26482 , n25655 );
and ( n26483 , n26482 , n25516 );
xor ( n26484 , n25516 , n25232 );
and ( n26485 , n26450 , n26451 );
xor ( n26486 , n26484 , n26485 );
and ( n26487 , n26486 , n25655 );
or ( n26488 , n26483 , n26487 );
buf ( n26489 , n26488 );
buf ( n26490 , n26489 );
and ( n26491 , n26456 , n26457 );
xor ( n26492 , n26490 , n26491 );
buf ( n26493 , n26492 );
and ( n26494 , n26493 , n25851 );
buf ( n26495 , RI2107f520_453);
and ( n26496 , n26495 , n25855 );
buf ( n26497 , RI21081b90_437);
and ( n26498 , n26497 , n25858 );
buf ( n26499 , RI210b73f8_342);
and ( n26500 , n26499 , n25861 );
or ( n26501 , n26494 , n26496 , n26498 , n26500 );
buf ( n26502 , n26501 );
and ( n26503 , n26481 , n26502 );
not ( n26504 , n26502 );
and ( n26505 , n26470 , n26471 );
xor ( n26506 , n26504 , n26505 );
and ( n26507 , n26506 , n25877 );
or ( n26508 , n26503 , n26507 );
buf ( n26509 , n26508 );
not ( n26510 , n26509 );
buf ( n26511 , n26510 );
buf ( n26512 , n26511 );
not ( n26513 , n26512 );
or ( n26514 , n26480 , n26513 );
not ( n26515 , n25877 );
not ( n26516 , n25655 );
and ( n26517 , n26516 , n25531 );
xor ( n26518 , n25531 , n25232 );
and ( n26519 , n26484 , n26485 );
xor ( n26520 , n26518 , n26519 );
and ( n26521 , n26520 , n25655 );
or ( n26522 , n26517 , n26521 );
buf ( n26523 , n26522 );
buf ( n26524 , n26523 );
and ( n26525 , n26490 , n26491 );
xor ( n26526 , n26524 , n26525 );
buf ( n26527 , n26526 );
and ( n26528 , n26527 , n25851 );
buf ( n26529 , RI2107f430_455);
and ( n26530 , n26529 , n25855 );
buf ( n26531 , RI210b4338_361);
and ( n26532 , n26531 , n25858 );
buf ( n26533 , RI210b6b10_344);
and ( n26534 , n26533 , n25861 );
or ( n26535 , n26528 , n26530 , n26532 , n26534 );
buf ( n26536 , n26535 );
and ( n26537 , n26515 , n26536 );
not ( n26538 , n26536 );
and ( n26539 , n26504 , n26505 );
xor ( n26540 , n26538 , n26539 );
and ( n26541 , n26540 , n25877 );
or ( n26542 , n26537 , n26541 );
buf ( n26543 , n26542 );
not ( n26544 , n26543 );
buf ( n26545 , n26544 );
buf ( n26546 , n26545 );
not ( n26547 , n26546 );
or ( n26548 , n26514 , n26547 );
not ( n26549 , n25877 );
not ( n26550 , n25655 );
and ( n26551 , n26550 , n25546 );
xor ( n26552 , n25546 , n25232 );
and ( n26553 , n26518 , n26519 );
xor ( n26554 , n26552 , n26553 );
and ( n26555 , n26554 , n25655 );
or ( n26556 , n26551 , n26555 );
buf ( n26557 , n26556 );
buf ( n26558 , n26557 );
and ( n26559 , n26524 , n26525 );
xor ( n26560 , n26558 , n26559 );
buf ( n26561 , n26560 );
and ( n26562 , n26561 , n25851 );
buf ( n26563 , RI210b1bd8_377);
and ( n26564 , n26563 , n25855 );
buf ( n26565 , RI210b42c0_362);
and ( n26566 , n26565 , n25858 );
buf ( n26567 , RI210b6a98_345);
and ( n26568 , n26567 , n25861 );
or ( n26569 , n26562 , n26564 , n26566 , n26568 );
buf ( n26570 , n26569 );
and ( n26571 , n26549 , n26570 );
not ( n26572 , n26570 );
and ( n26573 , n26538 , n26539 );
xor ( n26574 , n26572 , n26573 );
and ( n26575 , n26574 , n25877 );
or ( n26576 , n26571 , n26575 );
buf ( n26577 , n26576 );
not ( n26578 , n26577 );
buf ( n26579 , n26578 );
buf ( n26580 , n26579 );
not ( n26581 , n26580 );
or ( n26582 , n26548 , n26581 );
not ( n26583 , n25877 );
not ( n26584 , n25655 );
and ( n26585 , n26584 , n25561 );
xor ( n26586 , n25561 , n25232 );
and ( n26587 , n26552 , n26553 );
xor ( n26588 , n26586 , n26587 );
and ( n26589 , n26588 , n25655 );
or ( n26590 , n26585 , n26589 );
buf ( n26591 , n26590 );
buf ( n26592 , n26591 );
and ( n26593 , n26558 , n26559 );
xor ( n26594 , n26592 , n26593 );
buf ( n26595 , n26594 );
and ( n26596 , n26595 , n25851 );
buf ( n26597 , RI210b1b60_378);
and ( n26598 , n26597 , n25855 );
buf ( n26599 , RI210b3a50_363);
and ( n26600 , n26599 , n25858 );
buf ( n26601 , RI210b6a20_346);
and ( n26602 , n26601 , n25861 );
or ( n26603 , n26596 , n26598 , n26600 , n26602 );
buf ( n26604 , n26603 );
and ( n26605 , n26583 , n26604 );
not ( n26606 , n26604 );
and ( n26607 , n26572 , n26573 );
xor ( n26608 , n26606 , n26607 );
and ( n26609 , n26608 , n25877 );
or ( n26610 , n26605 , n26609 );
buf ( n26611 , n26610 );
not ( n26612 , n26611 );
buf ( n26613 , n26612 );
buf ( n26614 , n26613 );
not ( n26615 , n26614 );
or ( n26616 , n26582 , n26615 );
not ( n26617 , n25877 );
not ( n26618 , n25655 );
and ( n26619 , n26618 , n25576 );
xor ( n26620 , n25576 , n25232 );
and ( n26621 , n26586 , n26587 );
xor ( n26622 , n26620 , n26621 );
and ( n26623 , n26622 , n25655 );
or ( n26624 , n26619 , n26623 );
buf ( n26625 , n26624 );
buf ( n26626 , n26625 );
and ( n26627 , n26592 , n26593 );
xor ( n26628 , n26626 , n26627 );
buf ( n26629 , n26628 );
and ( n26630 , n26629 , n25851 );
buf ( n26631 , RI210b12f0_379);
and ( n26632 , n26631 , n25855 );
buf ( n26633 , RI210b39d8_364);
and ( n26634 , n26633 , n25858 );
buf ( n26635 , RI210b61b0_347);
and ( n26636 , n26635 , n25861 );
or ( n26637 , n26630 , n26632 , n26634 , n26636 );
buf ( n26638 , n26637 );
and ( n26639 , n26617 , n26638 );
not ( n26640 , n26638 );
and ( n26641 , n26606 , n26607 );
xor ( n26642 , n26640 , n26641 );
and ( n26643 , n26642 , n25877 );
or ( n26644 , n26639 , n26643 );
buf ( n26645 , n26644 );
not ( n26646 , n26645 );
buf ( n26647 , n26646 );
buf ( n26648 , n26647 );
not ( n26649 , n26648 );
or ( n26650 , n26616 , n26649 );
not ( n26651 , n25877 );
not ( n26652 , n25655 );
and ( n26653 , n26652 , n25591 );
xor ( n26654 , n25591 , n25232 );
and ( n26655 , n26620 , n26621 );
xor ( n26656 , n26654 , n26655 );
and ( n26657 , n26656 , n25655 );
or ( n26658 , n26653 , n26657 );
buf ( n26659 , n26658 );
buf ( n26660 , n26659 );
and ( n26661 , n26626 , n26627 );
xor ( n26662 , n26660 , n26661 );
buf ( n26663 , n26662 );
and ( n26664 , n26663 , n25851 );
buf ( n26665 , RI210b1278_380);
and ( n26666 , n26665 , n25855 );
buf ( n26667 , RI210b3960_365);
and ( n26668 , n26667 , n25858 );
buf ( n26669 , RI210b6138_348);
and ( n26670 , n26669 , n25861 );
or ( n26671 , n26664 , n26666 , n26668 , n26670 );
buf ( n26672 , n26671 );
and ( n26673 , n26651 , n26672 );
not ( n26674 , n26672 );
and ( n26675 , n26640 , n26641 );
xor ( n26676 , n26674 , n26675 );
and ( n26677 , n26676 , n25877 );
or ( n26678 , n26673 , n26677 );
buf ( n26679 , n26678 );
not ( n26680 , n26679 );
buf ( n26681 , n26680 );
buf ( n26682 , n26681 );
not ( n26683 , n26682 );
or ( n26684 , n26650 , n26683 );
not ( n26685 , n25877 );
not ( n26686 , n25655 );
and ( n26687 , n26686 , n25606 );
xor ( n26688 , n25606 , n25232 );
and ( n26689 , n26654 , n26655 );
xor ( n26690 , n26688 , n26689 );
and ( n26691 , n26690 , n25655 );
or ( n26692 , n26687 , n26691 );
buf ( n26693 , n26692 );
buf ( n26694 , n26693 );
and ( n26695 , n26660 , n26661 );
xor ( n26696 , n26694 , n26695 );
buf ( n26697 , n26696 );
and ( n26698 , n26697 , n25851 );
buf ( n26699 , RI210b1200_381);
and ( n26700 , n26699 , n25855 );
buf ( n26701 , RI210b38e8_366);
and ( n26702 , n26701 , n25858 );
buf ( n26703 , RI210b60c0_349);
and ( n26704 , n26703 , n25861 );
or ( n26705 , n26698 , n26700 , n26702 , n26704 );
buf ( n26706 , n26705 );
and ( n26707 , n26685 , n26706 );
not ( n26708 , n26706 );
and ( n26709 , n26674 , n26675 );
xor ( n26710 , n26708 , n26709 );
and ( n26711 , n26710 , n25877 );
or ( n26712 , n26707 , n26711 );
buf ( n26713 , n26712 );
not ( n26714 , n26713 );
buf ( n26715 , n26714 );
buf ( n26716 , n26715 );
not ( n26717 , n26716 );
or ( n26718 , n26684 , n26717 );
not ( n26719 , n25877 );
not ( n26720 , n25655 );
and ( n26721 , n26720 , n25621 );
xor ( n26722 , n25621 , n25232 );
and ( n26723 , n26688 , n26689 );
xor ( n26724 , n26722 , n26723 );
and ( n26725 , n26724 , n25655 );
or ( n26726 , n26721 , n26725 );
buf ( n26727 , n26726 );
buf ( n26728 , n26727 );
and ( n26729 , n26694 , n26695 );
xor ( n26730 , n26728 , n26729 );
buf ( n26731 , n26730 );
and ( n26732 , n26731 , n25851 );
buf ( n26733 , RI210b1188_382);
and ( n26734 , n26733 , n25855 );
buf ( n26735 , RI210b3078_367);
and ( n26736 , n26735 , n25858 );
buf ( n26737 , RI210b6048_350);
and ( n26738 , n26737 , n25861 );
or ( n26739 , n26732 , n26734 , n26736 , n26738 );
buf ( n26740 , n26739 );
and ( n26741 , n26719 , n26740 );
not ( n26742 , n26740 );
and ( n26743 , n26708 , n26709 );
xor ( n26744 , n26742 , n26743 );
and ( n26745 , n26744 , n25877 );
or ( n26746 , n26741 , n26745 );
buf ( n26747 , n26746 );
not ( n26748 , n26747 );
buf ( n26749 , n26748 );
buf ( n26750 , n26749 );
not ( n26751 , n26750 );
or ( n26752 , n26718 , n26751 );
not ( n26753 , n25877 );
not ( n26754 , n25655 );
and ( n26755 , n26754 , n25636 );
xor ( n26756 , n25636 , n25232 );
and ( n26757 , n26722 , n26723 );
xor ( n26758 , n26756 , n26757 );
and ( n26759 , n26758 , n25655 );
or ( n26760 , n26755 , n26759 );
buf ( n26761 , n26760 );
buf ( n26762 , n26761 );
and ( n26763 , n26728 , n26729 );
xor ( n26764 , n26762 , n26763 );
buf ( n26765 , n26764 );
and ( n26766 , n26765 , n25851 );
buf ( n26767 , RI210b0918_383);
and ( n26768 , n26767 , n25855 );
buf ( n26769 , RI210b3000_368);
and ( n26770 , n26769 , n25858 );
buf ( n26771 , RI210b57d8_351);
and ( n26772 , n26771 , n25861 );
or ( n26773 , n26766 , n26768 , n26770 , n26772 );
buf ( n26774 , n26773 );
and ( n26775 , n26753 , n26774 );
not ( n26776 , n26774 );
and ( n26777 , n26742 , n26743 );
xor ( n26778 , n26776 , n26777 );
and ( n26779 , n26778 , n25877 );
or ( n26780 , n26775 , n26779 );
buf ( n26781 , n26780 );
not ( n26782 , n26781 );
buf ( n26783 , n26782 );
buf ( n26784 , n26783 );
not ( n26785 , n26784 );
or ( n26786 , n26752 , n26785 );
not ( n26787 , n25877 );
not ( n26788 , n25655 );
and ( n26789 , n26788 , n25651 );
xor ( n26790 , n25651 , n25232 );
and ( n26791 , n26756 , n26757 );
xor ( n26792 , n26790 , n26791 );
and ( n26793 , n26792 , n25655 );
or ( n26794 , n26789 , n26793 );
buf ( n26795 , n26794 );
buf ( n26796 , n26795 );
and ( n26797 , n26762 , n26763 );
xor ( n26798 , n26796 , n26797 );
buf ( n26799 , n26798 );
and ( n26800 , n26799 , n25851 );
buf ( n26801 , RI210b08a0_384);
and ( n26802 , n26801 , n25855 );
buf ( n26803 , RI210b2f88_369);
and ( n26804 , n26803 , n25858 );
buf ( n26805 , RI210b5760_352);
and ( n26806 , n26805 , n25861 );
or ( n26807 , n26800 , n26802 , n26804 , n26806 );
buf ( n26808 , n26807 );
and ( n26809 , n26787 , n26808 );
not ( n26810 , n26808 );
and ( n26811 , n26776 , n26777 );
xor ( n26812 , n26810 , n26811 );
and ( n26813 , n26812 , n25877 );
or ( n26814 , n26809 , n26813 );
buf ( n26815 , n26814 );
not ( n26816 , n26815 );
buf ( n26817 , n26816 );
buf ( n26818 , n26817 );
not ( n26819 , n26818 );
or ( n26820 , n26786 , n26819 );
buf ( n26821 , n26820 );
buf ( n26822 , n26821 );
and ( n26823 , n26822 , n25877 );
not ( n26824 , n26823 );
and ( n26825 , n26824 , n25869 );
xor ( n26826 , n25869 , n25877 );
xor ( n26827 , n26826 , n25877 );
and ( n26828 , n26827 , n26823 );
or ( n26829 , n26825 , n26828 );
buf ( n26830 , n26829 );
buf ( n26831 , n24061 );
not ( n26832 , n26831 );
buf ( n26833 , n24349 );
and ( n26834 , n26832 , n26833 );
not ( n26835 , n26833 );
buf ( n26836 , n24357 );
not ( n26837 , n26836 );
buf ( n26838 , n24365 );
not ( n26839 , n26838 );
buf ( n26840 , n24373 );
not ( n26841 , n26840 );
buf ( n26842 , n24069 );
not ( n26843 , n26842 );
buf ( n26844 , n24078 );
not ( n26845 , n26844 );
buf ( n26846 , n24086 );
not ( n26847 , n26846 );
buf ( n26848 , n24094 );
not ( n26849 , n26848 );
buf ( n26850 , n24102 );
not ( n26851 , n26850 );
buf ( n26852 , n24110 );
not ( n26853 , n26852 );
buf ( n26854 , n24118 );
not ( n26855 , n26854 );
buf ( n26856 , n24126 );
not ( n26857 , n26856 );
buf ( n26858 , n24134 );
not ( n26859 , n26858 );
buf ( n26860 , n24142 );
not ( n26861 , n26860 );
buf ( n26862 , n24150 );
not ( n26863 , n26862 );
buf ( n26864 , n24158 );
not ( n26865 , n26864 );
buf ( n26866 , n24166 );
not ( n26867 , n26866 );
buf ( n26868 , n24174 );
not ( n26869 , n26868 );
buf ( n26870 , n24182 );
not ( n26871 , n26870 );
buf ( n26872 , n24190 );
not ( n26873 , n26872 );
buf ( n26874 , n24198 );
not ( n26875 , n26874 );
buf ( n26876 , n24206 );
not ( n26877 , n26876 );
buf ( n26878 , n24214 );
not ( n26879 , n26878 );
buf ( n26880 , n24222 );
not ( n26881 , n26880 );
buf ( n26882 , n24230 );
not ( n26883 , n26882 );
buf ( n26884 , n24238 );
not ( n26885 , n26884 );
buf ( n26886 , n24246 );
not ( n26887 , n26886 );
buf ( n26888 , n24249 );
not ( n26889 , n26888 );
and ( n26890 , n26887 , n26889 );
and ( n26891 , n26885 , n26890 );
and ( n26892 , n26883 , n26891 );
and ( n26893 , n26881 , n26892 );
and ( n26894 , n26879 , n26893 );
and ( n26895 , n26877 , n26894 );
and ( n26896 , n26875 , n26895 );
and ( n26897 , n26873 , n26896 );
and ( n26898 , n26871 , n26897 );
and ( n26899 , n26869 , n26898 );
and ( n26900 , n26867 , n26899 );
and ( n26901 , n26865 , n26900 );
and ( n26902 , n26863 , n26901 );
and ( n26903 , n26861 , n26902 );
and ( n26904 , n26859 , n26903 );
and ( n26905 , n26857 , n26904 );
and ( n26906 , n26855 , n26905 );
and ( n26907 , n26853 , n26906 );
and ( n26908 , n26851 , n26907 );
and ( n26909 , n26849 , n26908 );
and ( n26910 , n26847 , n26909 );
and ( n26911 , n26845 , n26910 );
and ( n26912 , n26843 , n26911 );
and ( n26913 , n26841 , n26912 );
and ( n26914 , n26839 , n26913 );
and ( n26915 , n26837 , n26914 );
xor ( n26916 , n26835 , n26915 );
and ( n26917 , n26916 , n26831 );
or ( n26918 , n26834 , n26917 );
buf ( n26919 , n26918 );
not ( n26920 , n26919 );
buf ( n26921 , n26920 );
buf ( n26922 , n26921 );
not ( n26923 , n26922 );
buf ( n26924 , n26923 );
buf ( n26925 , n26924 );
buf ( n26926 , n26925 );
not ( n26927 , n26926 );
buf ( n26928 , n26927 );
buf ( n26929 , n26928 );
not ( n26930 , n26929 );
not ( n26931 , n26831 );
buf ( n26932 , n24325 );
not ( n26933 , n26932 );
buf ( n26934 , n24333 );
not ( n26935 , n26934 );
buf ( n26936 , n24341 );
not ( n26937 , n26936 );
and ( n26938 , n26835 , n26915 );
and ( n26939 , n26937 , n26938 );
and ( n26940 , n26935 , n26939 );
and ( n26941 , n26933 , n26940 );
xor ( n26942 , n26931 , n26941 );
buf ( n26943 , n26831 );
and ( n26944 , n26942 , n26943 );
or ( n26945 , C0 , n26944 );
buf ( n26946 , n26945 );
not ( n26947 , n26946 );
buf ( n26948 , n26947 );
buf ( n26949 , n26948 );
not ( n26950 , n26949 );
buf ( n26951 , n26950 );
not ( n26952 , n26951 );
buf ( n26953 , n26952 );
not ( n26954 , n26831 );
and ( n26955 , n26954 , n26932 );
xor ( n26956 , n26933 , n26940 );
and ( n26957 , n26956 , n26831 );
or ( n26958 , n26955 , n26957 );
buf ( n26959 , n26958 );
not ( n26960 , n26959 );
buf ( n26961 , n26960 );
buf ( n26962 , n26961 );
not ( n26963 , n26962 );
buf ( n26964 , n26963 );
not ( n26965 , n26964 );
buf ( n26966 , n26965 );
not ( n26967 , n26831 );
and ( n26968 , n26967 , n26934 );
xor ( n26969 , n26935 , n26939 );
and ( n26970 , n26969 , n26831 );
or ( n26971 , n26968 , n26970 );
buf ( n26972 , n26971 );
not ( n26973 , n26972 );
buf ( n26974 , n26973 );
buf ( n26975 , n26974 );
not ( n26976 , n26975 );
buf ( n26977 , n26976 );
not ( n26978 , n26977 );
buf ( n26979 , n26978 );
not ( n26980 , n26831 );
and ( n26981 , n26980 , n26936 );
xor ( n26982 , n26937 , n26938 );
and ( n26983 , n26982 , n26831 );
or ( n26984 , n26981 , n26983 );
buf ( n26985 , n26984 );
not ( n26986 , n26985 );
buf ( n26987 , n26986 );
buf ( n26988 , n26987 );
not ( n26989 , n26988 );
buf ( n26990 , n26989 );
not ( n26991 , n26990 );
buf ( n26992 , n26991 );
not ( n26993 , n26924 );
buf ( n26994 , n26993 );
and ( n26995 , n26992 , n26994 );
and ( n26996 , n26979 , n26995 );
and ( n26997 , n26966 , n26996 );
and ( n26998 , n26953 , n26997 );
not ( n26999 , n26998 );
buf ( n27000 , n26999 );
buf ( n27001 , n26831 );
and ( n27002 , n27000 , n27001 );
or ( n27003 , C0 , n27002 );
buf ( n27004 , n27003 );
buf ( n27005 , n27004 );
not ( n27006 , n27005 );
not ( n27007 , n27001 );
buf ( n27008 , n26990 );
and ( n27009 , n27007 , n27008 );
xor ( n27010 , n26992 , n26994 );
buf ( n27011 , n27010 );
and ( n27012 , n27011 , n27001 );
or ( n27013 , n27009 , n27012 );
buf ( n27014 , n27013 );
buf ( n27015 , n27014 );
and ( n27016 , n27006 , n27015 );
not ( n27017 , n27015 );
not ( n27018 , n26925 );
xor ( n27019 , n27017 , n27018 );
and ( n27020 , n27019 , n27005 );
or ( n27021 , n27016 , n27020 );
buf ( n27022 , n27021 );
not ( n27023 , n27022 );
buf ( n27024 , n27023 );
buf ( n27025 , n27024 );
not ( n27026 , n27025 );
or ( n27027 , n26930 , n27026 );
buf ( n27028 , n27027 );
buf ( n27029 , n27028 );
and ( n27030 , n27029 , n27005 );
not ( n27031 , n27030 );
and ( n27032 , n27031 , n26930 );
xor ( n27033 , n26930 , n27005 );
xor ( n27034 , n27033 , n27005 );
and ( n27035 , n27034 , n27030 );
or ( n27036 , n27032 , n27035 );
buf ( n27037 , n27036 );
not ( n27038 , n27030 );
and ( n27039 , n27038 , n27026 );
xor ( n27040 , n27026 , n27005 );
and ( n27041 , n27033 , n27005 );
xor ( n27042 , n27040 , n27041 );
and ( n27043 , n27042 , n27030 );
or ( n27044 , n27039 , n27043 );
buf ( n27045 , n27044 );
and ( n27046 , n27037 , n27045 );
and ( n27047 , n26830 , n27046 );
not ( n27048 , n27037 );
and ( n27049 , n27048 , n27045 );
and ( n27050 , n26830 , n27049 );
buf ( n27051 , RI210cdec8_250);
not ( n27052 , n27051 );
buf ( n27053 , n25876 );
buf ( n27054 , n27053 );
not ( n27055 , n27054 );
not ( n27056 , n27053 );
buf ( n27057 , n25925 );
and ( n27058 , n27056 , n27057 );
not ( n27059 , n27057 );
buf ( n27060 , n25894 );
not ( n27061 , n27060 );
buf ( n27062 , n25863 );
not ( n27063 , n27062 );
and ( n27064 , n27061 , n27063 );
xor ( n27065 , n27059 , n27064 );
and ( n27066 , n27065 , n27053 );
or ( n27067 , n27058 , n27066 );
buf ( n27068 , n27067 );
not ( n27069 , n27068 );
buf ( n27070 , n27069 );
buf ( n27071 , n27070 );
and ( n27072 , C1 , n27071 );
and ( n27073 , C1 , n27072 );
and ( n27074 , C1 , n27073 );
and ( n27075 , C1 , n27074 );
and ( n27076 , C1 , n27075 );
and ( n27077 , C1 , n27076 );
and ( n27078 , C1 , n27077 );
and ( n27079 , C1 , n27078 );
and ( n27080 , C1 , n27079 );
and ( n27081 , C1 , n27080 );
and ( n27082 , C1 , n27081 );
and ( n27083 , C1 , n27082 );
and ( n27084 , C1 , n27083 );
and ( n27085 , C1 , n27084 );
and ( n27086 , C1 , n27085 );
and ( n27087 , C1 , n27086 );
and ( n27088 , C1 , n27087 );
and ( n27089 , C1 , n27088 );
and ( n27090 , C1 , n27089 );
and ( n27091 , C1 , n27090 );
and ( n27092 , C1 , n27091 );
and ( n27093 , C1 , n27092 );
and ( n27094 , C1 , n27093 );
and ( n27095 , C1 , n27094 );
and ( n27096 , C1 , n27095 );
and ( n27097 , C1 , n27096 );
and ( n27098 , C1 , n27097 );
and ( n27099 , C1 , n27098 );
buf ( n27100 , n27099 );
not ( n27101 , n27100 );
buf ( n27102 , n27101 );
buf ( n27103 , n27102 );
and ( n27104 , n27055 , n27103 );
not ( n27105 , n27102 );
buf ( n27106 , n27105 );
not ( n27107 , n27053 );
and ( n27108 , n27107 , n27060 );
xor ( n27109 , n27061 , n27063 );
and ( n27110 , n27109 , n27053 );
or ( n27111 , n27108 , n27110 );
buf ( n27112 , n27111 );
not ( n27113 , n27112 );
buf ( n27114 , n27113 );
buf ( n27115 , n27114 );
and ( n27116 , C1 , n27115 );
and ( n27117 , C1 , n27116 );
and ( n27118 , C1 , n27117 );
and ( n27119 , C1 , n27118 );
and ( n27120 , C1 , n27119 );
and ( n27121 , C1 , n27120 );
and ( n27122 , C1 , n27121 );
and ( n27123 , C1 , n27122 );
and ( n27124 , C1 , n27123 );
and ( n27125 , C1 , n27124 );
and ( n27126 , C1 , n27125 );
and ( n27127 , C1 , n27126 );
and ( n27128 , C1 , n27127 );
and ( n27129 , C1 , n27128 );
and ( n27130 , C1 , n27129 );
and ( n27131 , C1 , n27130 );
and ( n27132 , C1 , n27131 );
and ( n27133 , C1 , n27132 );
and ( n27134 , C1 , n27133 );
and ( n27135 , C1 , n27134 );
and ( n27136 , C1 , n27135 );
and ( n27137 , C1 , n27136 );
and ( n27138 , C1 , n27137 );
and ( n27139 , C1 , n27138 );
and ( n27140 , C1 , n27139 );
and ( n27141 , C1 , n27140 );
and ( n27142 , C1 , n27141 );
and ( n27143 , C1 , n27142 );
and ( n27144 , C1 , n27143 );
buf ( n27145 , n27144 );
not ( n27146 , n27145 );
buf ( n27147 , n27146 );
not ( n27148 , n27147 );
buf ( n27149 , n27148 );
xor ( n27150 , n27106 , n27149 );
buf ( n27151 , n27150 );
and ( n27152 , n27151 , n27054 );
or ( n27153 , n27104 , n27152 );
buf ( n27154 , n27153 );
and ( n27155 , n27052 , n27154 );
buf ( n27156 , n27147 );
buf ( n27157 , n27156 );
buf ( n27158 , n27157 );
not ( n27159 , n27158 );
buf ( n27160 , n27159 );
buf ( n27161 , n27160 );
not ( n27162 , n27161 );
not ( n27163 , n27053 );
and ( n27164 , n26790 , n26791 );
buf ( n27165 , n27164 );
and ( n27166 , n27165 , n25655 );
or ( n27167 , C0 , n27166 );
buf ( n27168 , n27167 );
buf ( n27169 , n27168 );
and ( n27170 , n26796 , n26797 );
and ( n27171 , n27169 , n27170 );
buf ( n27172 , n27171 );
buf ( n27173 , n27172 );
and ( n27174 , n27173 , n25851 );
buf ( n27175 , RI210aff40_387);
and ( n27176 , n27175 , n25855 );
buf ( n27177 , RI210b26a0_371);
and ( n27178 , n27177 , n25858 );
buf ( n27179 , RI210b4e00_355);
and ( n27180 , n27179 , n25861 );
or ( n27181 , n27174 , n27176 , n27178 , n27180 );
buf ( n27182 , n27181 );
not ( n27183 , n27182 );
xor ( n27184 , n27169 , n27170 );
buf ( n27185 , n27184 );
and ( n27186 , n27185 , n25851 );
buf ( n27187 , RI210b0828_385);
and ( n27188 , n27187 , n25855 );
buf ( n27189 , RI210b2f10_370);
and ( n27190 , n27189 , n25858 );
buf ( n27191 , RI210b56e8_353);
and ( n27192 , n27191 , n25861 );
or ( n27193 , n27186 , n27188 , n27190 , n27192 );
buf ( n27194 , n27193 );
not ( n27195 , n27194 );
buf ( n27196 , n26807 );
not ( n27197 , n27196 );
buf ( n27198 , n26773 );
not ( n27199 , n27198 );
buf ( n27200 , n26739 );
not ( n27201 , n27200 );
buf ( n27202 , n26705 );
not ( n27203 , n27202 );
buf ( n27204 , n26671 );
not ( n27205 , n27204 );
buf ( n27206 , n26637 );
not ( n27207 , n27206 );
buf ( n27208 , n26603 );
not ( n27209 , n27208 );
buf ( n27210 , n26569 );
not ( n27211 , n27210 );
buf ( n27212 , n26535 );
not ( n27213 , n27212 );
buf ( n27214 , n26501 );
not ( n27215 , n27214 );
buf ( n27216 , n26467 );
not ( n27217 , n27216 );
buf ( n27218 , n26433 );
not ( n27219 , n27218 );
buf ( n27220 , n26399 );
not ( n27221 , n27220 );
buf ( n27222 , n26365 );
not ( n27223 , n27222 );
buf ( n27224 , n26331 );
not ( n27225 , n27224 );
buf ( n27226 , n26297 );
not ( n27227 , n27226 );
buf ( n27228 , n26263 );
not ( n27229 , n27228 );
buf ( n27230 , n26229 );
not ( n27231 , n27230 );
buf ( n27232 , n26195 );
not ( n27233 , n27232 );
buf ( n27234 , n26161 );
not ( n27235 , n27234 );
buf ( n27236 , n26127 );
not ( n27237 , n27236 );
buf ( n27238 , n26093 );
not ( n27239 , n27238 );
buf ( n27240 , n26059 );
not ( n27241 , n27240 );
buf ( n27242 , n26025 );
not ( n27243 , n27242 );
buf ( n27244 , n25991 );
not ( n27245 , n27244 );
buf ( n27246 , n25958 );
not ( n27247 , n27246 );
and ( n27248 , n27059 , n27064 );
and ( n27249 , n27247 , n27248 );
and ( n27250 , n27245 , n27249 );
and ( n27251 , n27243 , n27250 );
and ( n27252 , n27241 , n27251 );
and ( n27253 , n27239 , n27252 );
and ( n27254 , n27237 , n27253 );
and ( n27255 , n27235 , n27254 );
and ( n27256 , n27233 , n27255 );
and ( n27257 , n27231 , n27256 );
and ( n27258 , n27229 , n27257 );
and ( n27259 , n27227 , n27258 );
and ( n27260 , n27225 , n27259 );
and ( n27261 , n27223 , n27260 );
and ( n27262 , n27221 , n27261 );
and ( n27263 , n27219 , n27262 );
and ( n27264 , n27217 , n27263 );
and ( n27265 , n27215 , n27264 );
and ( n27266 , n27213 , n27265 );
and ( n27267 , n27211 , n27266 );
and ( n27268 , n27209 , n27267 );
and ( n27269 , n27207 , n27268 );
and ( n27270 , n27205 , n27269 );
and ( n27271 , n27203 , n27270 );
and ( n27272 , n27201 , n27271 );
and ( n27273 , n27199 , n27272 );
and ( n27274 , n27197 , n27273 );
and ( n27275 , n27195 , n27274 );
and ( n27276 , n27183 , n27275 );
xor ( n27277 , n27163 , n27276 );
buf ( n27278 , n27053 );
and ( n27279 , n27277 , n27278 );
or ( n27280 , C0 , n27279 );
buf ( n27281 , n27280 );
not ( n27282 , n27281 );
buf ( n27283 , n27282 );
not ( n27284 , n27283 );
buf ( n27285 , n27284 );
not ( n27286 , n27285 );
buf ( n27287 , n27286 );
not ( n27288 , n27053 );
and ( n27289 , n27288 , n27182 );
xor ( n27290 , n27183 , n27275 );
and ( n27291 , n27290 , n27053 );
or ( n27292 , n27289 , n27291 );
buf ( n27293 , n27292 );
not ( n27294 , n27293 );
buf ( n27295 , n27294 );
buf ( n27296 , n27295 );
not ( n27297 , n27296 );
buf ( n27298 , n27297 );
not ( n27299 , n27298 );
buf ( n27300 , n27299 );
not ( n27301 , n27053 );
and ( n27302 , n27301 , n27194 );
xor ( n27303 , n27195 , n27274 );
and ( n27304 , n27303 , n27053 );
or ( n27305 , n27302 , n27304 );
buf ( n27306 , n27305 );
not ( n27307 , n27306 );
buf ( n27308 , n27307 );
buf ( n27309 , n27308 );
not ( n27310 , n27309 );
buf ( n27311 , n27310 );
not ( n27312 , n27311 );
buf ( n27313 , n27312 );
not ( n27314 , n27053 );
and ( n27315 , n27314 , n27196 );
xor ( n27316 , n27197 , n27273 );
and ( n27317 , n27316 , n27053 );
or ( n27318 , n27315 , n27317 );
buf ( n27319 , n27318 );
not ( n27320 , n27319 );
buf ( n27321 , n27320 );
buf ( n27322 , n27321 );
not ( n27323 , n27322 );
buf ( n27324 , n27323 );
not ( n27325 , n27324 );
buf ( n27326 , n27325 );
not ( n27327 , n27053 );
and ( n27328 , n27327 , n27198 );
xor ( n27329 , n27199 , n27272 );
and ( n27330 , n27329 , n27053 );
or ( n27331 , n27328 , n27330 );
buf ( n27332 , n27331 );
not ( n27333 , n27332 );
buf ( n27334 , n27333 );
buf ( n27335 , n27334 );
not ( n27336 , n27335 );
buf ( n27337 , n27336 );
not ( n27338 , n27337 );
buf ( n27339 , n27338 );
not ( n27340 , n27053 );
and ( n27341 , n27340 , n27200 );
xor ( n27342 , n27201 , n27271 );
and ( n27343 , n27342 , n27053 );
or ( n27344 , n27341 , n27343 );
buf ( n27345 , n27344 );
not ( n27346 , n27345 );
buf ( n27347 , n27346 );
buf ( n27348 , n27347 );
not ( n27349 , n27348 );
buf ( n27350 , n27349 );
not ( n27351 , n27350 );
buf ( n27352 , n27351 );
not ( n27353 , n27053 );
and ( n27354 , n27353 , n27202 );
xor ( n27355 , n27203 , n27270 );
and ( n27356 , n27355 , n27053 );
or ( n27357 , n27354 , n27356 );
buf ( n27358 , n27357 );
not ( n27359 , n27358 );
buf ( n27360 , n27359 );
buf ( n27361 , n27360 );
not ( n27362 , n27361 );
buf ( n27363 , n27362 );
not ( n27364 , n27363 );
buf ( n27365 , n27364 );
not ( n27366 , n27053 );
and ( n27367 , n27366 , n27204 );
xor ( n27368 , n27205 , n27269 );
and ( n27369 , n27368 , n27053 );
or ( n27370 , n27367 , n27369 );
buf ( n27371 , n27370 );
not ( n27372 , n27371 );
buf ( n27373 , n27372 );
buf ( n27374 , n27373 );
not ( n27375 , n27374 );
buf ( n27376 , n27375 );
not ( n27377 , n27376 );
buf ( n27378 , n27377 );
not ( n27379 , n27053 );
and ( n27380 , n27379 , n27206 );
xor ( n27381 , n27207 , n27268 );
and ( n27382 , n27381 , n27053 );
or ( n27383 , n27380 , n27382 );
buf ( n27384 , n27383 );
not ( n27385 , n27384 );
buf ( n27386 , n27385 );
buf ( n27387 , n27386 );
not ( n27388 , n27387 );
buf ( n27389 , n27388 );
not ( n27390 , n27389 );
buf ( n27391 , n27390 );
not ( n27392 , n27053 );
and ( n27393 , n27392 , n27208 );
xor ( n27394 , n27209 , n27267 );
and ( n27395 , n27394 , n27053 );
or ( n27396 , n27393 , n27395 );
buf ( n27397 , n27396 );
not ( n27398 , n27397 );
buf ( n27399 , n27398 );
buf ( n27400 , n27399 );
not ( n27401 , n27400 );
buf ( n27402 , n27401 );
not ( n27403 , n27402 );
buf ( n27404 , n27403 );
not ( n27405 , n27053 );
and ( n27406 , n27405 , n27210 );
xor ( n27407 , n27211 , n27266 );
and ( n27408 , n27407 , n27053 );
or ( n27409 , n27406 , n27408 );
buf ( n27410 , n27409 );
not ( n27411 , n27410 );
buf ( n27412 , n27411 );
buf ( n27413 , n27412 );
not ( n27414 , n27413 );
buf ( n27415 , n27414 );
not ( n27416 , n27415 );
buf ( n27417 , n27416 );
not ( n27418 , n27053 );
and ( n27419 , n27418 , n27212 );
xor ( n27420 , n27213 , n27265 );
and ( n27421 , n27420 , n27053 );
or ( n27422 , n27419 , n27421 );
buf ( n27423 , n27422 );
not ( n27424 , n27423 );
buf ( n27425 , n27424 );
buf ( n27426 , n27425 );
not ( n27427 , n27426 );
buf ( n27428 , n27427 );
not ( n27429 , n27428 );
buf ( n27430 , n27429 );
not ( n27431 , n27053 );
and ( n27432 , n27431 , n27214 );
xor ( n27433 , n27215 , n27264 );
and ( n27434 , n27433 , n27053 );
or ( n27435 , n27432 , n27434 );
buf ( n27436 , n27435 );
not ( n27437 , n27436 );
buf ( n27438 , n27437 );
buf ( n27439 , n27438 );
not ( n27440 , n27439 );
buf ( n27441 , n27440 );
not ( n27442 , n27441 );
buf ( n27443 , n27442 );
not ( n27444 , n27053 );
and ( n27445 , n27444 , n27216 );
xor ( n27446 , n27217 , n27263 );
and ( n27447 , n27446 , n27053 );
or ( n27448 , n27445 , n27447 );
buf ( n27449 , n27448 );
not ( n27450 , n27449 );
buf ( n27451 , n27450 );
buf ( n27452 , n27451 );
not ( n27453 , n27452 );
buf ( n27454 , n27453 );
not ( n27455 , n27454 );
buf ( n27456 , n27455 );
not ( n27457 , n27053 );
and ( n27458 , n27457 , n27218 );
xor ( n27459 , n27219 , n27262 );
and ( n27460 , n27459 , n27053 );
or ( n27461 , n27458 , n27460 );
buf ( n27462 , n27461 );
not ( n27463 , n27462 );
buf ( n27464 , n27463 );
buf ( n27465 , n27464 );
not ( n27466 , n27465 );
buf ( n27467 , n27466 );
not ( n27468 , n27467 );
buf ( n27469 , n27468 );
not ( n27470 , n27053 );
and ( n27471 , n27470 , n27220 );
xor ( n27472 , n27221 , n27261 );
and ( n27473 , n27472 , n27053 );
or ( n27474 , n27471 , n27473 );
buf ( n27475 , n27474 );
not ( n27476 , n27475 );
buf ( n27477 , n27476 );
buf ( n27478 , n27477 );
not ( n27479 , n27478 );
buf ( n27480 , n27479 );
not ( n27481 , n27480 );
buf ( n27482 , n27481 );
not ( n27483 , n27053 );
and ( n27484 , n27483 , n27222 );
xor ( n27485 , n27223 , n27260 );
and ( n27486 , n27485 , n27053 );
or ( n27487 , n27484 , n27486 );
buf ( n27488 , n27487 );
not ( n27489 , n27488 );
buf ( n27490 , n27489 );
buf ( n27491 , n27490 );
not ( n27492 , n27491 );
buf ( n27493 , n27492 );
not ( n27494 , n27493 );
buf ( n27495 , n27494 );
not ( n27496 , n27053 );
and ( n27497 , n27496 , n27224 );
xor ( n27498 , n27225 , n27259 );
and ( n27499 , n27498 , n27053 );
or ( n27500 , n27497 , n27499 );
buf ( n27501 , n27500 );
not ( n27502 , n27501 );
buf ( n27503 , n27502 );
buf ( n27504 , n27503 );
not ( n27505 , n27504 );
buf ( n27506 , n27505 );
not ( n27507 , n27506 );
buf ( n27508 , n27507 );
not ( n27509 , n27053 );
and ( n27510 , n27509 , n27226 );
xor ( n27511 , n27227 , n27258 );
and ( n27512 , n27511 , n27053 );
or ( n27513 , n27510 , n27512 );
buf ( n27514 , n27513 );
not ( n27515 , n27514 );
buf ( n27516 , n27515 );
buf ( n27517 , n27516 );
not ( n27518 , n27517 );
buf ( n27519 , n27518 );
not ( n27520 , n27519 );
buf ( n27521 , n27520 );
not ( n27522 , n27053 );
and ( n27523 , n27522 , n27228 );
xor ( n27524 , n27229 , n27257 );
and ( n27525 , n27524 , n27053 );
or ( n27526 , n27523 , n27525 );
buf ( n27527 , n27526 );
not ( n27528 , n27527 );
buf ( n27529 , n27528 );
buf ( n27530 , n27529 );
not ( n27531 , n27530 );
buf ( n27532 , n27531 );
not ( n27533 , n27532 );
buf ( n27534 , n27533 );
not ( n27535 , n27053 );
and ( n27536 , n27535 , n27230 );
xor ( n27537 , n27231 , n27256 );
and ( n27538 , n27537 , n27053 );
or ( n27539 , n27536 , n27538 );
buf ( n27540 , n27539 );
not ( n27541 , n27540 );
buf ( n27542 , n27541 );
buf ( n27543 , n27542 );
not ( n27544 , n27543 );
buf ( n27545 , n27544 );
not ( n27546 , n27545 );
buf ( n27547 , n27546 );
not ( n27548 , n27053 );
and ( n27549 , n27548 , n27232 );
xor ( n27550 , n27233 , n27255 );
and ( n27551 , n27550 , n27053 );
or ( n27552 , n27549 , n27551 );
buf ( n27553 , n27552 );
not ( n27554 , n27553 );
buf ( n27555 , n27554 );
buf ( n27556 , n27555 );
and ( n27557 , C1 , n27556 );
and ( n27558 , C1 , n27557 );
and ( n27559 , C1 , n27558 );
and ( n27560 , C1 , n27559 );
and ( n27561 , C1 , n27560 );
and ( n27562 , C1 , n27561 );
and ( n27563 , C1 , n27562 );
and ( n27564 , C1 , n27563 );
and ( n27565 , C1 , n27564 );
and ( n27566 , C1 , n27565 );
and ( n27567 , C1 , n27566 );
and ( n27568 , C1 , n27567 );
and ( n27569 , C1 , n27568 );
and ( n27570 , C1 , n27569 );
and ( n27571 , C1 , n27570 );
and ( n27572 , C1 , n27571 );
and ( n27573 , C1 , n27572 );
and ( n27574 , C1 , n27573 );
and ( n27575 , C1 , n27574 );
and ( n27576 , C1 , n27575 );
and ( n27577 , C1 , n27576 );
not ( n27578 , n27577 );
buf ( n27579 , n27578 );
not ( n27580 , n27579 );
buf ( n27581 , n27580 );
not ( n27582 , n27053 );
and ( n27583 , n27582 , n27234 );
xor ( n27584 , n27235 , n27254 );
and ( n27585 , n27584 , n27053 );
or ( n27586 , n27583 , n27585 );
buf ( n27587 , n27586 );
not ( n27588 , n27587 );
buf ( n27589 , n27588 );
buf ( n27590 , n27589 );
and ( n27591 , C1 , n27590 );
and ( n27592 , C1 , n27591 );
and ( n27593 , C1 , n27592 );
and ( n27594 , C1 , n27593 );
and ( n27595 , C1 , n27594 );
and ( n27596 , C1 , n27595 );
and ( n27597 , C1 , n27596 );
and ( n27598 , C1 , n27597 );
and ( n27599 , C1 , n27598 );
and ( n27600 , C1 , n27599 );
and ( n27601 , C1 , n27600 );
and ( n27602 , C1 , n27601 );
and ( n27603 , C1 , n27602 );
and ( n27604 , C1 , n27603 );
and ( n27605 , C1 , n27604 );
and ( n27606 , C1 , n27605 );
and ( n27607 , C1 , n27606 );
and ( n27608 , C1 , n27607 );
and ( n27609 , C1 , n27608 );
and ( n27610 , C1 , n27609 );
and ( n27611 , C1 , n27610 );
buf ( n27612 , n27611 );
not ( n27613 , n27612 );
buf ( n27614 , n27613 );
not ( n27615 , n27614 );
buf ( n27616 , n27615 );
not ( n27617 , n27053 );
and ( n27618 , n27617 , n27236 );
xor ( n27619 , n27237 , n27253 );
and ( n27620 , n27619 , n27053 );
or ( n27621 , n27618 , n27620 );
buf ( n27622 , n27621 );
not ( n27623 , n27622 );
buf ( n27624 , n27623 );
buf ( n27625 , n27624 );
and ( n27626 , C1 , n27625 );
and ( n27627 , C1 , n27626 );
and ( n27628 , C1 , n27627 );
and ( n27629 , C1 , n27628 );
and ( n27630 , C1 , n27629 );
and ( n27631 , C1 , n27630 );
and ( n27632 , C1 , n27631 );
and ( n27633 , C1 , n27632 );
and ( n27634 , C1 , n27633 );
and ( n27635 , C1 , n27634 );
and ( n27636 , C1 , n27635 );
and ( n27637 , C1 , n27636 );
and ( n27638 , C1 , n27637 );
and ( n27639 , C1 , n27638 );
and ( n27640 , C1 , n27639 );
and ( n27641 , C1 , n27640 );
and ( n27642 , C1 , n27641 );
and ( n27643 , C1 , n27642 );
and ( n27644 , C1 , n27643 );
and ( n27645 , C1 , n27644 );
and ( n27646 , C1 , n27645 );
and ( n27647 , C1 , n27646 );
buf ( n27648 , n27647 );
not ( n27649 , n27648 );
buf ( n27650 , n27649 );
not ( n27651 , n27650 );
buf ( n27652 , n27651 );
not ( n27653 , n27053 );
and ( n27654 , n27653 , n27238 );
xor ( n27655 , n27239 , n27252 );
and ( n27656 , n27655 , n27053 );
or ( n27657 , n27654 , n27656 );
buf ( n27658 , n27657 );
not ( n27659 , n27658 );
buf ( n27660 , n27659 );
buf ( n27661 , n27660 );
and ( n27662 , C1 , n27661 );
and ( n27663 , C1 , n27662 );
and ( n27664 , C1 , n27663 );
and ( n27665 , C1 , n27664 );
and ( n27666 , C1 , n27665 );
and ( n27667 , C1 , n27666 );
and ( n27668 , C1 , n27667 );
and ( n27669 , C1 , n27668 );
and ( n27670 , C1 , n27669 );
and ( n27671 , C1 , n27670 );
and ( n27672 , C1 , n27671 );
and ( n27673 , C1 , n27672 );
and ( n27674 , C1 , n27673 );
and ( n27675 , C1 , n27674 );
and ( n27676 , C1 , n27675 );
and ( n27677 , C1 , n27676 );
and ( n27678 , C1 , n27677 );
and ( n27679 , C1 , n27678 );
and ( n27680 , C1 , n27679 );
and ( n27681 , C1 , n27680 );
and ( n27682 , C1 , n27681 );
and ( n27683 , C1 , n27682 );
and ( n27684 , C1 , n27683 );
buf ( n27685 , n27684 );
not ( n27686 , n27685 );
buf ( n27687 , n27686 );
not ( n27688 , n27687 );
buf ( n27689 , n27688 );
not ( n27690 , n27053 );
and ( n27691 , n27690 , n27240 );
xor ( n27692 , n27241 , n27251 );
and ( n27693 , n27692 , n27053 );
or ( n27694 , n27691 , n27693 );
buf ( n27695 , n27694 );
not ( n27696 , n27695 );
buf ( n27697 , n27696 );
buf ( n27698 , n27697 );
and ( n27699 , C1 , n27698 );
and ( n27700 , C1 , n27699 );
and ( n27701 , C1 , n27700 );
and ( n27702 , C1 , n27701 );
and ( n27703 , C1 , n27702 );
and ( n27704 , C1 , n27703 );
and ( n27705 , C1 , n27704 );
and ( n27706 , C1 , n27705 );
and ( n27707 , C1 , n27706 );
and ( n27708 , C1 , n27707 );
and ( n27709 , C1 , n27708 );
and ( n27710 , C1 , n27709 );
and ( n27711 , C1 , n27710 );
and ( n27712 , C1 , n27711 );
and ( n27713 , C1 , n27712 );
and ( n27714 , C1 , n27713 );
and ( n27715 , C1 , n27714 );
and ( n27716 , C1 , n27715 );
and ( n27717 , C1 , n27716 );
and ( n27718 , C1 , n27717 );
and ( n27719 , C1 , n27718 );
and ( n27720 , C1 , n27719 );
and ( n27721 , C1 , n27720 );
and ( n27722 , C1 , n27721 );
buf ( n27723 , n27722 );
not ( n27724 , n27723 );
buf ( n27725 , n27724 );
not ( n27726 , n27725 );
buf ( n27727 , n27726 );
not ( n27728 , n27053 );
and ( n27729 , n27728 , n27242 );
xor ( n27730 , n27243 , n27250 );
and ( n27731 , n27730 , n27053 );
or ( n27732 , n27729 , n27731 );
buf ( n27733 , n27732 );
not ( n27734 , n27733 );
buf ( n27735 , n27734 );
buf ( n27736 , n27735 );
and ( n27737 , C1 , n27736 );
and ( n27738 , C1 , n27737 );
and ( n27739 , C1 , n27738 );
and ( n27740 , C1 , n27739 );
and ( n27741 , C1 , n27740 );
and ( n27742 , C1 , n27741 );
and ( n27743 , C1 , n27742 );
and ( n27744 , C1 , n27743 );
and ( n27745 , C1 , n27744 );
and ( n27746 , C1 , n27745 );
and ( n27747 , C1 , n27746 );
and ( n27748 , C1 , n27747 );
and ( n27749 , C1 , n27748 );
and ( n27750 , C1 , n27749 );
and ( n27751 , C1 , n27750 );
and ( n27752 , C1 , n27751 );
and ( n27753 , C1 , n27752 );
and ( n27754 , C1 , n27753 );
and ( n27755 , C1 , n27754 );
and ( n27756 , C1 , n27755 );
and ( n27757 , C1 , n27756 );
and ( n27758 , C1 , n27757 );
and ( n27759 , C1 , n27758 );
and ( n27760 , C1 , n27759 );
and ( n27761 , C1 , n27760 );
buf ( n27762 , n27761 );
not ( n27763 , n27762 );
buf ( n27764 , n27763 );
not ( n27765 , n27764 );
buf ( n27766 , n27765 );
not ( n27767 , n27053 );
and ( n27768 , n27767 , n27244 );
xor ( n27769 , n27245 , n27249 );
and ( n27770 , n27769 , n27053 );
or ( n27771 , n27768 , n27770 );
buf ( n27772 , n27771 );
not ( n27773 , n27772 );
buf ( n27774 , n27773 );
buf ( n27775 , n27774 );
and ( n27776 , C1 , n27775 );
and ( n27777 , C1 , n27776 );
and ( n27778 , C1 , n27777 );
and ( n27779 , C1 , n27778 );
and ( n27780 , C1 , n27779 );
and ( n27781 , C1 , n27780 );
and ( n27782 , C1 , n27781 );
and ( n27783 , C1 , n27782 );
and ( n27784 , C1 , n27783 );
and ( n27785 , C1 , n27784 );
and ( n27786 , C1 , n27785 );
and ( n27787 , C1 , n27786 );
and ( n27788 , C1 , n27787 );
and ( n27789 , C1 , n27788 );
and ( n27790 , C1 , n27789 );
and ( n27791 , C1 , n27790 );
and ( n27792 , C1 , n27791 );
and ( n27793 , C1 , n27792 );
and ( n27794 , C1 , n27793 );
and ( n27795 , C1 , n27794 );
and ( n27796 , C1 , n27795 );
and ( n27797 , C1 , n27796 );
and ( n27798 , C1 , n27797 );
and ( n27799 , C1 , n27798 );
and ( n27800 , C1 , n27799 );
and ( n27801 , C1 , n27800 );
buf ( n27802 , n27801 );
not ( n27803 , n27802 );
buf ( n27804 , n27803 );
not ( n27805 , n27804 );
buf ( n27806 , n27805 );
not ( n27807 , n27053 );
and ( n27808 , n27807 , n27246 );
xor ( n27809 , n27247 , n27248 );
and ( n27810 , n27809 , n27053 );
or ( n27811 , n27808 , n27810 );
buf ( n27812 , n27811 );
not ( n27813 , n27812 );
buf ( n27814 , n27813 );
buf ( n27815 , n27814 );
and ( n27816 , C1 , n27815 );
and ( n27817 , C1 , n27816 );
and ( n27818 , C1 , n27817 );
and ( n27819 , C1 , n27818 );
and ( n27820 , C1 , n27819 );
and ( n27821 , C1 , n27820 );
and ( n27822 , C1 , n27821 );
and ( n27823 , C1 , n27822 );
and ( n27824 , C1 , n27823 );
and ( n27825 , C1 , n27824 );
and ( n27826 , C1 , n27825 );
and ( n27827 , C1 , n27826 );
and ( n27828 , C1 , n27827 );
and ( n27829 , C1 , n27828 );
and ( n27830 , C1 , n27829 );
and ( n27831 , C1 , n27830 );
and ( n27832 , C1 , n27831 );
and ( n27833 , C1 , n27832 );
and ( n27834 , C1 , n27833 );
and ( n27835 , C1 , n27834 );
and ( n27836 , C1 , n27835 );
and ( n27837 , C1 , n27836 );
and ( n27838 , C1 , n27837 );
and ( n27839 , C1 , n27838 );
and ( n27840 , C1 , n27839 );
and ( n27841 , C1 , n27840 );
and ( n27842 , C1 , n27841 );
buf ( n27843 , n27842 );
not ( n27844 , n27843 );
buf ( n27845 , n27844 );
not ( n27846 , n27845 );
buf ( n27847 , n27846 );
and ( n27848 , n27106 , n27149 );
and ( n27849 , n27847 , n27848 );
and ( n27850 , n27806 , n27849 );
and ( n27851 , n27766 , n27850 );
and ( n27852 , n27727 , n27851 );
and ( n27853 , n27689 , n27852 );
and ( n27854 , n27652 , n27853 );
and ( n27855 , n27616 , n27854 );
and ( n27856 , n27581 , n27855 );
and ( n27857 , n27547 , n27856 );
and ( n27858 , n27534 , n27857 );
and ( n27859 , n27521 , n27858 );
and ( n27860 , n27508 , n27859 );
and ( n27861 , n27495 , n27860 );
and ( n27862 , n27482 , n27861 );
and ( n27863 , n27469 , n27862 );
and ( n27864 , n27456 , n27863 );
and ( n27865 , n27443 , n27864 );
and ( n27866 , n27430 , n27865 );
and ( n27867 , n27417 , n27866 );
and ( n27868 , n27404 , n27867 );
and ( n27869 , n27391 , n27868 );
and ( n27870 , n27378 , n27869 );
and ( n27871 , n27365 , n27870 );
and ( n27872 , n27352 , n27871 );
and ( n27873 , n27339 , n27872 );
and ( n27874 , n27326 , n27873 );
and ( n27875 , n27313 , n27874 );
and ( n27876 , n27300 , n27875 );
and ( n27877 , n27287 , n27876 );
not ( n27878 , n27877 );
buf ( n27879 , n27878 );
and ( n27880 , n27879 , n27054 );
or ( n27881 , C0 , n27880 );
buf ( n27882 , n27881 );
buf ( n27883 , n27882 );
not ( n27884 , n27883 );
buf ( n27885 , n27154 );
and ( n27886 , n27884 , n27885 );
not ( n27887 , n27885 );
not ( n27888 , n27157 );
xor ( n27889 , n27887 , n27888 );
and ( n27890 , n27889 , n27883 );
or ( n27891 , n27886 , n27890 );
buf ( n27892 , n27891 );
not ( n27893 , n27892 );
buf ( n27894 , n27893 );
buf ( n27895 , n27894 );
not ( n27896 , n27895 );
or ( n27897 , n27162 , n27896 );
not ( n27898 , n27883 );
not ( n27899 , n27054 );
buf ( n27900 , n27845 );
and ( n27901 , n27899 , n27900 );
xor ( n27902 , n27847 , n27848 );
buf ( n27903 , n27902 );
and ( n27904 , n27903 , n27054 );
or ( n27905 , n27901 , n27904 );
buf ( n27906 , n27905 );
buf ( n27907 , n27906 );
and ( n27908 , n27898 , n27907 );
not ( n27909 , n27907 );
and ( n27910 , n27887 , n27888 );
xor ( n27911 , n27909 , n27910 );
and ( n27912 , n27911 , n27883 );
or ( n27913 , n27908 , n27912 );
buf ( n27914 , n27913 );
not ( n27915 , n27914 );
buf ( n27916 , n27915 );
buf ( n27917 , n27916 );
not ( n27918 , n27917 );
or ( n27919 , n27897 , n27918 );
not ( n27920 , n27883 );
not ( n27921 , n27054 );
buf ( n27922 , n27804 );
and ( n27923 , n27921 , n27922 );
xor ( n27924 , n27806 , n27849 );
buf ( n27925 , n27924 );
and ( n27926 , n27925 , n27054 );
or ( n27927 , n27923 , n27926 );
buf ( n27928 , n27927 );
buf ( n27929 , n27928 );
and ( n27930 , n27920 , n27929 );
not ( n27931 , n27929 );
and ( n27932 , n27909 , n27910 );
xor ( n27933 , n27931 , n27932 );
and ( n27934 , n27933 , n27883 );
or ( n27935 , n27930 , n27934 );
buf ( n27936 , n27935 );
not ( n27937 , n27936 );
buf ( n27938 , n27937 );
buf ( n27939 , n27938 );
not ( n27940 , n27939 );
or ( n27941 , n27919 , n27940 );
not ( n27942 , n27883 );
not ( n27943 , n27054 );
buf ( n27944 , n27764 );
and ( n27945 , n27943 , n27944 );
xor ( n27946 , n27766 , n27850 );
buf ( n27947 , n27946 );
and ( n27948 , n27947 , n27054 );
or ( n27949 , n27945 , n27948 );
buf ( n27950 , n27949 );
buf ( n27951 , n27950 );
and ( n27952 , n27942 , n27951 );
not ( n27953 , n27951 );
and ( n27954 , n27931 , n27932 );
xor ( n27955 , n27953 , n27954 );
and ( n27956 , n27955 , n27883 );
or ( n27957 , n27952 , n27956 );
buf ( n27958 , n27957 );
not ( n27959 , n27958 );
buf ( n27960 , n27959 );
buf ( n27961 , n27960 );
not ( n27962 , n27961 );
or ( n27963 , n27941 , n27962 );
not ( n27964 , n27883 );
not ( n27965 , n27054 );
buf ( n27966 , n27725 );
and ( n27967 , n27965 , n27966 );
xor ( n27968 , n27727 , n27851 );
buf ( n27969 , n27968 );
and ( n27970 , n27969 , n27054 );
or ( n27971 , n27967 , n27970 );
buf ( n27972 , n27971 );
buf ( n27973 , n27972 );
and ( n27974 , n27964 , n27973 );
not ( n27975 , n27973 );
and ( n27976 , n27953 , n27954 );
xor ( n27977 , n27975 , n27976 );
and ( n27978 , n27977 , n27883 );
or ( n27979 , n27974 , n27978 );
buf ( n27980 , n27979 );
not ( n27981 , n27980 );
buf ( n27982 , n27981 );
buf ( n27983 , n27982 );
not ( n27984 , n27983 );
or ( n27985 , n27963 , n27984 );
not ( n27986 , n27883 );
not ( n27987 , n27054 );
buf ( n27988 , n27687 );
and ( n27989 , n27987 , n27988 );
xor ( n27990 , n27689 , n27852 );
buf ( n27991 , n27990 );
and ( n27992 , n27991 , n27054 );
or ( n27993 , n27989 , n27992 );
buf ( n27994 , n27993 );
buf ( n27995 , n27994 );
and ( n27996 , n27986 , n27995 );
not ( n27997 , n27995 );
and ( n27998 , n27975 , n27976 );
xor ( n27999 , n27997 , n27998 );
and ( n28000 , n27999 , n27883 );
or ( n28001 , n27996 , n28000 );
buf ( n28002 , n28001 );
not ( n28003 , n28002 );
buf ( n28004 , n28003 );
buf ( n28005 , n28004 );
not ( n28006 , n28005 );
or ( n28007 , n27985 , n28006 );
not ( n28008 , n27883 );
not ( n28009 , n27054 );
buf ( n28010 , n27650 );
and ( n28011 , n28009 , n28010 );
xor ( n28012 , n27652 , n27853 );
buf ( n28013 , n28012 );
and ( n28014 , n28013 , n27054 );
or ( n28015 , n28011 , n28014 );
buf ( n28016 , n28015 );
buf ( n28017 , n28016 );
and ( n28018 , n28008 , n28017 );
not ( n28019 , n28017 );
and ( n28020 , n27997 , n27998 );
xor ( n28021 , n28019 , n28020 );
and ( n28022 , n28021 , n27883 );
or ( n28023 , n28018 , n28022 );
buf ( n28024 , n28023 );
not ( n28025 , n28024 );
buf ( n28026 , n28025 );
buf ( n28027 , n28026 );
not ( n28028 , n28027 );
or ( n28029 , n28007 , n28028 );
not ( n28030 , n27883 );
not ( n28031 , n27054 );
buf ( n28032 , n27614 );
and ( n28033 , n28031 , n28032 );
xor ( n28034 , n27616 , n27854 );
buf ( n28035 , n28034 );
and ( n28036 , n28035 , n27054 );
or ( n28037 , n28033 , n28036 );
buf ( n28038 , n28037 );
buf ( n28039 , n28038 );
and ( n28040 , n28030 , n28039 );
not ( n28041 , n28039 );
and ( n28042 , n28019 , n28020 );
xor ( n28043 , n28041 , n28042 );
and ( n28044 , n28043 , n27883 );
or ( n28045 , n28040 , n28044 );
buf ( n28046 , n28045 );
not ( n28047 , n28046 );
buf ( n28048 , n28047 );
buf ( n28049 , n28048 );
not ( n28050 , n28049 );
or ( n28051 , n28029 , n28050 );
not ( n28052 , n27883 );
not ( n28053 , n27054 );
buf ( n28054 , n27579 );
and ( n28055 , n28053 , n28054 );
xor ( n28056 , n27581 , n27855 );
buf ( n28057 , n28056 );
and ( n28058 , n28057 , n27054 );
or ( n28059 , n28055 , n28058 );
buf ( n28060 , n28059 );
buf ( n28061 , n28060 );
and ( n28062 , n28052 , n28061 );
not ( n28063 , n28061 );
and ( n28064 , n28041 , n28042 );
xor ( n28065 , n28063 , n28064 );
and ( n28066 , n28065 , n27883 );
or ( n28067 , n28062 , n28066 );
buf ( n28068 , n28067 );
not ( n28069 , n28068 );
buf ( n28070 , n28069 );
buf ( n28071 , n28070 );
not ( n28072 , n28071 );
or ( n28073 , n28051 , n28072 );
not ( n28074 , n27883 );
not ( n28075 , n27054 );
buf ( n28076 , n27545 );
and ( n28077 , n28075 , n28076 );
xor ( n28078 , n27547 , n27856 );
buf ( n28079 , n28078 );
and ( n28080 , n28079 , n27054 );
or ( n28081 , n28077 , n28080 );
buf ( n28082 , n28081 );
buf ( n28083 , n28082 );
and ( n28084 , n28074 , n28083 );
not ( n28085 , n28083 );
and ( n28086 , n28063 , n28064 );
xor ( n28087 , n28085 , n28086 );
and ( n28088 , n28087 , n27883 );
or ( n28089 , n28084 , n28088 );
buf ( n28090 , n28089 );
not ( n28091 , n28090 );
buf ( n28092 , n28091 );
buf ( n28093 , n28092 );
not ( n28094 , n28093 );
or ( n28095 , n28073 , n28094 );
not ( n28096 , n27883 );
not ( n28097 , n27054 );
buf ( n28098 , n27532 );
and ( n28099 , n28097 , n28098 );
xor ( n28100 , n27534 , n27857 );
buf ( n28101 , n28100 );
and ( n28102 , n28101 , n27054 );
or ( n28103 , n28099 , n28102 );
buf ( n28104 , n28103 );
buf ( n28105 , n28104 );
and ( n28106 , n28096 , n28105 );
not ( n28107 , n28105 );
and ( n28108 , n28085 , n28086 );
xor ( n28109 , n28107 , n28108 );
and ( n28110 , n28109 , n27883 );
or ( n28111 , n28106 , n28110 );
buf ( n28112 , n28111 );
not ( n28113 , n28112 );
buf ( n28114 , n28113 );
buf ( n28115 , n28114 );
not ( n28116 , n28115 );
or ( n28117 , n28095 , n28116 );
not ( n28118 , n27883 );
not ( n28119 , n27054 );
buf ( n28120 , n27519 );
and ( n28121 , n28119 , n28120 );
xor ( n28122 , n27521 , n27858 );
buf ( n28123 , n28122 );
and ( n28124 , n28123 , n27054 );
or ( n28125 , n28121 , n28124 );
buf ( n28126 , n28125 );
buf ( n28127 , n28126 );
and ( n28128 , n28118 , n28127 );
not ( n28129 , n28127 );
and ( n28130 , n28107 , n28108 );
xor ( n28131 , n28129 , n28130 );
and ( n28132 , n28131 , n27883 );
or ( n28133 , n28128 , n28132 );
buf ( n28134 , n28133 );
not ( n28135 , n28134 );
buf ( n28136 , n28135 );
buf ( n28137 , n28136 );
not ( n28138 , n28137 );
or ( n28139 , n28117 , n28138 );
not ( n28140 , n27883 );
not ( n28141 , n27054 );
buf ( n28142 , n27506 );
and ( n28143 , n28141 , n28142 );
xor ( n28144 , n27508 , n27859 );
buf ( n28145 , n28144 );
and ( n28146 , n28145 , n27054 );
or ( n28147 , n28143 , n28146 );
buf ( n28148 , n28147 );
buf ( n28149 , n28148 );
and ( n28150 , n28140 , n28149 );
not ( n28151 , n28149 );
and ( n28152 , n28129 , n28130 );
xor ( n28153 , n28151 , n28152 );
and ( n28154 , n28153 , n27883 );
or ( n28155 , n28150 , n28154 );
buf ( n28156 , n28155 );
not ( n28157 , n28156 );
buf ( n28158 , n28157 );
buf ( n28159 , n28158 );
not ( n28160 , n28159 );
or ( n28161 , n28139 , n28160 );
not ( n28162 , n27883 );
not ( n28163 , n27054 );
buf ( n28164 , n27493 );
and ( n28165 , n28163 , n28164 );
xor ( n28166 , n27495 , n27860 );
buf ( n28167 , n28166 );
and ( n28168 , n28167 , n27054 );
or ( n28169 , n28165 , n28168 );
buf ( n28170 , n28169 );
buf ( n28171 , n28170 );
and ( n28172 , n28162 , n28171 );
not ( n28173 , n28171 );
and ( n28174 , n28151 , n28152 );
xor ( n28175 , n28173 , n28174 );
and ( n28176 , n28175 , n27883 );
or ( n28177 , n28172 , n28176 );
buf ( n28178 , n28177 );
not ( n28179 , n28178 );
buf ( n28180 , n28179 );
buf ( n28181 , n28180 );
not ( n28182 , n28181 );
or ( n28183 , n28161 , n28182 );
not ( n28184 , n27883 );
not ( n28185 , n27054 );
buf ( n28186 , n27480 );
and ( n28187 , n28185 , n28186 );
xor ( n28188 , n27482 , n27861 );
buf ( n28189 , n28188 );
and ( n28190 , n28189 , n27054 );
or ( n28191 , n28187 , n28190 );
buf ( n28192 , n28191 );
buf ( n28193 , n28192 );
and ( n28194 , n28184 , n28193 );
not ( n28195 , n28193 );
and ( n28196 , n28173 , n28174 );
xor ( n28197 , n28195 , n28196 );
and ( n28198 , n28197 , n27883 );
or ( n28199 , n28194 , n28198 );
buf ( n28200 , n28199 );
not ( n28201 , n28200 );
buf ( n28202 , n28201 );
buf ( n28203 , n28202 );
not ( n28204 , n28203 );
or ( n28205 , n28183 , n28204 );
not ( n28206 , n27883 );
not ( n28207 , n27054 );
buf ( n28208 , n27467 );
and ( n28209 , n28207 , n28208 );
xor ( n28210 , n27469 , n27862 );
buf ( n28211 , n28210 );
and ( n28212 , n28211 , n27054 );
or ( n28213 , n28209 , n28212 );
buf ( n28214 , n28213 );
buf ( n28215 , n28214 );
and ( n28216 , n28206 , n28215 );
not ( n28217 , n28215 );
and ( n28218 , n28195 , n28196 );
xor ( n28219 , n28217 , n28218 );
and ( n28220 , n28219 , n27883 );
or ( n28221 , n28216 , n28220 );
buf ( n28222 , n28221 );
not ( n28223 , n28222 );
buf ( n28224 , n28223 );
buf ( n28225 , n28224 );
not ( n28226 , n28225 );
or ( n28227 , n28205 , n28226 );
not ( n28228 , n27883 );
not ( n28229 , n27054 );
buf ( n28230 , n27454 );
and ( n28231 , n28229 , n28230 );
xor ( n28232 , n27456 , n27863 );
buf ( n28233 , n28232 );
and ( n28234 , n28233 , n27054 );
or ( n28235 , n28231 , n28234 );
buf ( n28236 , n28235 );
buf ( n28237 , n28236 );
and ( n28238 , n28228 , n28237 );
not ( n28239 , n28237 );
and ( n28240 , n28217 , n28218 );
xor ( n28241 , n28239 , n28240 );
and ( n28242 , n28241 , n27883 );
or ( n28243 , n28238 , n28242 );
buf ( n28244 , n28243 );
not ( n28245 , n28244 );
buf ( n28246 , n28245 );
buf ( n28247 , n28246 );
not ( n28248 , n28247 );
or ( n28249 , n28227 , n28248 );
not ( n28250 , n27883 );
not ( n28251 , n27054 );
buf ( n28252 , n27441 );
and ( n28253 , n28251 , n28252 );
xor ( n28254 , n27443 , n27864 );
buf ( n28255 , n28254 );
and ( n28256 , n28255 , n27054 );
or ( n28257 , n28253 , n28256 );
buf ( n28258 , n28257 );
buf ( n28259 , n28258 );
and ( n28260 , n28250 , n28259 );
not ( n28261 , n28259 );
and ( n28262 , n28239 , n28240 );
xor ( n28263 , n28261 , n28262 );
and ( n28264 , n28263 , n27883 );
or ( n28265 , n28260 , n28264 );
buf ( n28266 , n28265 );
not ( n28267 , n28266 );
buf ( n28268 , n28267 );
buf ( n28269 , n28268 );
not ( n28270 , n28269 );
or ( n28271 , n28249 , n28270 );
not ( n28272 , n27883 );
not ( n28273 , n27054 );
buf ( n28274 , n27428 );
and ( n28275 , n28273 , n28274 );
xor ( n28276 , n27430 , n27865 );
buf ( n28277 , n28276 );
and ( n28278 , n28277 , n27054 );
or ( n28279 , n28275 , n28278 );
buf ( n28280 , n28279 );
buf ( n28281 , n28280 );
and ( n28282 , n28272 , n28281 );
not ( n28283 , n28281 );
and ( n28284 , n28261 , n28262 );
xor ( n28285 , n28283 , n28284 );
and ( n28286 , n28285 , n27883 );
or ( n28287 , n28282 , n28286 );
buf ( n28288 , n28287 );
not ( n28289 , n28288 );
buf ( n28290 , n28289 );
buf ( n28291 , n28290 );
not ( n28292 , n28291 );
or ( n28293 , n28271 , n28292 );
not ( n28294 , n27883 );
not ( n28295 , n27054 );
buf ( n28296 , n27415 );
and ( n28297 , n28295 , n28296 );
xor ( n28298 , n27417 , n27866 );
buf ( n28299 , n28298 );
and ( n28300 , n28299 , n27054 );
or ( n28301 , n28297 , n28300 );
buf ( n28302 , n28301 );
buf ( n28303 , n28302 );
and ( n28304 , n28294 , n28303 );
not ( n28305 , n28303 );
and ( n28306 , n28283 , n28284 );
xor ( n28307 , n28305 , n28306 );
and ( n28308 , n28307 , n27883 );
or ( n28309 , n28304 , n28308 );
buf ( n28310 , n28309 );
not ( n28311 , n28310 );
buf ( n28312 , n28311 );
buf ( n28313 , n28312 );
not ( n28314 , n28313 );
or ( n28315 , n28293 , n28314 );
not ( n28316 , n27883 );
not ( n28317 , n27054 );
buf ( n28318 , n27402 );
and ( n28319 , n28317 , n28318 );
xor ( n28320 , n27404 , n27867 );
buf ( n28321 , n28320 );
and ( n28322 , n28321 , n27054 );
or ( n28323 , n28319 , n28322 );
buf ( n28324 , n28323 );
buf ( n28325 , n28324 );
and ( n28326 , n28316 , n28325 );
not ( n28327 , n28325 );
and ( n28328 , n28305 , n28306 );
xor ( n28329 , n28327 , n28328 );
and ( n28330 , n28329 , n27883 );
or ( n28331 , n28326 , n28330 );
buf ( n28332 , n28331 );
not ( n28333 , n28332 );
buf ( n28334 , n28333 );
buf ( n28335 , n28334 );
not ( n28336 , n28335 );
or ( n28337 , n28315 , n28336 );
not ( n28338 , n27883 );
not ( n28339 , n27054 );
buf ( n28340 , n27389 );
and ( n28341 , n28339 , n28340 );
xor ( n28342 , n27391 , n27868 );
buf ( n28343 , n28342 );
and ( n28344 , n28343 , n27054 );
or ( n28345 , n28341 , n28344 );
buf ( n28346 , n28345 );
buf ( n28347 , n28346 );
and ( n28348 , n28338 , n28347 );
not ( n28349 , n28347 );
and ( n28350 , n28327 , n28328 );
xor ( n28351 , n28349 , n28350 );
and ( n28352 , n28351 , n27883 );
or ( n28353 , n28348 , n28352 );
buf ( n28354 , n28353 );
not ( n28355 , n28354 );
buf ( n28356 , n28355 );
buf ( n28357 , n28356 );
not ( n28358 , n28357 );
or ( n28359 , n28337 , n28358 );
not ( n28360 , n27883 );
not ( n28361 , n27054 );
buf ( n28362 , n27376 );
and ( n28363 , n28361 , n28362 );
xor ( n28364 , n27378 , n27869 );
buf ( n28365 , n28364 );
and ( n28366 , n28365 , n27054 );
or ( n28367 , n28363 , n28366 );
buf ( n28368 , n28367 );
buf ( n28369 , n28368 );
and ( n28370 , n28360 , n28369 );
not ( n28371 , n28369 );
and ( n28372 , n28349 , n28350 );
xor ( n28373 , n28371 , n28372 );
and ( n28374 , n28373 , n27883 );
or ( n28375 , n28370 , n28374 );
buf ( n28376 , n28375 );
not ( n28377 , n28376 );
buf ( n28378 , n28377 );
buf ( n28379 , n28378 );
not ( n28380 , n28379 );
or ( n28381 , n28359 , n28380 );
not ( n28382 , n27883 );
not ( n28383 , n27054 );
buf ( n28384 , n27363 );
and ( n28385 , n28383 , n28384 );
xor ( n28386 , n27365 , n27870 );
buf ( n28387 , n28386 );
and ( n28388 , n28387 , n27054 );
or ( n28389 , n28385 , n28388 );
buf ( n28390 , n28389 );
buf ( n28391 , n28390 );
and ( n28392 , n28382 , n28391 );
not ( n28393 , n28391 );
and ( n28394 , n28371 , n28372 );
xor ( n28395 , n28393 , n28394 );
and ( n28396 , n28395 , n27883 );
or ( n28397 , n28392 , n28396 );
buf ( n28398 , n28397 );
not ( n28399 , n28398 );
buf ( n28400 , n28399 );
buf ( n28401 , n28400 );
not ( n28402 , n28401 );
or ( n28403 , n28381 , n28402 );
not ( n28404 , n27883 );
not ( n28405 , n27054 );
buf ( n28406 , n27350 );
and ( n28407 , n28405 , n28406 );
xor ( n28408 , n27352 , n27871 );
buf ( n28409 , n28408 );
and ( n28410 , n28409 , n27054 );
or ( n28411 , n28407 , n28410 );
buf ( n28412 , n28411 );
buf ( n28413 , n28412 );
and ( n28414 , n28404 , n28413 );
not ( n28415 , n28413 );
and ( n28416 , n28393 , n28394 );
xor ( n28417 , n28415 , n28416 );
and ( n28418 , n28417 , n27883 );
or ( n28419 , n28414 , n28418 );
buf ( n28420 , n28419 );
not ( n28421 , n28420 );
buf ( n28422 , n28421 );
buf ( n28423 , n28422 );
not ( n28424 , n28423 );
or ( n28425 , n28403 , n28424 );
not ( n28426 , n27883 );
not ( n28427 , n27054 );
buf ( n28428 , n27337 );
and ( n28429 , n28427 , n28428 );
xor ( n28430 , n27339 , n27872 );
buf ( n28431 , n28430 );
and ( n28432 , n28431 , n27054 );
or ( n28433 , n28429 , n28432 );
buf ( n28434 , n28433 );
buf ( n28435 , n28434 );
and ( n28436 , n28426 , n28435 );
not ( n28437 , n28435 );
and ( n28438 , n28415 , n28416 );
xor ( n28439 , n28437 , n28438 );
and ( n28440 , n28439 , n27883 );
or ( n28441 , n28436 , n28440 );
buf ( n28442 , n28441 );
not ( n28443 , n28442 );
buf ( n28444 , n28443 );
buf ( n28445 , n28444 );
not ( n28446 , n28445 );
or ( n28447 , n28425 , n28446 );
not ( n28448 , n27883 );
not ( n28449 , n27054 );
buf ( n28450 , n27324 );
and ( n28451 , n28449 , n28450 );
xor ( n28452 , n27326 , n27873 );
buf ( n28453 , n28452 );
and ( n28454 , n28453 , n27054 );
or ( n28455 , n28451 , n28454 );
buf ( n28456 , n28455 );
buf ( n28457 , n28456 );
and ( n28458 , n28448 , n28457 );
not ( n28459 , n28457 );
and ( n28460 , n28437 , n28438 );
xor ( n28461 , n28459 , n28460 );
and ( n28462 , n28461 , n27883 );
or ( n28463 , n28458 , n28462 );
buf ( n28464 , n28463 );
not ( n28465 , n28464 );
buf ( n28466 , n28465 );
buf ( n28467 , n28466 );
not ( n28468 , n28467 );
or ( n28469 , n28447 , n28468 );
not ( n28470 , n27883 );
not ( n28471 , n27054 );
buf ( n28472 , n27311 );
and ( n28473 , n28471 , n28472 );
xor ( n28474 , n27313 , n27874 );
buf ( n28475 , n28474 );
and ( n28476 , n28475 , n27054 );
or ( n28477 , n28473 , n28476 );
buf ( n28478 , n28477 );
buf ( n28479 , n28478 );
and ( n28480 , n28470 , n28479 );
not ( n28481 , n28479 );
and ( n28482 , n28459 , n28460 );
xor ( n28483 , n28481 , n28482 );
and ( n28484 , n28483 , n27883 );
or ( n28485 , n28480 , n28484 );
buf ( n28486 , n28485 );
not ( n28487 , n28486 );
buf ( n28488 , n28487 );
buf ( n28489 , n28488 );
not ( n28490 , n28489 );
or ( n28491 , n28469 , n28490 );
buf ( n28492 , n28491 );
buf ( n28493 , n28492 );
and ( n28494 , n28493 , n27883 );
not ( n28495 , n28494 );
and ( n28496 , n28495 , n27896 );
xor ( n28497 , n27896 , n27883 );
xor ( n28498 , n27162 , n27883 );
and ( n28499 , n28498 , n27883 );
xor ( n28500 , n28497 , n28499 );
and ( n28501 , n28500 , n28494 );
or ( n28502 , n28496 , n28501 );
buf ( n28503 , n28502 );
and ( n28504 , n28503 , n27051 );
or ( n28505 , n27155 , n28504 );
nor ( n28506 , n27048 , n27045 );
and ( n28507 , n28505 , n28506 );
nor ( n28508 , n27037 , n27045 );
and ( n28509 , n27154 , n28508 );
or ( n28510 , n27047 , n27050 , n28507 , n28509 );
not ( n28511 , n24782 );
not ( n28512 , n24798 );
nor ( n28513 , n28511 , n24790 , n28512 );
not ( n28514 , n28513 );
nor ( n28515 , n24782 , n24790 , n28512 );
not ( n28516 , n28515 );
and ( n28517 , n24782 , n24790 , n28512 );
not ( n28518 , n28517 );
and ( n28519 , n28511 , n24790 , n28512 );
not ( n28520 , n28519 );
nor ( n28521 , n28511 , n24790 , n24798 );
not ( n28522 , n28521 );
nor ( n28523 , n24782 , n24790 , n24798 );
not ( n28524 , n28523 );
buf ( n28525 , RI210bd668_302);
and ( n28526 , n28524 , n28525 );
or ( n28527 , n28526 , C0 );
and ( n28528 , n28522 , n28527 );
and ( n28529 , C1 , n28521 );
or ( n28530 , n28528 , n28529 );
and ( n28531 , n28520 , n28530 );
or ( n28532 , n28531 , C0 );
and ( n28533 , n28518 , n28532 );
and ( n28534 , C1 , n28517 );
or ( n28535 , n28533 , n28534 );
and ( n28536 , n28516 , n28535 );
not ( n28537 , n27051 );
and ( n28538 , n28537 , n28525 );
and ( n28539 , C1 , n27051 );
or ( n28540 , n28538 , n28539 );
and ( n28541 , n28540 , n28515 );
or ( n28542 , n28536 , n28541 );
and ( n28543 , n28514 , n28542 );
not ( n28544 , n27051 );
not ( n28545 , n28544 );
and ( n28546 , n28545 , n28525 );
and ( n28547 , C1 , n28544 );
or ( n28548 , n28546 , n28547 );
and ( n28549 , n28548 , n28513 );
or ( n28550 , n28543 , n28549 );
not ( n28551 , n28513 );
not ( n28552 , n28515 );
not ( n28553 , n28517 );
not ( n28554 , n28519 );
not ( n28555 , n28521 );
not ( n28556 , n28523 );
buf ( n28557 , RI210bcdf8_303);
and ( n28558 , n28556 , n28557 );
or ( n28559 , n28558 , C0 );
and ( n28560 , n28555 , n28559 );
or ( n28561 , n28560 , C0 );
and ( n28562 , n28554 , n28561 );
and ( n28563 , C1 , n28519 );
or ( n28564 , n28562 , n28563 );
and ( n28565 , n28553 , n28564 );
and ( n28566 , C1 , n28517 );
or ( n28567 , n28565 , n28566 );
and ( n28568 , n28552 , n28567 );
not ( n28569 , n27051 );
and ( n28570 , n28569 , n28557 );
and ( n28571 , C1 , n27051 );
or ( n28572 , n28570 , n28571 );
and ( n28573 , n28572 , n28515 );
or ( n28574 , n28568 , n28573 );
and ( n28575 , n28551 , n28574 );
not ( n28576 , n28544 );
and ( n28577 , n28576 , n28557 );
and ( n28578 , C1 , n28544 );
or ( n28579 , n28577 , n28578 );
and ( n28580 , n28579 , n28513 );
or ( n28581 , n28575 , n28580 );
not ( n28582 , n28581 );
nor ( n28583 , n28550 , n28582 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n28584 , n28510 , n28583 );
not ( n28585 , n28550 );
nor ( n28586 , n28585 , n28581 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
nor ( n28587 , n28550 , n28581 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
or ( n28588 , n28586 , n28587 );
nor ( n28589 , n28585 , n28582 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
or ( n28590 , n28588 , n28589 );
or ( n28591 , n28590 , C0 );
and ( n28592 , n24802 , n28591 );
or ( n28593 , n28584 , n28592 );
and ( n28594 , n25218 , n25200 , n25208 , n25216 );
and ( n28595 , n28593 , n28594 );
buf ( n28596 , n25863 );
not ( n28597 , n14641 );
buf ( n28598 , n14831 );
buf ( n28599 , n15852 );
xor ( n28600 , n28598 , n28599 );
buf ( n28601 , n28600 );
and ( n28602 , n28597 , n28601 );
and ( n28603 , n14831 , n14641 );
or ( n28604 , n28602 , n28603 );
or ( n28605 , n28506 , n27049 );
or ( n28606 , n28605 , n27046 );
and ( n28607 , n28604 , n28606 );
buf ( n28608 , n24249 );
buf ( n28609 , n28608 );
not ( n28610 , n28609 );
buf ( n28611 , n28610 );
buf ( n28612 , n28611 );
not ( n28613 , n28612 );
buf ( n28614 , n24061 );
not ( n28615 , n28614 );
buf ( n28616 , n24246 );
and ( n28617 , n28615 , n28616 );
not ( n28618 , n28616 );
not ( n28619 , n28608 );
xor ( n28620 , n28618 , n28619 );
and ( n28621 , n28620 , n28614 );
or ( n28622 , n28617 , n28621 );
buf ( n28623 , n28622 );
not ( n28624 , n28623 );
buf ( n28625 , n28624 );
buf ( n28626 , n28625 );
not ( n28627 , n28626 );
or ( n28628 , n28613 , n28627 );
not ( n28629 , n28614 );
buf ( n28630 , n24238 );
and ( n28631 , n28629 , n28630 );
not ( n28632 , n28630 );
and ( n28633 , n28618 , n28619 );
xor ( n28634 , n28632 , n28633 );
and ( n28635 , n28634 , n28614 );
or ( n28636 , n28631 , n28635 );
buf ( n28637 , n28636 );
not ( n28638 , n28637 );
buf ( n28639 , n28638 );
buf ( n28640 , n28639 );
not ( n28641 , n28640 );
or ( n28642 , n28628 , n28641 );
not ( n28643 , n28614 );
buf ( n28644 , n24230 );
and ( n28645 , n28643 , n28644 );
not ( n28646 , n28644 );
and ( n28647 , n28632 , n28633 );
xor ( n28648 , n28646 , n28647 );
and ( n28649 , n28648 , n28614 );
or ( n28650 , n28645 , n28649 );
buf ( n28651 , n28650 );
not ( n28652 , n28651 );
buf ( n28653 , n28652 );
buf ( n28654 , n28653 );
not ( n28655 , n28654 );
or ( n28656 , n28642 , n28655 );
not ( n28657 , n28614 );
buf ( n28658 , n24222 );
and ( n28659 , n28657 , n28658 );
not ( n28660 , n28658 );
and ( n28661 , n28646 , n28647 );
xor ( n28662 , n28660 , n28661 );
and ( n28663 , n28662 , n28614 );
or ( n28664 , n28659 , n28663 );
buf ( n28665 , n28664 );
not ( n28666 , n28665 );
buf ( n28667 , n28666 );
buf ( n28668 , n28667 );
not ( n28669 , n28668 );
or ( n28670 , n28656 , n28669 );
not ( n28671 , n28614 );
buf ( n28672 , n24214 );
and ( n28673 , n28671 , n28672 );
not ( n28674 , n28672 );
and ( n28675 , n28660 , n28661 );
xor ( n28676 , n28674 , n28675 );
and ( n28677 , n28676 , n28614 );
or ( n28678 , n28673 , n28677 );
buf ( n28679 , n28678 );
not ( n28680 , n28679 );
buf ( n28681 , n28680 );
buf ( n28682 , n28681 );
not ( n28683 , n28682 );
or ( n28684 , n28670 , n28683 );
not ( n28685 , n28614 );
buf ( n28686 , n24206 );
and ( n28687 , n28685 , n28686 );
not ( n28688 , n28686 );
and ( n28689 , n28674 , n28675 );
xor ( n28690 , n28688 , n28689 );
and ( n28691 , n28690 , n28614 );
or ( n28692 , n28687 , n28691 );
buf ( n28693 , n28692 );
not ( n28694 , n28693 );
buf ( n28695 , n28694 );
buf ( n28696 , n28695 );
not ( n28697 , n28696 );
or ( n28698 , n28684 , n28697 );
not ( n28699 , n28614 );
buf ( n28700 , n24198 );
and ( n28701 , n28699 , n28700 );
not ( n28702 , n28700 );
and ( n28703 , n28688 , n28689 );
xor ( n28704 , n28702 , n28703 );
and ( n28705 , n28704 , n28614 );
or ( n28706 , n28701 , n28705 );
buf ( n28707 , n28706 );
not ( n28708 , n28707 );
buf ( n28709 , n28708 );
buf ( n28710 , n28709 );
not ( n28711 , n28710 );
or ( n28712 , n28698 , n28711 );
not ( n28713 , n28614 );
buf ( n28714 , n24190 );
and ( n28715 , n28713 , n28714 );
not ( n28716 , n28714 );
and ( n28717 , n28702 , n28703 );
xor ( n28718 , n28716 , n28717 );
and ( n28719 , n28718 , n28614 );
or ( n28720 , n28715 , n28719 );
buf ( n28721 , n28720 );
not ( n28722 , n28721 );
buf ( n28723 , n28722 );
buf ( n28724 , n28723 );
not ( n28725 , n28724 );
or ( n28726 , n28712 , n28725 );
not ( n28727 , n28614 );
buf ( n28728 , n24182 );
and ( n28729 , n28727 , n28728 );
not ( n28730 , n28728 );
and ( n28731 , n28716 , n28717 );
xor ( n28732 , n28730 , n28731 );
and ( n28733 , n28732 , n28614 );
or ( n28734 , n28729 , n28733 );
buf ( n28735 , n28734 );
not ( n28736 , n28735 );
buf ( n28737 , n28736 );
buf ( n28738 , n28737 );
not ( n28739 , n28738 );
or ( n28740 , n28726 , n28739 );
not ( n28741 , n28614 );
buf ( n28742 , n24174 );
and ( n28743 , n28741 , n28742 );
not ( n28744 , n28742 );
and ( n28745 , n28730 , n28731 );
xor ( n28746 , n28744 , n28745 );
and ( n28747 , n28746 , n28614 );
or ( n28748 , n28743 , n28747 );
buf ( n28749 , n28748 );
not ( n28750 , n28749 );
buf ( n28751 , n28750 );
buf ( n28752 , n28751 );
not ( n28753 , n28752 );
or ( n28754 , n28740 , n28753 );
not ( n28755 , n28614 );
buf ( n28756 , n24166 );
and ( n28757 , n28755 , n28756 );
not ( n28758 , n28756 );
and ( n28759 , n28744 , n28745 );
xor ( n28760 , n28758 , n28759 );
and ( n28761 , n28760 , n28614 );
or ( n28762 , n28757 , n28761 );
buf ( n28763 , n28762 );
not ( n28764 , n28763 );
buf ( n28765 , n28764 );
buf ( n28766 , n28765 );
not ( n28767 , n28766 );
or ( n28768 , n28754 , n28767 );
not ( n28769 , n28614 );
buf ( n28770 , n24158 );
and ( n28771 , n28769 , n28770 );
not ( n28772 , n28770 );
and ( n28773 , n28758 , n28759 );
xor ( n28774 , n28772 , n28773 );
and ( n28775 , n28774 , n28614 );
or ( n28776 , n28771 , n28775 );
buf ( n28777 , n28776 );
not ( n28778 , n28777 );
buf ( n28779 , n28778 );
buf ( n28780 , n28779 );
not ( n28781 , n28780 );
or ( n28782 , n28768 , n28781 );
not ( n28783 , n28614 );
buf ( n28784 , n24150 );
and ( n28785 , n28783 , n28784 );
not ( n28786 , n28784 );
and ( n28787 , n28772 , n28773 );
xor ( n28788 , n28786 , n28787 );
and ( n28789 , n28788 , n28614 );
or ( n28790 , n28785 , n28789 );
buf ( n28791 , n28790 );
not ( n28792 , n28791 );
buf ( n28793 , n28792 );
buf ( n28794 , n28793 );
not ( n28795 , n28794 );
or ( n28796 , n28782 , n28795 );
not ( n28797 , n28614 );
buf ( n28798 , n24142 );
and ( n28799 , n28797 , n28798 );
not ( n28800 , n28798 );
and ( n28801 , n28786 , n28787 );
xor ( n28802 , n28800 , n28801 );
and ( n28803 , n28802 , n28614 );
or ( n28804 , n28799 , n28803 );
buf ( n28805 , n28804 );
not ( n28806 , n28805 );
buf ( n28807 , n28806 );
buf ( n28808 , n28807 );
not ( n28809 , n28808 );
or ( n28810 , n28796 , n28809 );
not ( n28811 , n28614 );
buf ( n28812 , n24134 );
and ( n28813 , n28811 , n28812 );
not ( n28814 , n28812 );
and ( n28815 , n28800 , n28801 );
xor ( n28816 , n28814 , n28815 );
and ( n28817 , n28816 , n28614 );
or ( n28818 , n28813 , n28817 );
buf ( n28819 , n28818 );
not ( n28820 , n28819 );
buf ( n28821 , n28820 );
buf ( n28822 , n28821 );
not ( n28823 , n28822 );
or ( n28824 , n28810 , n28823 );
not ( n28825 , n28614 );
buf ( n28826 , n24126 );
and ( n28827 , n28825 , n28826 );
not ( n28828 , n28826 );
and ( n28829 , n28814 , n28815 );
xor ( n28830 , n28828 , n28829 );
and ( n28831 , n28830 , n28614 );
or ( n28832 , n28827 , n28831 );
buf ( n28833 , n28832 );
not ( n28834 , n28833 );
buf ( n28835 , n28834 );
buf ( n28836 , n28835 );
not ( n28837 , n28836 );
or ( n28838 , n28824 , n28837 );
not ( n28839 , n28614 );
buf ( n28840 , n24118 );
and ( n28841 , n28839 , n28840 );
not ( n28842 , n28840 );
and ( n28843 , n28828 , n28829 );
xor ( n28844 , n28842 , n28843 );
and ( n28845 , n28844 , n28614 );
or ( n28846 , n28841 , n28845 );
buf ( n28847 , n28846 );
not ( n28848 , n28847 );
buf ( n28849 , n28848 );
buf ( n28850 , n28849 );
not ( n28851 , n28850 );
or ( n28852 , n28838 , n28851 );
not ( n28853 , n28614 );
buf ( n28854 , n24110 );
and ( n28855 , n28853 , n28854 );
not ( n28856 , n28854 );
and ( n28857 , n28842 , n28843 );
xor ( n28858 , n28856 , n28857 );
and ( n28859 , n28858 , n28614 );
or ( n28860 , n28855 , n28859 );
buf ( n28861 , n28860 );
not ( n28862 , n28861 );
buf ( n28863 , n28862 );
buf ( n28864 , n28863 );
not ( n28865 , n28864 );
or ( n28866 , n28852 , n28865 );
not ( n28867 , n28614 );
buf ( n28868 , n24102 );
and ( n28869 , n28867 , n28868 );
not ( n28870 , n28868 );
and ( n28871 , n28856 , n28857 );
xor ( n28872 , n28870 , n28871 );
and ( n28873 , n28872 , n28614 );
or ( n28874 , n28869 , n28873 );
buf ( n28875 , n28874 );
not ( n28876 , n28875 );
buf ( n28877 , n28876 );
buf ( n28878 , n28877 );
not ( n28879 , n28878 );
or ( n28880 , n28866 , n28879 );
buf ( n28881 , n28880 );
buf ( n28882 , n28881 );
and ( n28883 , n28882 , n28614 );
not ( n28884 , n28883 );
and ( n28885 , n28884 , n28613 );
xor ( n28886 , n28613 , n28614 );
xor ( n28887 , n28886 , n28614 );
and ( n28888 , n28887 , n28883 );
or ( n28889 , n28885 , n28888 );
buf ( n28890 , n28889 );
and ( n28891 , n28890 , n28508 );
or ( n28892 , n28607 , n28891 );
buf ( n28893 , n28892 );
xor ( n28894 , n28596 , n28893 );
buf ( n28895 , n28894 );
buf ( n28896 , n28895 );
buf ( n28897 , n28896 );
not ( n28898 , n28897 );
buf ( n28899 , n28898 );
buf ( n28900 , n28899 );
not ( n28901 , n28900 );
buf ( n28902 , n25876 );
not ( n28903 , n14641 );
buf ( n28904 , n14645 );
buf ( n28905 , n14643 );
xor ( n28906 , n28904 , n28905 );
buf ( n28907 , n14651 );
buf ( n28908 , n14944 );
and ( n28909 , n28907 , n28908 );
buf ( n28910 , n14657 );
buf ( n28911 , n14969 );
and ( n28912 , n28910 , n28911 );
buf ( n28913 , n14663 );
buf ( n28914 , n14984 );
and ( n28915 , n28913 , n28914 );
buf ( n28916 , n14669 );
buf ( n28917 , n14999 );
and ( n28918 , n28916 , n28917 );
buf ( n28919 , n14675 );
buf ( n28920 , n15014 );
and ( n28921 , n28919 , n28920 );
buf ( n28922 , n14681 );
buf ( n28923 , n15029 );
and ( n28924 , n28922 , n28923 );
buf ( n28925 , n14687 );
buf ( n28926 , n15044 );
and ( n28927 , n28925 , n28926 );
buf ( n28928 , n14693 );
buf ( n28929 , n15059 );
and ( n28930 , n28928 , n28929 );
buf ( n28931 , n14699 );
buf ( n28932 , n15074 );
and ( n28933 , n28931 , n28932 );
buf ( n28934 , n14705 );
buf ( n28935 , n15089 );
and ( n28936 , n28934 , n28935 );
buf ( n28937 , n14711 );
buf ( n28938 , n15104 );
and ( n28939 , n28937 , n28938 );
buf ( n28940 , n14717 );
buf ( n28941 , n15119 );
and ( n28942 , n28940 , n28941 );
buf ( n28943 , n14723 );
buf ( n28944 , n15456 );
and ( n28945 , n28943 , n28944 );
buf ( n28946 , n14729 );
buf ( n28947 , n15478 );
and ( n28948 , n28946 , n28947 );
buf ( n28949 , n14735 );
buf ( n28950 , n15500 );
and ( n28951 , n28949 , n28950 );
buf ( n28952 , n14741 );
buf ( n28953 , n15522 );
and ( n28954 , n28952 , n28953 );
buf ( n28955 , n14747 );
buf ( n28956 , n15544 );
and ( n28957 , n28955 , n28956 );
buf ( n28958 , n14753 );
buf ( n28959 , n15566 );
and ( n28960 , n28958 , n28959 );
buf ( n28961 , n14759 );
buf ( n28962 , n15588 );
and ( n28963 , n28961 , n28962 );
buf ( n28964 , n14765 );
buf ( n28965 , n15610 );
and ( n28966 , n28964 , n28965 );
buf ( n28967 , n14771 );
buf ( n28968 , n15632 );
and ( n28969 , n28967 , n28968 );
buf ( n28970 , n14777 );
buf ( n28971 , n15654 );
and ( n28972 , n28970 , n28971 );
buf ( n28973 , n14783 );
buf ( n28974 , n15676 );
and ( n28975 , n28973 , n28974 );
buf ( n28976 , n14789 );
buf ( n28977 , n15698 );
and ( n28978 , n28976 , n28977 );
buf ( n28979 , n14795 );
buf ( n28980 , n15720 );
and ( n28981 , n28979 , n28980 );
buf ( n28982 , n14801 );
buf ( n28983 , n15742 );
and ( n28984 , n28982 , n28983 );
buf ( n28985 , n14807 );
buf ( n28986 , n15764 );
and ( n28987 , n28985 , n28986 );
buf ( n28988 , n14813 );
buf ( n28989 , n15786 );
and ( n28990 , n28988 , n28989 );
buf ( n28991 , n14819 );
buf ( n28992 , n15808 );
and ( n28993 , n28991 , n28992 );
buf ( n28994 , n14825 );
buf ( n28995 , n15830 );
and ( n28996 , n28994 , n28995 );
and ( n28997 , n28598 , n28599 );
and ( n28998 , n28995 , n28997 );
and ( n28999 , n28994 , n28997 );
or ( n29000 , n28996 , n28998 , n28999 );
and ( n29001 , n28992 , n29000 );
and ( n29002 , n28991 , n29000 );
or ( n29003 , n28993 , n29001 , n29002 );
and ( n29004 , n28989 , n29003 );
and ( n29005 , n28988 , n29003 );
or ( n29006 , n28990 , n29004 , n29005 );
and ( n29007 , n28986 , n29006 );
and ( n29008 , n28985 , n29006 );
or ( n29009 , n28987 , n29007 , n29008 );
and ( n29010 , n28983 , n29009 );
and ( n29011 , n28982 , n29009 );
or ( n29012 , n28984 , n29010 , n29011 );
and ( n29013 , n28980 , n29012 );
and ( n29014 , n28979 , n29012 );
or ( n29015 , n28981 , n29013 , n29014 );
and ( n29016 , n28977 , n29015 );
and ( n29017 , n28976 , n29015 );
or ( n29018 , n28978 , n29016 , n29017 );
and ( n29019 , n28974 , n29018 );
and ( n29020 , n28973 , n29018 );
or ( n29021 , n28975 , n29019 , n29020 );
and ( n29022 , n28971 , n29021 );
and ( n29023 , n28970 , n29021 );
or ( n29024 , n28972 , n29022 , n29023 );
and ( n29025 , n28968 , n29024 );
and ( n29026 , n28967 , n29024 );
or ( n29027 , n28969 , n29025 , n29026 );
and ( n29028 , n28965 , n29027 );
and ( n29029 , n28964 , n29027 );
or ( n29030 , n28966 , n29028 , n29029 );
and ( n29031 , n28962 , n29030 );
and ( n29032 , n28961 , n29030 );
or ( n29033 , n28963 , n29031 , n29032 );
and ( n29034 , n28959 , n29033 );
and ( n29035 , n28958 , n29033 );
or ( n29036 , n28960 , n29034 , n29035 );
and ( n29037 , n28956 , n29036 );
and ( n29038 , n28955 , n29036 );
or ( n29039 , n28957 , n29037 , n29038 );
and ( n29040 , n28953 , n29039 );
and ( n29041 , n28952 , n29039 );
or ( n29042 , n28954 , n29040 , n29041 );
and ( n29043 , n28950 , n29042 );
and ( n29044 , n28949 , n29042 );
or ( n29045 , n28951 , n29043 , n29044 );
and ( n29046 , n28947 , n29045 );
and ( n29047 , n28946 , n29045 );
or ( n29048 , n28948 , n29046 , n29047 );
and ( n29049 , n28944 , n29048 );
and ( n29050 , n28943 , n29048 );
or ( n29051 , n28945 , n29049 , n29050 );
and ( n29052 , n28941 , n29051 );
and ( n29053 , n28940 , n29051 );
or ( n29054 , n28942 , n29052 , n29053 );
and ( n29055 , n28938 , n29054 );
and ( n29056 , n28937 , n29054 );
or ( n29057 , n28939 , n29055 , n29056 );
and ( n29058 , n28935 , n29057 );
and ( n29059 , n28934 , n29057 );
or ( n29060 , n28936 , n29058 , n29059 );
and ( n29061 , n28932 , n29060 );
and ( n29062 , n28931 , n29060 );
or ( n29063 , n28933 , n29061 , n29062 );
and ( n29064 , n28929 , n29063 );
and ( n29065 , n28928 , n29063 );
or ( n29066 , n28930 , n29064 , n29065 );
and ( n29067 , n28926 , n29066 );
and ( n29068 , n28925 , n29066 );
or ( n29069 , n28927 , n29067 , n29068 );
and ( n29070 , n28923 , n29069 );
and ( n29071 , n28922 , n29069 );
or ( n29072 , n28924 , n29070 , n29071 );
and ( n29073 , n28920 , n29072 );
and ( n29074 , n28919 , n29072 );
or ( n29075 , n28921 , n29073 , n29074 );
and ( n29076 , n28917 , n29075 );
and ( n29077 , n28916 , n29075 );
or ( n29078 , n28918 , n29076 , n29077 );
and ( n29079 , n28914 , n29078 );
and ( n29080 , n28913 , n29078 );
or ( n29081 , n28915 , n29079 , n29080 );
and ( n29082 , n28911 , n29081 );
and ( n29083 , n28910 , n29081 );
or ( n29084 , n28912 , n29082 , n29083 );
and ( n29085 , n28908 , n29084 );
and ( n29086 , n28907 , n29084 );
or ( n29087 , n28909 , n29085 , n29086 );
xor ( n29088 , n28906 , n29087 );
buf ( n29089 , n29088 );
and ( n29090 , n28903 , n29089 );
and ( n29091 , n14645 , n14641 );
or ( n29092 , n29090 , n29091 );
and ( n29093 , n29092 , n28606 );
buf ( n29094 , n29093 );
buf ( n29095 , n29094 );
not ( n29096 , n29095 );
xor ( n29097 , n28902 , n29096 );
buf ( n29098 , n27181 );
not ( n29099 , n14641 );
xor ( n29100 , n28907 , n28908 );
xor ( n29101 , n29100 , n29084 );
buf ( n29102 , n29101 );
and ( n29103 , n29099 , n29102 );
and ( n29104 , n14651 , n14641 );
or ( n29105 , n29103 , n29104 );
and ( n29106 , n29105 , n28606 );
buf ( n29107 , n29106 );
buf ( n29108 , n29107 );
not ( n29109 , n29108 );
and ( n29110 , n29098 , n29109 );
buf ( n29111 , n27193 );
not ( n29112 , n14641 );
xor ( n29113 , n28910 , n28911 );
xor ( n29114 , n29113 , n29081 );
buf ( n29115 , n29114 );
and ( n29116 , n29112 , n29115 );
and ( n29117 , n14657 , n14641 );
or ( n29118 , n29116 , n29117 );
and ( n29119 , n29118 , n28606 );
buf ( n29120 , n29119 );
buf ( n29121 , n29120 );
not ( n29122 , n29121 );
and ( n29123 , n29111 , n29122 );
buf ( n29124 , n26807 );
not ( n29125 , n14641 );
xor ( n29126 , n28913 , n28914 );
xor ( n29127 , n29126 , n29078 );
buf ( n29128 , n29127 );
and ( n29129 , n29125 , n29128 );
and ( n29130 , n14663 , n14641 );
or ( n29131 , n29129 , n29130 );
and ( n29132 , n29131 , n28606 );
buf ( n29133 , n29132 );
buf ( n29134 , n29133 );
not ( n29135 , n29134 );
and ( n29136 , n29124 , n29135 );
buf ( n29137 , n26773 );
not ( n29138 , n14641 );
xor ( n29139 , n28916 , n28917 );
xor ( n29140 , n29139 , n29075 );
buf ( n29141 , n29140 );
and ( n29142 , n29138 , n29141 );
and ( n29143 , n14669 , n14641 );
or ( n29144 , n29142 , n29143 );
and ( n29145 , n29144 , n28606 );
buf ( n29146 , n29145 );
buf ( n29147 , n29146 );
not ( n29148 , n29147 );
and ( n29149 , n29137 , n29148 );
buf ( n29150 , n26739 );
not ( n29151 , n14641 );
xor ( n29152 , n28919 , n28920 );
xor ( n29153 , n29152 , n29072 );
buf ( n29154 , n29153 );
and ( n29155 , n29151 , n29154 );
and ( n29156 , n14675 , n14641 );
or ( n29157 , n29155 , n29156 );
and ( n29158 , n29157 , n28606 );
buf ( n29159 , n29158 );
buf ( n29160 , n29159 );
not ( n29161 , n29160 );
and ( n29162 , n29150 , n29161 );
buf ( n29163 , n26705 );
not ( n29164 , n14641 );
xor ( n29165 , n28922 , n28923 );
xor ( n29166 , n29165 , n29069 );
buf ( n29167 , n29166 );
and ( n29168 , n29164 , n29167 );
and ( n29169 , n14681 , n14641 );
or ( n29170 , n29168 , n29169 );
and ( n29171 , n29170 , n28606 );
buf ( n29172 , n29171 );
buf ( n29173 , n29172 );
not ( n29174 , n29173 );
and ( n29175 , n29163 , n29174 );
buf ( n29176 , n26671 );
not ( n29177 , n14641 );
xor ( n29178 , n28925 , n28926 );
xor ( n29179 , n29178 , n29066 );
buf ( n29180 , n29179 );
and ( n29181 , n29177 , n29180 );
and ( n29182 , n14687 , n14641 );
or ( n29183 , n29181 , n29182 );
and ( n29184 , n29183 , n28606 );
buf ( n29185 , n29184 );
buf ( n29186 , n29185 );
not ( n29187 , n29186 );
and ( n29188 , n29176 , n29187 );
buf ( n29189 , n26637 );
not ( n29190 , n14641 );
xor ( n29191 , n28928 , n28929 );
xor ( n29192 , n29191 , n29063 );
buf ( n29193 , n29192 );
and ( n29194 , n29190 , n29193 );
and ( n29195 , n14693 , n14641 );
or ( n29196 , n29194 , n29195 );
and ( n29197 , n29196 , n28606 );
buf ( n29198 , n29197 );
buf ( n29199 , n29198 );
not ( n29200 , n29199 );
and ( n29201 , n29189 , n29200 );
buf ( n29202 , n26603 );
not ( n29203 , n14641 );
xor ( n29204 , n28931 , n28932 );
xor ( n29205 , n29204 , n29060 );
buf ( n29206 , n29205 );
and ( n29207 , n29203 , n29206 );
and ( n29208 , n14699 , n14641 );
or ( n29209 , n29207 , n29208 );
and ( n29210 , n29209 , n28606 );
buf ( n29211 , n29210 );
buf ( n29212 , n29211 );
not ( n29213 , n29212 );
and ( n29214 , n29202 , n29213 );
buf ( n29215 , n26569 );
not ( n29216 , n14641 );
xor ( n29217 , n28934 , n28935 );
xor ( n29218 , n29217 , n29057 );
buf ( n29219 , n29218 );
and ( n29220 , n29216 , n29219 );
and ( n29221 , n14705 , n14641 );
or ( n29222 , n29220 , n29221 );
and ( n29223 , n29222 , n28606 );
buf ( n29224 , n29223 );
buf ( n29225 , n29224 );
not ( n29226 , n29225 );
and ( n29227 , n29215 , n29226 );
buf ( n29228 , n26535 );
not ( n29229 , n14641 );
xor ( n29230 , n28937 , n28938 );
xor ( n29231 , n29230 , n29054 );
buf ( n29232 , n29231 );
and ( n29233 , n29229 , n29232 );
and ( n29234 , n14711 , n14641 );
or ( n29235 , n29233 , n29234 );
and ( n29236 , n29235 , n28606 );
buf ( n29237 , n29236 );
buf ( n29238 , n29237 );
not ( n29239 , n29238 );
and ( n29240 , n29228 , n29239 );
buf ( n29241 , n26501 );
not ( n29242 , n14641 );
xor ( n29243 , n28940 , n28941 );
xor ( n29244 , n29243 , n29051 );
buf ( n29245 , n29244 );
and ( n29246 , n29242 , n29245 );
and ( n29247 , n14717 , n14641 );
or ( n29248 , n29246 , n29247 );
and ( n29249 , n29248 , n28606 );
not ( n29250 , n28883 );
and ( n29251 , n29250 , n28879 );
xor ( n29252 , n28879 , n28614 );
xor ( n29253 , n28865 , n28614 );
xor ( n29254 , n28851 , n28614 );
xor ( n29255 , n28837 , n28614 );
xor ( n29256 , n28823 , n28614 );
xor ( n29257 , n28809 , n28614 );
xor ( n29258 , n28795 , n28614 );
xor ( n29259 , n28781 , n28614 );
xor ( n29260 , n28767 , n28614 );
xor ( n29261 , n28753 , n28614 );
xor ( n29262 , n28739 , n28614 );
xor ( n29263 , n28725 , n28614 );
xor ( n29264 , n28711 , n28614 );
xor ( n29265 , n28697 , n28614 );
xor ( n29266 , n28683 , n28614 );
xor ( n29267 , n28669 , n28614 );
xor ( n29268 , n28655 , n28614 );
xor ( n29269 , n28641 , n28614 );
xor ( n29270 , n28627 , n28614 );
and ( n29271 , n28886 , n28614 );
and ( n29272 , n29270 , n29271 );
and ( n29273 , n29269 , n29272 );
and ( n29274 , n29268 , n29273 );
and ( n29275 , n29267 , n29274 );
and ( n29276 , n29266 , n29275 );
and ( n29277 , n29265 , n29276 );
and ( n29278 , n29264 , n29277 );
and ( n29279 , n29263 , n29278 );
and ( n29280 , n29262 , n29279 );
and ( n29281 , n29261 , n29280 );
and ( n29282 , n29260 , n29281 );
and ( n29283 , n29259 , n29282 );
and ( n29284 , n29258 , n29283 );
and ( n29285 , n29257 , n29284 );
and ( n29286 , n29256 , n29285 );
and ( n29287 , n29255 , n29286 );
and ( n29288 , n29254 , n29287 );
and ( n29289 , n29253 , n29288 );
xor ( n29290 , n29252 , n29289 );
and ( n29291 , n29290 , n28883 );
or ( n29292 , n29251 , n29291 );
buf ( n29293 , n29292 );
and ( n29294 , n29293 , n28508 );
or ( n29295 , n29249 , n29294 );
buf ( n29296 , n29295 );
not ( n29297 , n29296 );
and ( n29298 , n29241 , n29297 );
buf ( n29299 , n26467 );
not ( n29300 , n14641 );
xor ( n29301 , n28943 , n28944 );
xor ( n29302 , n29301 , n29048 );
buf ( n29303 , n29302 );
and ( n29304 , n29300 , n29303 );
and ( n29305 , n14723 , n14641 );
or ( n29306 , n29304 , n29305 );
and ( n29307 , n29306 , n28606 );
not ( n29308 , n28883 );
and ( n29309 , n29308 , n28865 );
xor ( n29310 , n29253 , n29288 );
and ( n29311 , n29310 , n28883 );
or ( n29312 , n29309 , n29311 );
buf ( n29313 , n29312 );
and ( n29314 , n29313 , n28508 );
or ( n29315 , n29307 , n29314 );
buf ( n29316 , n29315 );
not ( n29317 , n29316 );
and ( n29318 , n29299 , n29317 );
buf ( n29319 , n26433 );
not ( n29320 , n14641 );
xor ( n29321 , n28946 , n28947 );
xor ( n29322 , n29321 , n29045 );
buf ( n29323 , n29322 );
and ( n29324 , n29320 , n29323 );
and ( n29325 , n14729 , n14641 );
or ( n29326 , n29324 , n29325 );
and ( n29327 , n29326 , n28606 );
not ( n29328 , n28883 );
and ( n29329 , n29328 , n28851 );
xor ( n29330 , n29254 , n29287 );
and ( n29331 , n29330 , n28883 );
or ( n29332 , n29329 , n29331 );
buf ( n29333 , n29332 );
and ( n29334 , n29333 , n28508 );
or ( n29335 , n29327 , n29334 );
buf ( n29336 , n29335 );
not ( n29337 , n29336 );
and ( n29338 , n29319 , n29337 );
buf ( n29339 , n26399 );
not ( n29340 , n14641 );
xor ( n29341 , n28949 , n28950 );
xor ( n29342 , n29341 , n29042 );
buf ( n29343 , n29342 );
and ( n29344 , n29340 , n29343 );
and ( n29345 , n14735 , n14641 );
or ( n29346 , n29344 , n29345 );
and ( n29347 , n29346 , n28606 );
not ( n29348 , n28883 );
and ( n29349 , n29348 , n28837 );
xor ( n29350 , n29255 , n29286 );
and ( n29351 , n29350 , n28883 );
or ( n29352 , n29349 , n29351 );
buf ( n29353 , n29352 );
and ( n29354 , n29353 , n28508 );
or ( n29355 , n29347 , n29354 );
buf ( n29356 , n29355 );
not ( n29357 , n29356 );
and ( n29358 , n29339 , n29357 );
buf ( n29359 , n26365 );
not ( n29360 , n14641 );
xor ( n29361 , n28952 , n28953 );
xor ( n29362 , n29361 , n29039 );
buf ( n29363 , n29362 );
and ( n29364 , n29360 , n29363 );
and ( n29365 , n14741 , n14641 );
or ( n29366 , n29364 , n29365 );
and ( n29367 , n29366 , n28606 );
not ( n29368 , n28883 );
and ( n29369 , n29368 , n28823 );
xor ( n29370 , n29256 , n29285 );
and ( n29371 , n29370 , n28883 );
or ( n29372 , n29369 , n29371 );
buf ( n29373 , n29372 );
and ( n29374 , n29373 , n28508 );
or ( n29375 , n29367 , n29374 );
buf ( n29376 , n29375 );
not ( n29377 , n29376 );
and ( n29378 , n29359 , n29377 );
buf ( n29379 , n26331 );
not ( n29380 , n14641 );
xor ( n29381 , n28955 , n28956 );
xor ( n29382 , n29381 , n29036 );
buf ( n29383 , n29382 );
and ( n29384 , n29380 , n29383 );
and ( n29385 , n14747 , n14641 );
or ( n29386 , n29384 , n29385 );
and ( n29387 , n29386 , n28606 );
not ( n29388 , n28883 );
and ( n29389 , n29388 , n28809 );
xor ( n29390 , n29257 , n29284 );
and ( n29391 , n29390 , n28883 );
or ( n29392 , n29389 , n29391 );
buf ( n29393 , n29392 );
and ( n29394 , n29393 , n28508 );
or ( n29395 , n29387 , n29394 );
buf ( n29396 , n29395 );
not ( n29397 , n29396 );
and ( n29398 , n29379 , n29397 );
buf ( n29399 , n26297 );
not ( n29400 , n14641 );
xor ( n29401 , n28958 , n28959 );
xor ( n29402 , n29401 , n29033 );
buf ( n29403 , n29402 );
and ( n29404 , n29400 , n29403 );
and ( n29405 , n14753 , n14641 );
or ( n29406 , n29404 , n29405 );
and ( n29407 , n29406 , n28606 );
not ( n29408 , n28883 );
and ( n29409 , n29408 , n28795 );
xor ( n29410 , n29258 , n29283 );
and ( n29411 , n29410 , n28883 );
or ( n29412 , n29409 , n29411 );
buf ( n29413 , n29412 );
and ( n29414 , n29413 , n28508 );
or ( n29415 , n29407 , n29414 );
buf ( n29416 , n29415 );
not ( n29417 , n29416 );
and ( n29418 , n29399 , n29417 );
buf ( n29419 , n26263 );
not ( n29420 , n14641 );
xor ( n29421 , n28961 , n28962 );
xor ( n29422 , n29421 , n29030 );
buf ( n29423 , n29422 );
and ( n29424 , n29420 , n29423 );
and ( n29425 , n14759 , n14641 );
or ( n29426 , n29424 , n29425 );
and ( n29427 , n29426 , n28606 );
not ( n29428 , n28883 );
and ( n29429 , n29428 , n28781 );
xor ( n29430 , n29259 , n29282 );
and ( n29431 , n29430 , n28883 );
or ( n29432 , n29429 , n29431 );
buf ( n29433 , n29432 );
and ( n29434 , n29433 , n28508 );
or ( n29435 , n29427 , n29434 );
buf ( n29436 , n29435 );
not ( n29437 , n29436 );
and ( n29438 , n29419 , n29437 );
buf ( n29439 , n26229 );
not ( n29440 , n14641 );
xor ( n29441 , n28964 , n28965 );
xor ( n29442 , n29441 , n29027 );
buf ( n29443 , n29442 );
and ( n29444 , n29440 , n29443 );
and ( n29445 , n14765 , n14641 );
or ( n29446 , n29444 , n29445 );
and ( n29447 , n29446 , n28606 );
not ( n29448 , n28883 );
and ( n29449 , n29448 , n28767 );
xor ( n29450 , n29260 , n29281 );
and ( n29451 , n29450 , n28883 );
or ( n29452 , n29449 , n29451 );
buf ( n29453 , n29452 );
and ( n29454 , n29453 , n28508 );
or ( n29455 , n29447 , n29454 );
buf ( n29456 , n29455 );
not ( n29457 , n29456 );
and ( n29458 , n29439 , n29457 );
buf ( n29459 , n26195 );
not ( n29460 , n14641 );
xor ( n29461 , n28967 , n28968 );
xor ( n29462 , n29461 , n29024 );
buf ( n29463 , n29462 );
and ( n29464 , n29460 , n29463 );
and ( n29465 , n14771 , n14641 );
or ( n29466 , n29464 , n29465 );
and ( n29467 , n29466 , n28606 );
not ( n29468 , n28883 );
and ( n29469 , n29468 , n28753 );
xor ( n29470 , n29261 , n29280 );
and ( n29471 , n29470 , n28883 );
or ( n29472 , n29469 , n29471 );
buf ( n29473 , n29472 );
and ( n29474 , n29473 , n28508 );
or ( n29475 , n29467 , n29474 );
buf ( n29476 , n29475 );
not ( n29477 , n29476 );
and ( n29478 , n29459 , n29477 );
buf ( n29479 , n26161 );
not ( n29480 , n14641 );
xor ( n29481 , n28970 , n28971 );
xor ( n29482 , n29481 , n29021 );
buf ( n29483 , n29482 );
and ( n29484 , n29480 , n29483 );
and ( n29485 , n14777 , n14641 );
or ( n29486 , n29484 , n29485 );
and ( n29487 , n29486 , n28606 );
not ( n29488 , n28883 );
and ( n29489 , n29488 , n28739 );
xor ( n29490 , n29262 , n29279 );
and ( n29491 , n29490 , n28883 );
or ( n29492 , n29489 , n29491 );
buf ( n29493 , n29492 );
and ( n29494 , n29493 , n28508 );
or ( n29495 , n29487 , n29494 );
buf ( n29496 , n29495 );
not ( n29497 , n29496 );
and ( n29498 , n29479 , n29497 );
buf ( n29499 , n26127 );
not ( n29500 , n14641 );
xor ( n29501 , n28973 , n28974 );
xor ( n29502 , n29501 , n29018 );
buf ( n29503 , n29502 );
and ( n29504 , n29500 , n29503 );
and ( n29505 , n14783 , n14641 );
or ( n29506 , n29504 , n29505 );
and ( n29507 , n29506 , n28606 );
not ( n29508 , n28883 );
and ( n29509 , n29508 , n28725 );
xor ( n29510 , n29263 , n29278 );
and ( n29511 , n29510 , n28883 );
or ( n29512 , n29509 , n29511 );
buf ( n29513 , n29512 );
and ( n29514 , n29513 , n28508 );
or ( n29515 , n29507 , n29514 );
buf ( n29516 , n29515 );
not ( n29517 , n29516 );
and ( n29518 , n29499 , n29517 );
buf ( n29519 , n26093 );
not ( n29520 , n14641 );
xor ( n29521 , n28976 , n28977 );
xor ( n29522 , n29521 , n29015 );
buf ( n29523 , n29522 );
and ( n29524 , n29520 , n29523 );
and ( n29525 , n14789 , n14641 );
or ( n29526 , n29524 , n29525 );
and ( n29527 , n29526 , n28606 );
not ( n29528 , n28883 );
and ( n29529 , n29528 , n28711 );
xor ( n29530 , n29264 , n29277 );
and ( n29531 , n29530 , n28883 );
or ( n29532 , n29529 , n29531 );
buf ( n29533 , n29532 );
and ( n29534 , n29533 , n28508 );
or ( n29535 , n29527 , n29534 );
buf ( n29536 , n29535 );
not ( n29537 , n29536 );
and ( n29538 , n29519 , n29537 );
buf ( n29539 , n26059 );
not ( n29540 , n14641 );
xor ( n29541 , n28979 , n28980 );
xor ( n29542 , n29541 , n29012 );
buf ( n29543 , n29542 );
and ( n29544 , n29540 , n29543 );
and ( n29545 , n14795 , n14641 );
or ( n29546 , n29544 , n29545 );
and ( n29547 , n29546 , n28606 );
not ( n29548 , n28883 );
and ( n29549 , n29548 , n28697 );
xor ( n29550 , n29265 , n29276 );
and ( n29551 , n29550 , n28883 );
or ( n29552 , n29549 , n29551 );
buf ( n29553 , n29552 );
and ( n29554 , n29553 , n28508 );
or ( n29555 , n29547 , n29554 );
buf ( n29556 , n29555 );
not ( n29557 , n29556 );
and ( n29558 , n29539 , n29557 );
buf ( n29559 , n26025 );
not ( n29560 , n14641 );
xor ( n29561 , n28982 , n28983 );
xor ( n29562 , n29561 , n29009 );
buf ( n29563 , n29562 );
and ( n29564 , n29560 , n29563 );
and ( n29565 , n14801 , n14641 );
or ( n29566 , n29564 , n29565 );
and ( n29567 , n29566 , n28606 );
not ( n29568 , n28883 );
and ( n29569 , n29568 , n28683 );
xor ( n29570 , n29266 , n29275 );
and ( n29571 , n29570 , n28883 );
or ( n29572 , n29569 , n29571 );
buf ( n29573 , n29572 );
and ( n29574 , n29573 , n28508 );
or ( n29575 , n29567 , n29574 );
buf ( n29576 , n29575 );
not ( n29577 , n29576 );
and ( n29578 , n29559 , n29577 );
buf ( n29579 , n25991 );
not ( n29580 , n14641 );
xor ( n29581 , n28985 , n28986 );
xor ( n29582 , n29581 , n29006 );
buf ( n29583 , n29582 );
and ( n29584 , n29580 , n29583 );
and ( n29585 , n14807 , n14641 );
or ( n29586 , n29584 , n29585 );
and ( n29587 , n29586 , n28606 );
not ( n29588 , n28883 );
and ( n29589 , n29588 , n28669 );
xor ( n29590 , n29267 , n29274 );
and ( n29591 , n29590 , n28883 );
or ( n29592 , n29589 , n29591 );
buf ( n29593 , n29592 );
and ( n29594 , n29593 , n28508 );
or ( n29595 , n29587 , n29594 );
buf ( n29596 , n29595 );
not ( n29597 , n29596 );
and ( n29598 , n29579 , n29597 );
buf ( n29599 , n25958 );
not ( n29600 , n14641 );
xor ( n29601 , n28988 , n28989 );
xor ( n29602 , n29601 , n29003 );
buf ( n29603 , n29602 );
and ( n29604 , n29600 , n29603 );
and ( n29605 , n14813 , n14641 );
or ( n29606 , n29604 , n29605 );
and ( n29607 , n29606 , n28606 );
not ( n29608 , n28883 );
and ( n29609 , n29608 , n28655 );
xor ( n29610 , n29268 , n29273 );
and ( n29611 , n29610 , n28883 );
or ( n29612 , n29609 , n29611 );
buf ( n29613 , n29612 );
and ( n29614 , n29613 , n28508 );
or ( n29615 , n29607 , n29614 );
buf ( n29616 , n29615 );
not ( n29617 , n29616 );
and ( n29618 , n29599 , n29617 );
buf ( n29619 , n25925 );
not ( n29620 , n14641 );
xor ( n29621 , n28991 , n28992 );
xor ( n29622 , n29621 , n29000 );
buf ( n29623 , n29622 );
and ( n29624 , n29620 , n29623 );
and ( n29625 , n14819 , n14641 );
or ( n29626 , n29624 , n29625 );
and ( n29627 , n29626 , n28606 );
not ( n29628 , n28883 );
and ( n29629 , n29628 , n28641 );
xor ( n29630 , n29269 , n29272 );
and ( n29631 , n29630 , n28883 );
or ( n29632 , n29629 , n29631 );
buf ( n29633 , n29632 );
and ( n29634 , n29633 , n28508 );
or ( n29635 , n29627 , n29634 );
buf ( n29636 , n29635 );
not ( n29637 , n29636 );
and ( n29638 , n29619 , n29637 );
buf ( n29639 , n25894 );
not ( n29640 , n14641 );
xor ( n29641 , n28994 , n28995 );
xor ( n29642 , n29641 , n28997 );
buf ( n29643 , n29642 );
and ( n29644 , n29640 , n29643 );
and ( n29645 , n14825 , n14641 );
or ( n29646 , n29644 , n29645 );
and ( n29647 , n29646 , n28606 );
not ( n29648 , n28883 );
and ( n29649 , n29648 , n28627 );
xor ( n29650 , n29270 , n29271 );
and ( n29651 , n29650 , n28883 );
or ( n29652 , n29649 , n29651 );
buf ( n29653 , n29652 );
and ( n29654 , n29653 , n28508 );
or ( n29655 , n29647 , n29654 );
buf ( n29656 , n29655 );
not ( n29657 , n29656 );
and ( n29658 , n29639 , n29657 );
not ( n29659 , n28893 );
or ( n29660 , n28596 , n29659 );
and ( n29661 , n29657 , n29660 );
and ( n29662 , n29639 , n29660 );
or ( n29663 , n29658 , n29661 , n29662 );
and ( n29664 , n29637 , n29663 );
and ( n29665 , n29619 , n29663 );
or ( n29666 , n29638 , n29664 , n29665 );
and ( n29667 , n29617 , n29666 );
and ( n29668 , n29599 , n29666 );
or ( n29669 , n29618 , n29667 , n29668 );
and ( n29670 , n29597 , n29669 );
and ( n29671 , n29579 , n29669 );
or ( n29672 , n29598 , n29670 , n29671 );
and ( n29673 , n29577 , n29672 );
and ( n29674 , n29559 , n29672 );
or ( n29675 , n29578 , n29673 , n29674 );
and ( n29676 , n29557 , n29675 );
and ( n29677 , n29539 , n29675 );
or ( n29678 , n29558 , n29676 , n29677 );
and ( n29679 , n29537 , n29678 );
and ( n29680 , n29519 , n29678 );
or ( n29681 , n29538 , n29679 , n29680 );
and ( n29682 , n29517 , n29681 );
and ( n29683 , n29499 , n29681 );
or ( n29684 , n29518 , n29682 , n29683 );
and ( n29685 , n29497 , n29684 );
and ( n29686 , n29479 , n29684 );
or ( n29687 , n29498 , n29685 , n29686 );
and ( n29688 , n29477 , n29687 );
and ( n29689 , n29459 , n29687 );
or ( n29690 , n29478 , n29688 , n29689 );
and ( n29691 , n29457 , n29690 );
and ( n29692 , n29439 , n29690 );
or ( n29693 , n29458 , n29691 , n29692 );
and ( n29694 , n29437 , n29693 );
and ( n29695 , n29419 , n29693 );
or ( n29696 , n29438 , n29694 , n29695 );
and ( n29697 , n29417 , n29696 );
and ( n29698 , n29399 , n29696 );
or ( n29699 , n29418 , n29697 , n29698 );
and ( n29700 , n29397 , n29699 );
and ( n29701 , n29379 , n29699 );
or ( n29702 , n29398 , n29700 , n29701 );
and ( n29703 , n29377 , n29702 );
and ( n29704 , n29359 , n29702 );
or ( n29705 , n29378 , n29703 , n29704 );
and ( n29706 , n29357 , n29705 );
and ( n29707 , n29339 , n29705 );
or ( n29708 , n29358 , n29706 , n29707 );
and ( n29709 , n29337 , n29708 );
and ( n29710 , n29319 , n29708 );
or ( n29711 , n29338 , n29709 , n29710 );
and ( n29712 , n29317 , n29711 );
and ( n29713 , n29299 , n29711 );
or ( n29714 , n29318 , n29712 , n29713 );
and ( n29715 , n29297 , n29714 );
and ( n29716 , n29241 , n29714 );
or ( n29717 , n29298 , n29715 , n29716 );
and ( n29718 , n29239 , n29717 );
and ( n29719 , n29228 , n29717 );
or ( n29720 , n29240 , n29718 , n29719 );
and ( n29721 , n29226 , n29720 );
and ( n29722 , n29215 , n29720 );
or ( n29723 , n29227 , n29721 , n29722 );
and ( n29724 , n29213 , n29723 );
and ( n29725 , n29202 , n29723 );
or ( n29726 , n29214 , n29724 , n29725 );
and ( n29727 , n29200 , n29726 );
and ( n29728 , n29189 , n29726 );
or ( n29729 , n29201 , n29727 , n29728 );
and ( n29730 , n29187 , n29729 );
and ( n29731 , n29176 , n29729 );
or ( n29732 , n29188 , n29730 , n29731 );
and ( n29733 , n29174 , n29732 );
and ( n29734 , n29163 , n29732 );
or ( n29735 , n29175 , n29733 , n29734 );
and ( n29736 , n29161 , n29735 );
and ( n29737 , n29150 , n29735 );
or ( n29738 , n29162 , n29736 , n29737 );
and ( n29739 , n29148 , n29738 );
and ( n29740 , n29137 , n29738 );
or ( n29741 , n29149 , n29739 , n29740 );
and ( n29742 , n29135 , n29741 );
and ( n29743 , n29124 , n29741 );
or ( n29744 , n29136 , n29742 , n29743 );
and ( n29745 , n29122 , n29744 );
and ( n29746 , n29111 , n29744 );
or ( n29747 , n29123 , n29745 , n29746 );
and ( n29748 , n29109 , n29747 );
and ( n29749 , n29098 , n29747 );
or ( n29750 , n29110 , n29748 , n29749 );
xor ( n29751 , n29097 , n29750 );
buf ( n29752 , n29751 );
buf ( n29753 , n29752 );
not ( n29754 , n29753 );
xor ( n29755 , n29639 , n29657 );
xor ( n29756 , n29755 , n29660 );
buf ( n29757 , n29756 );
buf ( n29758 , n29757 );
and ( n29759 , n29754 , n29758 );
not ( n29760 , n29758 );
not ( n29761 , n28896 );
xor ( n29762 , n29760 , n29761 );
and ( n29763 , n29762 , n29753 );
or ( n29764 , n29759 , n29763 );
buf ( n29765 , n29764 );
not ( n29766 , n29765 );
buf ( n29767 , n29766 );
buf ( n29768 , n29767 );
not ( n29769 , n29768 );
or ( n29770 , n28901 , n29769 );
not ( n29771 , n29753 );
xor ( n29772 , n29619 , n29637 );
xor ( n29773 , n29772 , n29663 );
buf ( n29774 , n29773 );
buf ( n29775 , n29774 );
and ( n29776 , n29771 , n29775 );
not ( n29777 , n29775 );
and ( n29778 , n29760 , n29761 );
xor ( n29779 , n29777 , n29778 );
and ( n29780 , n29779 , n29753 );
or ( n29781 , n29776 , n29780 );
buf ( n29782 , n29781 );
not ( n29783 , n29782 );
buf ( n29784 , n29783 );
buf ( n29785 , n29784 );
not ( n29786 , n29785 );
or ( n29787 , n29770 , n29786 );
not ( n29788 , n29753 );
xor ( n29789 , n29599 , n29617 );
xor ( n29790 , n29789 , n29666 );
buf ( n29791 , n29790 );
buf ( n29792 , n29791 );
and ( n29793 , n29788 , n29792 );
not ( n29794 , n29792 );
and ( n29795 , n29777 , n29778 );
xor ( n29796 , n29794 , n29795 );
and ( n29797 , n29796 , n29753 );
or ( n29798 , n29793 , n29797 );
buf ( n29799 , n29798 );
not ( n29800 , n29799 );
buf ( n29801 , n29800 );
buf ( n29802 , n29801 );
not ( n29803 , n29802 );
or ( n29804 , n29787 , n29803 );
not ( n29805 , n29753 );
xor ( n29806 , n29579 , n29597 );
xor ( n29807 , n29806 , n29669 );
buf ( n29808 , n29807 );
buf ( n29809 , n29808 );
and ( n29810 , n29805 , n29809 );
not ( n29811 , n29809 );
and ( n29812 , n29794 , n29795 );
xor ( n29813 , n29811 , n29812 );
and ( n29814 , n29813 , n29753 );
or ( n29815 , n29810 , n29814 );
buf ( n29816 , n29815 );
not ( n29817 , n29816 );
buf ( n29818 , n29817 );
buf ( n29819 , n29818 );
not ( n29820 , n29819 );
or ( n29821 , n29804 , n29820 );
not ( n29822 , n29753 );
xor ( n29823 , n29559 , n29577 );
xor ( n29824 , n29823 , n29672 );
buf ( n29825 , n29824 );
buf ( n29826 , n29825 );
and ( n29827 , n29822 , n29826 );
not ( n29828 , n29826 );
and ( n29829 , n29811 , n29812 );
xor ( n29830 , n29828 , n29829 );
and ( n29831 , n29830 , n29753 );
or ( n29832 , n29827 , n29831 );
buf ( n29833 , n29832 );
not ( n29834 , n29833 );
buf ( n29835 , n29834 );
buf ( n29836 , n29835 );
not ( n29837 , n29836 );
or ( n29838 , n29821 , n29837 );
not ( n29839 , n29753 );
xor ( n29840 , n29539 , n29557 );
xor ( n29841 , n29840 , n29675 );
buf ( n29842 , n29841 );
buf ( n29843 , n29842 );
and ( n29844 , n29839 , n29843 );
not ( n29845 , n29843 );
and ( n29846 , n29828 , n29829 );
xor ( n29847 , n29845 , n29846 );
and ( n29848 , n29847 , n29753 );
or ( n29849 , n29844 , n29848 );
buf ( n29850 , n29849 );
not ( n29851 , n29850 );
buf ( n29852 , n29851 );
buf ( n29853 , n29852 );
not ( n29854 , n29853 );
or ( n29855 , n29838 , n29854 );
not ( n29856 , n29753 );
xor ( n29857 , n29519 , n29537 );
xor ( n29858 , n29857 , n29678 );
buf ( n29859 , n29858 );
buf ( n29860 , n29859 );
and ( n29861 , n29856 , n29860 );
not ( n29862 , n29860 );
and ( n29863 , n29845 , n29846 );
xor ( n29864 , n29862 , n29863 );
and ( n29865 , n29864 , n29753 );
or ( n29866 , n29861 , n29865 );
buf ( n29867 , n29866 );
not ( n29868 , n29867 );
buf ( n29869 , n29868 );
buf ( n29870 , n29869 );
not ( n29871 , n29870 );
or ( n29872 , n29855 , n29871 );
not ( n29873 , n29753 );
xor ( n29874 , n29499 , n29517 );
xor ( n29875 , n29874 , n29681 );
buf ( n29876 , n29875 );
buf ( n29877 , n29876 );
and ( n29878 , n29873 , n29877 );
not ( n29879 , n29877 );
and ( n29880 , n29862 , n29863 );
xor ( n29881 , n29879 , n29880 );
and ( n29882 , n29881 , n29753 );
or ( n29883 , n29878 , n29882 );
buf ( n29884 , n29883 );
not ( n29885 , n29884 );
buf ( n29886 , n29885 );
buf ( n29887 , n29886 );
not ( n29888 , n29887 );
or ( n29889 , n29872 , n29888 );
not ( n29890 , n29753 );
xor ( n29891 , n29479 , n29497 );
xor ( n29892 , n29891 , n29684 );
buf ( n29893 , n29892 );
buf ( n29894 , n29893 );
and ( n29895 , n29890 , n29894 );
not ( n29896 , n29894 );
and ( n29897 , n29879 , n29880 );
xor ( n29898 , n29896 , n29897 );
and ( n29899 , n29898 , n29753 );
or ( n29900 , n29895 , n29899 );
buf ( n29901 , n29900 );
not ( n29902 , n29901 );
buf ( n29903 , n29902 );
buf ( n29904 , n29903 );
not ( n29905 , n29904 );
or ( n29906 , n29889 , n29905 );
not ( n29907 , n29753 );
xor ( n29908 , n29459 , n29477 );
xor ( n29909 , n29908 , n29687 );
buf ( n29910 , n29909 );
buf ( n29911 , n29910 );
and ( n29912 , n29907 , n29911 );
not ( n29913 , n29911 );
and ( n29914 , n29896 , n29897 );
xor ( n29915 , n29913 , n29914 );
and ( n29916 , n29915 , n29753 );
or ( n29917 , n29912 , n29916 );
buf ( n29918 , n29917 );
not ( n29919 , n29918 );
buf ( n29920 , n29919 );
buf ( n29921 , n29920 );
not ( n29922 , n29921 );
or ( n29923 , n29906 , n29922 );
not ( n29924 , n29753 );
xor ( n29925 , n29439 , n29457 );
xor ( n29926 , n29925 , n29690 );
buf ( n29927 , n29926 );
buf ( n29928 , n29927 );
and ( n29929 , n29924 , n29928 );
not ( n29930 , n29928 );
and ( n29931 , n29913 , n29914 );
xor ( n29932 , n29930 , n29931 );
and ( n29933 , n29932 , n29753 );
or ( n29934 , n29929 , n29933 );
buf ( n29935 , n29934 );
not ( n29936 , n29935 );
buf ( n29937 , n29936 );
buf ( n29938 , n29937 );
not ( n29939 , n29938 );
or ( n29940 , n29923 , n29939 );
not ( n29941 , n29753 );
xor ( n29942 , n29419 , n29437 );
xor ( n29943 , n29942 , n29693 );
buf ( n29944 , n29943 );
buf ( n29945 , n29944 );
and ( n29946 , n29941 , n29945 );
not ( n29947 , n29945 );
and ( n29948 , n29930 , n29931 );
xor ( n29949 , n29947 , n29948 );
and ( n29950 , n29949 , n29753 );
or ( n29951 , n29946 , n29950 );
buf ( n29952 , n29951 );
not ( n29953 , n29952 );
buf ( n29954 , n29953 );
buf ( n29955 , n29954 );
not ( n29956 , n29955 );
or ( n29957 , n29940 , n29956 );
not ( n29958 , n29753 );
xor ( n29959 , n29399 , n29417 );
xor ( n29960 , n29959 , n29696 );
buf ( n29961 , n29960 );
buf ( n29962 , n29961 );
and ( n29963 , n29958 , n29962 );
not ( n29964 , n29962 );
and ( n29965 , n29947 , n29948 );
xor ( n29966 , n29964 , n29965 );
and ( n29967 , n29966 , n29753 );
or ( n29968 , n29963 , n29967 );
buf ( n29969 , n29968 );
not ( n29970 , n29969 );
buf ( n29971 , n29970 );
buf ( n29972 , n29971 );
not ( n29973 , n29972 );
or ( n29974 , n29957 , n29973 );
not ( n29975 , n29753 );
xor ( n29976 , n29379 , n29397 );
xor ( n29977 , n29976 , n29699 );
buf ( n29978 , n29977 );
buf ( n29979 , n29978 );
and ( n29980 , n29975 , n29979 );
not ( n29981 , n29979 );
and ( n29982 , n29964 , n29965 );
xor ( n29983 , n29981 , n29982 );
and ( n29984 , n29983 , n29753 );
or ( n29985 , n29980 , n29984 );
buf ( n29986 , n29985 );
not ( n29987 , n29986 );
buf ( n29988 , n29987 );
buf ( n29989 , n29988 );
not ( n29990 , n29989 );
or ( n29991 , n29974 , n29990 );
not ( n29992 , n29753 );
xor ( n29993 , n29359 , n29377 );
xor ( n29994 , n29993 , n29702 );
buf ( n29995 , n29994 );
buf ( n29996 , n29995 );
and ( n29997 , n29992 , n29996 );
not ( n29998 , n29996 );
and ( n29999 , n29981 , n29982 );
xor ( n30000 , n29998 , n29999 );
and ( n30001 , n30000 , n29753 );
or ( n30002 , n29997 , n30001 );
buf ( n30003 , n30002 );
not ( n30004 , n30003 );
buf ( n30005 , n30004 );
buf ( n30006 , n30005 );
not ( n30007 , n30006 );
or ( n30008 , n29991 , n30007 );
not ( n30009 , n29753 );
xor ( n30010 , n29339 , n29357 );
xor ( n30011 , n30010 , n29705 );
buf ( n30012 , n30011 );
buf ( n30013 , n30012 );
and ( n30014 , n30009 , n30013 );
not ( n30015 , n30013 );
and ( n30016 , n29998 , n29999 );
xor ( n30017 , n30015 , n30016 );
and ( n30018 , n30017 , n29753 );
or ( n30019 , n30014 , n30018 );
buf ( n30020 , n30019 );
not ( n30021 , n30020 );
buf ( n30022 , n30021 );
buf ( n30023 , n30022 );
not ( n30024 , n30023 );
or ( n30025 , n30008 , n30024 );
not ( n30026 , n29753 );
xor ( n30027 , n29319 , n29337 );
xor ( n30028 , n30027 , n29708 );
buf ( n30029 , n30028 );
buf ( n30030 , n30029 );
and ( n30031 , n30026 , n30030 );
not ( n30032 , n30030 );
and ( n30033 , n30015 , n30016 );
xor ( n30034 , n30032 , n30033 );
and ( n30035 , n30034 , n29753 );
or ( n30036 , n30031 , n30035 );
buf ( n30037 , n30036 );
not ( n30038 , n30037 );
buf ( n30039 , n30038 );
buf ( n30040 , n30039 );
not ( n30041 , n30040 );
or ( n30042 , n30025 , n30041 );
not ( n30043 , n29753 );
xor ( n30044 , n29299 , n29317 );
xor ( n30045 , n30044 , n29711 );
buf ( n30046 , n30045 );
buf ( n30047 , n30046 );
and ( n30048 , n30043 , n30047 );
not ( n30049 , n30047 );
and ( n30050 , n30032 , n30033 );
xor ( n30051 , n30049 , n30050 );
and ( n30052 , n30051 , n29753 );
or ( n30053 , n30048 , n30052 );
buf ( n30054 , n30053 );
not ( n30055 , n30054 );
buf ( n30056 , n30055 );
buf ( n30057 , n30056 );
not ( n30058 , n30057 );
or ( n30059 , n30042 , n30058 );
not ( n30060 , n29753 );
xor ( n30061 , n29241 , n29297 );
xor ( n30062 , n30061 , n29714 );
buf ( n30063 , n30062 );
buf ( n30064 , n30063 );
and ( n30065 , n30060 , n30064 );
not ( n30066 , n30064 );
and ( n30067 , n30049 , n30050 );
xor ( n30068 , n30066 , n30067 );
and ( n30069 , n30068 , n29753 );
or ( n30070 , n30065 , n30069 );
buf ( n30071 , n30070 );
not ( n30072 , n30071 );
buf ( n30073 , n30072 );
buf ( n30074 , n30073 );
not ( n30075 , n30074 );
or ( n30076 , n30059 , n30075 );
not ( n30077 , n29753 );
xor ( n30078 , n29228 , n29239 );
xor ( n30079 , n30078 , n29717 );
buf ( n30080 , n30079 );
buf ( n30081 , n30080 );
and ( n30082 , n30077 , n30081 );
not ( n30083 , n30081 );
and ( n30084 , n30066 , n30067 );
xor ( n30085 , n30083 , n30084 );
and ( n30086 , n30085 , n29753 );
or ( n30087 , n30082 , n30086 );
buf ( n30088 , n30087 );
not ( n30089 , n30088 );
buf ( n30090 , n30089 );
buf ( n30091 , n30090 );
not ( n30092 , n30091 );
or ( n30093 , n30076 , n30092 );
not ( n30094 , n29753 );
xor ( n30095 , n29215 , n29226 );
xor ( n30096 , n30095 , n29720 );
buf ( n30097 , n30096 );
buf ( n30098 , n30097 );
and ( n30099 , n30094 , n30098 );
not ( n30100 , n30098 );
and ( n30101 , n30083 , n30084 );
xor ( n30102 , n30100 , n30101 );
and ( n30103 , n30102 , n29753 );
or ( n30104 , n30099 , n30103 );
buf ( n30105 , n30104 );
not ( n30106 , n30105 );
buf ( n30107 , n30106 );
buf ( n30108 , n30107 );
not ( n30109 , n30108 );
or ( n30110 , n30093 , n30109 );
not ( n30111 , n29753 );
xor ( n30112 , n29202 , n29213 );
xor ( n30113 , n30112 , n29723 );
buf ( n30114 , n30113 );
buf ( n30115 , n30114 );
and ( n30116 , n30111 , n30115 );
not ( n30117 , n30115 );
and ( n30118 , n30100 , n30101 );
xor ( n30119 , n30117 , n30118 );
and ( n30120 , n30119 , n29753 );
or ( n30121 , n30116 , n30120 );
buf ( n30122 , n30121 );
not ( n30123 , n30122 );
buf ( n30124 , n30123 );
buf ( n30125 , n30124 );
not ( n30126 , n30125 );
or ( n30127 , n30110 , n30126 );
not ( n30128 , n29753 );
xor ( n30129 , n29189 , n29200 );
xor ( n30130 , n30129 , n29726 );
buf ( n30131 , n30130 );
buf ( n30132 , n30131 );
and ( n30133 , n30128 , n30132 );
not ( n30134 , n30132 );
and ( n30135 , n30117 , n30118 );
xor ( n30136 , n30134 , n30135 );
and ( n30137 , n30136 , n29753 );
or ( n30138 , n30133 , n30137 );
buf ( n30139 , n30138 );
not ( n30140 , n30139 );
buf ( n30141 , n30140 );
buf ( n30142 , n30141 );
not ( n30143 , n30142 );
or ( n30144 , n30127 , n30143 );
not ( n30145 , n29753 );
xor ( n30146 , n29176 , n29187 );
xor ( n30147 , n30146 , n29729 );
buf ( n30148 , n30147 );
buf ( n30149 , n30148 );
and ( n30150 , n30145 , n30149 );
not ( n30151 , n30149 );
and ( n30152 , n30134 , n30135 );
xor ( n30153 , n30151 , n30152 );
and ( n30154 , n30153 , n29753 );
or ( n30155 , n30150 , n30154 );
buf ( n30156 , n30155 );
not ( n30157 , n30156 );
buf ( n30158 , n30157 );
buf ( n30159 , n30158 );
not ( n30160 , n30159 );
or ( n30161 , n30144 , n30160 );
not ( n30162 , n29753 );
xor ( n30163 , n29163 , n29174 );
xor ( n30164 , n30163 , n29732 );
buf ( n30165 , n30164 );
buf ( n30166 , n30165 );
and ( n30167 , n30162 , n30166 );
not ( n30168 , n30166 );
and ( n30169 , n30151 , n30152 );
xor ( n30170 , n30168 , n30169 );
and ( n30171 , n30170 , n29753 );
or ( n30172 , n30167 , n30171 );
buf ( n30173 , n30172 );
not ( n30174 , n30173 );
buf ( n30175 , n30174 );
buf ( n30176 , n30175 );
not ( n30177 , n30176 );
or ( n30178 , n30161 , n30177 );
not ( n30179 , n29753 );
xor ( n30180 , n29150 , n29161 );
xor ( n30181 , n30180 , n29735 );
buf ( n30182 , n30181 );
buf ( n30183 , n30182 );
and ( n30184 , n30179 , n30183 );
not ( n30185 , n30183 );
and ( n30186 , n30168 , n30169 );
xor ( n30187 , n30185 , n30186 );
and ( n30188 , n30187 , n29753 );
or ( n30189 , n30184 , n30188 );
buf ( n30190 , n30189 );
not ( n30191 , n30190 );
buf ( n30192 , n30191 );
buf ( n30193 , n30192 );
not ( n30194 , n30193 );
or ( n30195 , n30178 , n30194 );
not ( n30196 , n29753 );
xor ( n30197 , n29137 , n29148 );
xor ( n30198 , n30197 , n29738 );
buf ( n30199 , n30198 );
buf ( n30200 , n30199 );
and ( n30201 , n30196 , n30200 );
not ( n30202 , n30200 );
and ( n30203 , n30185 , n30186 );
xor ( n30204 , n30202 , n30203 );
and ( n30205 , n30204 , n29753 );
or ( n30206 , n30201 , n30205 );
buf ( n30207 , n30206 );
not ( n30208 , n30207 );
buf ( n30209 , n30208 );
buf ( n30210 , n30209 );
not ( n30211 , n30210 );
or ( n30212 , n30195 , n30211 );
not ( n30213 , n29753 );
xor ( n30214 , n29124 , n29135 );
xor ( n30215 , n30214 , n29741 );
buf ( n30216 , n30215 );
buf ( n30217 , n30216 );
and ( n30218 , n30213 , n30217 );
not ( n30219 , n30217 );
and ( n30220 , n30202 , n30203 );
xor ( n30221 , n30219 , n30220 );
and ( n30222 , n30221 , n29753 );
or ( n30223 , n30218 , n30222 );
buf ( n30224 , n30223 );
not ( n30225 , n30224 );
buf ( n30226 , n30225 );
buf ( n30227 , n30226 );
not ( n30228 , n30227 );
or ( n30229 , n30212 , n30228 );
not ( n30230 , n29753 );
xor ( n30231 , n29111 , n29122 );
xor ( n30232 , n30231 , n29744 );
buf ( n30233 , n30232 );
buf ( n30234 , n30233 );
and ( n30235 , n30230 , n30234 );
not ( n30236 , n30234 );
and ( n30237 , n30219 , n30220 );
xor ( n30238 , n30236 , n30237 );
and ( n30239 , n30238 , n29753 );
or ( n30240 , n30235 , n30239 );
buf ( n30241 , n30240 );
not ( n30242 , n30241 );
buf ( n30243 , n30242 );
buf ( n30244 , n30243 );
not ( n30245 , n30244 );
or ( n30246 , n30229 , n30245 );
buf ( n30247 , n30246 );
buf ( n30248 , n30247 );
and ( n30249 , n30248 , n29753 );
not ( n30250 , n30249 );
and ( n30251 , n30250 , n29769 );
xor ( n30252 , n29769 , n29753 );
xor ( n30253 , n28901 , n29753 );
and ( n30254 , n30253 , n29753 );
xor ( n30255 , n30252 , n30254 );
and ( n30256 , n30255 , n30249 );
or ( n30257 , n30251 , n30256 );
buf ( n30258 , n30257 );
and ( n30259 , n30258 , n28583 );
and ( n30260 , n24802 , n28591 );
or ( n30261 , n30259 , n30260 );
not ( n30262 , n25216 );
and ( n30263 , n25218 , n25199 , n25208 , n30262 );
and ( n30264 , n25191 , n25199 , n25208 , n30262 );
or ( n30265 , n30263 , n30264 );
nor ( n30266 , n25218 , n25199 , n25208 , n30262 );
or ( n30267 , n30265 , n30266 );
nor ( n30268 , n25218 , n25200 , n25208 , n30262 );
or ( n30269 , n30267 , n30268 );
and ( n30270 , n30261 , n30269 );
buf ( n30271 , n25863 );
buf ( n30272 , n28892 );
xor ( n30273 , n30271 , n30272 );
buf ( n30274 , n30273 );
buf ( n30275 , n30274 );
buf ( n30276 , n30275 );
not ( n30277 , n30276 );
buf ( n30278 , n30277 );
buf ( n30279 , n30278 );
not ( n30280 , n30279 );
buf ( n30281 , n25876 );
buf ( n30282 , n29094 );
xor ( n30283 , n30281 , n30282 );
buf ( n30284 , n27181 );
buf ( n30285 , n29107 );
and ( n30286 , n30284 , n30285 );
buf ( n30287 , n27193 );
buf ( n30288 , n29120 );
and ( n30289 , n30287 , n30288 );
buf ( n30290 , n26807 );
buf ( n30291 , n29133 );
and ( n30292 , n30290 , n30291 );
buf ( n30293 , n26773 );
buf ( n30294 , n29146 );
and ( n30295 , n30293 , n30294 );
buf ( n30296 , n26739 );
buf ( n30297 , n29159 );
and ( n30298 , n30296 , n30297 );
buf ( n30299 , n26705 );
buf ( n30300 , n29172 );
and ( n30301 , n30299 , n30300 );
buf ( n30302 , n26671 );
buf ( n30303 , n29185 );
and ( n30304 , n30302 , n30303 );
buf ( n30305 , n26637 );
buf ( n30306 , n29198 );
and ( n30307 , n30305 , n30306 );
buf ( n30308 , n26603 );
buf ( n30309 , n29211 );
and ( n30310 , n30308 , n30309 );
buf ( n30311 , n26569 );
buf ( n30312 , n29224 );
and ( n30313 , n30311 , n30312 );
buf ( n30314 , n26535 );
buf ( n30315 , n29237 );
and ( n30316 , n30314 , n30315 );
buf ( n30317 , n26501 );
buf ( n30318 , n29295 );
and ( n30319 , n30317 , n30318 );
buf ( n30320 , n26467 );
buf ( n30321 , n29315 );
and ( n30322 , n30320 , n30321 );
buf ( n30323 , n26433 );
buf ( n30324 , n29335 );
and ( n30325 , n30323 , n30324 );
buf ( n30326 , n26399 );
buf ( n30327 , n29355 );
and ( n30328 , n30326 , n30327 );
buf ( n30329 , n26365 );
buf ( n30330 , n29375 );
and ( n30331 , n30329 , n30330 );
buf ( n30332 , n26331 );
buf ( n30333 , n29395 );
and ( n30334 , n30332 , n30333 );
buf ( n30335 , n26297 );
buf ( n30336 , n29415 );
and ( n30337 , n30335 , n30336 );
buf ( n30338 , n26263 );
buf ( n30339 , n29435 );
and ( n30340 , n30338 , n30339 );
buf ( n30341 , n26229 );
buf ( n30342 , n29455 );
and ( n30343 , n30341 , n30342 );
buf ( n30344 , n26195 );
buf ( n30345 , n29475 );
and ( n30346 , n30344 , n30345 );
buf ( n30347 , n26161 );
buf ( n30348 , n29495 );
and ( n30349 , n30347 , n30348 );
buf ( n30350 , n26127 );
buf ( n30351 , n29515 );
and ( n30352 , n30350 , n30351 );
buf ( n30353 , n26093 );
buf ( n30354 , n29535 );
and ( n30355 , n30353 , n30354 );
buf ( n30356 , n26059 );
buf ( n30357 , n29555 );
and ( n30358 , n30356 , n30357 );
buf ( n30359 , n26025 );
buf ( n30360 , n29575 );
and ( n30361 , n30359 , n30360 );
buf ( n30362 , n25991 );
buf ( n30363 , n29595 );
and ( n30364 , n30362 , n30363 );
buf ( n30365 , n25958 );
buf ( n30366 , n29615 );
and ( n30367 , n30365 , n30366 );
buf ( n30368 , n25925 );
buf ( n30369 , n29635 );
and ( n30370 , n30368 , n30369 );
buf ( n30371 , n25894 );
buf ( n30372 , n29655 );
and ( n30373 , n30371 , n30372 );
and ( n30374 , n30271 , n30272 );
and ( n30375 , n30372 , n30374 );
and ( n30376 , n30371 , n30374 );
or ( n30377 , n30373 , n30375 , n30376 );
and ( n30378 , n30369 , n30377 );
and ( n30379 , n30368 , n30377 );
or ( n30380 , n30370 , n30378 , n30379 );
and ( n30381 , n30366 , n30380 );
and ( n30382 , n30365 , n30380 );
or ( n30383 , n30367 , n30381 , n30382 );
and ( n30384 , n30363 , n30383 );
and ( n30385 , n30362 , n30383 );
or ( n30386 , n30364 , n30384 , n30385 );
and ( n30387 , n30360 , n30386 );
and ( n30388 , n30359 , n30386 );
or ( n30389 , n30361 , n30387 , n30388 );
and ( n30390 , n30357 , n30389 );
and ( n30391 , n30356 , n30389 );
or ( n30392 , n30358 , n30390 , n30391 );
and ( n30393 , n30354 , n30392 );
and ( n30394 , n30353 , n30392 );
or ( n30395 , n30355 , n30393 , n30394 );
and ( n30396 , n30351 , n30395 );
and ( n30397 , n30350 , n30395 );
or ( n30398 , n30352 , n30396 , n30397 );
and ( n30399 , n30348 , n30398 );
and ( n30400 , n30347 , n30398 );
or ( n30401 , n30349 , n30399 , n30400 );
and ( n30402 , n30345 , n30401 );
and ( n30403 , n30344 , n30401 );
or ( n30404 , n30346 , n30402 , n30403 );
and ( n30405 , n30342 , n30404 );
and ( n30406 , n30341 , n30404 );
or ( n30407 , n30343 , n30405 , n30406 );
and ( n30408 , n30339 , n30407 );
and ( n30409 , n30338 , n30407 );
or ( n30410 , n30340 , n30408 , n30409 );
and ( n30411 , n30336 , n30410 );
and ( n30412 , n30335 , n30410 );
or ( n30413 , n30337 , n30411 , n30412 );
and ( n30414 , n30333 , n30413 );
and ( n30415 , n30332 , n30413 );
or ( n30416 , n30334 , n30414 , n30415 );
and ( n30417 , n30330 , n30416 );
and ( n30418 , n30329 , n30416 );
or ( n30419 , n30331 , n30417 , n30418 );
and ( n30420 , n30327 , n30419 );
and ( n30421 , n30326 , n30419 );
or ( n30422 , n30328 , n30420 , n30421 );
and ( n30423 , n30324 , n30422 );
and ( n30424 , n30323 , n30422 );
or ( n30425 , n30325 , n30423 , n30424 );
and ( n30426 , n30321 , n30425 );
and ( n30427 , n30320 , n30425 );
or ( n30428 , n30322 , n30426 , n30427 );
and ( n30429 , n30318 , n30428 );
and ( n30430 , n30317 , n30428 );
or ( n30431 , n30319 , n30429 , n30430 );
and ( n30432 , n30315 , n30431 );
and ( n30433 , n30314 , n30431 );
or ( n30434 , n30316 , n30432 , n30433 );
and ( n30435 , n30312 , n30434 );
and ( n30436 , n30311 , n30434 );
or ( n30437 , n30313 , n30435 , n30436 );
and ( n30438 , n30309 , n30437 );
and ( n30439 , n30308 , n30437 );
or ( n30440 , n30310 , n30438 , n30439 );
and ( n30441 , n30306 , n30440 );
and ( n30442 , n30305 , n30440 );
or ( n30443 , n30307 , n30441 , n30442 );
and ( n30444 , n30303 , n30443 );
and ( n30445 , n30302 , n30443 );
or ( n30446 , n30304 , n30444 , n30445 );
and ( n30447 , n30300 , n30446 );
and ( n30448 , n30299 , n30446 );
or ( n30449 , n30301 , n30447 , n30448 );
and ( n30450 , n30297 , n30449 );
and ( n30451 , n30296 , n30449 );
or ( n30452 , n30298 , n30450 , n30451 );
and ( n30453 , n30294 , n30452 );
and ( n30454 , n30293 , n30452 );
or ( n30455 , n30295 , n30453 , n30454 );
and ( n30456 , n30291 , n30455 );
and ( n30457 , n30290 , n30455 );
or ( n30458 , n30292 , n30456 , n30457 );
and ( n30459 , n30288 , n30458 );
and ( n30460 , n30287 , n30458 );
or ( n30461 , n30289 , n30459 , n30460 );
and ( n30462 , n30285 , n30461 );
and ( n30463 , n30284 , n30461 );
or ( n30464 , n30286 , n30462 , n30463 );
xor ( n30465 , n30283 , n30464 );
buf ( n30466 , n30465 );
buf ( n30467 , n30466 );
not ( n30468 , n30467 );
xor ( n30469 , n30371 , n30372 );
xor ( n30470 , n30469 , n30374 );
buf ( n30471 , n30470 );
buf ( n30472 , n30471 );
and ( n30473 , n30468 , n30472 );
not ( n30474 , n30472 );
not ( n30475 , n30275 );
xor ( n30476 , n30474 , n30475 );
and ( n30477 , n30476 , n30467 );
or ( n30478 , n30473 , n30477 );
buf ( n30479 , n30478 );
not ( n30480 , n30479 );
buf ( n30481 , n30480 );
buf ( n30482 , n30481 );
not ( n30483 , n30482 );
or ( n30484 , n30280 , n30483 );
not ( n30485 , n30467 );
xor ( n30486 , n30368 , n30369 );
xor ( n30487 , n30486 , n30377 );
buf ( n30488 , n30487 );
buf ( n30489 , n30488 );
and ( n30490 , n30485 , n30489 );
not ( n30491 , n30489 );
and ( n30492 , n30474 , n30475 );
xor ( n30493 , n30491 , n30492 );
and ( n30494 , n30493 , n30467 );
or ( n30495 , n30490 , n30494 );
buf ( n30496 , n30495 );
not ( n30497 , n30496 );
buf ( n30498 , n30497 );
buf ( n30499 , n30498 );
not ( n30500 , n30499 );
or ( n30501 , n30484 , n30500 );
not ( n30502 , n30467 );
xor ( n30503 , n30365 , n30366 );
xor ( n30504 , n30503 , n30380 );
buf ( n30505 , n30504 );
buf ( n30506 , n30505 );
and ( n30507 , n30502 , n30506 );
not ( n30508 , n30506 );
and ( n30509 , n30491 , n30492 );
xor ( n30510 , n30508 , n30509 );
and ( n30511 , n30510 , n30467 );
or ( n30512 , n30507 , n30511 );
buf ( n30513 , n30512 );
not ( n30514 , n30513 );
buf ( n30515 , n30514 );
buf ( n30516 , n30515 );
not ( n30517 , n30516 );
or ( n30518 , n30501 , n30517 );
not ( n30519 , n30467 );
xor ( n30520 , n30362 , n30363 );
xor ( n30521 , n30520 , n30383 );
buf ( n30522 , n30521 );
buf ( n30523 , n30522 );
and ( n30524 , n30519 , n30523 );
not ( n30525 , n30523 );
and ( n30526 , n30508 , n30509 );
xor ( n30527 , n30525 , n30526 );
and ( n30528 , n30527 , n30467 );
or ( n30529 , n30524 , n30528 );
buf ( n30530 , n30529 );
not ( n30531 , n30530 );
buf ( n30532 , n30531 );
buf ( n30533 , n30532 );
not ( n30534 , n30533 );
or ( n30535 , n30518 , n30534 );
not ( n30536 , n30467 );
xor ( n30537 , n30359 , n30360 );
xor ( n30538 , n30537 , n30386 );
buf ( n30539 , n30538 );
buf ( n30540 , n30539 );
and ( n30541 , n30536 , n30540 );
not ( n30542 , n30540 );
and ( n30543 , n30525 , n30526 );
xor ( n30544 , n30542 , n30543 );
and ( n30545 , n30544 , n30467 );
or ( n30546 , n30541 , n30545 );
buf ( n30547 , n30546 );
not ( n30548 , n30547 );
buf ( n30549 , n30548 );
buf ( n30550 , n30549 );
not ( n30551 , n30550 );
or ( n30552 , n30535 , n30551 );
not ( n30553 , n30467 );
xor ( n30554 , n30356 , n30357 );
xor ( n30555 , n30554 , n30389 );
buf ( n30556 , n30555 );
buf ( n30557 , n30556 );
and ( n30558 , n30553 , n30557 );
not ( n30559 , n30557 );
and ( n30560 , n30542 , n30543 );
xor ( n30561 , n30559 , n30560 );
and ( n30562 , n30561 , n30467 );
or ( n30563 , n30558 , n30562 );
buf ( n30564 , n30563 );
not ( n30565 , n30564 );
buf ( n30566 , n30565 );
buf ( n30567 , n30566 );
not ( n30568 , n30567 );
or ( n30569 , n30552 , n30568 );
not ( n30570 , n30467 );
xor ( n30571 , n30353 , n30354 );
xor ( n30572 , n30571 , n30392 );
buf ( n30573 , n30572 );
buf ( n30574 , n30573 );
and ( n30575 , n30570 , n30574 );
not ( n30576 , n30574 );
and ( n30577 , n30559 , n30560 );
xor ( n30578 , n30576 , n30577 );
and ( n30579 , n30578 , n30467 );
or ( n30580 , n30575 , n30579 );
buf ( n30581 , n30580 );
not ( n30582 , n30581 );
buf ( n30583 , n30582 );
buf ( n30584 , n30583 );
not ( n30585 , n30584 );
or ( n30586 , n30569 , n30585 );
not ( n30587 , n30467 );
xor ( n30588 , n30350 , n30351 );
xor ( n30589 , n30588 , n30395 );
buf ( n30590 , n30589 );
buf ( n30591 , n30590 );
and ( n30592 , n30587 , n30591 );
not ( n30593 , n30591 );
and ( n30594 , n30576 , n30577 );
xor ( n30595 , n30593 , n30594 );
and ( n30596 , n30595 , n30467 );
or ( n30597 , n30592 , n30596 );
buf ( n30598 , n30597 );
not ( n30599 , n30598 );
buf ( n30600 , n30599 );
buf ( n30601 , n30600 );
not ( n30602 , n30601 );
or ( n30603 , n30586 , n30602 );
not ( n30604 , n30467 );
xor ( n30605 , n30347 , n30348 );
xor ( n30606 , n30605 , n30398 );
buf ( n30607 , n30606 );
buf ( n30608 , n30607 );
and ( n30609 , n30604 , n30608 );
not ( n30610 , n30608 );
and ( n30611 , n30593 , n30594 );
xor ( n30612 , n30610 , n30611 );
and ( n30613 , n30612 , n30467 );
or ( n30614 , n30609 , n30613 );
buf ( n30615 , n30614 );
not ( n30616 , n30615 );
buf ( n30617 , n30616 );
buf ( n30618 , n30617 );
not ( n30619 , n30618 );
or ( n30620 , n30603 , n30619 );
not ( n30621 , n30467 );
xor ( n30622 , n30344 , n30345 );
xor ( n30623 , n30622 , n30401 );
buf ( n30624 , n30623 );
buf ( n30625 , n30624 );
and ( n30626 , n30621 , n30625 );
not ( n30627 , n30625 );
and ( n30628 , n30610 , n30611 );
xor ( n30629 , n30627 , n30628 );
and ( n30630 , n30629 , n30467 );
or ( n30631 , n30626 , n30630 );
buf ( n30632 , n30631 );
not ( n30633 , n30632 );
buf ( n30634 , n30633 );
buf ( n30635 , n30634 );
not ( n30636 , n30635 );
or ( n30637 , n30620 , n30636 );
not ( n30638 , n30467 );
xor ( n30639 , n30341 , n30342 );
xor ( n30640 , n30639 , n30404 );
buf ( n30641 , n30640 );
buf ( n30642 , n30641 );
and ( n30643 , n30638 , n30642 );
not ( n30644 , n30642 );
and ( n30645 , n30627 , n30628 );
xor ( n30646 , n30644 , n30645 );
and ( n30647 , n30646 , n30467 );
or ( n30648 , n30643 , n30647 );
buf ( n30649 , n30648 );
not ( n30650 , n30649 );
buf ( n30651 , n30650 );
buf ( n30652 , n30651 );
not ( n30653 , n30652 );
or ( n30654 , n30637 , n30653 );
not ( n30655 , n30467 );
xor ( n30656 , n30338 , n30339 );
xor ( n30657 , n30656 , n30407 );
buf ( n30658 , n30657 );
buf ( n30659 , n30658 );
and ( n30660 , n30655 , n30659 );
not ( n30661 , n30659 );
and ( n30662 , n30644 , n30645 );
xor ( n30663 , n30661 , n30662 );
and ( n30664 , n30663 , n30467 );
or ( n30665 , n30660 , n30664 );
buf ( n30666 , n30665 );
not ( n30667 , n30666 );
buf ( n30668 , n30667 );
buf ( n30669 , n30668 );
not ( n30670 , n30669 );
or ( n30671 , n30654 , n30670 );
not ( n30672 , n30467 );
xor ( n30673 , n30335 , n30336 );
xor ( n30674 , n30673 , n30410 );
buf ( n30675 , n30674 );
buf ( n30676 , n30675 );
and ( n30677 , n30672 , n30676 );
not ( n30678 , n30676 );
and ( n30679 , n30661 , n30662 );
xor ( n30680 , n30678 , n30679 );
and ( n30681 , n30680 , n30467 );
or ( n30682 , n30677 , n30681 );
buf ( n30683 , n30682 );
not ( n30684 , n30683 );
buf ( n30685 , n30684 );
buf ( n30686 , n30685 );
not ( n30687 , n30686 );
or ( n30688 , n30671 , n30687 );
not ( n30689 , n30467 );
xor ( n30690 , n30332 , n30333 );
xor ( n30691 , n30690 , n30413 );
buf ( n30692 , n30691 );
buf ( n30693 , n30692 );
and ( n30694 , n30689 , n30693 );
not ( n30695 , n30693 );
and ( n30696 , n30678 , n30679 );
xor ( n30697 , n30695 , n30696 );
and ( n30698 , n30697 , n30467 );
or ( n30699 , n30694 , n30698 );
buf ( n30700 , n30699 );
not ( n30701 , n30700 );
buf ( n30702 , n30701 );
buf ( n30703 , n30702 );
not ( n30704 , n30703 );
or ( n30705 , n30688 , n30704 );
not ( n30706 , n30467 );
xor ( n30707 , n30329 , n30330 );
xor ( n30708 , n30707 , n30416 );
buf ( n30709 , n30708 );
buf ( n30710 , n30709 );
and ( n30711 , n30706 , n30710 );
not ( n30712 , n30710 );
and ( n30713 , n30695 , n30696 );
xor ( n30714 , n30712 , n30713 );
and ( n30715 , n30714 , n30467 );
or ( n30716 , n30711 , n30715 );
buf ( n30717 , n30716 );
not ( n30718 , n30717 );
buf ( n30719 , n30718 );
buf ( n30720 , n30719 );
not ( n30721 , n30720 );
or ( n30722 , n30705 , n30721 );
not ( n30723 , n30467 );
xor ( n30724 , n30326 , n30327 );
xor ( n30725 , n30724 , n30419 );
buf ( n30726 , n30725 );
buf ( n30727 , n30726 );
and ( n30728 , n30723 , n30727 );
not ( n30729 , n30727 );
and ( n30730 , n30712 , n30713 );
xor ( n30731 , n30729 , n30730 );
and ( n30732 , n30731 , n30467 );
or ( n30733 , n30728 , n30732 );
buf ( n30734 , n30733 );
not ( n30735 , n30734 );
buf ( n30736 , n30735 );
buf ( n30737 , n30736 );
not ( n30738 , n30737 );
or ( n30739 , n30722 , n30738 );
not ( n30740 , n30467 );
xor ( n30741 , n30323 , n30324 );
xor ( n30742 , n30741 , n30422 );
buf ( n30743 , n30742 );
buf ( n30744 , n30743 );
and ( n30745 , n30740 , n30744 );
not ( n30746 , n30744 );
and ( n30747 , n30729 , n30730 );
xor ( n30748 , n30746 , n30747 );
and ( n30749 , n30748 , n30467 );
or ( n30750 , n30745 , n30749 );
buf ( n30751 , n30750 );
not ( n30752 , n30751 );
buf ( n30753 , n30752 );
buf ( n30754 , n30753 );
not ( n30755 , n30754 );
or ( n30756 , n30739 , n30755 );
not ( n30757 , n30467 );
xor ( n30758 , n30320 , n30321 );
xor ( n30759 , n30758 , n30425 );
buf ( n30760 , n30759 );
buf ( n30761 , n30760 );
and ( n30762 , n30757 , n30761 );
not ( n30763 , n30761 );
and ( n30764 , n30746 , n30747 );
xor ( n30765 , n30763 , n30764 );
and ( n30766 , n30765 , n30467 );
or ( n30767 , n30762 , n30766 );
buf ( n30768 , n30767 );
not ( n30769 , n30768 );
buf ( n30770 , n30769 );
buf ( n30771 , n30770 );
not ( n30772 , n30771 );
or ( n30773 , n30756 , n30772 );
not ( n30774 , n30467 );
xor ( n30775 , n30317 , n30318 );
xor ( n30776 , n30775 , n30428 );
buf ( n30777 , n30776 );
buf ( n30778 , n30777 );
and ( n30779 , n30774 , n30778 );
not ( n30780 , n30778 );
and ( n30781 , n30763 , n30764 );
xor ( n30782 , n30780 , n30781 );
and ( n30783 , n30782 , n30467 );
or ( n30784 , n30779 , n30783 );
buf ( n30785 , n30784 );
not ( n30786 , n30785 );
buf ( n30787 , n30786 );
buf ( n30788 , n30787 );
not ( n30789 , n30788 );
or ( n30790 , n30773 , n30789 );
not ( n30791 , n30467 );
xor ( n30792 , n30314 , n30315 );
xor ( n30793 , n30792 , n30431 );
buf ( n30794 , n30793 );
buf ( n30795 , n30794 );
and ( n30796 , n30791 , n30795 );
not ( n30797 , n30795 );
and ( n30798 , n30780 , n30781 );
xor ( n30799 , n30797 , n30798 );
and ( n30800 , n30799 , n30467 );
or ( n30801 , n30796 , n30800 );
buf ( n30802 , n30801 );
not ( n30803 , n30802 );
buf ( n30804 , n30803 );
buf ( n30805 , n30804 );
not ( n30806 , n30805 );
or ( n30807 , n30790 , n30806 );
not ( n30808 , n30467 );
xor ( n30809 , n30311 , n30312 );
xor ( n30810 , n30809 , n30434 );
buf ( n30811 , n30810 );
buf ( n30812 , n30811 );
and ( n30813 , n30808 , n30812 );
not ( n30814 , n30812 );
and ( n30815 , n30797 , n30798 );
xor ( n30816 , n30814 , n30815 );
and ( n30817 , n30816 , n30467 );
or ( n30818 , n30813 , n30817 );
buf ( n30819 , n30818 );
not ( n30820 , n30819 );
buf ( n30821 , n30820 );
buf ( n30822 , n30821 );
not ( n30823 , n30822 );
or ( n30824 , n30807 , n30823 );
not ( n30825 , n30467 );
xor ( n30826 , n30308 , n30309 );
xor ( n30827 , n30826 , n30437 );
buf ( n30828 , n30827 );
buf ( n30829 , n30828 );
and ( n30830 , n30825 , n30829 );
not ( n30831 , n30829 );
and ( n30832 , n30814 , n30815 );
xor ( n30833 , n30831 , n30832 );
and ( n30834 , n30833 , n30467 );
or ( n30835 , n30830 , n30834 );
buf ( n30836 , n30835 );
not ( n30837 , n30836 );
buf ( n30838 , n30837 );
buf ( n30839 , n30838 );
not ( n30840 , n30839 );
or ( n30841 , n30824 , n30840 );
not ( n30842 , n30467 );
xor ( n30843 , n30305 , n30306 );
xor ( n30844 , n30843 , n30440 );
buf ( n30845 , n30844 );
buf ( n30846 , n30845 );
and ( n30847 , n30842 , n30846 );
not ( n30848 , n30846 );
and ( n30849 , n30831 , n30832 );
xor ( n30850 , n30848 , n30849 );
and ( n30851 , n30850 , n30467 );
or ( n30852 , n30847 , n30851 );
buf ( n30853 , n30852 );
not ( n30854 , n30853 );
buf ( n30855 , n30854 );
buf ( n30856 , n30855 );
not ( n30857 , n30856 );
or ( n30858 , n30841 , n30857 );
not ( n30859 , n30467 );
xor ( n30860 , n30302 , n30303 );
xor ( n30861 , n30860 , n30443 );
buf ( n30862 , n30861 );
buf ( n30863 , n30862 );
and ( n30864 , n30859 , n30863 );
not ( n30865 , n30863 );
and ( n30866 , n30848 , n30849 );
xor ( n30867 , n30865 , n30866 );
and ( n30868 , n30867 , n30467 );
or ( n30869 , n30864 , n30868 );
buf ( n30870 , n30869 );
not ( n30871 , n30870 );
buf ( n30872 , n30871 );
buf ( n30873 , n30872 );
not ( n30874 , n30873 );
or ( n30875 , n30858 , n30874 );
not ( n30876 , n30467 );
xor ( n30877 , n30299 , n30300 );
xor ( n30878 , n30877 , n30446 );
buf ( n30879 , n30878 );
buf ( n30880 , n30879 );
and ( n30881 , n30876 , n30880 );
not ( n30882 , n30880 );
and ( n30883 , n30865 , n30866 );
xor ( n30884 , n30882 , n30883 );
and ( n30885 , n30884 , n30467 );
or ( n30886 , n30881 , n30885 );
buf ( n30887 , n30886 );
not ( n30888 , n30887 );
buf ( n30889 , n30888 );
buf ( n30890 , n30889 );
not ( n30891 , n30890 );
or ( n30892 , n30875 , n30891 );
not ( n30893 , n30467 );
xor ( n30894 , n30296 , n30297 );
xor ( n30895 , n30894 , n30449 );
buf ( n30896 , n30895 );
buf ( n30897 , n30896 );
and ( n30898 , n30893 , n30897 );
not ( n30899 , n30897 );
and ( n30900 , n30882 , n30883 );
xor ( n30901 , n30899 , n30900 );
and ( n30902 , n30901 , n30467 );
or ( n30903 , n30898 , n30902 );
buf ( n30904 , n30903 );
not ( n30905 , n30904 );
buf ( n30906 , n30905 );
buf ( n30907 , n30906 );
not ( n30908 , n30907 );
or ( n30909 , n30892 , n30908 );
not ( n30910 , n30467 );
xor ( n30911 , n30293 , n30294 );
xor ( n30912 , n30911 , n30452 );
buf ( n30913 , n30912 );
buf ( n30914 , n30913 );
and ( n30915 , n30910 , n30914 );
not ( n30916 , n30914 );
and ( n30917 , n30899 , n30900 );
xor ( n30918 , n30916 , n30917 );
and ( n30919 , n30918 , n30467 );
or ( n30920 , n30915 , n30919 );
buf ( n30921 , n30920 );
not ( n30922 , n30921 );
buf ( n30923 , n30922 );
buf ( n30924 , n30923 );
not ( n30925 , n30924 );
or ( n30926 , n30909 , n30925 );
not ( n30927 , n30467 );
xor ( n30928 , n30290 , n30291 );
xor ( n30929 , n30928 , n30455 );
buf ( n30930 , n30929 );
buf ( n30931 , n30930 );
and ( n30932 , n30927 , n30931 );
not ( n30933 , n30931 );
and ( n30934 , n30916 , n30917 );
xor ( n30935 , n30933 , n30934 );
and ( n30936 , n30935 , n30467 );
or ( n30937 , n30932 , n30936 );
buf ( n30938 , n30937 );
not ( n30939 , n30938 );
buf ( n30940 , n30939 );
buf ( n30941 , n30940 );
not ( n30942 , n30941 );
or ( n30943 , n30926 , n30942 );
not ( n30944 , n30467 );
xor ( n30945 , n30287 , n30288 );
xor ( n30946 , n30945 , n30458 );
buf ( n30947 , n30946 );
buf ( n30948 , n30947 );
and ( n30949 , n30944 , n30948 );
not ( n30950 , n30948 );
and ( n30951 , n30933 , n30934 );
xor ( n30952 , n30950 , n30951 );
and ( n30953 , n30952 , n30467 );
or ( n30954 , n30949 , n30953 );
buf ( n30955 , n30954 );
not ( n30956 , n30955 );
buf ( n30957 , n30956 );
buf ( n30958 , n30957 );
not ( n30959 , n30958 );
or ( n30960 , n30943 , n30959 );
buf ( n30961 , n30960 );
buf ( n30962 , n30961 );
and ( n30963 , n30962 , n30467 );
not ( n30964 , n30963 );
and ( n30965 , n30964 , n30483 );
xor ( n30966 , n30483 , n30467 );
xor ( n30967 , n30280 , n30467 );
and ( n30968 , n30967 , n30467 );
xor ( n30969 , n30966 , n30968 );
and ( n30970 , n30969 , n30963 );
or ( n30971 , n30965 , n30970 );
buf ( n30972 , n30971 );
and ( n30973 , n30972 , n28583 );
and ( n30974 , n24802 , n28591 );
or ( n30975 , n30973 , n30974 );
and ( n30976 , n25218 , n25200 , n25208 , n30262 );
and ( n30977 , n25191 , n25200 , n25208 , n30262 );
or ( n30978 , n30976 , n30977 );
nor ( n30979 , n25191 , n25199 , n25208 , n30262 );
or ( n30980 , n30978 , n30979 );
nor ( n30981 , n25191 , n25200 , n25208 , n30262 );
or ( n30982 , n30980 , n30981 );
and ( n30983 , n30975 , n30982 );
and ( n30984 , n29655 , n28583 );
and ( n30985 , n24802 , n28591 );
or ( n30986 , n30984 , n30985 );
nor ( n30987 , n25191 , n25200 , n25208 , n25216 );
nor ( n30988 , n25218 , n25200 , n25208 , n25216 );
or ( n30989 , n30987 , n30988 );
and ( n30990 , n30986 , n30989 );
nor ( n30991 , n25218 , n25199 , n25208 , n25216 );
and ( n30992 , n25887 , n30991 );
buf ( n30993 , n29655 );
not ( n30994 , n30993 );
buf ( n30995 , n28892 );
not ( n30996 , n30995 );
xor ( n30997 , n30994 , n30996 );
buf ( n30998 , n30997 );
and ( n30999 , n30998 , n28583 );
and ( n31000 , n24802 , n28591 );
or ( n31001 , n30999 , n31000 );
nor ( n31002 , n25191 , n25199 , n25208 , n25216 );
and ( n31003 , n31001 , n31002 );
or ( n31004 , n25223 , n28595 , n30270 , n30983 , n30990 , n30992 , n31003 );
and ( n31005 , n24801 , n31004 );
and ( n31006 , n24802 , n24800 );
or ( n31007 , n31005 , n31006 );
buf ( n31008 , n10617 );
and ( n31009 , n31007 , n31008 );
and ( n31010 , n24802 , n10618 );
or ( n31011 , n31009 , n31010 );
buf ( n31012 , n31011 );
buf ( n31013 , n31012 );
not ( n31014 , n24800 );
and ( n31015 , n26187 , n25222 );
not ( n31016 , n26823 );
and ( n31017 , n31016 , n26173 );
xor ( n31018 , n26173 , n25877 );
xor ( n31019 , n26139 , n25877 );
xor ( n31020 , n26105 , n25877 );
xor ( n31021 , n26071 , n25877 );
xor ( n31022 , n26037 , n25877 );
xor ( n31023 , n26003 , n25877 );
xor ( n31024 , n25970 , n25877 );
xor ( n31025 , n25937 , n25877 );
xor ( n31026 , n25906 , n25877 );
and ( n31027 , n26826 , n25877 );
and ( n31028 , n31026 , n31027 );
and ( n31029 , n31025 , n31028 );
and ( n31030 , n31024 , n31029 );
and ( n31031 , n31023 , n31030 );
and ( n31032 , n31022 , n31031 );
and ( n31033 , n31021 , n31032 );
and ( n31034 , n31020 , n31033 );
and ( n31035 , n31019 , n31034 );
xor ( n31036 , n31018 , n31035 );
and ( n31037 , n31036 , n26823 );
or ( n31038 , n31017 , n31037 );
buf ( n31039 , n31038 );
and ( n31040 , n31039 , n27046 );
and ( n31041 , n31039 , n27049 );
not ( n31042 , n27051 );
and ( n31043 , n31042 , n28082 );
not ( n31044 , n28494 );
and ( n31045 , n31044 , n28094 );
xor ( n31046 , n28094 , n27883 );
xor ( n31047 , n28072 , n27883 );
xor ( n31048 , n28050 , n27883 );
xor ( n31049 , n28028 , n27883 );
xor ( n31050 , n28006 , n27883 );
xor ( n31051 , n27984 , n27883 );
xor ( n31052 , n27962 , n27883 );
xor ( n31053 , n27940 , n27883 );
xor ( n31054 , n27918 , n27883 );
and ( n31055 , n28497 , n28499 );
and ( n31056 , n31054 , n31055 );
and ( n31057 , n31053 , n31056 );
and ( n31058 , n31052 , n31057 );
and ( n31059 , n31051 , n31058 );
and ( n31060 , n31050 , n31059 );
and ( n31061 , n31049 , n31060 );
and ( n31062 , n31048 , n31061 );
and ( n31063 , n31047 , n31062 );
xor ( n31064 , n31046 , n31063 );
and ( n31065 , n31064 , n28494 );
or ( n31066 , n31045 , n31065 );
buf ( n31067 , n31066 );
and ( n31068 , n31067 , n27051 );
or ( n31069 , n31043 , n31068 );
and ( n31070 , n31069 , n28506 );
and ( n31071 , n28082 , n28508 );
or ( n31072 , n31040 , n31041 , n31070 , n31071 );
and ( n31073 , n31072 , n28589 );
or ( n31074 , n28588 , n28583 );
or ( n31075 , n31074 , C0 );
and ( n31076 , n26187 , n31075 );
or ( n31077 , n31073 , n31076 );
and ( n31078 , n31077 , n28594 );
not ( n31079 , n30249 );
and ( n31080 , n31079 , n29922 );
xor ( n31081 , n29922 , n29753 );
xor ( n31082 , n29905 , n29753 );
xor ( n31083 , n29888 , n29753 );
xor ( n31084 , n29871 , n29753 );
xor ( n31085 , n29854 , n29753 );
xor ( n31086 , n29837 , n29753 );
xor ( n31087 , n29820 , n29753 );
xor ( n31088 , n29803 , n29753 );
xor ( n31089 , n29786 , n29753 );
and ( n31090 , n30252 , n30254 );
and ( n31091 , n31089 , n31090 );
and ( n31092 , n31088 , n31091 );
and ( n31093 , n31087 , n31092 );
and ( n31094 , n31086 , n31093 );
and ( n31095 , n31085 , n31094 );
and ( n31096 , n31084 , n31095 );
and ( n31097 , n31083 , n31096 );
and ( n31098 , n31082 , n31097 );
xor ( n31099 , n31081 , n31098 );
and ( n31100 , n31099 , n30249 );
or ( n31101 , n31080 , n31100 );
buf ( n31102 , n31101 );
and ( n31103 , n31102 , n28589 );
and ( n31104 , n26187 , n31075 );
or ( n31105 , n31103 , n31104 );
and ( n31106 , n31105 , n30269 );
not ( n31107 , n30963 );
and ( n31108 , n31107 , n30636 );
xor ( n31109 , n30636 , n30467 );
xor ( n31110 , n30619 , n30467 );
xor ( n31111 , n30602 , n30467 );
xor ( n31112 , n30585 , n30467 );
xor ( n31113 , n30568 , n30467 );
xor ( n31114 , n30551 , n30467 );
xor ( n31115 , n30534 , n30467 );
xor ( n31116 , n30517 , n30467 );
xor ( n31117 , n30500 , n30467 );
and ( n31118 , n30966 , n30968 );
and ( n31119 , n31117 , n31118 );
and ( n31120 , n31116 , n31119 );
and ( n31121 , n31115 , n31120 );
and ( n31122 , n31114 , n31121 );
and ( n31123 , n31113 , n31122 );
and ( n31124 , n31112 , n31123 );
and ( n31125 , n31111 , n31124 );
and ( n31126 , n31110 , n31125 );
xor ( n31127 , n31109 , n31126 );
and ( n31128 , n31127 , n30963 );
or ( n31129 , n31108 , n31128 );
buf ( n31130 , n31129 );
and ( n31131 , n31130 , n28589 );
and ( n31132 , n26187 , n31075 );
or ( n31133 , n31131 , n31132 );
and ( n31134 , n31133 , n30982 );
and ( n31135 , n29475 , n28589 );
and ( n31136 , n26187 , n31075 );
or ( n31137 , n31135 , n31136 );
and ( n31138 , n31137 , n30989 );
and ( n31139 , n29475 , n30991 );
buf ( n31140 , n29475 );
not ( n31141 , n31140 );
buf ( n31142 , n29495 );
not ( n31143 , n31142 );
buf ( n31144 , n29515 );
not ( n31145 , n31144 );
buf ( n31146 , n29535 );
not ( n31147 , n31146 );
buf ( n31148 , n29555 );
not ( n31149 , n31148 );
buf ( n31150 , n29575 );
not ( n31151 , n31150 );
buf ( n31152 , n29595 );
not ( n31153 , n31152 );
buf ( n31154 , n29615 );
not ( n31155 , n31154 );
buf ( n31156 , n29635 );
not ( n31157 , n31156 );
and ( n31158 , n30994 , n30996 );
and ( n31159 , n31157 , n31158 );
and ( n31160 , n31155 , n31159 );
and ( n31161 , n31153 , n31160 );
and ( n31162 , n31151 , n31161 );
and ( n31163 , n31149 , n31162 );
and ( n31164 , n31147 , n31163 );
and ( n31165 , n31145 , n31164 );
and ( n31166 , n31143 , n31165 );
xor ( n31167 , n31141 , n31166 );
buf ( n31168 , n31167 );
and ( n31169 , n31168 , n28589 );
and ( n31170 , n26187 , n31075 );
or ( n31171 , n31169 , n31170 );
and ( n31172 , n31171 , n31002 );
or ( n31173 , n31015 , n31078 , n31106 , n31134 , n31138 , n31139 , n31172 );
and ( n31174 , n31014 , n31173 );
and ( n31175 , n26187 , n24800 );
or ( n31176 , n31174 , n31175 );
and ( n31177 , n31176 , n31008 );
and ( n31178 , n25369 , n10618 );
or ( n31179 , n31177 , n31178 );
buf ( n31180 , n31179 );
buf ( n31181 , n31180 );
buf ( n31182 , n10615 );
buf ( n31183 , n10613 );
buf ( n31184 , n10615 );
not ( n31185 , n11954 );
not ( n31186 , n12243 );
or ( n31187 , n14562 , n14592 );
and ( n31188 , n10628 , n31187 );
buf ( n31189 , n15864 );
buf ( n31190 , n13508 );
xor ( n31191 , n31189 , n31190 );
buf ( n31192 , n31191 );
buf ( n31193 , n31192 );
buf ( n31194 , n31193 );
not ( n31195 , n31194 );
buf ( n31196 , n31195 );
buf ( n31197 , n31196 );
not ( n31198 , n31197 );
buf ( n31199 , n13140 );
not ( n31200 , n31199 );
buf ( n31201 , n14605 );
not ( n31202 , n31201 );
buf ( n31203 , n14958 );
not ( n31204 , n31203 );
buf ( n31205 , n13156 );
not ( n31206 , n31205 );
buf ( n31207 , n13169 );
not ( n31208 , n31207 );
buf ( n31209 , n13181 );
not ( n31210 , n31209 );
buf ( n31211 , n13193 );
not ( n31212 , n31211 );
buf ( n31213 , n13205 );
not ( n31214 , n31213 );
buf ( n31215 , n13217 );
not ( n31216 , n31215 );
buf ( n31217 , n13229 );
not ( n31218 , n31217 );
buf ( n31219 , n13241 );
not ( n31220 , n31219 );
buf ( n31221 , n13253 );
not ( n31222 , n31221 );
buf ( n31223 , n15447 );
buf ( n31224 , n13265 );
not ( n31225 , n31224 );
and ( n31226 , n31223 , n31225 );
buf ( n31227 , n15469 );
buf ( n31228 , n13277 );
not ( n31229 , n31228 );
and ( n31230 , n31227 , n31229 );
buf ( n31231 , n15491 );
buf ( n31232 , n13289 );
not ( n31233 , n31232 );
and ( n31234 , n31231 , n31233 );
buf ( n31235 , n15513 );
buf ( n31236 , n13301 );
not ( n31237 , n31236 );
and ( n31238 , n31235 , n31237 );
buf ( n31239 , n15535 );
buf ( n31240 , n13313 );
not ( n31241 , n31240 );
and ( n31242 , n31239 , n31241 );
buf ( n31243 , n15557 );
buf ( n31244 , n13325 );
not ( n31245 , n31244 );
and ( n31246 , n31243 , n31245 );
buf ( n31247 , n15579 );
buf ( n31248 , n13337 );
not ( n31249 , n31248 );
and ( n31250 , n31247 , n31249 );
buf ( n31251 , n15601 );
buf ( n31252 , n13349 );
not ( n31253 , n31252 );
and ( n31254 , n31251 , n31253 );
buf ( n31255 , n15623 );
buf ( n31256 , n13361 );
not ( n31257 , n31256 );
and ( n31258 , n31255 , n31257 );
buf ( n31259 , n15645 );
buf ( n31260 , n13373 );
not ( n31261 , n31260 );
and ( n31262 , n31259 , n31261 );
buf ( n31263 , n15667 );
buf ( n31264 , n13385 );
not ( n31265 , n31264 );
and ( n31266 , n31263 , n31265 );
buf ( n31267 , n15689 );
buf ( n31268 , n13397 );
not ( n31269 , n31268 );
and ( n31270 , n31267 , n31269 );
buf ( n31271 , n15711 );
buf ( n31272 , n13409 );
not ( n31273 , n31272 );
and ( n31274 , n31271 , n31273 );
buf ( n31275 , n15733 );
buf ( n31276 , n13421 );
not ( n31277 , n31276 );
and ( n31278 , n31275 , n31277 );
buf ( n31279 , n15755 );
buf ( n31280 , n13433 );
not ( n31281 , n31280 );
and ( n31282 , n31279 , n31281 );
buf ( n31283 , n15777 );
buf ( n31284 , n13445 );
not ( n31285 , n31284 );
and ( n31286 , n31283 , n31285 );
buf ( n31287 , n15799 );
buf ( n31288 , n13457 );
not ( n31289 , n31288 );
and ( n31290 , n31287 , n31289 );
buf ( n31291 , n15821 );
buf ( n31292 , n13474 );
not ( n31293 , n31292 );
and ( n31294 , n31291 , n31293 );
buf ( n31295 , n15843 );
buf ( n31296 , n13491 );
not ( n31297 , n31296 );
and ( n31298 , n31295 , n31297 );
not ( n31299 , n31190 );
or ( n31300 , n31189 , n31299 );
and ( n31301 , n31297 , n31300 );
and ( n31302 , n31295 , n31300 );
or ( n31303 , n31298 , n31301 , n31302 );
and ( n31304 , n31293 , n31303 );
and ( n31305 , n31291 , n31303 );
or ( n31306 , n31294 , n31304 , n31305 );
and ( n31307 , n31289 , n31306 );
and ( n31308 , n31287 , n31306 );
or ( n31309 , n31290 , n31307 , n31308 );
and ( n31310 , n31285 , n31309 );
and ( n31311 , n31283 , n31309 );
or ( n31312 , n31286 , n31310 , n31311 );
and ( n31313 , n31281 , n31312 );
and ( n31314 , n31279 , n31312 );
or ( n31315 , n31282 , n31313 , n31314 );
and ( n31316 , n31277 , n31315 );
and ( n31317 , n31275 , n31315 );
or ( n31318 , n31278 , n31316 , n31317 );
and ( n31319 , n31273 , n31318 );
and ( n31320 , n31271 , n31318 );
or ( n31321 , n31274 , n31319 , n31320 );
and ( n31322 , n31269 , n31321 );
and ( n31323 , n31267 , n31321 );
or ( n31324 , n31270 , n31322 , n31323 );
and ( n31325 , n31265 , n31324 );
and ( n31326 , n31263 , n31324 );
or ( n31327 , n31266 , n31325 , n31326 );
and ( n31328 , n31261 , n31327 );
and ( n31329 , n31259 , n31327 );
or ( n31330 , n31262 , n31328 , n31329 );
and ( n31331 , n31257 , n31330 );
and ( n31332 , n31255 , n31330 );
or ( n31333 , n31258 , n31331 , n31332 );
and ( n31334 , n31253 , n31333 );
and ( n31335 , n31251 , n31333 );
or ( n31336 , n31254 , n31334 , n31335 );
and ( n31337 , n31249 , n31336 );
and ( n31338 , n31247 , n31336 );
or ( n31339 , n31250 , n31337 , n31338 );
and ( n31340 , n31245 , n31339 );
and ( n31341 , n31243 , n31339 );
or ( n31342 , n31246 , n31340 , n31341 );
and ( n31343 , n31241 , n31342 );
and ( n31344 , n31239 , n31342 );
or ( n31345 , n31242 , n31343 , n31344 );
and ( n31346 , n31237 , n31345 );
and ( n31347 , n31235 , n31345 );
or ( n31348 , n31238 , n31346 , n31347 );
and ( n31349 , n31233 , n31348 );
and ( n31350 , n31231 , n31348 );
or ( n31351 , n31234 , n31349 , n31350 );
and ( n31352 , n31229 , n31351 );
and ( n31353 , n31227 , n31351 );
or ( n31354 , n31230 , n31352 , n31353 );
and ( n31355 , n31225 , n31354 );
and ( n31356 , n31223 , n31354 );
or ( n31357 , n31226 , n31355 , n31356 );
and ( n31358 , n31222 , n31357 );
and ( n31359 , n31220 , n31358 );
and ( n31360 , n31218 , n31359 );
and ( n31361 , n31216 , n31360 );
and ( n31362 , n31214 , n31361 );
and ( n31363 , n31212 , n31362 );
and ( n31364 , n31210 , n31363 );
and ( n31365 , n31208 , n31364 );
and ( n31366 , n31206 , n31365 );
and ( n31367 , n31204 , n31366 );
and ( n31368 , n31202 , n31367 );
xor ( n31369 , n31200 , n31368 );
buf ( n31370 , n31369 );
buf ( n31371 , n31370 );
not ( n31372 , n31371 );
xor ( n31373 , n31295 , n31297 );
xor ( n31374 , n31373 , n31300 );
buf ( n31375 , n31374 );
buf ( n31376 , n31375 );
and ( n31377 , n31372 , n31376 );
not ( n31378 , n31376 );
not ( n31379 , n31193 );
xor ( n31380 , n31378 , n31379 );
and ( n31381 , n31380 , n31371 );
or ( n31382 , n31377 , n31381 );
buf ( n31383 , n31382 );
not ( n31384 , n31383 );
buf ( n31385 , n31384 );
buf ( n31386 , n31385 );
not ( n31387 , n31386 );
or ( n31388 , n31198 , n31387 );
not ( n31389 , n31371 );
xor ( n31390 , n31291 , n31293 );
xor ( n31391 , n31390 , n31303 );
buf ( n31392 , n31391 );
buf ( n31393 , n31392 );
and ( n31394 , n31389 , n31393 );
not ( n31395 , n31393 );
and ( n31396 , n31378 , n31379 );
xor ( n31397 , n31395 , n31396 );
and ( n31398 , n31397 , n31371 );
or ( n31399 , n31394 , n31398 );
buf ( n31400 , n31399 );
not ( n31401 , n31400 );
buf ( n31402 , n31401 );
buf ( n31403 , n31402 );
not ( n31404 , n31403 );
or ( n31405 , n31388 , n31404 );
not ( n31406 , n31371 );
xor ( n31407 , n31287 , n31289 );
xor ( n31408 , n31407 , n31306 );
buf ( n31409 , n31408 );
buf ( n31410 , n31409 );
and ( n31411 , n31406 , n31410 );
not ( n31412 , n31410 );
and ( n31413 , n31395 , n31396 );
xor ( n31414 , n31412 , n31413 );
and ( n31415 , n31414 , n31371 );
or ( n31416 , n31411 , n31415 );
buf ( n31417 , n31416 );
not ( n31418 , n31417 );
buf ( n31419 , n31418 );
buf ( n31420 , n31419 );
not ( n31421 , n31420 );
or ( n31422 , n31405 , n31421 );
not ( n31423 , n31371 );
xor ( n31424 , n31283 , n31285 );
xor ( n31425 , n31424 , n31309 );
buf ( n31426 , n31425 );
buf ( n31427 , n31426 );
and ( n31428 , n31423 , n31427 );
not ( n31429 , n31427 );
and ( n31430 , n31412 , n31413 );
xor ( n31431 , n31429 , n31430 );
and ( n31432 , n31431 , n31371 );
or ( n31433 , n31428 , n31432 );
buf ( n31434 , n31433 );
not ( n31435 , n31434 );
buf ( n31436 , n31435 );
buf ( n31437 , n31436 );
not ( n31438 , n31437 );
or ( n31439 , n31422 , n31438 );
not ( n31440 , n31371 );
xor ( n31441 , n31279 , n31281 );
xor ( n31442 , n31441 , n31312 );
buf ( n31443 , n31442 );
buf ( n31444 , n31443 );
and ( n31445 , n31440 , n31444 );
not ( n31446 , n31444 );
and ( n31447 , n31429 , n31430 );
xor ( n31448 , n31446 , n31447 );
and ( n31449 , n31448 , n31371 );
or ( n31450 , n31445 , n31449 );
buf ( n31451 , n31450 );
not ( n31452 , n31451 );
buf ( n31453 , n31452 );
buf ( n31454 , n31453 );
not ( n31455 , n31454 );
or ( n31456 , n31439 , n31455 );
not ( n31457 , n31371 );
xor ( n31458 , n31275 , n31277 );
xor ( n31459 , n31458 , n31315 );
buf ( n31460 , n31459 );
buf ( n31461 , n31460 );
and ( n31462 , n31457 , n31461 );
not ( n31463 , n31461 );
and ( n31464 , n31446 , n31447 );
xor ( n31465 , n31463 , n31464 );
and ( n31466 , n31465 , n31371 );
or ( n31467 , n31462 , n31466 );
buf ( n31468 , n31467 );
not ( n31469 , n31468 );
buf ( n31470 , n31469 );
buf ( n31471 , n31470 );
not ( n31472 , n31471 );
or ( n31473 , n31456 , n31472 );
not ( n31474 , n31371 );
xor ( n31475 , n31271 , n31273 );
xor ( n31476 , n31475 , n31318 );
buf ( n31477 , n31476 );
buf ( n31478 , n31477 );
and ( n31479 , n31474 , n31478 );
not ( n31480 , n31478 );
and ( n31481 , n31463 , n31464 );
xor ( n31482 , n31480 , n31481 );
and ( n31483 , n31482 , n31371 );
or ( n31484 , n31479 , n31483 );
buf ( n31485 , n31484 );
not ( n31486 , n31485 );
buf ( n31487 , n31486 );
buf ( n31488 , n31487 );
not ( n31489 , n31488 );
or ( n31490 , n31473 , n31489 );
not ( n31491 , n31371 );
xor ( n31492 , n31267 , n31269 );
xor ( n31493 , n31492 , n31321 );
buf ( n31494 , n31493 );
buf ( n31495 , n31494 );
and ( n31496 , n31491 , n31495 );
not ( n31497 , n31495 );
and ( n31498 , n31480 , n31481 );
xor ( n31499 , n31497 , n31498 );
and ( n31500 , n31499 , n31371 );
or ( n31501 , n31496 , n31500 );
buf ( n31502 , n31501 );
not ( n31503 , n31502 );
buf ( n31504 , n31503 );
buf ( n31505 , n31504 );
not ( n31506 , n31505 );
or ( n31507 , n31490 , n31506 );
not ( n31508 , n31371 );
xor ( n31509 , n31263 , n31265 );
xor ( n31510 , n31509 , n31324 );
buf ( n31511 , n31510 );
buf ( n31512 , n31511 );
and ( n31513 , n31508 , n31512 );
not ( n31514 , n31512 );
and ( n31515 , n31497 , n31498 );
xor ( n31516 , n31514 , n31515 );
and ( n31517 , n31516 , n31371 );
or ( n31518 , n31513 , n31517 );
buf ( n31519 , n31518 );
not ( n31520 , n31519 );
buf ( n31521 , n31520 );
buf ( n31522 , n31521 );
not ( n31523 , n31522 );
or ( n31524 , n31507 , n31523 );
not ( n31525 , n31371 );
xor ( n31526 , n31259 , n31261 );
xor ( n31527 , n31526 , n31327 );
buf ( n31528 , n31527 );
buf ( n31529 , n31528 );
and ( n31530 , n31525 , n31529 );
not ( n31531 , n31529 );
and ( n31532 , n31514 , n31515 );
xor ( n31533 , n31531 , n31532 );
and ( n31534 , n31533 , n31371 );
or ( n31535 , n31530 , n31534 );
buf ( n31536 , n31535 );
not ( n31537 , n31536 );
buf ( n31538 , n31537 );
buf ( n31539 , n31538 );
not ( n31540 , n31539 );
or ( n31541 , n31524 , n31540 );
not ( n31542 , n31371 );
xor ( n31543 , n31255 , n31257 );
xor ( n31544 , n31543 , n31330 );
buf ( n31545 , n31544 );
buf ( n31546 , n31545 );
and ( n31547 , n31542 , n31546 );
not ( n31548 , n31546 );
and ( n31549 , n31531 , n31532 );
xor ( n31550 , n31548 , n31549 );
and ( n31551 , n31550 , n31371 );
or ( n31552 , n31547 , n31551 );
buf ( n31553 , n31552 );
not ( n31554 , n31553 );
buf ( n31555 , n31554 );
buf ( n31556 , n31555 );
not ( n31557 , n31556 );
or ( n31558 , n31541 , n31557 );
not ( n31559 , n31371 );
xor ( n31560 , n31251 , n31253 );
xor ( n31561 , n31560 , n31333 );
buf ( n31562 , n31561 );
buf ( n31563 , n31562 );
and ( n31564 , n31559 , n31563 );
not ( n31565 , n31563 );
and ( n31566 , n31548 , n31549 );
xor ( n31567 , n31565 , n31566 );
and ( n31568 , n31567 , n31371 );
or ( n31569 , n31564 , n31568 );
buf ( n31570 , n31569 );
not ( n31571 , n31570 );
buf ( n31572 , n31571 );
buf ( n31573 , n31572 );
not ( n31574 , n31573 );
or ( n31575 , n31558 , n31574 );
not ( n31576 , n31371 );
xor ( n31577 , n31247 , n31249 );
xor ( n31578 , n31577 , n31336 );
buf ( n31579 , n31578 );
buf ( n31580 , n31579 );
and ( n31581 , n31576 , n31580 );
not ( n31582 , n31580 );
and ( n31583 , n31565 , n31566 );
xor ( n31584 , n31582 , n31583 );
and ( n31585 , n31584 , n31371 );
or ( n31586 , n31581 , n31585 );
buf ( n31587 , n31586 );
not ( n31588 , n31587 );
buf ( n31589 , n31588 );
buf ( n31590 , n31589 );
not ( n31591 , n31590 );
or ( n31592 , n31575 , n31591 );
not ( n31593 , n31371 );
xor ( n31594 , n31243 , n31245 );
xor ( n31595 , n31594 , n31339 );
buf ( n31596 , n31595 );
buf ( n31597 , n31596 );
and ( n31598 , n31593 , n31597 );
not ( n31599 , n31597 );
and ( n31600 , n31582 , n31583 );
xor ( n31601 , n31599 , n31600 );
and ( n31602 , n31601 , n31371 );
or ( n31603 , n31598 , n31602 );
buf ( n31604 , n31603 );
not ( n31605 , n31604 );
buf ( n31606 , n31605 );
buf ( n31607 , n31606 );
not ( n31608 , n31607 );
or ( n31609 , n31592 , n31608 );
not ( n31610 , n31371 );
xor ( n31611 , n31239 , n31241 );
xor ( n31612 , n31611 , n31342 );
buf ( n31613 , n31612 );
buf ( n31614 , n31613 );
and ( n31615 , n31610 , n31614 );
not ( n31616 , n31614 );
and ( n31617 , n31599 , n31600 );
xor ( n31618 , n31616 , n31617 );
and ( n31619 , n31618 , n31371 );
or ( n31620 , n31615 , n31619 );
buf ( n31621 , n31620 );
not ( n31622 , n31621 );
buf ( n31623 , n31622 );
buf ( n31624 , n31623 );
not ( n31625 , n31624 );
or ( n31626 , n31609 , n31625 );
not ( n31627 , n31371 );
xor ( n31628 , n31235 , n31237 );
xor ( n31629 , n31628 , n31345 );
buf ( n31630 , n31629 );
buf ( n31631 , n31630 );
and ( n31632 , n31627 , n31631 );
not ( n31633 , n31631 );
and ( n31634 , n31616 , n31617 );
xor ( n31635 , n31633 , n31634 );
and ( n31636 , n31635 , n31371 );
or ( n31637 , n31632 , n31636 );
buf ( n31638 , n31637 );
not ( n31639 , n31638 );
buf ( n31640 , n31639 );
buf ( n31641 , n31640 );
not ( n31642 , n31641 );
or ( n31643 , n31626 , n31642 );
not ( n31644 , n31371 );
xor ( n31645 , n31231 , n31233 );
xor ( n31646 , n31645 , n31348 );
buf ( n31647 , n31646 );
buf ( n31648 , n31647 );
and ( n31649 , n31644 , n31648 );
not ( n31650 , n31648 );
and ( n31651 , n31633 , n31634 );
xor ( n31652 , n31650 , n31651 );
and ( n31653 , n31652 , n31371 );
or ( n31654 , n31649 , n31653 );
buf ( n31655 , n31654 );
not ( n31656 , n31655 );
buf ( n31657 , n31656 );
buf ( n31658 , n31657 );
not ( n31659 , n31658 );
or ( n31660 , n31643 , n31659 );
not ( n31661 , n31371 );
xor ( n31662 , n31227 , n31229 );
xor ( n31663 , n31662 , n31351 );
buf ( n31664 , n31663 );
buf ( n31665 , n31664 );
and ( n31666 , n31661 , n31665 );
not ( n31667 , n31665 );
and ( n31668 , n31650 , n31651 );
xor ( n31669 , n31667 , n31668 );
and ( n31670 , n31669 , n31371 );
or ( n31671 , n31666 , n31670 );
buf ( n31672 , n31671 );
not ( n31673 , n31672 );
buf ( n31674 , n31673 );
buf ( n31675 , n31674 );
not ( n31676 , n31675 );
or ( n31677 , n31660 , n31676 );
not ( n31678 , n31371 );
xor ( n31679 , n31223 , n31225 );
xor ( n31680 , n31679 , n31354 );
buf ( n31681 , n31680 );
buf ( n31682 , n31681 );
and ( n31683 , n31678 , n31682 );
not ( n31684 , n31682 );
and ( n31685 , n31667 , n31668 );
xor ( n31686 , n31684 , n31685 );
and ( n31687 , n31686 , n31371 );
or ( n31688 , n31683 , n31687 );
buf ( n31689 , n31688 );
not ( n31690 , n31689 );
buf ( n31691 , n31690 );
buf ( n31692 , n31691 );
not ( n31693 , n31692 );
or ( n31694 , n31677 , n31693 );
buf ( n31695 , n31694 );
buf ( n31696 , n31695 );
and ( n31697 , n31696 , n31371 );
not ( n31698 , n31697 );
and ( n31699 , n31698 , n31198 );
xor ( n31700 , n31198 , n31371 );
xor ( n31701 , n31700 , n31371 );
and ( n31702 , n31701 , n31697 );
or ( n31703 , n31699 , n31702 );
buf ( n31704 , n31703 );
and ( n31705 , n31704 , n14140 );
buf ( n31706 , n15864 );
buf ( n31707 , n13510 );
xor ( n31708 , n31706 , n31707 );
buf ( n31709 , n31708 );
buf ( n31710 , n31709 );
buf ( n31711 , n31710 );
not ( n31712 , n31711 );
buf ( n31713 , n31712 );
buf ( n31714 , n31713 );
not ( n31715 , n31714 );
buf ( n31716 , n13144 );
not ( n31717 , n31716 );
buf ( n31718 , n14607 );
not ( n31719 , n31718 );
buf ( n31720 , n14960 );
not ( n31721 , n31720 );
buf ( n31722 , n13158 );
not ( n31723 , n31722 );
buf ( n31724 , n13171 );
not ( n31725 , n31724 );
buf ( n31726 , n13183 );
not ( n31727 , n31726 );
buf ( n31728 , n13195 );
not ( n31729 , n31728 );
buf ( n31730 , n13207 );
not ( n31731 , n31730 );
buf ( n31732 , n13219 );
not ( n31733 , n31732 );
buf ( n31734 , n13231 );
not ( n31735 , n31734 );
buf ( n31736 , n13243 );
not ( n31737 , n31736 );
buf ( n31738 , n13255 );
not ( n31739 , n31738 );
buf ( n31740 , n15447 );
buf ( n31741 , n13267 );
not ( n31742 , n31741 );
and ( n31743 , n31740 , n31742 );
buf ( n31744 , n15469 );
buf ( n31745 , n13279 );
not ( n31746 , n31745 );
and ( n31747 , n31744 , n31746 );
buf ( n31748 , n15491 );
buf ( n31749 , n13291 );
not ( n31750 , n31749 );
and ( n31751 , n31748 , n31750 );
buf ( n31752 , n15513 );
buf ( n31753 , n13303 );
not ( n31754 , n31753 );
and ( n31755 , n31752 , n31754 );
buf ( n31756 , n15535 );
buf ( n31757 , n13315 );
not ( n31758 , n31757 );
and ( n31759 , n31756 , n31758 );
buf ( n31760 , n15557 );
buf ( n31761 , n13327 );
not ( n31762 , n31761 );
and ( n31763 , n31760 , n31762 );
buf ( n31764 , n15579 );
buf ( n31765 , n13339 );
not ( n31766 , n31765 );
and ( n31767 , n31764 , n31766 );
buf ( n31768 , n15601 );
buf ( n31769 , n13351 );
not ( n31770 , n31769 );
and ( n31771 , n31768 , n31770 );
buf ( n31772 , n15623 );
buf ( n31773 , n13363 );
not ( n31774 , n31773 );
and ( n31775 , n31772 , n31774 );
buf ( n31776 , n15645 );
buf ( n31777 , n13375 );
not ( n31778 , n31777 );
and ( n31779 , n31776 , n31778 );
buf ( n31780 , n15667 );
buf ( n31781 , n13387 );
not ( n31782 , n31781 );
and ( n31783 , n31780 , n31782 );
buf ( n31784 , n15689 );
buf ( n31785 , n13399 );
not ( n31786 , n31785 );
and ( n31787 , n31784 , n31786 );
buf ( n31788 , n15711 );
buf ( n31789 , n13411 );
not ( n31790 , n31789 );
and ( n31791 , n31788 , n31790 );
buf ( n31792 , n15733 );
buf ( n31793 , n13423 );
not ( n31794 , n31793 );
and ( n31795 , n31792 , n31794 );
buf ( n31796 , n15755 );
buf ( n31797 , n13435 );
not ( n31798 , n31797 );
and ( n31799 , n31796 , n31798 );
buf ( n31800 , n15777 );
buf ( n31801 , n13447 );
not ( n31802 , n31801 );
and ( n31803 , n31800 , n31802 );
buf ( n31804 , n15799 );
buf ( n31805 , n13459 );
not ( n31806 , n31805 );
and ( n31807 , n31804 , n31806 );
buf ( n31808 , n15821 );
buf ( n31809 , n13476 );
not ( n31810 , n31809 );
and ( n31811 , n31808 , n31810 );
buf ( n31812 , n15843 );
buf ( n31813 , n13493 );
not ( n31814 , n31813 );
and ( n31815 , n31812 , n31814 );
not ( n31816 , n31707 );
or ( n31817 , n31706 , n31816 );
and ( n31818 , n31814 , n31817 );
and ( n31819 , n31812 , n31817 );
or ( n31820 , n31815 , n31818 , n31819 );
and ( n31821 , n31810 , n31820 );
and ( n31822 , n31808 , n31820 );
or ( n31823 , n31811 , n31821 , n31822 );
and ( n31824 , n31806 , n31823 );
and ( n31825 , n31804 , n31823 );
or ( n31826 , n31807 , n31824 , n31825 );
and ( n31827 , n31802 , n31826 );
and ( n31828 , n31800 , n31826 );
or ( n31829 , n31803 , n31827 , n31828 );
and ( n31830 , n31798 , n31829 );
and ( n31831 , n31796 , n31829 );
or ( n31832 , n31799 , n31830 , n31831 );
and ( n31833 , n31794 , n31832 );
and ( n31834 , n31792 , n31832 );
or ( n31835 , n31795 , n31833 , n31834 );
and ( n31836 , n31790 , n31835 );
and ( n31837 , n31788 , n31835 );
or ( n31838 , n31791 , n31836 , n31837 );
and ( n31839 , n31786 , n31838 );
and ( n31840 , n31784 , n31838 );
or ( n31841 , n31787 , n31839 , n31840 );
and ( n31842 , n31782 , n31841 );
and ( n31843 , n31780 , n31841 );
or ( n31844 , n31783 , n31842 , n31843 );
and ( n31845 , n31778 , n31844 );
and ( n31846 , n31776 , n31844 );
or ( n31847 , n31779 , n31845 , n31846 );
and ( n31848 , n31774 , n31847 );
and ( n31849 , n31772 , n31847 );
or ( n31850 , n31775 , n31848 , n31849 );
and ( n31851 , n31770 , n31850 );
and ( n31852 , n31768 , n31850 );
or ( n31853 , n31771 , n31851 , n31852 );
and ( n31854 , n31766 , n31853 );
and ( n31855 , n31764 , n31853 );
or ( n31856 , n31767 , n31854 , n31855 );
and ( n31857 , n31762 , n31856 );
and ( n31858 , n31760 , n31856 );
or ( n31859 , n31763 , n31857 , n31858 );
and ( n31860 , n31758 , n31859 );
and ( n31861 , n31756 , n31859 );
or ( n31862 , n31759 , n31860 , n31861 );
and ( n31863 , n31754 , n31862 );
and ( n31864 , n31752 , n31862 );
or ( n31865 , n31755 , n31863 , n31864 );
and ( n31866 , n31750 , n31865 );
and ( n31867 , n31748 , n31865 );
or ( n31868 , n31751 , n31866 , n31867 );
and ( n31869 , n31746 , n31868 );
and ( n31870 , n31744 , n31868 );
or ( n31871 , n31747 , n31869 , n31870 );
and ( n31872 , n31742 , n31871 );
and ( n31873 , n31740 , n31871 );
or ( n31874 , n31743 , n31872 , n31873 );
and ( n31875 , n31739 , n31874 );
and ( n31876 , n31737 , n31875 );
and ( n31877 , n31735 , n31876 );
and ( n31878 , n31733 , n31877 );
and ( n31879 , n31731 , n31878 );
and ( n31880 , n31729 , n31879 );
and ( n31881 , n31727 , n31880 );
and ( n31882 , n31725 , n31881 );
and ( n31883 , n31723 , n31882 );
and ( n31884 , n31721 , n31883 );
and ( n31885 , n31719 , n31884 );
xor ( n31886 , n31717 , n31885 );
buf ( n31887 , n31886 );
buf ( n31888 , n31887 );
not ( n31889 , n31888 );
xor ( n31890 , n31812 , n31814 );
xor ( n31891 , n31890 , n31817 );
buf ( n31892 , n31891 );
buf ( n31893 , n31892 );
and ( n31894 , n31889 , n31893 );
not ( n31895 , n31893 );
not ( n31896 , n31710 );
xor ( n31897 , n31895 , n31896 );
and ( n31898 , n31897 , n31888 );
or ( n31899 , n31894 , n31898 );
buf ( n31900 , n31899 );
not ( n31901 , n31900 );
buf ( n31902 , n31901 );
buf ( n31903 , n31902 );
not ( n31904 , n31903 );
or ( n31905 , n31715 , n31904 );
not ( n31906 , n31888 );
xor ( n31907 , n31808 , n31810 );
xor ( n31908 , n31907 , n31820 );
buf ( n31909 , n31908 );
buf ( n31910 , n31909 );
and ( n31911 , n31906 , n31910 );
not ( n31912 , n31910 );
and ( n31913 , n31895 , n31896 );
xor ( n31914 , n31912 , n31913 );
and ( n31915 , n31914 , n31888 );
or ( n31916 , n31911 , n31915 );
buf ( n31917 , n31916 );
not ( n31918 , n31917 );
buf ( n31919 , n31918 );
buf ( n31920 , n31919 );
not ( n31921 , n31920 );
or ( n31922 , n31905 , n31921 );
not ( n31923 , n31888 );
xor ( n31924 , n31804 , n31806 );
xor ( n31925 , n31924 , n31823 );
buf ( n31926 , n31925 );
buf ( n31927 , n31926 );
and ( n31928 , n31923 , n31927 );
not ( n31929 , n31927 );
and ( n31930 , n31912 , n31913 );
xor ( n31931 , n31929 , n31930 );
and ( n31932 , n31931 , n31888 );
or ( n31933 , n31928 , n31932 );
buf ( n31934 , n31933 );
not ( n31935 , n31934 );
buf ( n31936 , n31935 );
buf ( n31937 , n31936 );
not ( n31938 , n31937 );
or ( n31939 , n31922 , n31938 );
not ( n31940 , n31888 );
xor ( n31941 , n31800 , n31802 );
xor ( n31942 , n31941 , n31826 );
buf ( n31943 , n31942 );
buf ( n31944 , n31943 );
and ( n31945 , n31940 , n31944 );
not ( n31946 , n31944 );
and ( n31947 , n31929 , n31930 );
xor ( n31948 , n31946 , n31947 );
and ( n31949 , n31948 , n31888 );
or ( n31950 , n31945 , n31949 );
buf ( n31951 , n31950 );
not ( n31952 , n31951 );
buf ( n31953 , n31952 );
buf ( n31954 , n31953 );
not ( n31955 , n31954 );
or ( n31956 , n31939 , n31955 );
not ( n31957 , n31888 );
xor ( n31958 , n31796 , n31798 );
xor ( n31959 , n31958 , n31829 );
buf ( n31960 , n31959 );
buf ( n31961 , n31960 );
and ( n31962 , n31957 , n31961 );
not ( n31963 , n31961 );
and ( n31964 , n31946 , n31947 );
xor ( n31965 , n31963 , n31964 );
and ( n31966 , n31965 , n31888 );
or ( n31967 , n31962 , n31966 );
buf ( n31968 , n31967 );
not ( n31969 , n31968 );
buf ( n31970 , n31969 );
buf ( n31971 , n31970 );
not ( n31972 , n31971 );
or ( n31973 , n31956 , n31972 );
not ( n31974 , n31888 );
xor ( n31975 , n31792 , n31794 );
xor ( n31976 , n31975 , n31832 );
buf ( n31977 , n31976 );
buf ( n31978 , n31977 );
and ( n31979 , n31974 , n31978 );
not ( n31980 , n31978 );
and ( n31981 , n31963 , n31964 );
xor ( n31982 , n31980 , n31981 );
and ( n31983 , n31982 , n31888 );
or ( n31984 , n31979 , n31983 );
buf ( n31985 , n31984 );
not ( n31986 , n31985 );
buf ( n31987 , n31986 );
buf ( n31988 , n31987 );
not ( n31989 , n31988 );
or ( n31990 , n31973 , n31989 );
not ( n31991 , n31888 );
xor ( n31992 , n31788 , n31790 );
xor ( n31993 , n31992 , n31835 );
buf ( n31994 , n31993 );
buf ( n31995 , n31994 );
and ( n31996 , n31991 , n31995 );
not ( n31997 , n31995 );
and ( n31998 , n31980 , n31981 );
xor ( n31999 , n31997 , n31998 );
and ( n32000 , n31999 , n31888 );
or ( n32001 , n31996 , n32000 );
buf ( n32002 , n32001 );
not ( n32003 , n32002 );
buf ( n32004 , n32003 );
buf ( n32005 , n32004 );
not ( n32006 , n32005 );
or ( n32007 , n31990 , n32006 );
not ( n32008 , n31888 );
xor ( n32009 , n31784 , n31786 );
xor ( n32010 , n32009 , n31838 );
buf ( n32011 , n32010 );
buf ( n32012 , n32011 );
and ( n32013 , n32008 , n32012 );
not ( n32014 , n32012 );
and ( n32015 , n31997 , n31998 );
xor ( n32016 , n32014 , n32015 );
and ( n32017 , n32016 , n31888 );
or ( n32018 , n32013 , n32017 );
buf ( n32019 , n32018 );
not ( n32020 , n32019 );
buf ( n32021 , n32020 );
buf ( n32022 , n32021 );
not ( n32023 , n32022 );
or ( n32024 , n32007 , n32023 );
not ( n32025 , n31888 );
xor ( n32026 , n31780 , n31782 );
xor ( n32027 , n32026 , n31841 );
buf ( n32028 , n32027 );
buf ( n32029 , n32028 );
and ( n32030 , n32025 , n32029 );
not ( n32031 , n32029 );
and ( n32032 , n32014 , n32015 );
xor ( n32033 , n32031 , n32032 );
and ( n32034 , n32033 , n31888 );
or ( n32035 , n32030 , n32034 );
buf ( n32036 , n32035 );
not ( n32037 , n32036 );
buf ( n32038 , n32037 );
buf ( n32039 , n32038 );
not ( n32040 , n32039 );
or ( n32041 , n32024 , n32040 );
not ( n32042 , n31888 );
xor ( n32043 , n31776 , n31778 );
xor ( n32044 , n32043 , n31844 );
buf ( n32045 , n32044 );
buf ( n32046 , n32045 );
and ( n32047 , n32042 , n32046 );
not ( n32048 , n32046 );
and ( n32049 , n32031 , n32032 );
xor ( n32050 , n32048 , n32049 );
and ( n32051 , n32050 , n31888 );
or ( n32052 , n32047 , n32051 );
buf ( n32053 , n32052 );
not ( n32054 , n32053 );
buf ( n32055 , n32054 );
buf ( n32056 , n32055 );
not ( n32057 , n32056 );
or ( n32058 , n32041 , n32057 );
not ( n32059 , n31888 );
xor ( n32060 , n31772 , n31774 );
xor ( n32061 , n32060 , n31847 );
buf ( n32062 , n32061 );
buf ( n32063 , n32062 );
and ( n32064 , n32059 , n32063 );
not ( n32065 , n32063 );
and ( n32066 , n32048 , n32049 );
xor ( n32067 , n32065 , n32066 );
and ( n32068 , n32067 , n31888 );
or ( n32069 , n32064 , n32068 );
buf ( n32070 , n32069 );
not ( n32071 , n32070 );
buf ( n32072 , n32071 );
buf ( n32073 , n32072 );
not ( n32074 , n32073 );
or ( n32075 , n32058 , n32074 );
not ( n32076 , n31888 );
xor ( n32077 , n31768 , n31770 );
xor ( n32078 , n32077 , n31850 );
buf ( n32079 , n32078 );
buf ( n32080 , n32079 );
and ( n32081 , n32076 , n32080 );
not ( n32082 , n32080 );
and ( n32083 , n32065 , n32066 );
xor ( n32084 , n32082 , n32083 );
and ( n32085 , n32084 , n31888 );
or ( n32086 , n32081 , n32085 );
buf ( n32087 , n32086 );
not ( n32088 , n32087 );
buf ( n32089 , n32088 );
buf ( n32090 , n32089 );
not ( n32091 , n32090 );
or ( n32092 , n32075 , n32091 );
not ( n32093 , n31888 );
xor ( n32094 , n31764 , n31766 );
xor ( n32095 , n32094 , n31853 );
buf ( n32096 , n32095 );
buf ( n32097 , n32096 );
and ( n32098 , n32093 , n32097 );
not ( n32099 , n32097 );
and ( n32100 , n32082 , n32083 );
xor ( n32101 , n32099 , n32100 );
and ( n32102 , n32101 , n31888 );
or ( n32103 , n32098 , n32102 );
buf ( n32104 , n32103 );
not ( n32105 , n32104 );
buf ( n32106 , n32105 );
buf ( n32107 , n32106 );
not ( n32108 , n32107 );
or ( n32109 , n32092 , n32108 );
not ( n32110 , n31888 );
xor ( n32111 , n31760 , n31762 );
xor ( n32112 , n32111 , n31856 );
buf ( n32113 , n32112 );
buf ( n32114 , n32113 );
and ( n32115 , n32110 , n32114 );
not ( n32116 , n32114 );
and ( n32117 , n32099 , n32100 );
xor ( n32118 , n32116 , n32117 );
and ( n32119 , n32118 , n31888 );
or ( n32120 , n32115 , n32119 );
buf ( n32121 , n32120 );
not ( n32122 , n32121 );
buf ( n32123 , n32122 );
buf ( n32124 , n32123 );
not ( n32125 , n32124 );
or ( n32126 , n32109 , n32125 );
not ( n32127 , n31888 );
xor ( n32128 , n31756 , n31758 );
xor ( n32129 , n32128 , n31859 );
buf ( n32130 , n32129 );
buf ( n32131 , n32130 );
and ( n32132 , n32127 , n32131 );
not ( n32133 , n32131 );
and ( n32134 , n32116 , n32117 );
xor ( n32135 , n32133 , n32134 );
and ( n32136 , n32135 , n31888 );
or ( n32137 , n32132 , n32136 );
buf ( n32138 , n32137 );
not ( n32139 , n32138 );
buf ( n32140 , n32139 );
buf ( n32141 , n32140 );
not ( n32142 , n32141 );
or ( n32143 , n32126 , n32142 );
not ( n32144 , n31888 );
xor ( n32145 , n31752 , n31754 );
xor ( n32146 , n32145 , n31862 );
buf ( n32147 , n32146 );
buf ( n32148 , n32147 );
and ( n32149 , n32144 , n32148 );
not ( n32150 , n32148 );
and ( n32151 , n32133 , n32134 );
xor ( n32152 , n32150 , n32151 );
and ( n32153 , n32152 , n31888 );
or ( n32154 , n32149 , n32153 );
buf ( n32155 , n32154 );
not ( n32156 , n32155 );
buf ( n32157 , n32156 );
buf ( n32158 , n32157 );
not ( n32159 , n32158 );
or ( n32160 , n32143 , n32159 );
not ( n32161 , n31888 );
xor ( n32162 , n31748 , n31750 );
xor ( n32163 , n32162 , n31865 );
buf ( n32164 , n32163 );
buf ( n32165 , n32164 );
and ( n32166 , n32161 , n32165 );
not ( n32167 , n32165 );
and ( n32168 , n32150 , n32151 );
xor ( n32169 , n32167 , n32168 );
and ( n32170 , n32169 , n31888 );
or ( n32171 , n32166 , n32170 );
buf ( n32172 , n32171 );
not ( n32173 , n32172 );
buf ( n32174 , n32173 );
buf ( n32175 , n32174 );
not ( n32176 , n32175 );
or ( n32177 , n32160 , n32176 );
not ( n32178 , n31888 );
xor ( n32179 , n31744 , n31746 );
xor ( n32180 , n32179 , n31868 );
buf ( n32181 , n32180 );
buf ( n32182 , n32181 );
and ( n32183 , n32178 , n32182 );
not ( n32184 , n32182 );
and ( n32185 , n32167 , n32168 );
xor ( n32186 , n32184 , n32185 );
and ( n32187 , n32186 , n31888 );
or ( n32188 , n32183 , n32187 );
buf ( n32189 , n32188 );
not ( n32190 , n32189 );
buf ( n32191 , n32190 );
buf ( n32192 , n32191 );
not ( n32193 , n32192 );
or ( n32194 , n32177 , n32193 );
not ( n32195 , n31888 );
xor ( n32196 , n31740 , n31742 );
xor ( n32197 , n32196 , n31871 );
buf ( n32198 , n32197 );
buf ( n32199 , n32198 );
and ( n32200 , n32195 , n32199 );
not ( n32201 , n32199 );
and ( n32202 , n32184 , n32185 );
xor ( n32203 , n32201 , n32202 );
and ( n32204 , n32203 , n31888 );
or ( n32205 , n32200 , n32204 );
buf ( n32206 , n32205 );
not ( n32207 , n32206 );
buf ( n32208 , n32207 );
buf ( n32209 , n32208 );
not ( n32210 , n32209 );
or ( n32211 , n32194 , n32210 );
buf ( n32212 , n32211 );
buf ( n32213 , n32212 );
and ( n32214 , n32213 , n31888 );
not ( n32215 , n32214 );
and ( n32216 , n32215 , n31715 );
xor ( n32217 , n31715 , n31888 );
xor ( n32218 , n32217 , n31888 );
and ( n32219 , n32218 , n32214 );
or ( n32220 , n32216 , n32219 );
buf ( n32221 , n32220 );
and ( n32222 , n32221 , n14137 );
and ( n32223 , n15864 , n14143 );
and ( n32224 , n10628 , n14141 );
or ( n32225 , n31705 , n32222 , n32223 , n32224 );
or ( n32226 , n14565 , n14564 );
or ( n32227 , n32226 , n14567 );
or ( n32228 , n32227 , n14569 );
or ( n32229 , n32228 , n14572 );
or ( n32230 , n32229 , n14574 );
or ( n32231 , n32230 , n14576 );
or ( n32232 , n32231 , n14578 );
or ( n32233 , n32232 , n14580 );
or ( n32234 , n32233 , n14582 );
or ( n32235 , n32234 , n14584 );
or ( n32236 , n32235 , n14586 );
and ( n32237 , n32225 , n32236 );
or ( n32238 , n31188 , n32237 );
and ( n32239 , n31186 , n32238 );
buf ( n32240 , n13508 );
buf ( n32241 , n32240 );
not ( n32242 , n32241 );
buf ( n32243 , n32242 );
buf ( n32244 , n32243 );
not ( n32245 , n32244 );
buf ( n32246 , n13140 );
not ( n32247 , n32246 );
buf ( n32248 , n13491 );
and ( n32249 , n32247 , n32248 );
not ( n32250 , n32248 );
not ( n32251 , n32240 );
xor ( n32252 , n32250 , n32251 );
and ( n32253 , n32252 , n32246 );
or ( n32254 , n32249 , n32253 );
buf ( n32255 , n32254 );
not ( n32256 , n32255 );
buf ( n32257 , n32256 );
buf ( n32258 , n32257 );
not ( n32259 , n32258 );
or ( n32260 , n32245 , n32259 );
not ( n32261 , n32246 );
buf ( n32262 , n13474 );
and ( n32263 , n32261 , n32262 );
not ( n32264 , n32262 );
and ( n32265 , n32250 , n32251 );
xor ( n32266 , n32264 , n32265 );
and ( n32267 , n32266 , n32246 );
or ( n32268 , n32263 , n32267 );
buf ( n32269 , n32268 );
not ( n32270 , n32269 );
buf ( n32271 , n32270 );
buf ( n32272 , n32271 );
not ( n32273 , n32272 );
or ( n32274 , n32260 , n32273 );
not ( n32275 , n32246 );
buf ( n32276 , n13457 );
and ( n32277 , n32275 , n32276 );
not ( n32278 , n32276 );
and ( n32279 , n32264 , n32265 );
xor ( n32280 , n32278 , n32279 );
and ( n32281 , n32280 , n32246 );
or ( n32282 , n32277 , n32281 );
buf ( n32283 , n32282 );
not ( n32284 , n32283 );
buf ( n32285 , n32284 );
buf ( n32286 , n32285 );
not ( n32287 , n32286 );
or ( n32288 , n32274 , n32287 );
not ( n32289 , n32246 );
buf ( n32290 , n13445 );
and ( n32291 , n32289 , n32290 );
not ( n32292 , n32290 );
and ( n32293 , n32278 , n32279 );
xor ( n32294 , n32292 , n32293 );
and ( n32295 , n32294 , n32246 );
or ( n32296 , n32291 , n32295 );
buf ( n32297 , n32296 );
not ( n32298 , n32297 );
buf ( n32299 , n32298 );
buf ( n32300 , n32299 );
not ( n32301 , n32300 );
or ( n32302 , n32288 , n32301 );
not ( n32303 , n32246 );
buf ( n32304 , n13433 );
and ( n32305 , n32303 , n32304 );
not ( n32306 , n32304 );
and ( n32307 , n32292 , n32293 );
xor ( n32308 , n32306 , n32307 );
and ( n32309 , n32308 , n32246 );
or ( n32310 , n32305 , n32309 );
buf ( n32311 , n32310 );
not ( n32312 , n32311 );
buf ( n32313 , n32312 );
buf ( n32314 , n32313 );
not ( n32315 , n32314 );
or ( n32316 , n32302 , n32315 );
not ( n32317 , n32246 );
buf ( n32318 , n13421 );
and ( n32319 , n32317 , n32318 );
not ( n32320 , n32318 );
and ( n32321 , n32306 , n32307 );
xor ( n32322 , n32320 , n32321 );
and ( n32323 , n32322 , n32246 );
or ( n32324 , n32319 , n32323 );
buf ( n32325 , n32324 );
not ( n32326 , n32325 );
buf ( n32327 , n32326 );
buf ( n32328 , n32327 );
not ( n32329 , n32328 );
or ( n32330 , n32316 , n32329 );
not ( n32331 , n32246 );
buf ( n32332 , n13409 );
and ( n32333 , n32331 , n32332 );
not ( n32334 , n32332 );
and ( n32335 , n32320 , n32321 );
xor ( n32336 , n32334 , n32335 );
and ( n32337 , n32336 , n32246 );
or ( n32338 , n32333 , n32337 );
buf ( n32339 , n32338 );
not ( n32340 , n32339 );
buf ( n32341 , n32340 );
buf ( n32342 , n32341 );
not ( n32343 , n32342 );
or ( n32344 , n32330 , n32343 );
not ( n32345 , n32246 );
buf ( n32346 , n13397 );
and ( n32347 , n32345 , n32346 );
not ( n32348 , n32346 );
and ( n32349 , n32334 , n32335 );
xor ( n32350 , n32348 , n32349 );
and ( n32351 , n32350 , n32246 );
or ( n32352 , n32347 , n32351 );
buf ( n32353 , n32352 );
not ( n32354 , n32353 );
buf ( n32355 , n32354 );
buf ( n32356 , n32355 );
not ( n32357 , n32356 );
or ( n32358 , n32344 , n32357 );
not ( n32359 , n32246 );
buf ( n32360 , n13385 );
and ( n32361 , n32359 , n32360 );
not ( n32362 , n32360 );
and ( n32363 , n32348 , n32349 );
xor ( n32364 , n32362 , n32363 );
and ( n32365 , n32364 , n32246 );
or ( n32366 , n32361 , n32365 );
buf ( n32367 , n32366 );
not ( n32368 , n32367 );
buf ( n32369 , n32368 );
buf ( n32370 , n32369 );
not ( n32371 , n32370 );
or ( n32372 , n32358 , n32371 );
not ( n32373 , n32246 );
buf ( n32374 , n13373 );
and ( n32375 , n32373 , n32374 );
not ( n32376 , n32374 );
and ( n32377 , n32362 , n32363 );
xor ( n32378 , n32376 , n32377 );
and ( n32379 , n32378 , n32246 );
or ( n32380 , n32375 , n32379 );
buf ( n32381 , n32380 );
not ( n32382 , n32381 );
buf ( n32383 , n32382 );
buf ( n32384 , n32383 );
not ( n32385 , n32384 );
or ( n32386 , n32372 , n32385 );
not ( n32387 , n32246 );
buf ( n32388 , n13361 );
and ( n32389 , n32387 , n32388 );
not ( n32390 , n32388 );
and ( n32391 , n32376 , n32377 );
xor ( n32392 , n32390 , n32391 );
and ( n32393 , n32392 , n32246 );
or ( n32394 , n32389 , n32393 );
buf ( n32395 , n32394 );
not ( n32396 , n32395 );
buf ( n32397 , n32396 );
buf ( n32398 , n32397 );
not ( n32399 , n32398 );
or ( n32400 , n32386 , n32399 );
not ( n32401 , n32246 );
buf ( n32402 , n13349 );
and ( n32403 , n32401 , n32402 );
not ( n32404 , n32402 );
and ( n32405 , n32390 , n32391 );
xor ( n32406 , n32404 , n32405 );
and ( n32407 , n32406 , n32246 );
or ( n32408 , n32403 , n32407 );
buf ( n32409 , n32408 );
not ( n32410 , n32409 );
buf ( n32411 , n32410 );
buf ( n32412 , n32411 );
not ( n32413 , n32412 );
or ( n32414 , n32400 , n32413 );
not ( n32415 , n32246 );
buf ( n32416 , n13337 );
and ( n32417 , n32415 , n32416 );
not ( n32418 , n32416 );
and ( n32419 , n32404 , n32405 );
xor ( n32420 , n32418 , n32419 );
and ( n32421 , n32420 , n32246 );
or ( n32422 , n32417 , n32421 );
buf ( n32423 , n32422 );
not ( n32424 , n32423 );
buf ( n32425 , n32424 );
buf ( n32426 , n32425 );
not ( n32427 , n32426 );
or ( n32428 , n32414 , n32427 );
not ( n32429 , n32246 );
buf ( n32430 , n13325 );
and ( n32431 , n32429 , n32430 );
not ( n32432 , n32430 );
and ( n32433 , n32418 , n32419 );
xor ( n32434 , n32432 , n32433 );
and ( n32435 , n32434 , n32246 );
or ( n32436 , n32431 , n32435 );
buf ( n32437 , n32436 );
not ( n32438 , n32437 );
buf ( n32439 , n32438 );
buf ( n32440 , n32439 );
not ( n32441 , n32440 );
or ( n32442 , n32428 , n32441 );
not ( n32443 , n32246 );
buf ( n32444 , n13313 );
and ( n32445 , n32443 , n32444 );
not ( n32446 , n32444 );
and ( n32447 , n32432 , n32433 );
xor ( n32448 , n32446 , n32447 );
and ( n32449 , n32448 , n32246 );
or ( n32450 , n32445 , n32449 );
buf ( n32451 , n32450 );
not ( n32452 , n32451 );
buf ( n32453 , n32452 );
buf ( n32454 , n32453 );
not ( n32455 , n32454 );
or ( n32456 , n32442 , n32455 );
not ( n32457 , n32246 );
buf ( n32458 , n13301 );
and ( n32459 , n32457 , n32458 );
not ( n32460 , n32458 );
and ( n32461 , n32446 , n32447 );
xor ( n32462 , n32460 , n32461 );
and ( n32463 , n32462 , n32246 );
or ( n32464 , n32459 , n32463 );
buf ( n32465 , n32464 );
not ( n32466 , n32465 );
buf ( n32467 , n32466 );
buf ( n32468 , n32467 );
not ( n32469 , n32468 );
or ( n32470 , n32456 , n32469 );
not ( n32471 , n32246 );
buf ( n32472 , n13289 );
and ( n32473 , n32471 , n32472 );
not ( n32474 , n32472 );
and ( n32475 , n32460 , n32461 );
xor ( n32476 , n32474 , n32475 );
and ( n32477 , n32476 , n32246 );
or ( n32478 , n32473 , n32477 );
buf ( n32479 , n32478 );
not ( n32480 , n32479 );
buf ( n32481 , n32480 );
buf ( n32482 , n32481 );
not ( n32483 , n32482 );
or ( n32484 , n32470 , n32483 );
not ( n32485 , n32246 );
buf ( n32486 , n13277 );
and ( n32487 , n32485 , n32486 );
not ( n32488 , n32486 );
and ( n32489 , n32474 , n32475 );
xor ( n32490 , n32488 , n32489 );
and ( n32491 , n32490 , n32246 );
or ( n32492 , n32487 , n32491 );
buf ( n32493 , n32492 );
not ( n32494 , n32493 );
buf ( n32495 , n32494 );
buf ( n32496 , n32495 );
not ( n32497 , n32496 );
or ( n32498 , n32484 , n32497 );
not ( n32499 , n32246 );
buf ( n32500 , n13265 );
and ( n32501 , n32499 , n32500 );
not ( n32502 , n32500 );
and ( n32503 , n32488 , n32489 );
xor ( n32504 , n32502 , n32503 );
and ( n32505 , n32504 , n32246 );
or ( n32506 , n32501 , n32505 );
buf ( n32507 , n32506 );
not ( n32508 , n32507 );
buf ( n32509 , n32508 );
buf ( n32510 , n32509 );
not ( n32511 , n32510 );
or ( n32512 , n32498 , n32511 );
buf ( n32513 , n32512 );
buf ( n32514 , n32513 );
and ( n32515 , n32514 , n32246 );
not ( n32516 , n32515 );
and ( n32517 , n32516 , n32245 );
xor ( n32518 , n32245 , n32246 );
xor ( n32519 , n32518 , n32246 );
and ( n32520 , n32519 , n32515 );
or ( n32521 , n32517 , n32520 );
buf ( n32522 , n32521 );
buf ( n32523 , n32522 );
buf ( n32524 , n15864 );
not ( n32525 , n32524 );
buf ( n32526 , n32525 );
not ( n32527 , n32526 );
buf ( n32528 , n32527 );
buf ( n32529 , n32528 );
buf ( n32530 , n32529 );
xor ( n32531 , n32523 , n32530 );
buf ( n32532 , n32531 );
and ( n32533 , n32532 , n14143 );
buf ( n32534 , n13510 );
buf ( n32535 , n32534 );
not ( n32536 , n32535 );
buf ( n32537 , n32536 );
buf ( n32538 , n32537 );
not ( n32539 , n32538 );
buf ( n32540 , n13144 );
not ( n32541 , n32540 );
buf ( n32542 , n13493 );
and ( n32543 , n32541 , n32542 );
not ( n32544 , n32542 );
not ( n32545 , n32534 );
xor ( n32546 , n32544 , n32545 );
and ( n32547 , n32546 , n32540 );
or ( n32548 , n32543 , n32547 );
buf ( n32549 , n32548 );
not ( n32550 , n32549 );
buf ( n32551 , n32550 );
buf ( n32552 , n32551 );
not ( n32553 , n32552 );
or ( n32554 , n32539 , n32553 );
not ( n32555 , n32540 );
buf ( n32556 , n13476 );
and ( n32557 , n32555 , n32556 );
not ( n32558 , n32556 );
and ( n32559 , n32544 , n32545 );
xor ( n32560 , n32558 , n32559 );
and ( n32561 , n32560 , n32540 );
or ( n32562 , n32557 , n32561 );
buf ( n32563 , n32562 );
not ( n32564 , n32563 );
buf ( n32565 , n32564 );
buf ( n32566 , n32565 );
not ( n32567 , n32566 );
or ( n32568 , n32554 , n32567 );
not ( n32569 , n32540 );
buf ( n32570 , n13459 );
and ( n32571 , n32569 , n32570 );
not ( n32572 , n32570 );
and ( n32573 , n32558 , n32559 );
xor ( n32574 , n32572 , n32573 );
and ( n32575 , n32574 , n32540 );
or ( n32576 , n32571 , n32575 );
buf ( n32577 , n32576 );
not ( n32578 , n32577 );
buf ( n32579 , n32578 );
buf ( n32580 , n32579 );
not ( n32581 , n32580 );
or ( n32582 , n32568 , n32581 );
not ( n32583 , n32540 );
buf ( n32584 , n13447 );
and ( n32585 , n32583 , n32584 );
not ( n32586 , n32584 );
and ( n32587 , n32572 , n32573 );
xor ( n32588 , n32586 , n32587 );
and ( n32589 , n32588 , n32540 );
or ( n32590 , n32585 , n32589 );
buf ( n32591 , n32590 );
not ( n32592 , n32591 );
buf ( n32593 , n32592 );
buf ( n32594 , n32593 );
not ( n32595 , n32594 );
or ( n32596 , n32582 , n32595 );
not ( n32597 , n32540 );
buf ( n32598 , n13435 );
and ( n32599 , n32597 , n32598 );
not ( n32600 , n32598 );
and ( n32601 , n32586 , n32587 );
xor ( n32602 , n32600 , n32601 );
and ( n32603 , n32602 , n32540 );
or ( n32604 , n32599 , n32603 );
buf ( n32605 , n32604 );
not ( n32606 , n32605 );
buf ( n32607 , n32606 );
buf ( n32608 , n32607 );
not ( n32609 , n32608 );
or ( n32610 , n32596 , n32609 );
not ( n32611 , n32540 );
buf ( n32612 , n13423 );
and ( n32613 , n32611 , n32612 );
not ( n32614 , n32612 );
and ( n32615 , n32600 , n32601 );
xor ( n32616 , n32614 , n32615 );
and ( n32617 , n32616 , n32540 );
or ( n32618 , n32613 , n32617 );
buf ( n32619 , n32618 );
not ( n32620 , n32619 );
buf ( n32621 , n32620 );
buf ( n32622 , n32621 );
not ( n32623 , n32622 );
or ( n32624 , n32610 , n32623 );
not ( n32625 , n32540 );
buf ( n32626 , n13411 );
and ( n32627 , n32625 , n32626 );
not ( n32628 , n32626 );
and ( n32629 , n32614 , n32615 );
xor ( n32630 , n32628 , n32629 );
and ( n32631 , n32630 , n32540 );
or ( n32632 , n32627 , n32631 );
buf ( n32633 , n32632 );
not ( n32634 , n32633 );
buf ( n32635 , n32634 );
buf ( n32636 , n32635 );
not ( n32637 , n32636 );
or ( n32638 , n32624 , n32637 );
not ( n32639 , n32540 );
buf ( n32640 , n13399 );
and ( n32641 , n32639 , n32640 );
not ( n32642 , n32640 );
and ( n32643 , n32628 , n32629 );
xor ( n32644 , n32642 , n32643 );
and ( n32645 , n32644 , n32540 );
or ( n32646 , n32641 , n32645 );
buf ( n32647 , n32646 );
not ( n32648 , n32647 );
buf ( n32649 , n32648 );
buf ( n32650 , n32649 );
not ( n32651 , n32650 );
or ( n32652 , n32638 , n32651 );
not ( n32653 , n32540 );
buf ( n32654 , n13387 );
and ( n32655 , n32653 , n32654 );
not ( n32656 , n32654 );
and ( n32657 , n32642 , n32643 );
xor ( n32658 , n32656 , n32657 );
and ( n32659 , n32658 , n32540 );
or ( n32660 , n32655 , n32659 );
buf ( n32661 , n32660 );
not ( n32662 , n32661 );
buf ( n32663 , n32662 );
buf ( n32664 , n32663 );
not ( n32665 , n32664 );
or ( n32666 , n32652 , n32665 );
not ( n32667 , n32540 );
buf ( n32668 , n13375 );
and ( n32669 , n32667 , n32668 );
not ( n32670 , n32668 );
and ( n32671 , n32656 , n32657 );
xor ( n32672 , n32670 , n32671 );
and ( n32673 , n32672 , n32540 );
or ( n32674 , n32669 , n32673 );
buf ( n32675 , n32674 );
not ( n32676 , n32675 );
buf ( n32677 , n32676 );
buf ( n32678 , n32677 );
not ( n32679 , n32678 );
or ( n32680 , n32666 , n32679 );
not ( n32681 , n32540 );
buf ( n32682 , n13363 );
and ( n32683 , n32681 , n32682 );
not ( n32684 , n32682 );
and ( n32685 , n32670 , n32671 );
xor ( n32686 , n32684 , n32685 );
and ( n32687 , n32686 , n32540 );
or ( n32688 , n32683 , n32687 );
buf ( n32689 , n32688 );
not ( n32690 , n32689 );
buf ( n32691 , n32690 );
buf ( n32692 , n32691 );
not ( n32693 , n32692 );
or ( n32694 , n32680 , n32693 );
not ( n32695 , n32540 );
buf ( n32696 , n13351 );
and ( n32697 , n32695 , n32696 );
not ( n32698 , n32696 );
and ( n32699 , n32684 , n32685 );
xor ( n32700 , n32698 , n32699 );
and ( n32701 , n32700 , n32540 );
or ( n32702 , n32697 , n32701 );
buf ( n32703 , n32702 );
not ( n32704 , n32703 );
buf ( n32705 , n32704 );
buf ( n32706 , n32705 );
not ( n32707 , n32706 );
or ( n32708 , n32694 , n32707 );
not ( n32709 , n32540 );
buf ( n32710 , n13339 );
and ( n32711 , n32709 , n32710 );
not ( n32712 , n32710 );
and ( n32713 , n32698 , n32699 );
xor ( n32714 , n32712 , n32713 );
and ( n32715 , n32714 , n32540 );
or ( n32716 , n32711 , n32715 );
buf ( n32717 , n32716 );
not ( n32718 , n32717 );
buf ( n32719 , n32718 );
buf ( n32720 , n32719 );
not ( n32721 , n32720 );
or ( n32722 , n32708 , n32721 );
not ( n32723 , n32540 );
buf ( n32724 , n13327 );
and ( n32725 , n32723 , n32724 );
not ( n32726 , n32724 );
and ( n32727 , n32712 , n32713 );
xor ( n32728 , n32726 , n32727 );
and ( n32729 , n32728 , n32540 );
or ( n32730 , n32725 , n32729 );
buf ( n32731 , n32730 );
not ( n32732 , n32731 );
buf ( n32733 , n32732 );
buf ( n32734 , n32733 );
not ( n32735 , n32734 );
or ( n32736 , n32722 , n32735 );
not ( n32737 , n32540 );
buf ( n32738 , n13315 );
and ( n32739 , n32737 , n32738 );
not ( n32740 , n32738 );
and ( n32741 , n32726 , n32727 );
xor ( n32742 , n32740 , n32741 );
and ( n32743 , n32742 , n32540 );
or ( n32744 , n32739 , n32743 );
buf ( n32745 , n32744 );
not ( n32746 , n32745 );
buf ( n32747 , n32746 );
buf ( n32748 , n32747 );
not ( n32749 , n32748 );
or ( n32750 , n32736 , n32749 );
not ( n32751 , n32540 );
buf ( n32752 , n13303 );
and ( n32753 , n32751 , n32752 );
not ( n32754 , n32752 );
and ( n32755 , n32740 , n32741 );
xor ( n32756 , n32754 , n32755 );
and ( n32757 , n32756 , n32540 );
or ( n32758 , n32753 , n32757 );
buf ( n32759 , n32758 );
not ( n32760 , n32759 );
buf ( n32761 , n32760 );
buf ( n32762 , n32761 );
not ( n32763 , n32762 );
or ( n32764 , n32750 , n32763 );
not ( n32765 , n32540 );
buf ( n32766 , n13291 );
and ( n32767 , n32765 , n32766 );
not ( n32768 , n32766 );
and ( n32769 , n32754 , n32755 );
xor ( n32770 , n32768 , n32769 );
and ( n32771 , n32770 , n32540 );
or ( n32772 , n32767 , n32771 );
buf ( n32773 , n32772 );
not ( n32774 , n32773 );
buf ( n32775 , n32774 );
buf ( n32776 , n32775 );
not ( n32777 , n32776 );
or ( n32778 , n32764 , n32777 );
not ( n32779 , n32540 );
buf ( n32780 , n13279 );
and ( n32781 , n32779 , n32780 );
not ( n32782 , n32780 );
and ( n32783 , n32768 , n32769 );
xor ( n32784 , n32782 , n32783 );
and ( n32785 , n32784 , n32540 );
or ( n32786 , n32781 , n32785 );
buf ( n32787 , n32786 );
not ( n32788 , n32787 );
buf ( n32789 , n32788 );
buf ( n32790 , n32789 );
not ( n32791 , n32790 );
or ( n32792 , n32778 , n32791 );
not ( n32793 , n32540 );
buf ( n32794 , n13267 );
and ( n32795 , n32793 , n32794 );
not ( n32796 , n32794 );
and ( n32797 , n32782 , n32783 );
xor ( n32798 , n32796 , n32797 );
and ( n32799 , n32798 , n32540 );
or ( n32800 , n32795 , n32799 );
buf ( n32801 , n32800 );
not ( n32802 , n32801 );
buf ( n32803 , n32802 );
buf ( n32804 , n32803 );
not ( n32805 , n32804 );
or ( n32806 , n32792 , n32805 );
buf ( n32807 , n32806 );
buf ( n32808 , n32807 );
and ( n32809 , n32808 , n32540 );
not ( n32810 , n32809 );
and ( n32811 , n32810 , n32539 );
xor ( n32812 , n32539 , n32540 );
xor ( n32813 , n32812 , n32540 );
and ( n32814 , n32813 , n32809 );
or ( n32815 , n32811 , n32814 );
buf ( n32816 , n32815 );
buf ( n32817 , n32816 );
buf ( n32818 , n32529 );
xor ( n32819 , n32817 , n32818 );
buf ( n32820 , n32819 );
and ( n32821 , n32820 , n14141 );
or ( n32822 , n14140 , n14137 );
and ( n32823 , n15864 , n32822 );
or ( n32824 , n32533 , n32821 , n32823 );
buf ( n32825 , n32824 );
buf ( n32826 , n32825 );
not ( n32827 , n32826 );
buf ( n32828 , n32827 );
buf ( n32829 , n32828 );
not ( n32830 , n32829 );
xor ( n32831 , n32511 , n32246 );
xor ( n32832 , n32497 , n32246 );
xor ( n32833 , n32483 , n32246 );
xor ( n32834 , n32469 , n32246 );
xor ( n32835 , n32455 , n32246 );
xor ( n32836 , n32441 , n32246 );
xor ( n32837 , n32427 , n32246 );
xor ( n32838 , n32413 , n32246 );
xor ( n32839 , n32399 , n32246 );
xor ( n32840 , n32385 , n32246 );
xor ( n32841 , n32371 , n32246 );
xor ( n32842 , n32357 , n32246 );
xor ( n32843 , n32343 , n32246 );
xor ( n32844 , n32329 , n32246 );
xor ( n32845 , n32315 , n32246 );
xor ( n32846 , n32301 , n32246 );
xor ( n32847 , n32287 , n32246 );
xor ( n32848 , n32273 , n32246 );
xor ( n32849 , n32259 , n32246 );
and ( n32850 , n32518 , n32246 );
and ( n32851 , n32849 , n32850 );
and ( n32852 , n32848 , n32851 );
and ( n32853 , n32847 , n32852 );
and ( n32854 , n32846 , n32853 );
and ( n32855 , n32845 , n32854 );
and ( n32856 , n32844 , n32855 );
and ( n32857 , n32843 , n32856 );
and ( n32858 , n32842 , n32857 );
and ( n32859 , n32841 , n32858 );
and ( n32860 , n32840 , n32859 );
and ( n32861 , n32839 , n32860 );
and ( n32862 , n32838 , n32861 );
and ( n32863 , n32837 , n32862 );
and ( n32864 , n32836 , n32863 );
and ( n32865 , n32835 , n32864 );
and ( n32866 , n32834 , n32865 );
and ( n32867 , n32833 , n32866 );
and ( n32868 , n32832 , n32867 );
and ( n32869 , n32831 , n32868 );
buf ( n32870 , n32869 );
and ( n32871 , n32870 , n32515 );
or ( n32872 , C0 , n32871 );
buf ( n32873 , n32872 );
buf ( n32874 , n32873 );
not ( n32875 , n32515 );
and ( n32876 , n32875 , n32511 );
xor ( n32877 , n32831 , n32868 );
and ( n32878 , n32877 , n32515 );
or ( n32879 , n32876 , n32878 );
buf ( n32880 , n32879 );
buf ( n32881 , n32880 );
buf ( n32882 , n15447 );
not ( n32883 , n32882 );
buf ( n32884 , n32883 );
buf ( n32885 , n32884 );
not ( n32886 , n32885 );
buf ( n32887 , n32886 );
buf ( n32888 , n32887 );
buf ( n32889 , n32888 );
not ( n32890 , n32889 );
and ( n32891 , n32881 , n32890 );
not ( n32892 , n32515 );
and ( n32893 , n32892 , n32497 );
xor ( n32894 , n32832 , n32867 );
and ( n32895 , n32894 , n32515 );
or ( n32896 , n32893 , n32895 );
buf ( n32897 , n32896 );
buf ( n32898 , n32897 );
buf ( n32899 , n15469 );
not ( n32900 , n32899 );
buf ( n32901 , n32900 );
buf ( n32902 , n32901 );
not ( n32903 , n32902 );
buf ( n32904 , n32903 );
buf ( n32905 , n32904 );
buf ( n32906 , n32905 );
not ( n32907 , n32906 );
and ( n32908 , n32898 , n32907 );
not ( n32909 , n32515 );
and ( n32910 , n32909 , n32483 );
xor ( n32911 , n32833 , n32866 );
and ( n32912 , n32911 , n32515 );
or ( n32913 , n32910 , n32912 );
buf ( n32914 , n32913 );
buf ( n32915 , n32914 );
buf ( n32916 , n15491 );
not ( n32917 , n32916 );
buf ( n32918 , n32917 );
buf ( n32919 , n32918 );
not ( n32920 , n32919 );
buf ( n32921 , n32920 );
buf ( n32922 , n32921 );
buf ( n32923 , n32922 );
not ( n32924 , n32923 );
and ( n32925 , n32915 , n32924 );
not ( n32926 , n32515 );
and ( n32927 , n32926 , n32469 );
xor ( n32928 , n32834 , n32865 );
and ( n32929 , n32928 , n32515 );
or ( n32930 , n32927 , n32929 );
buf ( n32931 , n32930 );
buf ( n32932 , n32931 );
buf ( n32933 , n15513 );
not ( n32934 , n32933 );
buf ( n32935 , n32934 );
buf ( n32936 , n32935 );
not ( n32937 , n32936 );
buf ( n32938 , n32937 );
buf ( n32939 , n32938 );
buf ( n32940 , n32939 );
not ( n32941 , n32940 );
and ( n32942 , n32932 , n32941 );
not ( n32943 , n32515 );
and ( n32944 , n32943 , n32455 );
xor ( n32945 , n32835 , n32864 );
and ( n32946 , n32945 , n32515 );
or ( n32947 , n32944 , n32946 );
buf ( n32948 , n32947 );
buf ( n32949 , n32948 );
buf ( n32950 , n15535 );
not ( n32951 , n32950 );
buf ( n32952 , n32951 );
buf ( n32953 , n32952 );
not ( n32954 , n32953 );
buf ( n32955 , n32954 );
buf ( n32956 , n32955 );
buf ( n32957 , n32956 );
not ( n32958 , n32957 );
and ( n32959 , n32949 , n32958 );
not ( n32960 , n32515 );
and ( n32961 , n32960 , n32441 );
xor ( n32962 , n32836 , n32863 );
and ( n32963 , n32962 , n32515 );
or ( n32964 , n32961 , n32963 );
buf ( n32965 , n32964 );
buf ( n32966 , n32965 );
buf ( n32967 , n15557 );
not ( n32968 , n32967 );
buf ( n32969 , n32968 );
buf ( n32970 , n32969 );
not ( n32971 , n32970 );
buf ( n32972 , n32971 );
buf ( n32973 , n32972 );
buf ( n32974 , n32973 );
not ( n32975 , n32974 );
and ( n32976 , n32966 , n32975 );
not ( n32977 , n32515 );
and ( n32978 , n32977 , n32427 );
xor ( n32979 , n32837 , n32862 );
and ( n32980 , n32979 , n32515 );
or ( n32981 , n32978 , n32980 );
buf ( n32982 , n32981 );
buf ( n32983 , n32982 );
buf ( n32984 , n15579 );
not ( n32985 , n32984 );
buf ( n32986 , n32985 );
buf ( n32987 , n32986 );
not ( n32988 , n32987 );
buf ( n32989 , n32988 );
buf ( n32990 , n32989 );
buf ( n32991 , n32990 );
not ( n32992 , n32991 );
and ( n32993 , n32983 , n32992 );
not ( n32994 , n32515 );
and ( n32995 , n32994 , n32413 );
xor ( n32996 , n32838 , n32861 );
and ( n32997 , n32996 , n32515 );
or ( n32998 , n32995 , n32997 );
buf ( n32999 , n32998 );
buf ( n33000 , n32999 );
buf ( n33001 , n15601 );
not ( n33002 , n33001 );
buf ( n33003 , n33002 );
buf ( n33004 , n33003 );
not ( n33005 , n33004 );
buf ( n33006 , n33005 );
buf ( n33007 , n33006 );
buf ( n33008 , n33007 );
not ( n33009 , n33008 );
and ( n33010 , n33000 , n33009 );
not ( n33011 , n32515 );
and ( n33012 , n33011 , n32399 );
xor ( n33013 , n32839 , n32860 );
and ( n33014 , n33013 , n32515 );
or ( n33015 , n33012 , n33014 );
buf ( n33016 , n33015 );
buf ( n33017 , n33016 );
buf ( n33018 , n15623 );
not ( n33019 , n33018 );
buf ( n33020 , n33019 );
buf ( n33021 , n33020 );
not ( n33022 , n33021 );
buf ( n33023 , n33022 );
buf ( n33024 , n33023 );
buf ( n33025 , n33024 );
not ( n33026 , n33025 );
and ( n33027 , n33017 , n33026 );
not ( n33028 , n32515 );
and ( n33029 , n33028 , n32385 );
xor ( n33030 , n32840 , n32859 );
and ( n33031 , n33030 , n32515 );
or ( n33032 , n33029 , n33031 );
buf ( n33033 , n33032 );
buf ( n33034 , n33033 );
buf ( n33035 , n15645 );
not ( n33036 , n33035 );
buf ( n33037 , n33036 );
buf ( n33038 , n33037 );
not ( n33039 , n33038 );
buf ( n33040 , n33039 );
buf ( n33041 , n33040 );
buf ( n33042 , n33041 );
not ( n33043 , n33042 );
and ( n33044 , n33034 , n33043 );
not ( n33045 , n32515 );
and ( n33046 , n33045 , n32371 );
xor ( n33047 , n32841 , n32858 );
and ( n33048 , n33047 , n32515 );
or ( n33049 , n33046 , n33048 );
buf ( n33050 , n33049 );
buf ( n33051 , n33050 );
buf ( n33052 , n15667 );
not ( n33053 , n33052 );
buf ( n33054 , n33053 );
buf ( n33055 , n33054 );
not ( n33056 , n33055 );
buf ( n33057 , n33056 );
buf ( n33058 , n33057 );
buf ( n33059 , n33058 );
not ( n33060 , n33059 );
and ( n33061 , n33051 , n33060 );
not ( n33062 , n32515 );
and ( n33063 , n33062 , n32357 );
xor ( n33064 , n32842 , n32857 );
and ( n33065 , n33064 , n32515 );
or ( n33066 , n33063 , n33065 );
buf ( n33067 , n33066 );
buf ( n33068 , n33067 );
buf ( n33069 , n15689 );
not ( n33070 , n33069 );
buf ( n33071 , n33070 );
buf ( n33072 , n33071 );
not ( n33073 , n33072 );
buf ( n33074 , n33073 );
buf ( n33075 , n33074 );
buf ( n33076 , n33075 );
not ( n33077 , n33076 );
and ( n33078 , n33068 , n33077 );
not ( n33079 , n32515 );
and ( n33080 , n33079 , n32343 );
xor ( n33081 , n32843 , n32856 );
and ( n33082 , n33081 , n32515 );
or ( n33083 , n33080 , n33082 );
buf ( n33084 , n33083 );
buf ( n33085 , n33084 );
buf ( n33086 , n15711 );
not ( n33087 , n33086 );
buf ( n33088 , n33087 );
buf ( n33089 , n33088 );
not ( n33090 , n33089 );
buf ( n33091 , n33090 );
buf ( n33092 , n33091 );
buf ( n33093 , n33092 );
not ( n33094 , n33093 );
and ( n33095 , n33085 , n33094 );
not ( n33096 , n32515 );
and ( n33097 , n33096 , n32329 );
xor ( n33098 , n32844 , n32855 );
and ( n33099 , n33098 , n32515 );
or ( n33100 , n33097 , n33099 );
buf ( n33101 , n33100 );
buf ( n33102 , n33101 );
buf ( n33103 , n15733 );
not ( n33104 , n33103 );
buf ( n33105 , n33104 );
buf ( n33106 , n33105 );
not ( n33107 , n33106 );
buf ( n33108 , n33107 );
buf ( n33109 , n33108 );
buf ( n33110 , n33109 );
not ( n33111 , n33110 );
and ( n33112 , n33102 , n33111 );
not ( n33113 , n32515 );
and ( n33114 , n33113 , n32315 );
xor ( n33115 , n32845 , n32854 );
and ( n33116 , n33115 , n32515 );
or ( n33117 , n33114 , n33116 );
buf ( n33118 , n33117 );
buf ( n33119 , n33118 );
buf ( n33120 , n15755 );
not ( n33121 , n33120 );
buf ( n33122 , n33121 );
buf ( n33123 , n33122 );
not ( n33124 , n33123 );
buf ( n33125 , n33124 );
buf ( n33126 , n33125 );
buf ( n33127 , n33126 );
not ( n33128 , n33127 );
and ( n33129 , n33119 , n33128 );
not ( n33130 , n32515 );
and ( n33131 , n33130 , n32301 );
xor ( n33132 , n32846 , n32853 );
and ( n33133 , n33132 , n32515 );
or ( n33134 , n33131 , n33133 );
buf ( n33135 , n33134 );
buf ( n33136 , n33135 );
buf ( n33137 , n15777 );
not ( n33138 , n33137 );
buf ( n33139 , n33138 );
buf ( n33140 , n33139 );
not ( n33141 , n33140 );
buf ( n33142 , n33141 );
buf ( n33143 , n33142 );
buf ( n33144 , n33143 );
not ( n33145 , n33144 );
and ( n33146 , n33136 , n33145 );
not ( n33147 , n32515 );
and ( n33148 , n33147 , n32287 );
xor ( n33149 , n32847 , n32852 );
and ( n33150 , n33149 , n32515 );
or ( n33151 , n33148 , n33150 );
buf ( n33152 , n33151 );
buf ( n33153 , n33152 );
buf ( n33154 , n15799 );
not ( n33155 , n33154 );
buf ( n33156 , n33155 );
buf ( n33157 , n33156 );
not ( n33158 , n33157 );
buf ( n33159 , n33158 );
buf ( n33160 , n33159 );
buf ( n33161 , n33160 );
not ( n33162 , n33161 );
and ( n33163 , n33153 , n33162 );
not ( n33164 , n32515 );
and ( n33165 , n33164 , n32273 );
xor ( n33166 , n32848 , n32851 );
and ( n33167 , n33166 , n32515 );
or ( n33168 , n33165 , n33167 );
buf ( n33169 , n33168 );
buf ( n33170 , n33169 );
buf ( n33171 , n15821 );
not ( n33172 , n33171 );
buf ( n33173 , n33172 );
buf ( n33174 , n33173 );
not ( n33175 , n33174 );
buf ( n33176 , n33175 );
buf ( n33177 , n33176 );
buf ( n33178 , n33177 );
not ( n33179 , n33178 );
and ( n33180 , n33170 , n33179 );
not ( n33181 , n32515 );
and ( n33182 , n33181 , n32259 );
xor ( n33183 , n32849 , n32850 );
and ( n33184 , n33183 , n32515 );
or ( n33185 , n33182 , n33184 );
buf ( n33186 , n33185 );
buf ( n33187 , n33186 );
buf ( n33188 , n15843 );
not ( n33189 , n33188 );
buf ( n33190 , n33189 );
buf ( n33191 , n33190 );
not ( n33192 , n33191 );
buf ( n33193 , n33192 );
buf ( n33194 , n33193 );
buf ( n33195 , n33194 );
not ( n33196 , n33195 );
and ( n33197 , n33187 , n33196 );
not ( n33198 , n32530 );
or ( n33199 , n32523 , n33198 );
and ( n33200 , n33196 , n33199 );
and ( n33201 , n33187 , n33199 );
or ( n33202 , n33197 , n33200 , n33201 );
and ( n33203 , n33179 , n33202 );
and ( n33204 , n33170 , n33202 );
or ( n33205 , n33180 , n33203 , n33204 );
and ( n33206 , n33162 , n33205 );
and ( n33207 , n33153 , n33205 );
or ( n33208 , n33163 , n33206 , n33207 );
and ( n33209 , n33145 , n33208 );
and ( n33210 , n33136 , n33208 );
or ( n33211 , n33146 , n33209 , n33210 );
and ( n33212 , n33128 , n33211 );
and ( n33213 , n33119 , n33211 );
or ( n33214 , n33129 , n33212 , n33213 );
and ( n33215 , n33111 , n33214 );
and ( n33216 , n33102 , n33214 );
or ( n33217 , n33112 , n33215 , n33216 );
and ( n33218 , n33094 , n33217 );
and ( n33219 , n33085 , n33217 );
or ( n33220 , n33095 , n33218 , n33219 );
and ( n33221 , n33077 , n33220 );
and ( n33222 , n33068 , n33220 );
or ( n33223 , n33078 , n33221 , n33222 );
and ( n33224 , n33060 , n33223 );
and ( n33225 , n33051 , n33223 );
or ( n33226 , n33061 , n33224 , n33225 );
and ( n33227 , n33043 , n33226 );
and ( n33228 , n33034 , n33226 );
or ( n33229 , n33044 , n33227 , n33228 );
and ( n33230 , n33026 , n33229 );
and ( n33231 , n33017 , n33229 );
or ( n33232 , n33027 , n33230 , n33231 );
and ( n33233 , n33009 , n33232 );
and ( n33234 , n33000 , n33232 );
or ( n33235 , n33010 , n33233 , n33234 );
and ( n33236 , n32992 , n33235 );
and ( n33237 , n32983 , n33235 );
or ( n33238 , n32993 , n33236 , n33237 );
and ( n33239 , n32975 , n33238 );
and ( n33240 , n32966 , n33238 );
or ( n33241 , n32976 , n33239 , n33240 );
and ( n33242 , n32958 , n33241 );
and ( n33243 , n32949 , n33241 );
or ( n33244 , n32959 , n33242 , n33243 );
and ( n33245 , n32941 , n33244 );
and ( n33246 , n32932 , n33244 );
or ( n33247 , n32942 , n33245 , n33246 );
and ( n33248 , n32924 , n33247 );
and ( n33249 , n32915 , n33247 );
or ( n33250 , n32925 , n33248 , n33249 );
and ( n33251 , n32907 , n33250 );
and ( n33252 , n32898 , n33250 );
or ( n33253 , n32908 , n33251 , n33252 );
and ( n33254 , n32890 , n33253 );
and ( n33255 , n32881 , n33253 );
or ( n33256 , n32891 , n33254 , n33255 );
or ( n33257 , n32874 , n33256 );
buf ( n33258 , n33257 );
buf ( n33259 , n33258 );
or ( n33260 , C0 , n33259 );
or ( n33261 , C0 , n33260 );
or ( n33262 , C0 , n33261 );
or ( n33263 , C0 , n33262 );
or ( n33264 , C0 , n33263 );
or ( n33265 , C0 , n33264 );
or ( n33266 , C0 , n33265 );
or ( n33267 , C0 , n33266 );
xnor ( n33268 , C0 , n33267 );
buf ( n33269 , n33268 );
and ( n33270 , n33269 , n14143 );
xor ( n33271 , n32805 , n32540 );
xor ( n33272 , n32791 , n32540 );
xor ( n33273 , n32777 , n32540 );
xor ( n33274 , n32763 , n32540 );
xor ( n33275 , n32749 , n32540 );
xor ( n33276 , n32735 , n32540 );
xor ( n33277 , n32721 , n32540 );
xor ( n33278 , n32707 , n32540 );
xor ( n33279 , n32693 , n32540 );
xor ( n33280 , n32679 , n32540 );
xor ( n33281 , n32665 , n32540 );
xor ( n33282 , n32651 , n32540 );
xor ( n33283 , n32637 , n32540 );
xor ( n33284 , n32623 , n32540 );
xor ( n33285 , n32609 , n32540 );
xor ( n33286 , n32595 , n32540 );
xor ( n33287 , n32581 , n32540 );
xor ( n33288 , n32567 , n32540 );
xor ( n33289 , n32553 , n32540 );
and ( n33290 , n32812 , n32540 );
and ( n33291 , n33289 , n33290 );
and ( n33292 , n33288 , n33291 );
and ( n33293 , n33287 , n33292 );
and ( n33294 , n33286 , n33293 );
and ( n33295 , n33285 , n33294 );
and ( n33296 , n33284 , n33295 );
and ( n33297 , n33283 , n33296 );
and ( n33298 , n33282 , n33297 );
and ( n33299 , n33281 , n33298 );
and ( n33300 , n33280 , n33299 );
and ( n33301 , n33279 , n33300 );
and ( n33302 , n33278 , n33301 );
and ( n33303 , n33277 , n33302 );
and ( n33304 , n33276 , n33303 );
and ( n33305 , n33275 , n33304 );
and ( n33306 , n33274 , n33305 );
and ( n33307 , n33273 , n33306 );
and ( n33308 , n33272 , n33307 );
and ( n33309 , n33271 , n33308 );
buf ( n33310 , n33309 );
and ( n33311 , n33310 , n32809 );
or ( n33312 , C0 , n33311 );
buf ( n33313 , n33312 );
buf ( n33314 , n33313 );
not ( n33315 , n32809 );
and ( n33316 , n33315 , n32805 );
xor ( n33317 , n33271 , n33308 );
and ( n33318 , n33317 , n32809 );
or ( n33319 , n33316 , n33318 );
buf ( n33320 , n33319 );
buf ( n33321 , n33320 );
buf ( n33322 , n32888 );
not ( n33323 , n33322 );
and ( n33324 , n33321 , n33323 );
not ( n33325 , n32809 );
and ( n33326 , n33325 , n32791 );
xor ( n33327 , n33272 , n33307 );
and ( n33328 , n33327 , n32809 );
or ( n33329 , n33326 , n33328 );
buf ( n33330 , n33329 );
buf ( n33331 , n33330 );
buf ( n33332 , n32905 );
not ( n33333 , n33332 );
and ( n33334 , n33331 , n33333 );
not ( n33335 , n32809 );
and ( n33336 , n33335 , n32777 );
xor ( n33337 , n33273 , n33306 );
and ( n33338 , n33337 , n32809 );
or ( n33339 , n33336 , n33338 );
buf ( n33340 , n33339 );
buf ( n33341 , n33340 );
buf ( n33342 , n32922 );
not ( n33343 , n33342 );
and ( n33344 , n33341 , n33343 );
not ( n33345 , n32809 );
and ( n33346 , n33345 , n32763 );
xor ( n33347 , n33274 , n33305 );
and ( n33348 , n33347 , n32809 );
or ( n33349 , n33346 , n33348 );
buf ( n33350 , n33349 );
buf ( n33351 , n33350 );
buf ( n33352 , n32939 );
not ( n33353 , n33352 );
and ( n33354 , n33351 , n33353 );
not ( n33355 , n32809 );
and ( n33356 , n33355 , n32749 );
xor ( n33357 , n33275 , n33304 );
and ( n33358 , n33357 , n32809 );
or ( n33359 , n33356 , n33358 );
buf ( n33360 , n33359 );
buf ( n33361 , n33360 );
buf ( n33362 , n32956 );
not ( n33363 , n33362 );
and ( n33364 , n33361 , n33363 );
not ( n33365 , n32809 );
and ( n33366 , n33365 , n32735 );
xor ( n33367 , n33276 , n33303 );
and ( n33368 , n33367 , n32809 );
or ( n33369 , n33366 , n33368 );
buf ( n33370 , n33369 );
buf ( n33371 , n33370 );
buf ( n33372 , n32973 );
not ( n33373 , n33372 );
and ( n33374 , n33371 , n33373 );
not ( n33375 , n32809 );
and ( n33376 , n33375 , n32721 );
xor ( n33377 , n33277 , n33302 );
and ( n33378 , n33377 , n32809 );
or ( n33379 , n33376 , n33378 );
buf ( n33380 , n33379 );
buf ( n33381 , n33380 );
buf ( n33382 , n32990 );
not ( n33383 , n33382 );
and ( n33384 , n33381 , n33383 );
not ( n33385 , n32809 );
and ( n33386 , n33385 , n32707 );
xor ( n33387 , n33278 , n33301 );
and ( n33388 , n33387 , n32809 );
or ( n33389 , n33386 , n33388 );
buf ( n33390 , n33389 );
buf ( n33391 , n33390 );
buf ( n33392 , n33007 );
not ( n33393 , n33392 );
and ( n33394 , n33391 , n33393 );
not ( n33395 , n32809 );
and ( n33396 , n33395 , n32693 );
xor ( n33397 , n33279 , n33300 );
and ( n33398 , n33397 , n32809 );
or ( n33399 , n33396 , n33398 );
buf ( n33400 , n33399 );
buf ( n33401 , n33400 );
buf ( n33402 , n33024 );
not ( n33403 , n33402 );
and ( n33404 , n33401 , n33403 );
not ( n33405 , n32809 );
and ( n33406 , n33405 , n32679 );
xor ( n33407 , n33280 , n33299 );
and ( n33408 , n33407 , n32809 );
or ( n33409 , n33406 , n33408 );
buf ( n33410 , n33409 );
buf ( n33411 , n33410 );
buf ( n33412 , n33041 );
not ( n33413 , n33412 );
and ( n33414 , n33411 , n33413 );
not ( n33415 , n32809 );
and ( n33416 , n33415 , n32665 );
xor ( n33417 , n33281 , n33298 );
and ( n33418 , n33417 , n32809 );
or ( n33419 , n33416 , n33418 );
buf ( n33420 , n33419 );
buf ( n33421 , n33420 );
buf ( n33422 , n33058 );
not ( n33423 , n33422 );
and ( n33424 , n33421 , n33423 );
not ( n33425 , n32809 );
and ( n33426 , n33425 , n32651 );
xor ( n33427 , n33282 , n33297 );
and ( n33428 , n33427 , n32809 );
or ( n33429 , n33426 , n33428 );
buf ( n33430 , n33429 );
buf ( n33431 , n33430 );
buf ( n33432 , n33075 );
not ( n33433 , n33432 );
and ( n33434 , n33431 , n33433 );
not ( n33435 , n32809 );
and ( n33436 , n33435 , n32637 );
xor ( n33437 , n33283 , n33296 );
and ( n33438 , n33437 , n32809 );
or ( n33439 , n33436 , n33438 );
buf ( n33440 , n33439 );
buf ( n33441 , n33440 );
buf ( n33442 , n33092 );
not ( n33443 , n33442 );
and ( n33444 , n33441 , n33443 );
not ( n33445 , n32809 );
and ( n33446 , n33445 , n32623 );
xor ( n33447 , n33284 , n33295 );
and ( n33448 , n33447 , n32809 );
or ( n33449 , n33446 , n33448 );
buf ( n33450 , n33449 );
buf ( n33451 , n33450 );
buf ( n33452 , n33109 );
not ( n33453 , n33452 );
and ( n33454 , n33451 , n33453 );
not ( n33455 , n32809 );
and ( n33456 , n33455 , n32609 );
xor ( n33457 , n33285 , n33294 );
and ( n33458 , n33457 , n32809 );
or ( n33459 , n33456 , n33458 );
buf ( n33460 , n33459 );
buf ( n33461 , n33460 );
buf ( n33462 , n33126 );
not ( n33463 , n33462 );
and ( n33464 , n33461 , n33463 );
not ( n33465 , n32809 );
and ( n33466 , n33465 , n32595 );
xor ( n33467 , n33286 , n33293 );
and ( n33468 , n33467 , n32809 );
or ( n33469 , n33466 , n33468 );
buf ( n33470 , n33469 );
buf ( n33471 , n33470 );
buf ( n33472 , n33143 );
not ( n33473 , n33472 );
and ( n33474 , n33471 , n33473 );
not ( n33475 , n32809 );
and ( n33476 , n33475 , n32581 );
xor ( n33477 , n33287 , n33292 );
and ( n33478 , n33477 , n32809 );
or ( n33479 , n33476 , n33478 );
buf ( n33480 , n33479 );
buf ( n33481 , n33480 );
buf ( n33482 , n33160 );
not ( n33483 , n33482 );
and ( n33484 , n33481 , n33483 );
not ( n33485 , n32809 );
and ( n33486 , n33485 , n32567 );
xor ( n33487 , n33288 , n33291 );
and ( n33488 , n33487 , n32809 );
or ( n33489 , n33486 , n33488 );
buf ( n33490 , n33489 );
buf ( n33491 , n33490 );
buf ( n33492 , n33177 );
not ( n33493 , n33492 );
and ( n33494 , n33491 , n33493 );
not ( n33495 , n32809 );
and ( n33496 , n33495 , n32553 );
xor ( n33497 , n33289 , n33290 );
and ( n33498 , n33497 , n32809 );
or ( n33499 , n33496 , n33498 );
buf ( n33500 , n33499 );
buf ( n33501 , n33500 );
buf ( n33502 , n33194 );
not ( n33503 , n33502 );
and ( n33504 , n33501 , n33503 );
not ( n33505 , n32818 );
or ( n33506 , n32817 , n33505 );
and ( n33507 , n33503 , n33506 );
and ( n33508 , n33501 , n33506 );
or ( n33509 , n33504 , n33507 , n33508 );
and ( n33510 , n33493 , n33509 );
and ( n33511 , n33491 , n33509 );
or ( n33512 , n33494 , n33510 , n33511 );
and ( n33513 , n33483 , n33512 );
and ( n33514 , n33481 , n33512 );
or ( n33515 , n33484 , n33513 , n33514 );
and ( n33516 , n33473 , n33515 );
and ( n33517 , n33471 , n33515 );
or ( n33518 , n33474 , n33516 , n33517 );
and ( n33519 , n33463 , n33518 );
and ( n33520 , n33461 , n33518 );
or ( n33521 , n33464 , n33519 , n33520 );
and ( n33522 , n33453 , n33521 );
and ( n33523 , n33451 , n33521 );
or ( n33524 , n33454 , n33522 , n33523 );
and ( n33525 , n33443 , n33524 );
and ( n33526 , n33441 , n33524 );
or ( n33527 , n33444 , n33525 , n33526 );
and ( n33528 , n33433 , n33527 );
and ( n33529 , n33431 , n33527 );
or ( n33530 , n33434 , n33528 , n33529 );
and ( n33531 , n33423 , n33530 );
and ( n33532 , n33421 , n33530 );
or ( n33533 , n33424 , n33531 , n33532 );
and ( n33534 , n33413 , n33533 );
and ( n33535 , n33411 , n33533 );
or ( n33536 , n33414 , n33534 , n33535 );
and ( n33537 , n33403 , n33536 );
and ( n33538 , n33401 , n33536 );
or ( n33539 , n33404 , n33537 , n33538 );
and ( n33540 , n33393 , n33539 );
and ( n33541 , n33391 , n33539 );
or ( n33542 , n33394 , n33540 , n33541 );
and ( n33543 , n33383 , n33542 );
and ( n33544 , n33381 , n33542 );
or ( n33545 , n33384 , n33543 , n33544 );
and ( n33546 , n33373 , n33545 );
and ( n33547 , n33371 , n33545 );
or ( n33548 , n33374 , n33546 , n33547 );
and ( n33549 , n33363 , n33548 );
and ( n33550 , n33361 , n33548 );
or ( n33551 , n33364 , n33549 , n33550 );
and ( n33552 , n33353 , n33551 );
and ( n33553 , n33351 , n33551 );
or ( n33554 , n33354 , n33552 , n33553 );
and ( n33555 , n33343 , n33554 );
and ( n33556 , n33341 , n33554 );
or ( n33557 , n33344 , n33555 , n33556 );
and ( n33558 , n33333 , n33557 );
and ( n33559 , n33331 , n33557 );
or ( n33560 , n33334 , n33558 , n33559 );
and ( n33561 , n33323 , n33560 );
and ( n33562 , n33321 , n33560 );
or ( n33563 , n33324 , n33561 , n33562 );
or ( n33564 , n33314 , n33563 );
buf ( n33565 , n33564 );
buf ( n33566 , n33565 );
or ( n33567 , C0 , n33566 );
or ( n33568 , C0 , n33567 );
or ( n33569 , C0 , n33568 );
or ( n33570 , C0 , n33569 );
or ( n33571 , C0 , n33570 );
or ( n33572 , C0 , n33571 );
or ( n33573 , C0 , n33572 );
or ( n33574 , C0 , n33573 );
xnor ( n33575 , C0 , n33574 );
buf ( n33576 , n33575 );
and ( n33577 , n33576 , n14141 );
or ( n33578 , n33270 , n33577 , C0 );
buf ( n33579 , n33578 );
not ( n33580 , n33579 );
xor ( n33581 , n33187 , n33196 );
xor ( n33582 , n33581 , n33199 );
buf ( n33583 , n33582 );
and ( n33584 , n33583 , n14143 );
xor ( n33585 , n33501 , n33503 );
xor ( n33586 , n33585 , n33506 );
buf ( n33587 , n33586 );
and ( n33588 , n33587 , n14141 );
and ( n33589 , n15843 , n32822 );
or ( n33590 , n33584 , n33588 , n33589 );
buf ( n33591 , n33590 );
and ( n33592 , n33580 , n33591 );
not ( n33593 , n33591 );
not ( n33594 , n32825 );
xor ( n33595 , n33593 , n33594 );
and ( n33596 , n33595 , n33579 );
or ( n33597 , n33592 , n33596 );
buf ( n33598 , n33597 );
not ( n33599 , n33598 );
buf ( n33600 , n33599 );
buf ( n33601 , n33600 );
not ( n33602 , n33601 );
or ( n33603 , n32830 , n33602 );
not ( n33604 , n33579 );
xor ( n33605 , n33170 , n33179 );
xor ( n33606 , n33605 , n33202 );
buf ( n33607 , n33606 );
and ( n33608 , n33607 , n14143 );
xor ( n33609 , n33491 , n33493 );
xor ( n33610 , n33609 , n33509 );
buf ( n33611 , n33610 );
and ( n33612 , n33611 , n14141 );
and ( n33613 , n15821 , n32822 );
or ( n33614 , n33608 , n33612 , n33613 );
buf ( n33615 , n33614 );
and ( n33616 , n33604 , n33615 );
not ( n33617 , n33615 );
and ( n33618 , n33593 , n33594 );
xor ( n33619 , n33617 , n33618 );
and ( n33620 , n33619 , n33579 );
or ( n33621 , n33616 , n33620 );
buf ( n33622 , n33621 );
not ( n33623 , n33622 );
buf ( n33624 , n33623 );
buf ( n33625 , n33624 );
not ( n33626 , n33625 );
or ( n33627 , n33603 , n33626 );
not ( n33628 , n33579 );
xor ( n33629 , n33153 , n33162 );
xor ( n33630 , n33629 , n33205 );
buf ( n33631 , n33630 );
and ( n33632 , n33631 , n14143 );
xor ( n33633 , n33481 , n33483 );
xor ( n33634 , n33633 , n33512 );
buf ( n33635 , n33634 );
and ( n33636 , n33635 , n14141 );
and ( n33637 , n15799 , n32822 );
or ( n33638 , n33632 , n33636 , n33637 );
buf ( n33639 , n33638 );
and ( n33640 , n33628 , n33639 );
not ( n33641 , n33639 );
and ( n33642 , n33617 , n33618 );
xor ( n33643 , n33641 , n33642 );
and ( n33644 , n33643 , n33579 );
or ( n33645 , n33640 , n33644 );
buf ( n33646 , n33645 );
not ( n33647 , n33646 );
buf ( n33648 , n33647 );
buf ( n33649 , n33648 );
not ( n33650 , n33649 );
or ( n33651 , n33627 , n33650 );
not ( n33652 , n33579 );
xor ( n33653 , n33136 , n33145 );
xor ( n33654 , n33653 , n33208 );
buf ( n33655 , n33654 );
and ( n33656 , n33655 , n14143 );
xor ( n33657 , n33471 , n33473 );
xor ( n33658 , n33657 , n33515 );
buf ( n33659 , n33658 );
and ( n33660 , n33659 , n14141 );
and ( n33661 , n15777 , n32822 );
or ( n33662 , n33656 , n33660 , n33661 );
buf ( n33663 , n33662 );
and ( n33664 , n33652 , n33663 );
not ( n33665 , n33663 );
and ( n33666 , n33641 , n33642 );
xor ( n33667 , n33665 , n33666 );
and ( n33668 , n33667 , n33579 );
or ( n33669 , n33664 , n33668 );
buf ( n33670 , n33669 );
not ( n33671 , n33670 );
buf ( n33672 , n33671 );
buf ( n33673 , n33672 );
not ( n33674 , n33673 );
or ( n33675 , n33651 , n33674 );
not ( n33676 , n33579 );
xor ( n33677 , n33119 , n33128 );
xor ( n33678 , n33677 , n33211 );
buf ( n33679 , n33678 );
and ( n33680 , n33679 , n14143 );
xor ( n33681 , n33461 , n33463 );
xor ( n33682 , n33681 , n33518 );
buf ( n33683 , n33682 );
and ( n33684 , n33683 , n14141 );
and ( n33685 , n15755 , n32822 );
or ( n33686 , n33680 , n33684 , n33685 );
buf ( n33687 , n33686 );
and ( n33688 , n33676 , n33687 );
not ( n33689 , n33687 );
and ( n33690 , n33665 , n33666 );
xor ( n33691 , n33689 , n33690 );
and ( n33692 , n33691 , n33579 );
or ( n33693 , n33688 , n33692 );
buf ( n33694 , n33693 );
not ( n33695 , n33694 );
buf ( n33696 , n33695 );
buf ( n33697 , n33696 );
not ( n33698 , n33697 );
or ( n33699 , n33675 , n33698 );
not ( n33700 , n33579 );
xor ( n33701 , n33102 , n33111 );
xor ( n33702 , n33701 , n33214 );
buf ( n33703 , n33702 );
and ( n33704 , n33703 , n14143 );
xor ( n33705 , n33451 , n33453 );
xor ( n33706 , n33705 , n33521 );
buf ( n33707 , n33706 );
and ( n33708 , n33707 , n14141 );
and ( n33709 , n15733 , n32822 );
or ( n33710 , n33704 , n33708 , n33709 );
buf ( n33711 , n33710 );
and ( n33712 , n33700 , n33711 );
not ( n33713 , n33711 );
and ( n33714 , n33689 , n33690 );
xor ( n33715 , n33713 , n33714 );
and ( n33716 , n33715 , n33579 );
or ( n33717 , n33712 , n33716 );
buf ( n33718 , n33717 );
not ( n33719 , n33718 );
buf ( n33720 , n33719 );
buf ( n33721 , n33720 );
not ( n33722 , n33721 );
or ( n33723 , n33699 , n33722 );
not ( n33724 , n33579 );
xor ( n33725 , n33085 , n33094 );
xor ( n33726 , n33725 , n33217 );
buf ( n33727 , n33726 );
and ( n33728 , n33727 , n14143 );
xor ( n33729 , n33441 , n33443 );
xor ( n33730 , n33729 , n33524 );
buf ( n33731 , n33730 );
and ( n33732 , n33731 , n14141 );
and ( n33733 , n15711 , n32822 );
or ( n33734 , n33728 , n33732 , n33733 );
buf ( n33735 , n33734 );
and ( n33736 , n33724 , n33735 );
not ( n33737 , n33735 );
and ( n33738 , n33713 , n33714 );
xor ( n33739 , n33737 , n33738 );
and ( n33740 , n33739 , n33579 );
or ( n33741 , n33736 , n33740 );
buf ( n33742 , n33741 );
not ( n33743 , n33742 );
buf ( n33744 , n33743 );
buf ( n33745 , n33744 );
not ( n33746 , n33745 );
or ( n33747 , n33723 , n33746 );
not ( n33748 , n33579 );
xor ( n33749 , n33068 , n33077 );
xor ( n33750 , n33749 , n33220 );
buf ( n33751 , n33750 );
and ( n33752 , n33751 , n14143 );
xor ( n33753 , n33431 , n33433 );
xor ( n33754 , n33753 , n33527 );
buf ( n33755 , n33754 );
and ( n33756 , n33755 , n14141 );
and ( n33757 , n15689 , n32822 );
or ( n33758 , n33752 , n33756 , n33757 );
buf ( n33759 , n33758 );
and ( n33760 , n33748 , n33759 );
not ( n33761 , n33759 );
and ( n33762 , n33737 , n33738 );
xor ( n33763 , n33761 , n33762 );
and ( n33764 , n33763 , n33579 );
or ( n33765 , n33760 , n33764 );
buf ( n33766 , n33765 );
not ( n33767 , n33766 );
buf ( n33768 , n33767 );
buf ( n33769 , n33768 );
not ( n33770 , n33769 );
or ( n33771 , n33747 , n33770 );
not ( n33772 , n33579 );
xor ( n33773 , n33051 , n33060 );
xor ( n33774 , n33773 , n33223 );
buf ( n33775 , n33774 );
and ( n33776 , n33775 , n14143 );
xor ( n33777 , n33421 , n33423 );
xor ( n33778 , n33777 , n33530 );
buf ( n33779 , n33778 );
and ( n33780 , n33779 , n14141 );
and ( n33781 , n15667 , n32822 );
or ( n33782 , n33776 , n33780 , n33781 );
buf ( n33783 , n33782 );
and ( n33784 , n33772 , n33783 );
not ( n33785 , n33783 );
and ( n33786 , n33761 , n33762 );
xor ( n33787 , n33785 , n33786 );
and ( n33788 , n33787 , n33579 );
or ( n33789 , n33784 , n33788 );
buf ( n33790 , n33789 );
not ( n33791 , n33790 );
buf ( n33792 , n33791 );
buf ( n33793 , n33792 );
not ( n33794 , n33793 );
or ( n33795 , n33771 , n33794 );
not ( n33796 , n33579 );
xor ( n33797 , n33034 , n33043 );
xor ( n33798 , n33797 , n33226 );
buf ( n33799 , n33798 );
and ( n33800 , n33799 , n14143 );
xor ( n33801 , n33411 , n33413 );
xor ( n33802 , n33801 , n33533 );
buf ( n33803 , n33802 );
and ( n33804 , n33803 , n14141 );
and ( n33805 , n15645 , n32822 );
or ( n33806 , n33800 , n33804 , n33805 );
buf ( n33807 , n33806 );
and ( n33808 , n33796 , n33807 );
not ( n33809 , n33807 );
and ( n33810 , n33785 , n33786 );
xor ( n33811 , n33809 , n33810 );
and ( n33812 , n33811 , n33579 );
or ( n33813 , n33808 , n33812 );
buf ( n33814 , n33813 );
not ( n33815 , n33814 );
buf ( n33816 , n33815 );
buf ( n33817 , n33816 );
not ( n33818 , n33817 );
or ( n33819 , n33795 , n33818 );
not ( n33820 , n33579 );
xor ( n33821 , n33017 , n33026 );
xor ( n33822 , n33821 , n33229 );
buf ( n33823 , n33822 );
and ( n33824 , n33823 , n14143 );
xor ( n33825 , n33401 , n33403 );
xor ( n33826 , n33825 , n33536 );
buf ( n33827 , n33826 );
and ( n33828 , n33827 , n14141 );
and ( n33829 , n15623 , n32822 );
or ( n33830 , n33824 , n33828 , n33829 );
buf ( n33831 , n33830 );
and ( n33832 , n33820 , n33831 );
not ( n33833 , n33831 );
and ( n33834 , n33809 , n33810 );
xor ( n33835 , n33833 , n33834 );
and ( n33836 , n33835 , n33579 );
or ( n33837 , n33832 , n33836 );
buf ( n33838 , n33837 );
not ( n33839 , n33838 );
buf ( n33840 , n33839 );
buf ( n33841 , n33840 );
not ( n33842 , n33841 );
or ( n33843 , n33819 , n33842 );
not ( n33844 , n33579 );
xor ( n33845 , n33000 , n33009 );
xor ( n33846 , n33845 , n33232 );
buf ( n33847 , n33846 );
and ( n33848 , n33847 , n14143 );
xor ( n33849 , n33391 , n33393 );
xor ( n33850 , n33849 , n33539 );
buf ( n33851 , n33850 );
and ( n33852 , n33851 , n14141 );
and ( n33853 , n15601 , n32822 );
or ( n33854 , n33848 , n33852 , n33853 );
buf ( n33855 , n33854 );
and ( n33856 , n33844 , n33855 );
not ( n33857 , n33855 );
and ( n33858 , n33833 , n33834 );
xor ( n33859 , n33857 , n33858 );
and ( n33860 , n33859 , n33579 );
or ( n33861 , n33856 , n33860 );
buf ( n33862 , n33861 );
not ( n33863 , n33862 );
buf ( n33864 , n33863 );
buf ( n33865 , n33864 );
not ( n33866 , n33865 );
or ( n33867 , n33843 , n33866 );
not ( n33868 , n33579 );
xor ( n33869 , n32983 , n32992 );
xor ( n33870 , n33869 , n33235 );
buf ( n33871 , n33870 );
and ( n33872 , n33871 , n14143 );
xor ( n33873 , n33381 , n33383 );
xor ( n33874 , n33873 , n33542 );
buf ( n33875 , n33874 );
and ( n33876 , n33875 , n14141 );
and ( n33877 , n15579 , n32822 );
or ( n33878 , n33872 , n33876 , n33877 );
buf ( n33879 , n33878 );
and ( n33880 , n33868 , n33879 );
not ( n33881 , n33879 );
and ( n33882 , n33857 , n33858 );
xor ( n33883 , n33881 , n33882 );
and ( n33884 , n33883 , n33579 );
or ( n33885 , n33880 , n33884 );
buf ( n33886 , n33885 );
not ( n33887 , n33886 );
buf ( n33888 , n33887 );
buf ( n33889 , n33888 );
not ( n33890 , n33889 );
or ( n33891 , n33867 , n33890 );
not ( n33892 , n33579 );
xor ( n33893 , n32966 , n32975 );
xor ( n33894 , n33893 , n33238 );
buf ( n33895 , n33894 );
and ( n33896 , n33895 , n14143 );
xor ( n33897 , n33371 , n33373 );
xor ( n33898 , n33897 , n33545 );
buf ( n33899 , n33898 );
and ( n33900 , n33899 , n14141 );
and ( n33901 , n15557 , n32822 );
or ( n33902 , n33896 , n33900 , n33901 );
buf ( n33903 , n33902 );
and ( n33904 , n33892 , n33903 );
not ( n33905 , n33903 );
and ( n33906 , n33881 , n33882 );
xor ( n33907 , n33905 , n33906 );
and ( n33908 , n33907 , n33579 );
or ( n33909 , n33904 , n33908 );
buf ( n33910 , n33909 );
not ( n33911 , n33910 );
buf ( n33912 , n33911 );
buf ( n33913 , n33912 );
not ( n33914 , n33913 );
or ( n33915 , n33891 , n33914 );
not ( n33916 , n33579 );
xor ( n33917 , n32949 , n32958 );
xor ( n33918 , n33917 , n33241 );
buf ( n33919 , n33918 );
and ( n33920 , n33919 , n14143 );
xor ( n33921 , n33361 , n33363 );
xor ( n33922 , n33921 , n33548 );
buf ( n33923 , n33922 );
and ( n33924 , n33923 , n14141 );
and ( n33925 , n15535 , n32822 );
or ( n33926 , n33920 , n33924 , n33925 );
buf ( n33927 , n33926 );
and ( n33928 , n33916 , n33927 );
not ( n33929 , n33927 );
and ( n33930 , n33905 , n33906 );
xor ( n33931 , n33929 , n33930 );
and ( n33932 , n33931 , n33579 );
or ( n33933 , n33928 , n33932 );
buf ( n33934 , n33933 );
not ( n33935 , n33934 );
buf ( n33936 , n33935 );
buf ( n33937 , n33936 );
not ( n33938 , n33937 );
or ( n33939 , n33915 , n33938 );
not ( n33940 , n33579 );
xor ( n33941 , n32932 , n32941 );
xor ( n33942 , n33941 , n33244 );
buf ( n33943 , n33942 );
and ( n33944 , n33943 , n14143 );
xor ( n33945 , n33351 , n33353 );
xor ( n33946 , n33945 , n33551 );
buf ( n33947 , n33946 );
and ( n33948 , n33947 , n14141 );
and ( n33949 , n15513 , n32822 );
or ( n33950 , n33944 , n33948 , n33949 );
buf ( n33951 , n33950 );
and ( n33952 , n33940 , n33951 );
not ( n33953 , n33951 );
and ( n33954 , n33929 , n33930 );
xor ( n33955 , n33953 , n33954 );
and ( n33956 , n33955 , n33579 );
or ( n33957 , n33952 , n33956 );
buf ( n33958 , n33957 );
not ( n33959 , n33958 );
buf ( n33960 , n33959 );
buf ( n33961 , n33960 );
not ( n33962 , n33961 );
or ( n33963 , n33939 , n33962 );
not ( n33964 , n33579 );
xor ( n33965 , n32915 , n32924 );
xor ( n33966 , n33965 , n33247 );
buf ( n33967 , n33966 );
and ( n33968 , n33967 , n14143 );
xor ( n33969 , n33341 , n33343 );
xor ( n33970 , n33969 , n33554 );
buf ( n33971 , n33970 );
and ( n33972 , n33971 , n14141 );
and ( n33973 , n15491 , n32822 );
or ( n33974 , n33968 , n33972 , n33973 );
buf ( n33975 , n33974 );
and ( n33976 , n33964 , n33975 );
not ( n33977 , n33975 );
and ( n33978 , n33953 , n33954 );
xor ( n33979 , n33977 , n33978 );
and ( n33980 , n33979 , n33579 );
or ( n33981 , n33976 , n33980 );
buf ( n33982 , n33981 );
not ( n33983 , n33982 );
buf ( n33984 , n33983 );
buf ( n33985 , n33984 );
not ( n33986 , n33985 );
or ( n33987 , n33963 , n33986 );
not ( n33988 , n33579 );
xor ( n33989 , n32898 , n32907 );
xor ( n33990 , n33989 , n33250 );
buf ( n33991 , n33990 );
and ( n33992 , n33991 , n14143 );
xor ( n33993 , n33331 , n33333 );
xor ( n33994 , n33993 , n33557 );
buf ( n33995 , n33994 );
and ( n33996 , n33995 , n14141 );
and ( n33997 , n15469 , n32822 );
or ( n33998 , n33992 , n33996 , n33997 );
buf ( n33999 , n33998 );
and ( n34000 , n33988 , n33999 );
not ( n34001 , n33999 );
and ( n34002 , n33977 , n33978 );
xor ( n34003 , n34001 , n34002 );
and ( n34004 , n34003 , n33579 );
or ( n34005 , n34000 , n34004 );
buf ( n34006 , n34005 );
not ( n34007 , n34006 );
buf ( n34008 , n34007 );
buf ( n34009 , n34008 );
not ( n34010 , n34009 );
or ( n34011 , n33987 , n34010 );
not ( n34012 , n33579 );
xor ( n34013 , n32881 , n32890 );
xor ( n34014 , n34013 , n33253 );
buf ( n34015 , n34014 );
and ( n34016 , n34015 , n14143 );
xor ( n34017 , n33321 , n33323 );
xor ( n34018 , n34017 , n33560 );
buf ( n34019 , n34018 );
and ( n34020 , n34019 , n14141 );
and ( n34021 , n15447 , n32822 );
or ( n34022 , n34016 , n34020 , n34021 );
buf ( n34023 , n34022 );
and ( n34024 , n34012 , n34023 );
not ( n34025 , n34023 );
and ( n34026 , n34001 , n34002 );
xor ( n34027 , n34025 , n34026 );
and ( n34028 , n34027 , n33579 );
or ( n34029 , n34024 , n34028 );
buf ( n34030 , n34029 );
not ( n34031 , n34030 );
buf ( n34032 , n34031 );
buf ( n34033 , n34032 );
not ( n34034 , n34033 );
or ( n34035 , n34011 , n34034 );
buf ( n34036 , n34035 );
buf ( n34037 , n34036 );
and ( n34038 , n34037 , n33579 );
not ( n34039 , n34038 );
and ( n34040 , n34039 , n32830 );
xor ( n34041 , n32830 , n33579 );
xor ( n34042 , n34041 , n33579 );
and ( n34043 , n34042 , n34038 );
or ( n34044 , n34040 , n34043 );
buf ( n34045 , n34044 );
and ( n34046 , n34045 , n12243 );
or ( n34047 , n32239 , n34046 );
and ( n34048 , n31185 , n34047 );
and ( n34049 , n32225 , n11954 );
or ( n34050 , n34048 , n34049 );
and ( n34051 , n34050 , n16574 );
buf ( n34052 , n12333 );
buf ( n34053 , n34052 );
not ( n34054 , n34053 );
buf ( n34055 , n34054 );
buf ( n34056 , n34055 );
not ( n34057 , n34056 );
buf ( n34058 , n12245 );
not ( n34059 , n34058 );
buf ( n34060 , n12330 );
and ( n34061 , n34059 , n34060 );
not ( n34062 , n34060 );
not ( n34063 , n34052 );
xor ( n34064 , n34062 , n34063 );
and ( n34065 , n34064 , n34058 );
or ( n34066 , n34061 , n34065 );
buf ( n34067 , n34066 );
not ( n34068 , n34067 );
buf ( n34069 , n34068 );
buf ( n34070 , n34069 );
not ( n34071 , n34070 );
or ( n34072 , n34057 , n34071 );
not ( n34073 , n34058 );
buf ( n34074 , n12327 );
and ( n34075 , n34073 , n34074 );
not ( n34076 , n34074 );
and ( n34077 , n34062 , n34063 );
xor ( n34078 , n34076 , n34077 );
and ( n34079 , n34078 , n34058 );
or ( n34080 , n34075 , n34079 );
buf ( n34081 , n34080 );
not ( n34082 , n34081 );
buf ( n34083 , n34082 );
buf ( n34084 , n34083 );
not ( n34085 , n34084 );
or ( n34086 , n34072 , n34085 );
not ( n34087 , n34058 );
buf ( n34088 , n12324 );
and ( n34089 , n34087 , n34088 );
not ( n34090 , n34088 );
and ( n34091 , n34076 , n34077 );
xor ( n34092 , n34090 , n34091 );
and ( n34093 , n34092 , n34058 );
or ( n34094 , n34089 , n34093 );
buf ( n34095 , n34094 );
not ( n34096 , n34095 );
buf ( n34097 , n34096 );
buf ( n34098 , n34097 );
not ( n34099 , n34098 );
or ( n34100 , n34086 , n34099 );
not ( n34101 , n34058 );
buf ( n34102 , n12321 );
and ( n34103 , n34101 , n34102 );
not ( n34104 , n34102 );
and ( n34105 , n34090 , n34091 );
xor ( n34106 , n34104 , n34105 );
and ( n34107 , n34106 , n34058 );
or ( n34108 , n34103 , n34107 );
buf ( n34109 , n34108 );
not ( n34110 , n34109 );
buf ( n34111 , n34110 );
buf ( n34112 , n34111 );
not ( n34113 , n34112 );
or ( n34114 , n34100 , n34113 );
not ( n34115 , n34058 );
buf ( n34116 , n12318 );
and ( n34117 , n34115 , n34116 );
not ( n34118 , n34116 );
and ( n34119 , n34104 , n34105 );
xor ( n34120 , n34118 , n34119 );
and ( n34121 , n34120 , n34058 );
or ( n34122 , n34117 , n34121 );
buf ( n34123 , n34122 );
not ( n34124 , n34123 );
buf ( n34125 , n34124 );
buf ( n34126 , n34125 );
not ( n34127 , n34126 );
or ( n34128 , n34114 , n34127 );
not ( n34129 , n34058 );
buf ( n34130 , n12315 );
and ( n34131 , n34129 , n34130 );
not ( n34132 , n34130 );
and ( n34133 , n34118 , n34119 );
xor ( n34134 , n34132 , n34133 );
and ( n34135 , n34134 , n34058 );
or ( n34136 , n34131 , n34135 );
buf ( n34137 , n34136 );
not ( n34138 , n34137 );
buf ( n34139 , n34138 );
buf ( n34140 , n34139 );
not ( n34141 , n34140 );
or ( n34142 , n34128 , n34141 );
not ( n34143 , n34058 );
buf ( n34144 , n12312 );
and ( n34145 , n34143 , n34144 );
not ( n34146 , n34144 );
and ( n34147 , n34132 , n34133 );
xor ( n34148 , n34146 , n34147 );
and ( n34149 , n34148 , n34058 );
or ( n34150 , n34145 , n34149 );
buf ( n34151 , n34150 );
not ( n34152 , n34151 );
buf ( n34153 , n34152 );
buf ( n34154 , n34153 );
not ( n34155 , n34154 );
or ( n34156 , n34142 , n34155 );
not ( n34157 , n34058 );
buf ( n34158 , n12309 );
and ( n34159 , n34157 , n34158 );
not ( n34160 , n34158 );
and ( n34161 , n34146 , n34147 );
xor ( n34162 , n34160 , n34161 );
and ( n34163 , n34162 , n34058 );
or ( n34164 , n34159 , n34163 );
buf ( n34165 , n34164 );
not ( n34166 , n34165 );
buf ( n34167 , n34166 );
buf ( n34168 , n34167 );
not ( n34169 , n34168 );
or ( n34170 , n34156 , n34169 );
not ( n34171 , n34058 );
buf ( n34172 , n12306 );
and ( n34173 , n34171 , n34172 );
not ( n34174 , n34172 );
and ( n34175 , n34160 , n34161 );
xor ( n34176 , n34174 , n34175 );
and ( n34177 , n34176 , n34058 );
or ( n34178 , n34173 , n34177 );
buf ( n34179 , n34178 );
not ( n34180 , n34179 );
buf ( n34181 , n34180 );
buf ( n34182 , n34181 );
not ( n34183 , n34182 );
or ( n34184 , n34170 , n34183 );
not ( n34185 , n34058 );
buf ( n34186 , n12303 );
and ( n34187 , n34185 , n34186 );
not ( n34188 , n34186 );
and ( n34189 , n34174 , n34175 );
xor ( n34190 , n34188 , n34189 );
and ( n34191 , n34190 , n34058 );
or ( n34192 , n34187 , n34191 );
buf ( n34193 , n34192 );
not ( n34194 , n34193 );
buf ( n34195 , n34194 );
buf ( n34196 , n34195 );
not ( n34197 , n34196 );
or ( n34198 , n34184 , n34197 );
not ( n34199 , n34058 );
buf ( n34200 , n12300 );
and ( n34201 , n34199 , n34200 );
not ( n34202 , n34200 );
and ( n34203 , n34188 , n34189 );
xor ( n34204 , n34202 , n34203 );
and ( n34205 , n34204 , n34058 );
or ( n34206 , n34201 , n34205 );
buf ( n34207 , n34206 );
not ( n34208 , n34207 );
buf ( n34209 , n34208 );
buf ( n34210 , n34209 );
not ( n34211 , n34210 );
or ( n34212 , n34198 , n34211 );
not ( n34213 , n34058 );
buf ( n34214 , n12297 );
and ( n34215 , n34213 , n34214 );
not ( n34216 , n34214 );
and ( n34217 , n34202 , n34203 );
xor ( n34218 , n34216 , n34217 );
and ( n34219 , n34218 , n34058 );
or ( n34220 , n34215 , n34219 );
buf ( n34221 , n34220 );
not ( n34222 , n34221 );
buf ( n34223 , n34222 );
buf ( n34224 , n34223 );
not ( n34225 , n34224 );
or ( n34226 , n34212 , n34225 );
not ( n34227 , n34058 );
buf ( n34228 , n12294 );
and ( n34229 , n34227 , n34228 );
not ( n34230 , n34228 );
and ( n34231 , n34216 , n34217 );
xor ( n34232 , n34230 , n34231 );
and ( n34233 , n34232 , n34058 );
or ( n34234 , n34229 , n34233 );
buf ( n34235 , n34234 );
not ( n34236 , n34235 );
buf ( n34237 , n34236 );
buf ( n34238 , n34237 );
not ( n34239 , n34238 );
or ( n34240 , n34226 , n34239 );
not ( n34241 , n34058 );
buf ( n34242 , n12291 );
and ( n34243 , n34241 , n34242 );
not ( n34244 , n34242 );
and ( n34245 , n34230 , n34231 );
xor ( n34246 , n34244 , n34245 );
and ( n34247 , n34246 , n34058 );
or ( n34248 , n34243 , n34247 );
buf ( n34249 , n34248 );
not ( n34250 , n34249 );
buf ( n34251 , n34250 );
buf ( n34252 , n34251 );
not ( n34253 , n34252 );
or ( n34254 , n34240 , n34253 );
not ( n34255 , n34058 );
buf ( n34256 , n12288 );
and ( n34257 , n34255 , n34256 );
not ( n34258 , n34256 );
and ( n34259 , n34244 , n34245 );
xor ( n34260 , n34258 , n34259 );
and ( n34261 , n34260 , n34058 );
or ( n34262 , n34257 , n34261 );
buf ( n34263 , n34262 );
not ( n34264 , n34263 );
buf ( n34265 , n34264 );
buf ( n34266 , n34265 );
not ( n34267 , n34266 );
or ( n34268 , n34254 , n34267 );
not ( n34269 , n34058 );
buf ( n34270 , n12285 );
and ( n34271 , n34269 , n34270 );
not ( n34272 , n34270 );
and ( n34273 , n34258 , n34259 );
xor ( n34274 , n34272 , n34273 );
and ( n34275 , n34274 , n34058 );
or ( n34276 , n34271 , n34275 );
buf ( n34277 , n34276 );
not ( n34278 , n34277 );
buf ( n34279 , n34278 );
buf ( n34280 , n34279 );
not ( n34281 , n34280 );
or ( n34282 , n34268 , n34281 );
not ( n34283 , n34058 );
buf ( n34284 , n12282 );
and ( n34285 , n34283 , n34284 );
not ( n34286 , n34284 );
and ( n34287 , n34272 , n34273 );
xor ( n34288 , n34286 , n34287 );
and ( n34289 , n34288 , n34058 );
or ( n34290 , n34285 , n34289 );
buf ( n34291 , n34290 );
not ( n34292 , n34291 );
buf ( n34293 , n34292 );
buf ( n34294 , n34293 );
not ( n34295 , n34294 );
or ( n34296 , n34282 , n34295 );
not ( n34297 , n34058 );
buf ( n34298 , n12279 );
and ( n34299 , n34297 , n34298 );
not ( n34300 , n34298 );
and ( n34301 , n34286 , n34287 );
xor ( n34302 , n34300 , n34301 );
and ( n34303 , n34302 , n34058 );
or ( n34304 , n34299 , n34303 );
buf ( n34305 , n34304 );
not ( n34306 , n34305 );
buf ( n34307 , n34306 );
buf ( n34308 , n34307 );
not ( n34309 , n34308 );
or ( n34310 , n34296 , n34309 );
not ( n34311 , n34058 );
buf ( n34312 , n12276 );
and ( n34313 , n34311 , n34312 );
not ( n34314 , n34312 );
and ( n34315 , n34300 , n34301 );
xor ( n34316 , n34314 , n34315 );
and ( n34317 , n34316 , n34058 );
or ( n34318 , n34313 , n34317 );
buf ( n34319 , n34318 );
not ( n34320 , n34319 );
buf ( n34321 , n34320 );
buf ( n34322 , n34321 );
not ( n34323 , n34322 );
or ( n34324 , n34310 , n34323 );
buf ( n34325 , n34324 );
buf ( n34326 , n34325 );
and ( n34327 , n34326 , n34058 );
not ( n34328 , n34327 );
and ( n34329 , n34328 , n34057 );
xor ( n34330 , n34057 , n34058 );
xor ( n34331 , n34330 , n34058 );
and ( n34332 , n34331 , n34327 );
or ( n34333 , n34329 , n34332 );
buf ( n34334 , n34333 );
and ( n34335 , n34334 , n16576 );
or ( n34336 , n34051 , n34335 );
buf ( n34337 , n34336 );
buf ( n34338 , n34337 );
not ( n34339 , n17451 );
and ( n34340 , n18504 , n17873 );
not ( n34341 , n19750 );
and ( n34342 , n34341 , n20459 );
not ( n34343 , n21193 );
and ( n34344 , n34343 , n20465 );
xor ( n34345 , n21221 , n20582 );
and ( n34346 , n34345 , n21193 );
or ( n34347 , n34344 , n34346 );
buf ( n34348 , n34347 );
and ( n34349 , n34348 , n19750 );
or ( n34350 , n34342 , n34349 );
and ( n34351 , n34350 , n21253 );
and ( n34352 , n20459 , n21255 );
or ( n34353 , C0 , C0 , n34351 , n34352 );
and ( n34354 , n34353 , n21330 );
and ( n34355 , n18504 , n21338 );
or ( n34356 , n34354 , n34355 );
and ( n34357 , n34356 , n21341 );
not ( n34358 , n22996 );
and ( n34359 , n34358 , n21648 );
xor ( n34360 , n23024 , n22500 );
and ( n34361 , n34360 , n22996 );
or ( n34362 , n34359 , n34361 );
buf ( n34363 , n34362 );
and ( n34364 , n34363 , n21330 );
and ( n34365 , n18504 , n21338 );
or ( n34366 , n34364 , n34365 );
and ( n34367 , n34366 , n23064 );
not ( n34368 , n23758 );
and ( n34369 , n34368 , n23075 );
xor ( n34370 , n23786 , n23262 );
and ( n34371 , n34370 , n23758 );
or ( n34372 , n34369 , n34371 );
buf ( n34373 , n34372 );
and ( n34374 , n34373 , n21330 );
and ( n34375 , n18504 , n21338 );
or ( n34376 , n34374 , n34375 );
and ( n34377 , n34376 , n23825 );
and ( n34378 , n21639 , n21330 );
and ( n34379 , n18504 , n21338 );
or ( n34380 , n34378 , n34379 );
and ( n34381 , n34380 , n23832 );
and ( n34382 , n18314 , n23834 );
buf ( n34383 , n23886 );
and ( n34384 , n34383 , n21330 );
and ( n34385 , n18504 , n21338 );
or ( n34386 , n34384 , n34385 );
and ( n34387 , n34386 , n23917 );
or ( n34388 , n34340 , n34357 , n34367 , n34377 , n34381 , n34382 , n34387 );
and ( n34389 , n34339 , n34388 );
and ( n34390 , n18504 , n17451 );
or ( n34391 , n34389 , n34390 );
and ( n34392 , n34391 , n23924 );
and ( n34393 , n18504 , n23926 );
or ( n34394 , n34392 , n34393 );
buf ( n34395 , n34394 );
buf ( n34396 , n34395 );
buf ( n34397 , n10613 );
buf ( n34398 , n10613 );
not ( n34399 , n17451 );
and ( n34400 , n19215 , n17873 );
not ( n34401 , n19474 );
and ( n34402 , n34401 , n19199 );
xor ( n34403 , n19481 , n19521 );
and ( n34404 , n34403 , n19474 );
or ( n34405 , n34402 , n34404 );
buf ( n34406 , n34405 );
and ( n34407 , n34406 , n19745 );
and ( n34408 , n34406 , n19748 );
not ( n34409 , n19750 );
and ( n34410 , n34409 , n21031 );
not ( n34411 , n21193 );
and ( n34412 , n34411 , n21043 );
xor ( n34413 , n21200 , n21242 );
and ( n34414 , n34413 , n21193 );
or ( n34415 , n34412 , n34414 );
buf ( n34416 , n34415 );
and ( n34417 , n34416 , n19750 );
or ( n34418 , n34410 , n34417 );
and ( n34419 , n34418 , n21253 );
and ( n34420 , n21031 , n21255 );
or ( n34421 , n34407 , n34408 , n34419 , n34420 );
and ( n34422 , n34421 , n21330 );
and ( n34423 , n19215 , n21338 );
or ( n34424 , n34422 , n34423 );
and ( n34425 , n34424 , n21341 );
not ( n34426 , n22996 );
and ( n34427 , n34426 , n22856 );
xor ( n34428 , n23003 , n23045 );
and ( n34429 , n34428 , n22996 );
or ( n34430 , n34427 , n34429 );
buf ( n34431 , n34430 );
and ( n34432 , n34431 , n21330 );
and ( n34433 , n19215 , n21338 );
or ( n34434 , n34432 , n34433 );
and ( n34435 , n34434 , n23064 );
not ( n34436 , n23758 );
and ( n34437 , n34436 , n23618 );
xor ( n34438 , n23765 , n23807 );
and ( n34439 , n34438 , n23758 );
or ( n34440 , n34437 , n34439 );
buf ( n34441 , n34440 );
and ( n34442 , n34441 , n21330 );
and ( n34443 , n19215 , n21338 );
or ( n34444 , n34442 , n34443 );
and ( n34445 , n34444 , n23825 );
and ( n34446 , n21971 , n21330 );
and ( n34447 , n19215 , n21338 );
or ( n34448 , n34446 , n34447 );
and ( n34449 , n34448 , n23832 );
and ( n34450 , n19213 , n23834 );
xor ( n34451 , n23845 , n23907 );
buf ( n34452 , n34451 );
and ( n34453 , n34452 , n21330 );
and ( n34454 , n19215 , n21338 );
or ( n34455 , n34453 , n34454 );
and ( n34456 , n34455 , n23917 );
or ( n34457 , n34400 , n34425 , n34435 , n34445 , n34449 , n34450 , n34456 );
and ( n34458 , n34399 , n34457 );
and ( n34459 , n19215 , n17451 );
or ( n34460 , n34458 , n34459 );
and ( n34461 , n34460 , n23924 );
and ( n34462 , n19215 , n23926 );
or ( n34463 , n34461 , n34462 );
buf ( n34464 , n34463 );
buf ( n34465 , n34464 );
buf ( n34466 , n10615 );
not ( n34467 , n17451 );
not ( n34468 , n19474 );
and ( n34469 , n34468 , n18825 );
xor ( n34470 , n19492 , n19510 );
and ( n34471 , n34470 , n19474 );
or ( n34472 , n34469 , n34471 );
buf ( n34473 , n34472 );
and ( n34474 , n34473 , n19745 );
and ( n34475 , n34473 , n19748 );
not ( n34476 , n19750 );
and ( n34477 , n34476 , n20789 );
not ( n34478 , n21193 );
and ( n34479 , n34478 , n20801 );
xor ( n34480 , n21211 , n21231 );
and ( n34481 , n34480 , n21193 );
or ( n34482 , n34479 , n34481 );
buf ( n34483 , n34482 );
and ( n34484 , n34483 , n19750 );
or ( n34485 , n34477 , n34484 );
and ( n34486 , n34485 , n21253 );
and ( n34487 , n20789 , n21255 );
or ( n34488 , n34474 , n34475 , n34486 , n34487 );
and ( n34489 , n34488 , n21334 );
or ( n34490 , n21333 , n21330 );
or ( n34491 , n34490 , n21336 );
or ( n34492 , n34491 , C0 );
and ( n34493 , n18845 , n34492 );
or ( n34494 , n34489 , n34493 );
and ( n34495 , n34494 , n21341 );
not ( n34496 , n22996 );
and ( n34497 , n34496 , n22669 );
xor ( n34498 , n23014 , n23034 );
and ( n34499 , n34498 , n22996 );
or ( n34500 , n34497 , n34499 );
buf ( n34501 , n34500 );
and ( n34502 , n34501 , n21334 );
and ( n34503 , n18845 , n34492 );
or ( n34504 , n34502 , n34503 );
and ( n34505 , n34504 , n23064 );
not ( n34506 , n23758 );
and ( n34507 , n34506 , n23431 );
xor ( n34508 , n23776 , n23796 );
and ( n34509 , n34508 , n23758 );
or ( n34510 , n34507 , n34509 );
buf ( n34511 , n34510 );
and ( n34512 , n34511 , n21334 );
and ( n34513 , n18845 , n34492 );
or ( n34514 , n34512 , n34513 );
and ( n34515 , n34514 , n23825 );
and ( n34516 , n22222 , n21334 );
and ( n34517 , n18845 , n34492 );
or ( n34518 , n34516 , n34517 );
and ( n34519 , n34518 , n23832 );
xor ( n34520 , n23867 , n23896 );
buf ( n34521 , n34520 );
and ( n34522 , n34521 , n21334 );
and ( n34523 , n18845 , n34492 );
or ( n34524 , n34522 , n34523 );
and ( n34525 , n34524 , n23917 );
or ( n34526 , n23834 , n17873 );
and ( n34527 , n18845 , n34526 );
or ( n34528 , n34495 , n34505 , n34515 , n34519 , n34525 , n34527 );
and ( n34529 , n34467 , n34528 );
and ( n34530 , n18845 , n17451 );
or ( n34531 , n34529 , n34530 );
and ( n34532 , n34531 , n23924 );
and ( n34533 , n18845 , n23926 );
or ( n34534 , n34532 , n34533 );
buf ( n34535 , n34534 );
buf ( n34536 , n34535 );
not ( n34537 , n17450 );
or ( n34538 , n17162 , n34537 );
not ( n34539 , n34538 );
and ( n34540 , n17450 , n34539 );
and ( n34541 , n34540 , n23924 );
buf ( n34542 , n34541 );
buf ( n34543 , n34542 );
buf ( n34544 , n10613 );
buf ( n34545 , n10615 );
buf ( n34546 , n10615 );
buf ( n34547 , n10615 );
not ( n34548 , n24800 );
not ( n34549 , n26823 );
and ( n34550 , n34549 , n25906 );
xor ( n34551 , n31026 , n31027 );
and ( n34552 , n34551 , n26823 );
or ( n34553 , n34550 , n34552 );
buf ( n34554 , n34553 );
and ( n34555 , n34554 , n27046 );
and ( n34556 , n34554 , n27049 );
not ( n34557 , n27051 );
and ( n34558 , n34557 , n27906 );
not ( n34559 , n28494 );
and ( n34560 , n34559 , n27918 );
xor ( n34561 , n31054 , n31055 );
and ( n34562 , n34561 , n28494 );
or ( n34563 , n34560 , n34562 );
buf ( n34564 , n34563 );
and ( n34565 , n34564 , n27051 );
or ( n34566 , n34558 , n34565 );
and ( n34567 , n34566 , n28506 );
and ( n34568 , n27906 , n28508 );
or ( n34569 , n34555 , n34556 , n34567 , n34568 );
and ( n34570 , n34569 , n28586 );
or ( n34571 , n28587 , n28583 );
or ( n34572 , n34571 , n28589 );
or ( n34573 , n34572 , C0 );
and ( n34574 , n25921 , n34573 );
or ( n34575 , n34570 , n34574 );
and ( n34576 , n34575 , n28594 );
not ( n34577 , n30249 );
and ( n34578 , n34577 , n29786 );
xor ( n34579 , n31089 , n31090 );
and ( n34580 , n34579 , n30249 );
or ( n34581 , n34578 , n34580 );
buf ( n34582 , n34581 );
and ( n34583 , n34582 , n28586 );
and ( n34584 , n25921 , n34573 );
or ( n34585 , n34583 , n34584 );
and ( n34586 , n34585 , n30269 );
not ( n34587 , n30963 );
and ( n34588 , n34587 , n30500 );
xor ( n34589 , n31117 , n31118 );
and ( n34590 , n34589 , n30963 );
or ( n34591 , n34588 , n34590 );
buf ( n34592 , n34591 );
and ( n34593 , n34592 , n28586 );
and ( n34594 , n25921 , n34573 );
or ( n34595 , n34593 , n34594 );
and ( n34596 , n34595 , n30982 );
and ( n34597 , n29635 , n28586 );
and ( n34598 , n25921 , n34573 );
or ( n34599 , n34597 , n34598 );
and ( n34600 , n34599 , n30989 );
xor ( n34601 , n31157 , n31158 );
buf ( n34602 , n34601 );
and ( n34603 , n34602 , n28586 );
and ( n34604 , n25921 , n34573 );
or ( n34605 , n34603 , n34604 );
and ( n34606 , n34605 , n31002 );
or ( n34607 , n30991 , n25222 );
and ( n34608 , n25921 , n34607 );
or ( n34609 , n34576 , n34586 , n34596 , n34600 , n34606 , n34608 );
and ( n34610 , n34548 , n34609 );
and ( n34611 , n25921 , n24800 );
or ( n34612 , n34610 , n34611 );
and ( n34613 , n34612 , n31008 );
and ( n34614 , n25921 , n10618 );
or ( n34615 , n34613 , n34614 );
buf ( n34616 , n34615 );
buf ( n34617 , n34616 );
buf ( n34618 , n10613 );
not ( n34619 , n24800 );
not ( n34620 , n26823 );
and ( n34621 , n34620 , n26309 );
xor ( n34622 , n26309 , n25877 );
xor ( n34623 , n26275 , n25877 );
xor ( n34624 , n26241 , n25877 );
xor ( n34625 , n26207 , n25877 );
and ( n34626 , n31018 , n31035 );
and ( n34627 , n34625 , n34626 );
and ( n34628 , n34624 , n34627 );
and ( n34629 , n34623 , n34628 );
xor ( n34630 , n34622 , n34629 );
and ( n34631 , n34630 , n26823 );
or ( n34632 , n34621 , n34631 );
buf ( n34633 , n34632 );
and ( n34634 , n34633 , n27046 );
and ( n34635 , n34633 , n27049 );
not ( n34636 , n27051 );
and ( n34637 , n34636 , n28170 );
not ( n34638 , n28494 );
and ( n34639 , n34638 , n28182 );
xor ( n34640 , n28182 , n27883 );
xor ( n34641 , n28160 , n27883 );
xor ( n34642 , n28138 , n27883 );
xor ( n34643 , n28116 , n27883 );
and ( n34644 , n31046 , n31063 );
and ( n34645 , n34643 , n34644 );
and ( n34646 , n34642 , n34645 );
and ( n34647 , n34641 , n34646 );
xor ( n34648 , n34640 , n34647 );
and ( n34649 , n34648 , n28494 );
or ( n34650 , n34639 , n34649 );
buf ( n34651 , n34650 );
and ( n34652 , n34651 , n27051 );
or ( n34653 , n34637 , n34652 );
and ( n34654 , n34653 , n28506 );
and ( n34655 , n28170 , n28508 );
or ( n34656 , n34634 , n34635 , n34654 , n34655 );
and ( n34657 , n34656 , n28586 );
and ( n34658 , n26327 , n34573 );
or ( n34659 , n34657 , n34658 );
and ( n34660 , n34659 , n28594 );
not ( n34661 , n30249 );
and ( n34662 , n34661 , n29990 );
xor ( n34663 , n29990 , n29753 );
xor ( n34664 , n29973 , n29753 );
xor ( n34665 , n29956 , n29753 );
xor ( n34666 , n29939 , n29753 );
and ( n34667 , n31081 , n31098 );
and ( n34668 , n34666 , n34667 );
and ( n34669 , n34665 , n34668 );
and ( n34670 , n34664 , n34669 );
xor ( n34671 , n34663 , n34670 );
and ( n34672 , n34671 , n30249 );
or ( n34673 , n34662 , n34672 );
buf ( n34674 , n34673 );
and ( n34675 , n34674 , n28586 );
and ( n34676 , n26327 , n34573 );
or ( n34677 , n34675 , n34676 );
and ( n34678 , n34677 , n30269 );
not ( n34679 , n30963 );
and ( n34680 , n34679 , n30704 );
xor ( n34681 , n30704 , n30467 );
xor ( n34682 , n30687 , n30467 );
xor ( n34683 , n30670 , n30467 );
xor ( n34684 , n30653 , n30467 );
and ( n34685 , n31109 , n31126 );
and ( n34686 , n34684 , n34685 );
and ( n34687 , n34683 , n34686 );
and ( n34688 , n34682 , n34687 );
xor ( n34689 , n34681 , n34688 );
and ( n34690 , n34689 , n30963 );
or ( n34691 , n34680 , n34690 );
buf ( n34692 , n34691 );
and ( n34693 , n34692 , n28586 );
and ( n34694 , n26327 , n34573 );
or ( n34695 , n34693 , n34694 );
and ( n34696 , n34695 , n30982 );
and ( n34697 , n29395 , n28586 );
and ( n34698 , n26327 , n34573 );
or ( n34699 , n34697 , n34698 );
and ( n34700 , n34699 , n30989 );
buf ( n34701 , n29395 );
not ( n34702 , n34701 );
buf ( n34703 , n29415 );
not ( n34704 , n34703 );
buf ( n34705 , n29435 );
not ( n34706 , n34705 );
buf ( n34707 , n29455 );
not ( n34708 , n34707 );
and ( n34709 , n31141 , n31166 );
and ( n34710 , n34708 , n34709 );
and ( n34711 , n34706 , n34710 );
and ( n34712 , n34704 , n34711 );
xor ( n34713 , n34702 , n34712 );
buf ( n34714 , n34713 );
and ( n34715 , n34714 , n28586 );
and ( n34716 , n26327 , n34573 );
or ( n34717 , n34715 , n34716 );
and ( n34718 , n34717 , n31002 );
and ( n34719 , n26327 , n34607 );
or ( n34720 , n34660 , n34678 , n34696 , n34700 , n34718 , n34719 );
and ( n34721 , n34619 , n34720 );
and ( n34722 , n26327 , n24800 );
or ( n34723 , n34721 , n34722 );
and ( n34724 , n34723 , n31008 );
and ( n34725 , n26327 , n10618 );
or ( n34726 , n34724 , n34725 );
buf ( n34727 , n34726 );
buf ( n34728 , n34727 );
buf ( n34729 , n10615 );
buf ( n34730 , n10613 );
buf ( n34731 , n10613 );
buf ( n34732 , n10613 );
not ( n34733 , n17451 );
not ( n34734 , n19474 );
and ( n34735 , n34734 , n18520 );
xor ( n34736 , n19501 , n18528 );
and ( n34737 , n34736 , n19474 );
or ( n34738 , n34735 , n34737 );
buf ( n34739 , n34738 );
and ( n34740 , n34739 , n19745 );
and ( n34741 , n34739 , n19748 );
not ( n34742 , n19750 );
and ( n34743 , n34742 , n20591 );
not ( n34744 , n21193 );
and ( n34745 , n34744 , n20603 );
xor ( n34746 , n21220 , n21222 );
and ( n34747 , n34746 , n21193 );
or ( n34748 , n34745 , n34747 );
buf ( n34749 , n34748 );
and ( n34750 , n34749 , n19750 );
or ( n34751 , n34743 , n34750 );
and ( n34752 , n34751 , n21253 );
and ( n34753 , n20591 , n21255 );
or ( n34754 , n34740 , n34741 , n34752 , n34753 );
and ( n34755 , n34754 , n21333 );
or ( n34756 , n21334 , n21330 );
or ( n34757 , n34756 , n21336 );
or ( n34758 , n34757 , C0 );
and ( n34759 , n18542 , n34758 );
or ( n34760 , n34755 , n34759 );
and ( n34761 , n34760 , n21341 );
not ( n34762 , n22996 );
and ( n34763 , n34762 , n22516 );
xor ( n34764 , n23023 , n23025 );
and ( n34765 , n34764 , n22996 );
or ( n34766 , n34763 , n34765 );
buf ( n34767 , n34766 );
and ( n34768 , n34767 , n21333 );
and ( n34769 , n18542 , n34758 );
or ( n34770 , n34768 , n34769 );
and ( n34771 , n34770 , n23064 );
not ( n34772 , n23758 );
and ( n34773 , n34772 , n23278 );
xor ( n34774 , n23785 , n23787 );
and ( n34775 , n34774 , n23758 );
or ( n34776 , n34773 , n34775 );
buf ( n34777 , n34776 );
and ( n34778 , n34777 , n21333 );
and ( n34779 , n18542 , n34758 );
or ( n34780 , n34778 , n34779 );
and ( n34781 , n34780 , n23825 );
and ( n34782 , n22402 , n21333 );
and ( n34783 , n18542 , n34758 );
or ( n34784 , n34782 , n34783 );
and ( n34785 , n34784 , n23832 );
xor ( n34786 , n23885 , n23887 );
buf ( n34787 , n34786 );
and ( n34788 , n34787 , n21333 );
and ( n34789 , n18542 , n34758 );
or ( n34790 , n34788 , n34789 );
and ( n34791 , n34790 , n23917 );
and ( n34792 , n18542 , n34526 );
or ( n34793 , n34761 , n34771 , n34781 , n34785 , n34791 , n34792 );
and ( n34794 , n34733 , n34793 );
and ( n34795 , n18542 , n17451 );
or ( n34796 , n34794 , n34795 );
and ( n34797 , n34796 , n23924 );
and ( n34798 , n18542 , n23926 );
or ( n34799 , n34797 , n34798 );
buf ( n34800 , n34799 );
buf ( n34801 , n34800 );
buf ( n34802 , n10613 );
not ( n34803 , n24799 );
or ( n34804 , n24511 , n34803 );
not ( n34805 , n34804 );
and ( n34806 , n34805 , n26569 );
and ( n34807 , n14707 , n34804 );
or ( n34808 , n34806 , n34807 );
and ( n34809 , n34808 , n31008 );
and ( n34810 , n14707 , n10618 );
or ( n34811 , n34809 , n34810 );
buf ( n34812 , n34811 );
buf ( n34813 , n34812 );
buf ( n34814 , n10615 );
buf ( n34815 , n10613 );
buf ( n34816 , n10615 );
buf ( n34817 , n10613 );
buf ( n34818 , n10613 );
buf ( n34819 , n10613 );
buf ( n34820 , n10615 );
or ( n34821 , n11954 , n12243 );
not ( n34822 , n34821 );
not ( n34823 , n13916 );
and ( n34824 , n34823 , n13793 );
xor ( n34825 , n13794 , n13861 );
and ( n34826 , n34825 , n13916 );
or ( n34827 , n34824 , n34826 );
buf ( n34828 , n34827 );
and ( n34829 , n34828 , n14137 );
and ( n34830 , n34828 , n14143 );
not ( n34831 , n14139 );
buf ( n34832 , n13150 );
buf ( n34833 , n34832 );
not ( n34834 , n34833 );
not ( n34835 , n34832 );
buf ( n34836 , n13403 );
and ( n34837 , n34835 , n34836 );
not ( n34838 , n34836 );
buf ( n34839 , n13415 );
not ( n34840 , n34839 );
buf ( n34841 , n13427 );
not ( n34842 , n34841 );
buf ( n34843 , n13439 );
not ( n34844 , n34843 );
buf ( n34845 , n13451 );
not ( n34846 , n34845 );
buf ( n34847 , n13463 );
not ( n34848 , n34847 );
buf ( n34849 , n13480 );
not ( n34850 , n34849 );
buf ( n34851 , n13497 );
not ( n34852 , n34851 );
buf ( n34853 , n13514 );
not ( n34854 , n34853 );
and ( n34855 , n34852 , n34854 );
and ( n34856 , n34850 , n34855 );
and ( n34857 , n34848 , n34856 );
and ( n34858 , n34846 , n34857 );
and ( n34859 , n34844 , n34858 );
and ( n34860 , n34842 , n34859 );
and ( n34861 , n34840 , n34860 );
xor ( n34862 , n34838 , n34861 );
and ( n34863 , n34862 , n34832 );
or ( n34864 , n34837 , n34863 );
buf ( n34865 , n34864 );
not ( n34866 , n34865 );
buf ( n34867 , n34866 );
buf ( n34868 , n34867 );
and ( n34869 , C1 , n34868 );
and ( n34870 , C1 , n34869 );
and ( n34871 , C1 , n34870 );
and ( n34872 , C1 , n34871 );
and ( n34873 , C1 , n34872 );
and ( n34874 , C1 , n34873 );
and ( n34875 , C1 , n34874 );
and ( n34876 , C1 , n34875 );
and ( n34877 , C1 , n34876 );
and ( n34878 , C1 , n34877 );
and ( n34879 , C1 , n34878 );
and ( n34880 , C1 , n34879 );
and ( n34881 , C1 , n34880 );
and ( n34882 , C1 , n34881 );
and ( n34883 , C1 , n34882 );
and ( n34884 , C1 , n34883 );
and ( n34885 , C1 , n34884 );
and ( n34886 , C1 , n34885 );
and ( n34887 , C1 , n34886 );
and ( n34888 , C1 , n34887 );
and ( n34889 , C1 , n34888 );
and ( n34890 , C1 , n34889 );
buf ( n34891 , n34890 );
not ( n34892 , n34891 );
buf ( n34893 , n34892 );
buf ( n34894 , n34893 );
and ( n34895 , n34834 , n34894 );
not ( n34896 , n34893 );
buf ( n34897 , n34896 );
not ( n34898 , n34832 );
and ( n34899 , n34898 , n34839 );
xor ( n34900 , n34840 , n34860 );
and ( n34901 , n34900 , n34832 );
or ( n34902 , n34899 , n34901 );
buf ( n34903 , n34902 );
not ( n34904 , n34903 );
buf ( n34905 , n34904 );
buf ( n34906 , n34905 );
and ( n34907 , C1 , n34906 );
and ( n34908 , C1 , n34907 );
and ( n34909 , C1 , n34908 );
and ( n34910 , C1 , n34909 );
and ( n34911 , C1 , n34910 );
and ( n34912 , C1 , n34911 );
and ( n34913 , C1 , n34912 );
and ( n34914 , C1 , n34913 );
and ( n34915 , C1 , n34914 );
and ( n34916 , C1 , n34915 );
and ( n34917 , C1 , n34916 );
and ( n34918 , C1 , n34917 );
and ( n34919 , C1 , n34918 );
and ( n34920 , C1 , n34919 );
and ( n34921 , C1 , n34920 );
and ( n34922 , C1 , n34921 );
and ( n34923 , C1 , n34922 );
and ( n34924 , C1 , n34923 );
and ( n34925 , C1 , n34924 );
and ( n34926 , C1 , n34925 );
and ( n34927 , C1 , n34926 );
and ( n34928 , C1 , n34927 );
and ( n34929 , C1 , n34928 );
buf ( n34930 , n34929 );
not ( n34931 , n34930 );
buf ( n34932 , n34931 );
not ( n34933 , n34932 );
buf ( n34934 , n34933 );
not ( n34935 , n34832 );
and ( n34936 , n34935 , n34841 );
xor ( n34937 , n34842 , n34859 );
and ( n34938 , n34937 , n34832 );
or ( n34939 , n34936 , n34938 );
buf ( n34940 , n34939 );
not ( n34941 , n34940 );
buf ( n34942 , n34941 );
buf ( n34943 , n34942 );
and ( n34944 , C1 , n34943 );
and ( n34945 , C1 , n34944 );
and ( n34946 , C1 , n34945 );
and ( n34947 , C1 , n34946 );
and ( n34948 , C1 , n34947 );
and ( n34949 , C1 , n34948 );
and ( n34950 , C1 , n34949 );
and ( n34951 , C1 , n34950 );
and ( n34952 , C1 , n34951 );
and ( n34953 , C1 , n34952 );
and ( n34954 , C1 , n34953 );
and ( n34955 , C1 , n34954 );
and ( n34956 , C1 , n34955 );
and ( n34957 , C1 , n34956 );
and ( n34958 , C1 , n34957 );
and ( n34959 , C1 , n34958 );
and ( n34960 , C1 , n34959 );
and ( n34961 , C1 , n34960 );
and ( n34962 , C1 , n34961 );
and ( n34963 , C1 , n34962 );
and ( n34964 , C1 , n34963 );
and ( n34965 , C1 , n34964 );
and ( n34966 , C1 , n34965 );
and ( n34967 , C1 , n34966 );
buf ( n34968 , n34967 );
not ( n34969 , n34968 );
buf ( n34970 , n34969 );
not ( n34971 , n34970 );
buf ( n34972 , n34971 );
not ( n34973 , n34832 );
and ( n34974 , n34973 , n34843 );
xor ( n34975 , n34844 , n34858 );
and ( n34976 , n34975 , n34832 );
or ( n34977 , n34974 , n34976 );
buf ( n34978 , n34977 );
not ( n34979 , n34978 );
buf ( n34980 , n34979 );
buf ( n34981 , n34980 );
and ( n34982 , C1 , n34981 );
and ( n34983 , C1 , n34982 );
and ( n34984 , C1 , n34983 );
and ( n34985 , C1 , n34984 );
and ( n34986 , C1 , n34985 );
and ( n34987 , C1 , n34986 );
and ( n34988 , C1 , n34987 );
and ( n34989 , C1 , n34988 );
and ( n34990 , C1 , n34989 );
and ( n34991 , C1 , n34990 );
and ( n34992 , C1 , n34991 );
and ( n34993 , C1 , n34992 );
and ( n34994 , C1 , n34993 );
and ( n34995 , C1 , n34994 );
and ( n34996 , C1 , n34995 );
and ( n34997 , C1 , n34996 );
and ( n34998 , C1 , n34997 );
and ( n34999 , C1 , n34998 );
and ( n35000 , C1 , n34999 );
and ( n35001 , C1 , n35000 );
and ( n35002 , C1 , n35001 );
and ( n35003 , C1 , n35002 );
and ( n35004 , C1 , n35003 );
and ( n35005 , C1 , n35004 );
and ( n35006 , C1 , n35005 );
buf ( n35007 , n35006 );
not ( n35008 , n35007 );
buf ( n35009 , n35008 );
not ( n35010 , n35009 );
buf ( n35011 , n35010 );
not ( n35012 , n34832 );
and ( n35013 , n35012 , n34845 );
xor ( n35014 , n34846 , n34857 );
and ( n35015 , n35014 , n34832 );
or ( n35016 , n35013 , n35015 );
buf ( n35017 , n35016 );
not ( n35018 , n35017 );
buf ( n35019 , n35018 );
buf ( n35020 , n35019 );
and ( n35021 , C1 , n35020 );
and ( n35022 , C1 , n35021 );
and ( n35023 , C1 , n35022 );
and ( n35024 , C1 , n35023 );
and ( n35025 , C1 , n35024 );
and ( n35026 , C1 , n35025 );
and ( n35027 , C1 , n35026 );
and ( n35028 , C1 , n35027 );
and ( n35029 , C1 , n35028 );
and ( n35030 , C1 , n35029 );
and ( n35031 , C1 , n35030 );
and ( n35032 , C1 , n35031 );
and ( n35033 , C1 , n35032 );
and ( n35034 , C1 , n35033 );
and ( n35035 , C1 , n35034 );
and ( n35036 , C1 , n35035 );
and ( n35037 , C1 , n35036 );
and ( n35038 , C1 , n35037 );
and ( n35039 , C1 , n35038 );
and ( n35040 , C1 , n35039 );
and ( n35041 , C1 , n35040 );
and ( n35042 , C1 , n35041 );
and ( n35043 , C1 , n35042 );
and ( n35044 , C1 , n35043 );
and ( n35045 , C1 , n35044 );
and ( n35046 , C1 , n35045 );
buf ( n35047 , n35046 );
not ( n35048 , n35047 );
buf ( n35049 , n35048 );
not ( n35050 , n35049 );
buf ( n35051 , n35050 );
not ( n35052 , n34832 );
and ( n35053 , n35052 , n34847 );
xor ( n35054 , n34848 , n34856 );
and ( n35055 , n35054 , n34832 );
or ( n35056 , n35053 , n35055 );
buf ( n35057 , n35056 );
not ( n35058 , n35057 );
buf ( n35059 , n35058 );
buf ( n35060 , n35059 );
and ( n35061 , C1 , n35060 );
and ( n35062 , C1 , n35061 );
and ( n35063 , C1 , n35062 );
and ( n35064 , C1 , n35063 );
and ( n35065 , C1 , n35064 );
and ( n35066 , C1 , n35065 );
and ( n35067 , C1 , n35066 );
and ( n35068 , C1 , n35067 );
and ( n35069 , C1 , n35068 );
and ( n35070 , C1 , n35069 );
and ( n35071 , C1 , n35070 );
and ( n35072 , C1 , n35071 );
and ( n35073 , C1 , n35072 );
and ( n35074 , C1 , n35073 );
and ( n35075 , C1 , n35074 );
and ( n35076 , C1 , n35075 );
and ( n35077 , C1 , n35076 );
and ( n35078 , C1 , n35077 );
and ( n35079 , C1 , n35078 );
and ( n35080 , C1 , n35079 );
and ( n35081 , C1 , n35080 );
and ( n35082 , C1 , n35081 );
and ( n35083 , C1 , n35082 );
and ( n35084 , C1 , n35083 );
and ( n35085 , C1 , n35084 );
and ( n35086 , C1 , n35085 );
and ( n35087 , C1 , n35086 );
buf ( n35088 , n35087 );
not ( n35089 , n35088 );
buf ( n35090 , n35089 );
not ( n35091 , n35090 );
buf ( n35092 , n35091 );
not ( n35093 , n34832 );
and ( n35094 , n35093 , n34849 );
xor ( n35095 , n34850 , n34855 );
and ( n35096 , n35095 , n34832 );
or ( n35097 , n35094 , n35096 );
buf ( n35098 , n35097 );
not ( n35099 , n35098 );
buf ( n35100 , n35099 );
buf ( n35101 , n35100 );
and ( n35102 , C1 , n35101 );
and ( n35103 , C1 , n35102 );
and ( n35104 , C1 , n35103 );
and ( n35105 , C1 , n35104 );
and ( n35106 , C1 , n35105 );
and ( n35107 , C1 , n35106 );
and ( n35108 , C1 , n35107 );
and ( n35109 , C1 , n35108 );
and ( n35110 , C1 , n35109 );
and ( n35111 , C1 , n35110 );
and ( n35112 , C1 , n35111 );
and ( n35113 , C1 , n35112 );
and ( n35114 , C1 , n35113 );
and ( n35115 , C1 , n35114 );
and ( n35116 , C1 , n35115 );
and ( n35117 , C1 , n35116 );
and ( n35118 , C1 , n35117 );
and ( n35119 , C1 , n35118 );
and ( n35120 , C1 , n35119 );
and ( n35121 , C1 , n35120 );
and ( n35122 , C1 , n35121 );
and ( n35123 , C1 , n35122 );
and ( n35124 , C1 , n35123 );
and ( n35125 , C1 , n35124 );
and ( n35126 , C1 , n35125 );
and ( n35127 , C1 , n35126 );
and ( n35128 , C1 , n35127 );
and ( n35129 , C1 , n35128 );
buf ( n35130 , n35129 );
not ( n35131 , n35130 );
buf ( n35132 , n35131 );
not ( n35133 , n35132 );
buf ( n35134 , n35133 );
not ( n35135 , n34832 );
and ( n35136 , n35135 , n34851 );
xor ( n35137 , n34852 , n34854 );
and ( n35138 , n35137 , n34832 );
or ( n35139 , n35136 , n35138 );
buf ( n35140 , n35139 );
not ( n35141 , n35140 );
buf ( n35142 , n35141 );
buf ( n35143 , n35142 );
and ( n35144 , C1 , n35143 );
and ( n35145 , C1 , n35144 );
and ( n35146 , C1 , n35145 );
and ( n35147 , C1 , n35146 );
and ( n35148 , C1 , n35147 );
and ( n35149 , C1 , n35148 );
and ( n35150 , C1 , n35149 );
and ( n35151 , C1 , n35150 );
and ( n35152 , C1 , n35151 );
and ( n35153 , C1 , n35152 );
and ( n35154 , C1 , n35153 );
and ( n35155 , C1 , n35154 );
and ( n35156 , C1 , n35155 );
and ( n35157 , C1 , n35156 );
and ( n35158 , C1 , n35157 );
and ( n35159 , C1 , n35158 );
and ( n35160 , C1 , n35159 );
and ( n35161 , C1 , n35160 );
and ( n35162 , C1 , n35161 );
and ( n35163 , C1 , n35162 );
and ( n35164 , C1 , n35163 );
and ( n35165 , C1 , n35164 );
and ( n35166 , C1 , n35165 );
and ( n35167 , C1 , n35166 );
and ( n35168 , C1 , n35167 );
and ( n35169 , C1 , n35168 );
and ( n35170 , C1 , n35169 );
and ( n35171 , C1 , n35170 );
and ( n35172 , C1 , n35171 );
buf ( n35173 , n35172 );
not ( n35174 , n35173 );
buf ( n35175 , n35174 );
not ( n35176 , n35175 );
buf ( n35177 , n35176 );
and ( n35178 , n35134 , n35177 );
and ( n35179 , n35092 , n35178 );
and ( n35180 , n35051 , n35179 );
and ( n35181 , n35011 , n35180 );
and ( n35182 , n34972 , n35181 );
and ( n35183 , n34934 , n35182 );
xor ( n35184 , n34897 , n35183 );
buf ( n35185 , n35184 );
and ( n35186 , n35185 , n34833 );
or ( n35187 , n34895 , n35186 );
buf ( n35188 , n35187 );
and ( n35189 , n34831 , n35188 );
buf ( n35190 , n35175 );
buf ( n35191 , n35190 );
buf ( n35192 , n35191 );
not ( n35193 , n35192 );
buf ( n35194 , n35193 );
buf ( n35195 , n35194 );
not ( n35196 , n35195 );
not ( n35197 , n34832 );
buf ( n35198 , n14611 );
not ( n35199 , n35198 );
buf ( n35200 , n14964 );
not ( n35201 , n35200 );
buf ( n35202 , n13162 );
not ( n35203 , n35202 );
buf ( n35204 , n13175 );
not ( n35205 , n35204 );
buf ( n35206 , n13187 );
not ( n35207 , n35206 );
buf ( n35208 , n13199 );
not ( n35209 , n35208 );
buf ( n35210 , n13211 );
not ( n35211 , n35210 );
buf ( n35212 , n13223 );
not ( n35213 , n35212 );
buf ( n35214 , n13235 );
not ( n35215 , n35214 );
buf ( n35216 , n13247 );
not ( n35217 , n35216 );
buf ( n35218 , n13259 );
not ( n35219 , n35218 );
buf ( n35220 , n13271 );
not ( n35221 , n35220 );
buf ( n35222 , n13283 );
not ( n35223 , n35222 );
buf ( n35224 , n13295 );
not ( n35225 , n35224 );
buf ( n35226 , n13307 );
not ( n35227 , n35226 );
buf ( n35228 , n13319 );
not ( n35229 , n35228 );
buf ( n35230 , n13331 );
not ( n35231 , n35230 );
buf ( n35232 , n13343 );
not ( n35233 , n35232 );
buf ( n35234 , n13355 );
not ( n35235 , n35234 );
buf ( n35236 , n13367 );
not ( n35237 , n35236 );
buf ( n35238 , n13379 );
not ( n35239 , n35238 );
buf ( n35240 , n13391 );
not ( n35241 , n35240 );
and ( n35242 , n34838 , n34861 );
and ( n35243 , n35241 , n35242 );
and ( n35244 , n35239 , n35243 );
and ( n35245 , n35237 , n35244 );
and ( n35246 , n35235 , n35245 );
and ( n35247 , n35233 , n35246 );
and ( n35248 , n35231 , n35247 );
and ( n35249 , n35229 , n35248 );
and ( n35250 , n35227 , n35249 );
and ( n35251 , n35225 , n35250 );
and ( n35252 , n35223 , n35251 );
and ( n35253 , n35221 , n35252 );
and ( n35254 , n35219 , n35253 );
and ( n35255 , n35217 , n35254 );
and ( n35256 , n35215 , n35255 );
and ( n35257 , n35213 , n35256 );
and ( n35258 , n35211 , n35257 );
and ( n35259 , n35209 , n35258 );
and ( n35260 , n35207 , n35259 );
and ( n35261 , n35205 , n35260 );
and ( n35262 , n35203 , n35261 );
and ( n35263 , n35201 , n35262 );
and ( n35264 , n35199 , n35263 );
xor ( n35265 , n35197 , n35264 );
buf ( n35266 , n34832 );
and ( n35267 , n35265 , n35266 );
or ( n35268 , C0 , n35267 );
buf ( n35269 , n35268 );
not ( n35270 , n35269 );
buf ( n35271 , n35270 );
not ( n35272 , n35271 );
buf ( n35273 , n35272 );
not ( n35274 , n35273 );
buf ( n35275 , n35274 );
not ( n35276 , n34832 );
and ( n35277 , n35276 , n35198 );
xor ( n35278 , n35199 , n35263 );
and ( n35279 , n35278 , n34832 );
or ( n35280 , n35277 , n35279 );
buf ( n35281 , n35280 );
not ( n35282 , n35281 );
buf ( n35283 , n35282 );
buf ( n35284 , n35283 );
not ( n35285 , n35284 );
buf ( n35286 , n35285 );
not ( n35287 , n35286 );
buf ( n35288 , n35287 );
not ( n35289 , n34832 );
and ( n35290 , n35289 , n35200 );
xor ( n35291 , n35201 , n35262 );
and ( n35292 , n35291 , n34832 );
or ( n35293 , n35290 , n35292 );
buf ( n35294 , n35293 );
not ( n35295 , n35294 );
buf ( n35296 , n35295 );
buf ( n35297 , n35296 );
not ( n35298 , n35297 );
buf ( n35299 , n35298 );
not ( n35300 , n35299 );
buf ( n35301 , n35300 );
not ( n35302 , n34832 );
and ( n35303 , n35302 , n35202 );
xor ( n35304 , n35203 , n35261 );
and ( n35305 , n35304 , n34832 );
or ( n35306 , n35303 , n35305 );
buf ( n35307 , n35306 );
not ( n35308 , n35307 );
buf ( n35309 , n35308 );
buf ( n35310 , n35309 );
not ( n35311 , n35310 );
buf ( n35312 , n35311 );
not ( n35313 , n35312 );
buf ( n35314 , n35313 );
not ( n35315 , n34832 );
and ( n35316 , n35315 , n35204 );
xor ( n35317 , n35205 , n35260 );
and ( n35318 , n35317 , n34832 );
or ( n35319 , n35316 , n35318 );
buf ( n35320 , n35319 );
not ( n35321 , n35320 );
buf ( n35322 , n35321 );
buf ( n35323 , n35322 );
not ( n35324 , n35323 );
buf ( n35325 , n35324 );
not ( n35326 , n35325 );
buf ( n35327 , n35326 );
not ( n35328 , n34832 );
and ( n35329 , n35328 , n35206 );
xor ( n35330 , n35207 , n35259 );
and ( n35331 , n35330 , n34832 );
or ( n35332 , n35329 , n35331 );
buf ( n35333 , n35332 );
not ( n35334 , n35333 );
buf ( n35335 , n35334 );
buf ( n35336 , n35335 );
not ( n35337 , n35336 );
buf ( n35338 , n35337 );
not ( n35339 , n35338 );
buf ( n35340 , n35339 );
not ( n35341 , n34832 );
and ( n35342 , n35341 , n35208 );
xor ( n35343 , n35209 , n35258 );
and ( n35344 , n35343 , n34832 );
or ( n35345 , n35342 , n35344 );
buf ( n35346 , n35345 );
not ( n35347 , n35346 );
buf ( n35348 , n35347 );
buf ( n35349 , n35348 );
not ( n35350 , n35349 );
buf ( n35351 , n35350 );
not ( n35352 , n35351 );
buf ( n35353 , n35352 );
not ( n35354 , n34832 );
and ( n35355 , n35354 , n35210 );
xor ( n35356 , n35211 , n35257 );
and ( n35357 , n35356 , n34832 );
or ( n35358 , n35355 , n35357 );
buf ( n35359 , n35358 );
not ( n35360 , n35359 );
buf ( n35361 , n35360 );
buf ( n35362 , n35361 );
not ( n35363 , n35362 );
buf ( n35364 , n35363 );
not ( n35365 , n35364 );
buf ( n35366 , n35365 );
not ( n35367 , n34832 );
and ( n35368 , n35367 , n35212 );
xor ( n35369 , n35213 , n35256 );
and ( n35370 , n35369 , n34832 );
or ( n35371 , n35368 , n35370 );
buf ( n35372 , n35371 );
not ( n35373 , n35372 );
buf ( n35374 , n35373 );
buf ( n35375 , n35374 );
not ( n35376 , n35375 );
buf ( n35377 , n35376 );
not ( n35378 , n35377 );
buf ( n35379 , n35378 );
not ( n35380 , n34832 );
and ( n35381 , n35380 , n35214 );
xor ( n35382 , n35215 , n35255 );
and ( n35383 , n35382 , n34832 );
or ( n35384 , n35381 , n35383 );
buf ( n35385 , n35384 );
not ( n35386 , n35385 );
buf ( n35387 , n35386 );
buf ( n35388 , n35387 );
not ( n35389 , n35388 );
buf ( n35390 , n35389 );
not ( n35391 , n35390 );
buf ( n35392 , n35391 );
not ( n35393 , n34832 );
and ( n35394 , n35393 , n35216 );
xor ( n35395 , n35217 , n35254 );
and ( n35396 , n35395 , n34832 );
or ( n35397 , n35394 , n35396 );
buf ( n35398 , n35397 );
not ( n35399 , n35398 );
buf ( n35400 , n35399 );
buf ( n35401 , n35400 );
not ( n35402 , n35401 );
buf ( n35403 , n35402 );
not ( n35404 , n35403 );
buf ( n35405 , n35404 );
not ( n35406 , n34832 );
and ( n35407 , n35406 , n35218 );
xor ( n35408 , n35219 , n35253 );
and ( n35409 , n35408 , n34832 );
or ( n35410 , n35407 , n35409 );
buf ( n35411 , n35410 );
not ( n35412 , n35411 );
buf ( n35413 , n35412 );
buf ( n35414 , n35413 );
not ( n35415 , n35414 );
buf ( n35416 , n35415 );
not ( n35417 , n35416 );
buf ( n35418 , n35417 );
not ( n35419 , n34832 );
and ( n35420 , n35419 , n35220 );
xor ( n35421 , n35221 , n35252 );
and ( n35422 , n35421 , n34832 );
or ( n35423 , n35420 , n35422 );
buf ( n35424 , n35423 );
not ( n35425 , n35424 );
buf ( n35426 , n35425 );
buf ( n35427 , n35426 );
not ( n35428 , n35427 );
buf ( n35429 , n35428 );
not ( n35430 , n35429 );
buf ( n35431 , n35430 );
not ( n35432 , n34832 );
and ( n35433 , n35432 , n35222 );
xor ( n35434 , n35223 , n35251 );
and ( n35435 , n35434 , n34832 );
or ( n35436 , n35433 , n35435 );
buf ( n35437 , n35436 );
not ( n35438 , n35437 );
buf ( n35439 , n35438 );
buf ( n35440 , n35439 );
not ( n35441 , n35440 );
buf ( n35442 , n35441 );
not ( n35443 , n35442 );
buf ( n35444 , n35443 );
not ( n35445 , n34832 );
and ( n35446 , n35445 , n35224 );
xor ( n35447 , n35225 , n35250 );
and ( n35448 , n35447 , n34832 );
or ( n35449 , n35446 , n35448 );
buf ( n35450 , n35449 );
not ( n35451 , n35450 );
buf ( n35452 , n35451 );
buf ( n35453 , n35452 );
not ( n35454 , n35453 );
buf ( n35455 , n35454 );
not ( n35456 , n35455 );
buf ( n35457 , n35456 );
not ( n35458 , n34832 );
and ( n35459 , n35458 , n35226 );
xor ( n35460 , n35227 , n35249 );
and ( n35461 , n35460 , n34832 );
or ( n35462 , n35459 , n35461 );
buf ( n35463 , n35462 );
not ( n35464 , n35463 );
buf ( n35465 , n35464 );
buf ( n35466 , n35465 );
not ( n35467 , n35466 );
buf ( n35468 , n35467 );
not ( n35469 , n35468 );
buf ( n35470 , n35469 );
not ( n35471 , n34832 );
and ( n35472 , n35471 , n35228 );
xor ( n35473 , n35229 , n35248 );
and ( n35474 , n35473 , n34832 );
or ( n35475 , n35472 , n35474 );
buf ( n35476 , n35475 );
not ( n35477 , n35476 );
buf ( n35478 , n35477 );
buf ( n35479 , n35478 );
not ( n35480 , n35479 );
buf ( n35481 , n35480 );
not ( n35482 , n35481 );
buf ( n35483 , n35482 );
not ( n35484 , n34832 );
and ( n35485 , n35484 , n35230 );
xor ( n35486 , n35231 , n35247 );
and ( n35487 , n35486 , n34832 );
or ( n35488 , n35485 , n35487 );
buf ( n35489 , n35488 );
not ( n35490 , n35489 );
buf ( n35491 , n35490 );
buf ( n35492 , n35491 );
not ( n35493 , n35492 );
buf ( n35494 , n35493 );
not ( n35495 , n35494 );
buf ( n35496 , n35495 );
not ( n35497 , n34832 );
and ( n35498 , n35497 , n35232 );
xor ( n35499 , n35233 , n35246 );
and ( n35500 , n35499 , n34832 );
or ( n35501 , n35498 , n35500 );
buf ( n35502 , n35501 );
not ( n35503 , n35502 );
buf ( n35504 , n35503 );
buf ( n35505 , n35504 );
not ( n35506 , n35505 );
buf ( n35507 , n35506 );
not ( n35508 , n35507 );
buf ( n35509 , n35508 );
not ( n35510 , n34832 );
and ( n35511 , n35510 , n35234 );
xor ( n35512 , n35235 , n35245 );
and ( n35513 , n35512 , n34832 );
or ( n35514 , n35511 , n35513 );
buf ( n35515 , n35514 );
not ( n35516 , n35515 );
buf ( n35517 , n35516 );
buf ( n35518 , n35517 );
not ( n35519 , n35518 );
buf ( n35520 , n35519 );
not ( n35521 , n35520 );
buf ( n35522 , n35521 );
not ( n35523 , n34832 );
and ( n35524 , n35523 , n35236 );
xor ( n35525 , n35237 , n35244 );
and ( n35526 , n35525 , n34832 );
or ( n35527 , n35524 , n35526 );
buf ( n35528 , n35527 );
not ( n35529 , n35528 );
buf ( n35530 , n35529 );
buf ( n35531 , n35530 );
not ( n35532 , n35531 );
buf ( n35533 , n35532 );
not ( n35534 , n35533 );
buf ( n35535 , n35534 );
not ( n35536 , n34832 );
and ( n35537 , n35536 , n35238 );
xor ( n35538 , n35239 , n35243 );
and ( n35539 , n35538 , n34832 );
or ( n35540 , n35537 , n35539 );
buf ( n35541 , n35540 );
not ( n35542 , n35541 );
buf ( n35543 , n35542 );
buf ( n35544 , n35543 );
and ( n35545 , C1 , n35544 );
and ( n35546 , C1 , n35545 );
and ( n35547 , C1 , n35546 );
and ( n35548 , C1 , n35547 );
and ( n35549 , C1 , n35548 );
and ( n35550 , C1 , n35549 );
and ( n35551 , C1 , n35550 );
and ( n35552 , C1 , n35551 );
and ( n35553 , C1 , n35552 );
and ( n35554 , C1 , n35553 );
and ( n35555 , C1 , n35554 );
and ( n35556 , C1 , n35555 );
and ( n35557 , C1 , n35556 );
and ( n35558 , C1 , n35557 );
and ( n35559 , C1 , n35558 );
and ( n35560 , C1 , n35559 );
and ( n35561 , C1 , n35560 );
and ( n35562 , C1 , n35561 );
and ( n35563 , C1 , n35562 );
and ( n35564 , C1 , n35563 );
and ( n35565 , C1 , n35564 );
not ( n35566 , n35565 );
buf ( n35567 , n35566 );
not ( n35568 , n35567 );
buf ( n35569 , n35568 );
not ( n35570 , n34832 );
and ( n35571 , n35570 , n35240 );
xor ( n35572 , n35241 , n35242 );
and ( n35573 , n35572 , n34832 );
or ( n35574 , n35571 , n35573 );
buf ( n35575 , n35574 );
not ( n35576 , n35575 );
buf ( n35577 , n35576 );
buf ( n35578 , n35577 );
and ( n35579 , C1 , n35578 );
and ( n35580 , C1 , n35579 );
and ( n35581 , C1 , n35580 );
and ( n35582 , C1 , n35581 );
and ( n35583 , C1 , n35582 );
and ( n35584 , C1 , n35583 );
and ( n35585 , C1 , n35584 );
and ( n35586 , C1 , n35585 );
and ( n35587 , C1 , n35586 );
and ( n35588 , C1 , n35587 );
and ( n35589 , C1 , n35588 );
and ( n35590 , C1 , n35589 );
and ( n35591 , C1 , n35590 );
and ( n35592 , C1 , n35591 );
and ( n35593 , C1 , n35592 );
and ( n35594 , C1 , n35593 );
and ( n35595 , C1 , n35594 );
and ( n35596 , C1 , n35595 );
and ( n35597 , C1 , n35596 );
and ( n35598 , C1 , n35597 );
and ( n35599 , C1 , n35598 );
buf ( n35600 , n35599 );
not ( n35601 , n35600 );
buf ( n35602 , n35601 );
not ( n35603 , n35602 );
buf ( n35604 , n35603 );
and ( n35605 , n34897 , n35183 );
and ( n35606 , n35604 , n35605 );
and ( n35607 , n35569 , n35606 );
and ( n35608 , n35535 , n35607 );
and ( n35609 , n35522 , n35608 );
and ( n35610 , n35509 , n35609 );
and ( n35611 , n35496 , n35610 );
and ( n35612 , n35483 , n35611 );
and ( n35613 , n35470 , n35612 );
and ( n35614 , n35457 , n35613 );
and ( n35615 , n35444 , n35614 );
and ( n35616 , n35431 , n35615 );
and ( n35617 , n35418 , n35616 );
and ( n35618 , n35405 , n35617 );
and ( n35619 , n35392 , n35618 );
and ( n35620 , n35379 , n35619 );
and ( n35621 , n35366 , n35620 );
and ( n35622 , n35353 , n35621 );
and ( n35623 , n35340 , n35622 );
and ( n35624 , n35327 , n35623 );
and ( n35625 , n35314 , n35624 );
and ( n35626 , n35301 , n35625 );
and ( n35627 , n35288 , n35626 );
and ( n35628 , n35275 , n35627 );
not ( n35629 , n35628 );
buf ( n35630 , n35629 );
and ( n35631 , n35630 , n34833 );
or ( n35632 , C0 , n35631 );
buf ( n35633 , n35632 );
buf ( n35634 , n35633 );
not ( n35635 , n35634 );
not ( n35636 , n34833 );
buf ( n35637 , n35132 );
and ( n35638 , n35636 , n35637 );
xor ( n35639 , n35134 , n35177 );
buf ( n35640 , n35639 );
and ( n35641 , n35640 , n34833 );
or ( n35642 , n35638 , n35641 );
buf ( n35643 , n35642 );
buf ( n35644 , n35643 );
and ( n35645 , n35635 , n35644 );
not ( n35646 , n35644 );
not ( n35647 , n35191 );
xor ( n35648 , n35646 , n35647 );
and ( n35649 , n35648 , n35634 );
or ( n35650 , n35645 , n35649 );
buf ( n35651 , n35650 );
not ( n35652 , n35651 );
buf ( n35653 , n35652 );
buf ( n35654 , n35653 );
not ( n35655 , n35654 );
or ( n35656 , n35196 , n35655 );
not ( n35657 , n35634 );
not ( n35658 , n34833 );
buf ( n35659 , n35090 );
and ( n35660 , n35658 , n35659 );
xor ( n35661 , n35092 , n35178 );
buf ( n35662 , n35661 );
and ( n35663 , n35662 , n34833 );
or ( n35664 , n35660 , n35663 );
buf ( n35665 , n35664 );
buf ( n35666 , n35665 );
and ( n35667 , n35657 , n35666 );
not ( n35668 , n35666 );
and ( n35669 , n35646 , n35647 );
xor ( n35670 , n35668 , n35669 );
and ( n35671 , n35670 , n35634 );
or ( n35672 , n35667 , n35671 );
buf ( n35673 , n35672 );
not ( n35674 , n35673 );
buf ( n35675 , n35674 );
buf ( n35676 , n35675 );
not ( n35677 , n35676 );
or ( n35678 , n35656 , n35677 );
not ( n35679 , n35634 );
not ( n35680 , n34833 );
buf ( n35681 , n35049 );
and ( n35682 , n35680 , n35681 );
xor ( n35683 , n35051 , n35179 );
buf ( n35684 , n35683 );
and ( n35685 , n35684 , n34833 );
or ( n35686 , n35682 , n35685 );
buf ( n35687 , n35686 );
buf ( n35688 , n35687 );
and ( n35689 , n35679 , n35688 );
not ( n35690 , n35688 );
and ( n35691 , n35668 , n35669 );
xor ( n35692 , n35690 , n35691 );
and ( n35693 , n35692 , n35634 );
or ( n35694 , n35689 , n35693 );
buf ( n35695 , n35694 );
not ( n35696 , n35695 );
buf ( n35697 , n35696 );
buf ( n35698 , n35697 );
not ( n35699 , n35698 );
or ( n35700 , n35678 , n35699 );
not ( n35701 , n35634 );
not ( n35702 , n34833 );
buf ( n35703 , n35009 );
and ( n35704 , n35702 , n35703 );
xor ( n35705 , n35011 , n35180 );
buf ( n35706 , n35705 );
and ( n35707 , n35706 , n34833 );
or ( n35708 , n35704 , n35707 );
buf ( n35709 , n35708 );
buf ( n35710 , n35709 );
and ( n35711 , n35701 , n35710 );
not ( n35712 , n35710 );
and ( n35713 , n35690 , n35691 );
xor ( n35714 , n35712 , n35713 );
and ( n35715 , n35714 , n35634 );
or ( n35716 , n35711 , n35715 );
buf ( n35717 , n35716 );
not ( n35718 , n35717 );
buf ( n35719 , n35718 );
buf ( n35720 , n35719 );
not ( n35721 , n35720 );
or ( n35722 , n35700 , n35721 );
not ( n35723 , n35634 );
not ( n35724 , n34833 );
buf ( n35725 , n34970 );
and ( n35726 , n35724 , n35725 );
xor ( n35727 , n34972 , n35181 );
buf ( n35728 , n35727 );
and ( n35729 , n35728 , n34833 );
or ( n35730 , n35726 , n35729 );
buf ( n35731 , n35730 );
buf ( n35732 , n35731 );
and ( n35733 , n35723 , n35732 );
not ( n35734 , n35732 );
and ( n35735 , n35712 , n35713 );
xor ( n35736 , n35734 , n35735 );
and ( n35737 , n35736 , n35634 );
or ( n35738 , n35733 , n35737 );
buf ( n35739 , n35738 );
not ( n35740 , n35739 );
buf ( n35741 , n35740 );
buf ( n35742 , n35741 );
not ( n35743 , n35742 );
or ( n35744 , n35722 , n35743 );
not ( n35745 , n35634 );
not ( n35746 , n34833 );
buf ( n35747 , n34932 );
and ( n35748 , n35746 , n35747 );
xor ( n35749 , n34934 , n35182 );
buf ( n35750 , n35749 );
and ( n35751 , n35750 , n34833 );
or ( n35752 , n35748 , n35751 );
buf ( n35753 , n35752 );
buf ( n35754 , n35753 );
and ( n35755 , n35745 , n35754 );
not ( n35756 , n35754 );
and ( n35757 , n35734 , n35735 );
xor ( n35758 , n35756 , n35757 );
and ( n35759 , n35758 , n35634 );
or ( n35760 , n35755 , n35759 );
buf ( n35761 , n35760 );
not ( n35762 , n35761 );
buf ( n35763 , n35762 );
buf ( n35764 , n35763 );
not ( n35765 , n35764 );
or ( n35766 , n35744 , n35765 );
not ( n35767 , n35634 );
buf ( n35768 , n35188 );
and ( n35769 , n35767 , n35768 );
not ( n35770 , n35768 );
and ( n35771 , n35756 , n35757 );
xor ( n35772 , n35770 , n35771 );
and ( n35773 , n35772 , n35634 );
or ( n35774 , n35769 , n35773 );
buf ( n35775 , n35774 );
not ( n35776 , n35775 );
buf ( n35777 , n35776 );
buf ( n35778 , n35777 );
not ( n35779 , n35778 );
or ( n35780 , n35766 , n35779 );
not ( n35781 , n35634 );
not ( n35782 , n34833 );
buf ( n35783 , n35602 );
and ( n35784 , n35782 , n35783 );
xor ( n35785 , n35604 , n35605 );
buf ( n35786 , n35785 );
and ( n35787 , n35786 , n34833 );
or ( n35788 , n35784 , n35787 );
buf ( n35789 , n35788 );
buf ( n35790 , n35789 );
and ( n35791 , n35781 , n35790 );
not ( n35792 , n35790 );
and ( n35793 , n35770 , n35771 );
xor ( n35794 , n35792 , n35793 );
and ( n35795 , n35794 , n35634 );
or ( n35796 , n35791 , n35795 );
buf ( n35797 , n35796 );
not ( n35798 , n35797 );
buf ( n35799 , n35798 );
buf ( n35800 , n35799 );
not ( n35801 , n35800 );
or ( n35802 , n35780 , n35801 );
not ( n35803 , n35634 );
not ( n35804 , n34833 );
buf ( n35805 , n35567 );
and ( n35806 , n35804 , n35805 );
xor ( n35807 , n35569 , n35606 );
buf ( n35808 , n35807 );
and ( n35809 , n35808 , n34833 );
or ( n35810 , n35806 , n35809 );
buf ( n35811 , n35810 );
buf ( n35812 , n35811 );
and ( n35813 , n35803 , n35812 );
not ( n35814 , n35812 );
and ( n35815 , n35792 , n35793 );
xor ( n35816 , n35814 , n35815 );
and ( n35817 , n35816 , n35634 );
or ( n35818 , n35813 , n35817 );
buf ( n35819 , n35818 );
not ( n35820 , n35819 );
buf ( n35821 , n35820 );
buf ( n35822 , n35821 );
not ( n35823 , n35822 );
or ( n35824 , n35802 , n35823 );
not ( n35825 , n35634 );
not ( n35826 , n34833 );
buf ( n35827 , n35533 );
and ( n35828 , n35826 , n35827 );
xor ( n35829 , n35535 , n35607 );
buf ( n35830 , n35829 );
and ( n35831 , n35830 , n34833 );
or ( n35832 , n35828 , n35831 );
buf ( n35833 , n35832 );
buf ( n35834 , n35833 );
and ( n35835 , n35825 , n35834 );
not ( n35836 , n35834 );
and ( n35837 , n35814 , n35815 );
xor ( n35838 , n35836 , n35837 );
and ( n35839 , n35838 , n35634 );
or ( n35840 , n35835 , n35839 );
buf ( n35841 , n35840 );
not ( n35842 , n35841 );
buf ( n35843 , n35842 );
buf ( n35844 , n35843 );
not ( n35845 , n35844 );
or ( n35846 , n35824 , n35845 );
not ( n35847 , n35634 );
not ( n35848 , n34833 );
buf ( n35849 , n35520 );
and ( n35850 , n35848 , n35849 );
xor ( n35851 , n35522 , n35608 );
buf ( n35852 , n35851 );
and ( n35853 , n35852 , n34833 );
or ( n35854 , n35850 , n35853 );
buf ( n35855 , n35854 );
buf ( n35856 , n35855 );
and ( n35857 , n35847 , n35856 );
not ( n35858 , n35856 );
and ( n35859 , n35836 , n35837 );
xor ( n35860 , n35858 , n35859 );
and ( n35861 , n35860 , n35634 );
or ( n35862 , n35857 , n35861 );
buf ( n35863 , n35862 );
not ( n35864 , n35863 );
buf ( n35865 , n35864 );
buf ( n35866 , n35865 );
not ( n35867 , n35866 );
or ( n35868 , n35846 , n35867 );
not ( n35869 , n35634 );
not ( n35870 , n34833 );
buf ( n35871 , n35507 );
and ( n35872 , n35870 , n35871 );
xor ( n35873 , n35509 , n35609 );
buf ( n35874 , n35873 );
and ( n35875 , n35874 , n34833 );
or ( n35876 , n35872 , n35875 );
buf ( n35877 , n35876 );
buf ( n35878 , n35877 );
and ( n35879 , n35869 , n35878 );
not ( n35880 , n35878 );
and ( n35881 , n35858 , n35859 );
xor ( n35882 , n35880 , n35881 );
and ( n35883 , n35882 , n35634 );
or ( n35884 , n35879 , n35883 );
buf ( n35885 , n35884 );
not ( n35886 , n35885 );
buf ( n35887 , n35886 );
buf ( n35888 , n35887 );
not ( n35889 , n35888 );
or ( n35890 , n35868 , n35889 );
not ( n35891 , n35634 );
not ( n35892 , n34833 );
buf ( n35893 , n35494 );
and ( n35894 , n35892 , n35893 );
xor ( n35895 , n35496 , n35610 );
buf ( n35896 , n35895 );
and ( n35897 , n35896 , n34833 );
or ( n35898 , n35894 , n35897 );
buf ( n35899 , n35898 );
buf ( n35900 , n35899 );
and ( n35901 , n35891 , n35900 );
not ( n35902 , n35900 );
and ( n35903 , n35880 , n35881 );
xor ( n35904 , n35902 , n35903 );
and ( n35905 , n35904 , n35634 );
or ( n35906 , n35901 , n35905 );
buf ( n35907 , n35906 );
not ( n35908 , n35907 );
buf ( n35909 , n35908 );
buf ( n35910 , n35909 );
not ( n35911 , n35910 );
or ( n35912 , n35890 , n35911 );
not ( n35913 , n35634 );
not ( n35914 , n34833 );
buf ( n35915 , n35481 );
and ( n35916 , n35914 , n35915 );
xor ( n35917 , n35483 , n35611 );
buf ( n35918 , n35917 );
and ( n35919 , n35918 , n34833 );
or ( n35920 , n35916 , n35919 );
buf ( n35921 , n35920 );
buf ( n35922 , n35921 );
and ( n35923 , n35913 , n35922 );
not ( n35924 , n35922 );
and ( n35925 , n35902 , n35903 );
xor ( n35926 , n35924 , n35925 );
and ( n35927 , n35926 , n35634 );
or ( n35928 , n35923 , n35927 );
buf ( n35929 , n35928 );
not ( n35930 , n35929 );
buf ( n35931 , n35930 );
buf ( n35932 , n35931 );
not ( n35933 , n35932 );
or ( n35934 , n35912 , n35933 );
not ( n35935 , n35634 );
not ( n35936 , n34833 );
buf ( n35937 , n35468 );
and ( n35938 , n35936 , n35937 );
xor ( n35939 , n35470 , n35612 );
buf ( n35940 , n35939 );
and ( n35941 , n35940 , n34833 );
or ( n35942 , n35938 , n35941 );
buf ( n35943 , n35942 );
buf ( n35944 , n35943 );
and ( n35945 , n35935 , n35944 );
not ( n35946 , n35944 );
and ( n35947 , n35924 , n35925 );
xor ( n35948 , n35946 , n35947 );
and ( n35949 , n35948 , n35634 );
or ( n35950 , n35945 , n35949 );
buf ( n35951 , n35950 );
not ( n35952 , n35951 );
buf ( n35953 , n35952 );
buf ( n35954 , n35953 );
not ( n35955 , n35954 );
or ( n35956 , n35934 , n35955 );
not ( n35957 , n35634 );
not ( n35958 , n34833 );
buf ( n35959 , n35455 );
and ( n35960 , n35958 , n35959 );
xor ( n35961 , n35457 , n35613 );
buf ( n35962 , n35961 );
and ( n35963 , n35962 , n34833 );
or ( n35964 , n35960 , n35963 );
buf ( n35965 , n35964 );
buf ( n35966 , n35965 );
and ( n35967 , n35957 , n35966 );
not ( n35968 , n35966 );
and ( n35969 , n35946 , n35947 );
xor ( n35970 , n35968 , n35969 );
and ( n35971 , n35970 , n35634 );
or ( n35972 , n35967 , n35971 );
buf ( n35973 , n35972 );
not ( n35974 , n35973 );
buf ( n35975 , n35974 );
buf ( n35976 , n35975 );
not ( n35977 , n35976 );
or ( n35978 , n35956 , n35977 );
not ( n35979 , n35634 );
not ( n35980 , n34833 );
buf ( n35981 , n35442 );
and ( n35982 , n35980 , n35981 );
xor ( n35983 , n35444 , n35614 );
buf ( n35984 , n35983 );
and ( n35985 , n35984 , n34833 );
or ( n35986 , n35982 , n35985 );
buf ( n35987 , n35986 );
buf ( n35988 , n35987 );
and ( n35989 , n35979 , n35988 );
not ( n35990 , n35988 );
and ( n35991 , n35968 , n35969 );
xor ( n35992 , n35990 , n35991 );
and ( n35993 , n35992 , n35634 );
or ( n35994 , n35989 , n35993 );
buf ( n35995 , n35994 );
not ( n35996 , n35995 );
buf ( n35997 , n35996 );
buf ( n35998 , n35997 );
not ( n35999 , n35998 );
or ( n36000 , n35978 , n35999 );
not ( n36001 , n35634 );
not ( n36002 , n34833 );
buf ( n36003 , n35429 );
and ( n36004 , n36002 , n36003 );
xor ( n36005 , n35431 , n35615 );
buf ( n36006 , n36005 );
and ( n36007 , n36006 , n34833 );
or ( n36008 , n36004 , n36007 );
buf ( n36009 , n36008 );
buf ( n36010 , n36009 );
and ( n36011 , n36001 , n36010 );
not ( n36012 , n36010 );
and ( n36013 , n35990 , n35991 );
xor ( n36014 , n36012 , n36013 );
and ( n36015 , n36014 , n35634 );
or ( n36016 , n36011 , n36015 );
buf ( n36017 , n36016 );
not ( n36018 , n36017 );
buf ( n36019 , n36018 );
buf ( n36020 , n36019 );
not ( n36021 , n36020 );
or ( n36022 , n36000 , n36021 );
not ( n36023 , n35634 );
not ( n36024 , n34833 );
buf ( n36025 , n35416 );
and ( n36026 , n36024 , n36025 );
xor ( n36027 , n35418 , n35616 );
buf ( n36028 , n36027 );
and ( n36029 , n36028 , n34833 );
or ( n36030 , n36026 , n36029 );
buf ( n36031 , n36030 );
buf ( n36032 , n36031 );
and ( n36033 , n36023 , n36032 );
not ( n36034 , n36032 );
and ( n36035 , n36012 , n36013 );
xor ( n36036 , n36034 , n36035 );
and ( n36037 , n36036 , n35634 );
or ( n36038 , n36033 , n36037 );
buf ( n36039 , n36038 );
not ( n36040 , n36039 );
buf ( n36041 , n36040 );
buf ( n36042 , n36041 );
not ( n36043 , n36042 );
or ( n36044 , n36022 , n36043 );
not ( n36045 , n35634 );
not ( n36046 , n34833 );
buf ( n36047 , n35403 );
and ( n36048 , n36046 , n36047 );
xor ( n36049 , n35405 , n35617 );
buf ( n36050 , n36049 );
and ( n36051 , n36050 , n34833 );
or ( n36052 , n36048 , n36051 );
buf ( n36053 , n36052 );
buf ( n36054 , n36053 );
and ( n36055 , n36045 , n36054 );
not ( n36056 , n36054 );
and ( n36057 , n36034 , n36035 );
xor ( n36058 , n36056 , n36057 );
and ( n36059 , n36058 , n35634 );
or ( n36060 , n36055 , n36059 );
buf ( n36061 , n36060 );
not ( n36062 , n36061 );
buf ( n36063 , n36062 );
buf ( n36064 , n36063 );
not ( n36065 , n36064 );
or ( n36066 , n36044 , n36065 );
not ( n36067 , n35634 );
not ( n36068 , n34833 );
buf ( n36069 , n35390 );
and ( n36070 , n36068 , n36069 );
xor ( n36071 , n35392 , n35618 );
buf ( n36072 , n36071 );
and ( n36073 , n36072 , n34833 );
or ( n36074 , n36070 , n36073 );
buf ( n36075 , n36074 );
buf ( n36076 , n36075 );
and ( n36077 , n36067 , n36076 );
not ( n36078 , n36076 );
and ( n36079 , n36056 , n36057 );
xor ( n36080 , n36078 , n36079 );
and ( n36081 , n36080 , n35634 );
or ( n36082 , n36077 , n36081 );
buf ( n36083 , n36082 );
not ( n36084 , n36083 );
buf ( n36085 , n36084 );
buf ( n36086 , n36085 );
not ( n36087 , n36086 );
or ( n36088 , n36066 , n36087 );
not ( n36089 , n35634 );
not ( n36090 , n34833 );
buf ( n36091 , n35377 );
and ( n36092 , n36090 , n36091 );
xor ( n36093 , n35379 , n35619 );
buf ( n36094 , n36093 );
and ( n36095 , n36094 , n34833 );
or ( n36096 , n36092 , n36095 );
buf ( n36097 , n36096 );
buf ( n36098 , n36097 );
and ( n36099 , n36089 , n36098 );
not ( n36100 , n36098 );
and ( n36101 , n36078 , n36079 );
xor ( n36102 , n36100 , n36101 );
and ( n36103 , n36102 , n35634 );
or ( n36104 , n36099 , n36103 );
buf ( n36105 , n36104 );
not ( n36106 , n36105 );
buf ( n36107 , n36106 );
buf ( n36108 , n36107 );
not ( n36109 , n36108 );
or ( n36110 , n36088 , n36109 );
not ( n36111 , n35634 );
not ( n36112 , n34833 );
buf ( n36113 , n35364 );
and ( n36114 , n36112 , n36113 );
xor ( n36115 , n35366 , n35620 );
buf ( n36116 , n36115 );
and ( n36117 , n36116 , n34833 );
or ( n36118 , n36114 , n36117 );
buf ( n36119 , n36118 );
buf ( n36120 , n36119 );
and ( n36121 , n36111 , n36120 );
not ( n36122 , n36120 );
and ( n36123 , n36100 , n36101 );
xor ( n36124 , n36122 , n36123 );
and ( n36125 , n36124 , n35634 );
or ( n36126 , n36121 , n36125 );
buf ( n36127 , n36126 );
not ( n36128 , n36127 );
buf ( n36129 , n36128 );
buf ( n36130 , n36129 );
not ( n36131 , n36130 );
or ( n36132 , n36110 , n36131 );
not ( n36133 , n35634 );
not ( n36134 , n34833 );
buf ( n36135 , n35351 );
and ( n36136 , n36134 , n36135 );
xor ( n36137 , n35353 , n35621 );
buf ( n36138 , n36137 );
and ( n36139 , n36138 , n34833 );
or ( n36140 , n36136 , n36139 );
buf ( n36141 , n36140 );
buf ( n36142 , n36141 );
and ( n36143 , n36133 , n36142 );
not ( n36144 , n36142 );
and ( n36145 , n36122 , n36123 );
xor ( n36146 , n36144 , n36145 );
and ( n36147 , n36146 , n35634 );
or ( n36148 , n36143 , n36147 );
buf ( n36149 , n36148 );
not ( n36150 , n36149 );
buf ( n36151 , n36150 );
buf ( n36152 , n36151 );
not ( n36153 , n36152 );
or ( n36154 , n36132 , n36153 );
not ( n36155 , n35634 );
not ( n36156 , n34833 );
buf ( n36157 , n35338 );
and ( n36158 , n36156 , n36157 );
xor ( n36159 , n35340 , n35622 );
buf ( n36160 , n36159 );
and ( n36161 , n36160 , n34833 );
or ( n36162 , n36158 , n36161 );
buf ( n36163 , n36162 );
buf ( n36164 , n36163 );
and ( n36165 , n36155 , n36164 );
not ( n36166 , n36164 );
and ( n36167 , n36144 , n36145 );
xor ( n36168 , n36166 , n36167 );
and ( n36169 , n36168 , n35634 );
or ( n36170 , n36165 , n36169 );
buf ( n36171 , n36170 );
not ( n36172 , n36171 );
buf ( n36173 , n36172 );
buf ( n36174 , n36173 );
not ( n36175 , n36174 );
or ( n36176 , n36154 , n36175 );
not ( n36177 , n35634 );
not ( n36178 , n34833 );
buf ( n36179 , n35325 );
and ( n36180 , n36178 , n36179 );
xor ( n36181 , n35327 , n35623 );
buf ( n36182 , n36181 );
and ( n36183 , n36182 , n34833 );
or ( n36184 , n36180 , n36183 );
buf ( n36185 , n36184 );
buf ( n36186 , n36185 );
and ( n36187 , n36177 , n36186 );
not ( n36188 , n36186 );
and ( n36189 , n36166 , n36167 );
xor ( n36190 , n36188 , n36189 );
and ( n36191 , n36190 , n35634 );
or ( n36192 , n36187 , n36191 );
buf ( n36193 , n36192 );
not ( n36194 , n36193 );
buf ( n36195 , n36194 );
buf ( n36196 , n36195 );
not ( n36197 , n36196 );
or ( n36198 , n36176 , n36197 );
not ( n36199 , n35634 );
not ( n36200 , n34833 );
buf ( n36201 , n35312 );
and ( n36202 , n36200 , n36201 );
xor ( n36203 , n35314 , n35624 );
buf ( n36204 , n36203 );
and ( n36205 , n36204 , n34833 );
or ( n36206 , n36202 , n36205 );
buf ( n36207 , n36206 );
buf ( n36208 , n36207 );
and ( n36209 , n36199 , n36208 );
not ( n36210 , n36208 );
and ( n36211 , n36188 , n36189 );
xor ( n36212 , n36210 , n36211 );
and ( n36213 , n36212 , n35634 );
or ( n36214 , n36209 , n36213 );
buf ( n36215 , n36214 );
not ( n36216 , n36215 );
buf ( n36217 , n36216 );
buf ( n36218 , n36217 );
not ( n36219 , n36218 );
or ( n36220 , n36198 , n36219 );
not ( n36221 , n35634 );
not ( n36222 , n34833 );
buf ( n36223 , n35299 );
and ( n36224 , n36222 , n36223 );
xor ( n36225 , n35301 , n35625 );
buf ( n36226 , n36225 );
and ( n36227 , n36226 , n34833 );
or ( n36228 , n36224 , n36227 );
buf ( n36229 , n36228 );
buf ( n36230 , n36229 );
and ( n36231 , n36221 , n36230 );
not ( n36232 , n36230 );
and ( n36233 , n36210 , n36211 );
xor ( n36234 , n36232 , n36233 );
and ( n36235 , n36234 , n35634 );
or ( n36236 , n36231 , n36235 );
buf ( n36237 , n36236 );
not ( n36238 , n36237 );
buf ( n36239 , n36238 );
buf ( n36240 , n36239 );
not ( n36241 , n36240 );
or ( n36242 , n36220 , n36241 );
buf ( n36243 , n36242 );
buf ( n36244 , n36243 );
and ( n36245 , n36244 , n35634 );
not ( n36246 , n36245 );
and ( n36247 , n36246 , n35779 );
xor ( n36248 , n35779 , n35634 );
xor ( n36249 , n35765 , n35634 );
xor ( n36250 , n35743 , n35634 );
xor ( n36251 , n35721 , n35634 );
xor ( n36252 , n35699 , n35634 );
xor ( n36253 , n35677 , n35634 );
xor ( n36254 , n35655 , n35634 );
xor ( n36255 , n35196 , n35634 );
and ( n36256 , n36255 , n35634 );
and ( n36257 , n36254 , n36256 );
and ( n36258 , n36253 , n36257 );
and ( n36259 , n36252 , n36258 );
and ( n36260 , n36251 , n36259 );
and ( n36261 , n36250 , n36260 );
and ( n36262 , n36249 , n36261 );
xor ( n36263 , n36248 , n36262 );
and ( n36264 , n36263 , n36245 );
or ( n36265 , n36247 , n36264 );
buf ( n36266 , n36265 );
and ( n36267 , n36266 , n14139 );
or ( n36268 , n35189 , n36267 );
and ( n36269 , n36268 , n14140 );
and ( n36270 , n35188 , n14141 );
or ( n36271 , n34829 , n34830 , n36269 , n36270 );
not ( n36272 , n12226 );
not ( n36273 , n12242 );
nor ( n36274 , n36272 , n12234 , n36273 );
not ( n36275 , n36274 );
nor ( n36276 , n12226 , n12234 , n36273 );
not ( n36277 , n36276 );
and ( n36278 , n12226 , n12234 , n36273 );
not ( n36279 , n36278 );
and ( n36280 , n36272 , n12234 , n36273 );
not ( n36281 , n36280 );
nor ( n36282 , n36272 , n12234 , n12242 );
not ( n36283 , n36282 );
nor ( n36284 , n12226 , n12234 , n12242 );
not ( n36285 , n36284 );
buf ( n36286 , RI21077000_517);
and ( n36287 , n36285 , n36286 );
or ( n36288 , n36287 , C0 );
and ( n36289 , n36283 , n36288 );
and ( n36290 , C1 , n36282 );
or ( n36291 , n36289 , n36290 );
and ( n36292 , n36281 , n36291 );
or ( n36293 , n36292 , C0 );
and ( n36294 , n36279 , n36293 );
and ( n36295 , C1 , n36278 );
or ( n36296 , n36294 , n36295 );
and ( n36297 , n36277 , n36296 );
not ( n36298 , n14139 );
and ( n36299 , n36298 , n36286 );
and ( n36300 , C1 , n14139 );
or ( n36301 , n36299 , n36300 );
and ( n36302 , n36301 , n36276 );
or ( n36303 , n36297 , n36302 );
and ( n36304 , n36275 , n36303 );
not ( n36305 , n14139 );
not ( n36306 , n36305 );
and ( n36307 , n36306 , n36286 );
and ( n36308 , C1 , n36305 );
or ( n36309 , n36307 , n36308 );
and ( n36310 , n36309 , n36274 );
or ( n36311 , n36304 , n36310 );
not ( n36312 , n36311 );
not ( n36313 , n36274 );
not ( n36314 , n36276 );
not ( n36315 , n36278 );
not ( n36316 , n36280 );
not ( n36317 , n36282 );
not ( n36318 , n36284 );
buf ( n36319 , RI21076538_518);
and ( n36320 , n36318 , n36319 );
or ( n36321 , n36320 , C0 );
and ( n36322 , n36317 , n36321 );
or ( n36323 , n36322 , C0 );
and ( n36324 , n36316 , n36323 );
and ( n36325 , C1 , n36280 );
or ( n36326 , n36324 , n36325 );
and ( n36327 , n36315 , n36326 );
and ( n36328 , C1 , n36278 );
or ( n36329 , n36327 , n36328 );
and ( n36330 , n36314 , n36329 );
not ( n36331 , n14139 );
and ( n36332 , n36331 , n36319 );
and ( n36333 , C1 , n14139 );
or ( n36334 , n36332 , n36333 );
and ( n36335 , n36334 , n36276 );
or ( n36336 , n36330 , n36335 );
and ( n36337 , n36313 , n36336 );
not ( n36338 , n36305 );
and ( n36339 , n36338 , n36319 );
and ( n36340 , C1 , n36305 );
or ( n36341 , n36339 , n36340 );
and ( n36342 , n36341 , n36274 );
or ( n36343 , n36337 , n36342 );
not ( n36344 , n36343 );
nor ( n36345 , n36312 , n36344 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
and ( n36346 , n36271 , n36345 );
nor ( n36347 , n36311 , n36344 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
nor ( n36348 , n36312 , n36343 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
or ( n36349 , n36347 , n36348 );
nor ( n36350 , n36311 , n36343 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 , C0 );
or ( n36351 , n36349 , n36350 );
or ( n36352 , n36351 , C0 );
and ( n36353 , n13413 , n36352 );
or ( n36354 , n36346 , n36353 );
and ( n36355 , n36354 , n14562 );
buf ( n36356 , n13514 );
buf ( n36357 , n15866 );
xor ( n36358 , n36356 , n36357 );
buf ( n36359 , n36358 );
buf ( n36360 , n36359 );
buf ( n36361 , n36360 );
not ( n36362 , n36361 );
buf ( n36363 , n36362 );
buf ( n36364 , n36363 );
not ( n36365 , n36364 );
buf ( n36366 , n13150 );
buf ( n36367 , n14934 );
xor ( n36368 , n36366 , n36367 );
buf ( n36369 , n14611 );
buf ( n36370 , n14952 );
and ( n36371 , n36369 , n36370 );
buf ( n36372 , n14964 );
buf ( n36373 , n14977 );
and ( n36374 , n36372 , n36373 );
buf ( n36375 , n13162 );
buf ( n36376 , n14992 );
and ( n36377 , n36375 , n36376 );
buf ( n36378 , n13175 );
buf ( n36379 , n15007 );
and ( n36380 , n36378 , n36379 );
buf ( n36381 , n13187 );
buf ( n36382 , n15022 );
and ( n36383 , n36381 , n36382 );
buf ( n36384 , n13199 );
buf ( n36385 , n15037 );
and ( n36386 , n36384 , n36385 );
buf ( n36387 , n13211 );
buf ( n36388 , n15052 );
and ( n36389 , n36387 , n36388 );
buf ( n36390 , n13223 );
buf ( n36391 , n15067 );
and ( n36392 , n36390 , n36391 );
buf ( n36393 , n13235 );
buf ( n36394 , n15082 );
and ( n36395 , n36393 , n36394 );
buf ( n36396 , n13247 );
buf ( n36397 , n15097 );
and ( n36398 , n36396 , n36397 );
buf ( n36399 , n13259 );
buf ( n36400 , n15112 );
and ( n36401 , n36399 , n36400 );
buf ( n36402 , n13271 );
buf ( n36403 , n15449 );
and ( n36404 , n36402 , n36403 );
buf ( n36405 , n13283 );
buf ( n36406 , n15471 );
and ( n36407 , n36405 , n36406 );
buf ( n36408 , n13295 );
buf ( n36409 , n15493 );
and ( n36410 , n36408 , n36409 );
buf ( n36411 , n13307 );
buf ( n36412 , n15515 );
and ( n36413 , n36411 , n36412 );
buf ( n36414 , n13319 );
buf ( n36415 , n15537 );
and ( n36416 , n36414 , n36415 );
buf ( n36417 , n13331 );
buf ( n36418 , n15559 );
and ( n36419 , n36417 , n36418 );
buf ( n36420 , n13343 );
buf ( n36421 , n15581 );
and ( n36422 , n36420 , n36421 );
buf ( n36423 , n13355 );
buf ( n36424 , n15603 );
and ( n36425 , n36423 , n36424 );
buf ( n36426 , n13367 );
buf ( n36427 , n15625 );
and ( n36428 , n36426 , n36427 );
buf ( n36429 , n13379 );
buf ( n36430 , n15647 );
and ( n36431 , n36429 , n36430 );
buf ( n36432 , n13391 );
buf ( n36433 , n15669 );
and ( n36434 , n36432 , n36433 );
buf ( n36435 , n13403 );
buf ( n36436 , n15691 );
and ( n36437 , n36435 , n36436 );
buf ( n36438 , n13415 );
buf ( n36439 , n15713 );
and ( n36440 , n36438 , n36439 );
buf ( n36441 , n13427 );
buf ( n36442 , n15735 );
and ( n36443 , n36441 , n36442 );
buf ( n36444 , n13439 );
buf ( n36445 , n15757 );
and ( n36446 , n36444 , n36445 );
buf ( n36447 , n13451 );
buf ( n36448 , n15779 );
and ( n36449 , n36447 , n36448 );
buf ( n36450 , n13463 );
buf ( n36451 , n15801 );
and ( n36452 , n36450 , n36451 );
buf ( n36453 , n13480 );
buf ( n36454 , n15823 );
and ( n36455 , n36453 , n36454 );
buf ( n36456 , n13497 );
buf ( n36457 , n15845 );
and ( n36458 , n36456 , n36457 );
and ( n36459 , n36356 , n36357 );
and ( n36460 , n36457 , n36459 );
and ( n36461 , n36456 , n36459 );
or ( n36462 , n36458 , n36460 , n36461 );
and ( n36463 , n36454 , n36462 );
and ( n36464 , n36453 , n36462 );
or ( n36465 , n36455 , n36463 , n36464 );
and ( n36466 , n36451 , n36465 );
and ( n36467 , n36450 , n36465 );
or ( n36468 , n36452 , n36466 , n36467 );
and ( n36469 , n36448 , n36468 );
and ( n36470 , n36447 , n36468 );
or ( n36471 , n36449 , n36469 , n36470 );
and ( n36472 , n36445 , n36471 );
and ( n36473 , n36444 , n36471 );
or ( n36474 , n36446 , n36472 , n36473 );
and ( n36475 , n36442 , n36474 );
and ( n36476 , n36441 , n36474 );
or ( n36477 , n36443 , n36475 , n36476 );
and ( n36478 , n36439 , n36477 );
and ( n36479 , n36438 , n36477 );
or ( n36480 , n36440 , n36478 , n36479 );
and ( n36481 , n36436 , n36480 );
and ( n36482 , n36435 , n36480 );
or ( n36483 , n36437 , n36481 , n36482 );
and ( n36484 , n36433 , n36483 );
and ( n36485 , n36432 , n36483 );
or ( n36486 , n36434 , n36484 , n36485 );
and ( n36487 , n36430 , n36486 );
and ( n36488 , n36429 , n36486 );
or ( n36489 , n36431 , n36487 , n36488 );
and ( n36490 , n36427 , n36489 );
and ( n36491 , n36426 , n36489 );
or ( n36492 , n36428 , n36490 , n36491 );
and ( n36493 , n36424 , n36492 );
and ( n36494 , n36423 , n36492 );
or ( n36495 , n36425 , n36493 , n36494 );
and ( n36496 , n36421 , n36495 );
and ( n36497 , n36420 , n36495 );
or ( n36498 , n36422 , n36496 , n36497 );
and ( n36499 , n36418 , n36498 );
and ( n36500 , n36417 , n36498 );
or ( n36501 , n36419 , n36499 , n36500 );
and ( n36502 , n36415 , n36501 );
and ( n36503 , n36414 , n36501 );
or ( n36504 , n36416 , n36502 , n36503 );
and ( n36505 , n36412 , n36504 );
and ( n36506 , n36411 , n36504 );
or ( n36507 , n36413 , n36505 , n36506 );
and ( n36508 , n36409 , n36507 );
and ( n36509 , n36408 , n36507 );
or ( n36510 , n36410 , n36508 , n36509 );
and ( n36511 , n36406 , n36510 );
and ( n36512 , n36405 , n36510 );
or ( n36513 , n36407 , n36511 , n36512 );
and ( n36514 , n36403 , n36513 );
and ( n36515 , n36402 , n36513 );
or ( n36516 , n36404 , n36514 , n36515 );
and ( n36517 , n36400 , n36516 );
and ( n36518 , n36399 , n36516 );
or ( n36519 , n36401 , n36517 , n36518 );
and ( n36520 , n36397 , n36519 );
and ( n36521 , n36396 , n36519 );
or ( n36522 , n36398 , n36520 , n36521 );
and ( n36523 , n36394 , n36522 );
and ( n36524 , n36393 , n36522 );
or ( n36525 , n36395 , n36523 , n36524 );
and ( n36526 , n36391 , n36525 );
and ( n36527 , n36390 , n36525 );
or ( n36528 , n36392 , n36526 , n36527 );
and ( n36529 , n36388 , n36528 );
and ( n36530 , n36387 , n36528 );
or ( n36531 , n36389 , n36529 , n36530 );
and ( n36532 , n36385 , n36531 );
and ( n36533 , n36384 , n36531 );
or ( n36534 , n36386 , n36532 , n36533 );
and ( n36535 , n36382 , n36534 );
and ( n36536 , n36381 , n36534 );
or ( n36537 , n36383 , n36535 , n36536 );
and ( n36538 , n36379 , n36537 );
and ( n36539 , n36378 , n36537 );
or ( n36540 , n36380 , n36538 , n36539 );
and ( n36541 , n36376 , n36540 );
and ( n36542 , n36375 , n36540 );
or ( n36543 , n36377 , n36541 , n36542 );
and ( n36544 , n36373 , n36543 );
and ( n36545 , n36372 , n36543 );
or ( n36546 , n36374 , n36544 , n36545 );
and ( n36547 , n36370 , n36546 );
and ( n36548 , n36369 , n36546 );
or ( n36549 , n36371 , n36547 , n36548 );
xor ( n36550 , n36368 , n36549 );
buf ( n36551 , n36550 );
buf ( n36552 , n36551 );
not ( n36553 , n36552 );
xor ( n36554 , n36456 , n36457 );
xor ( n36555 , n36554 , n36459 );
buf ( n36556 , n36555 );
buf ( n36557 , n36556 );
and ( n36558 , n36553 , n36557 );
not ( n36559 , n36557 );
not ( n36560 , n36360 );
xor ( n36561 , n36559 , n36560 );
and ( n36562 , n36561 , n36552 );
or ( n36563 , n36558 , n36562 );
buf ( n36564 , n36563 );
not ( n36565 , n36564 );
buf ( n36566 , n36565 );
buf ( n36567 , n36566 );
not ( n36568 , n36567 );
or ( n36569 , n36365 , n36568 );
not ( n36570 , n36552 );
xor ( n36571 , n36453 , n36454 );
xor ( n36572 , n36571 , n36462 );
buf ( n36573 , n36572 );
buf ( n36574 , n36573 );
and ( n36575 , n36570 , n36574 );
not ( n36576 , n36574 );
and ( n36577 , n36559 , n36560 );
xor ( n36578 , n36576 , n36577 );
and ( n36579 , n36578 , n36552 );
or ( n36580 , n36575 , n36579 );
buf ( n36581 , n36580 );
not ( n36582 , n36581 );
buf ( n36583 , n36582 );
buf ( n36584 , n36583 );
not ( n36585 , n36584 );
or ( n36586 , n36569 , n36585 );
not ( n36587 , n36552 );
xor ( n36588 , n36450 , n36451 );
xor ( n36589 , n36588 , n36465 );
buf ( n36590 , n36589 );
buf ( n36591 , n36590 );
and ( n36592 , n36587 , n36591 );
not ( n36593 , n36591 );
and ( n36594 , n36576 , n36577 );
xor ( n36595 , n36593 , n36594 );
and ( n36596 , n36595 , n36552 );
or ( n36597 , n36592 , n36596 );
buf ( n36598 , n36597 );
not ( n36599 , n36598 );
buf ( n36600 , n36599 );
buf ( n36601 , n36600 );
not ( n36602 , n36601 );
or ( n36603 , n36586 , n36602 );
not ( n36604 , n36552 );
xor ( n36605 , n36447 , n36448 );
xor ( n36606 , n36605 , n36468 );
buf ( n36607 , n36606 );
buf ( n36608 , n36607 );
and ( n36609 , n36604 , n36608 );
not ( n36610 , n36608 );
and ( n36611 , n36593 , n36594 );
xor ( n36612 , n36610 , n36611 );
and ( n36613 , n36612 , n36552 );
or ( n36614 , n36609 , n36613 );
buf ( n36615 , n36614 );
not ( n36616 , n36615 );
buf ( n36617 , n36616 );
buf ( n36618 , n36617 );
not ( n36619 , n36618 );
or ( n36620 , n36603 , n36619 );
not ( n36621 , n36552 );
xor ( n36622 , n36444 , n36445 );
xor ( n36623 , n36622 , n36471 );
buf ( n36624 , n36623 );
buf ( n36625 , n36624 );
and ( n36626 , n36621 , n36625 );
not ( n36627 , n36625 );
and ( n36628 , n36610 , n36611 );
xor ( n36629 , n36627 , n36628 );
and ( n36630 , n36629 , n36552 );
or ( n36631 , n36626 , n36630 );
buf ( n36632 , n36631 );
not ( n36633 , n36632 );
buf ( n36634 , n36633 );
buf ( n36635 , n36634 );
not ( n36636 , n36635 );
or ( n36637 , n36620 , n36636 );
not ( n36638 , n36552 );
xor ( n36639 , n36441 , n36442 );
xor ( n36640 , n36639 , n36474 );
buf ( n36641 , n36640 );
buf ( n36642 , n36641 );
and ( n36643 , n36638 , n36642 );
not ( n36644 , n36642 );
and ( n36645 , n36627 , n36628 );
xor ( n36646 , n36644 , n36645 );
and ( n36647 , n36646 , n36552 );
or ( n36648 , n36643 , n36647 );
buf ( n36649 , n36648 );
not ( n36650 , n36649 );
buf ( n36651 , n36650 );
buf ( n36652 , n36651 );
not ( n36653 , n36652 );
or ( n36654 , n36637 , n36653 );
not ( n36655 , n36552 );
xor ( n36656 , n36438 , n36439 );
xor ( n36657 , n36656 , n36477 );
buf ( n36658 , n36657 );
buf ( n36659 , n36658 );
and ( n36660 , n36655 , n36659 );
not ( n36661 , n36659 );
and ( n36662 , n36644 , n36645 );
xor ( n36663 , n36661 , n36662 );
and ( n36664 , n36663 , n36552 );
or ( n36665 , n36660 , n36664 );
buf ( n36666 , n36665 );
not ( n36667 , n36666 );
buf ( n36668 , n36667 );
buf ( n36669 , n36668 );
not ( n36670 , n36669 );
or ( n36671 , n36654 , n36670 );
not ( n36672 , n36552 );
xor ( n36673 , n36435 , n36436 );
xor ( n36674 , n36673 , n36480 );
buf ( n36675 , n36674 );
buf ( n36676 , n36675 );
and ( n36677 , n36672 , n36676 );
not ( n36678 , n36676 );
and ( n36679 , n36661 , n36662 );
xor ( n36680 , n36678 , n36679 );
and ( n36681 , n36680 , n36552 );
or ( n36682 , n36677 , n36681 );
buf ( n36683 , n36682 );
not ( n36684 , n36683 );
buf ( n36685 , n36684 );
buf ( n36686 , n36685 );
not ( n36687 , n36686 );
or ( n36688 , n36671 , n36687 );
not ( n36689 , n36552 );
xor ( n36690 , n36432 , n36433 );
xor ( n36691 , n36690 , n36483 );
buf ( n36692 , n36691 );
buf ( n36693 , n36692 );
and ( n36694 , n36689 , n36693 );
not ( n36695 , n36693 );
and ( n36696 , n36678 , n36679 );
xor ( n36697 , n36695 , n36696 );
and ( n36698 , n36697 , n36552 );
or ( n36699 , n36694 , n36698 );
buf ( n36700 , n36699 );
not ( n36701 , n36700 );
buf ( n36702 , n36701 );
buf ( n36703 , n36702 );
not ( n36704 , n36703 );
or ( n36705 , n36688 , n36704 );
not ( n36706 , n36552 );
xor ( n36707 , n36429 , n36430 );
xor ( n36708 , n36707 , n36486 );
buf ( n36709 , n36708 );
buf ( n36710 , n36709 );
and ( n36711 , n36706 , n36710 );
not ( n36712 , n36710 );
and ( n36713 , n36695 , n36696 );
xor ( n36714 , n36712 , n36713 );
and ( n36715 , n36714 , n36552 );
or ( n36716 , n36711 , n36715 );
buf ( n36717 , n36716 );
not ( n36718 , n36717 );
buf ( n36719 , n36718 );
buf ( n36720 , n36719 );
not ( n36721 , n36720 );
or ( n36722 , n36705 , n36721 );
not ( n36723 , n36552 );
xor ( n36724 , n36426 , n36427 );
xor ( n36725 , n36724 , n36489 );
buf ( n36726 , n36725 );
buf ( n36727 , n36726 );
and ( n36728 , n36723 , n36727 );
not ( n36729 , n36727 );
and ( n36730 , n36712 , n36713 );
xor ( n36731 , n36729 , n36730 );
and ( n36732 , n36731 , n36552 );
or ( n36733 , n36728 , n36732 );
buf ( n36734 , n36733 );
not ( n36735 , n36734 );
buf ( n36736 , n36735 );
buf ( n36737 , n36736 );
not ( n36738 , n36737 );
or ( n36739 , n36722 , n36738 );
not ( n36740 , n36552 );
xor ( n36741 , n36423 , n36424 );
xor ( n36742 , n36741 , n36492 );
buf ( n36743 , n36742 );
buf ( n36744 , n36743 );
and ( n36745 , n36740 , n36744 );
not ( n36746 , n36744 );
and ( n36747 , n36729 , n36730 );
xor ( n36748 , n36746 , n36747 );
and ( n36749 , n36748 , n36552 );
or ( n36750 , n36745 , n36749 );
buf ( n36751 , n36750 );
not ( n36752 , n36751 );
buf ( n36753 , n36752 );
buf ( n36754 , n36753 );
not ( n36755 , n36754 );
or ( n36756 , n36739 , n36755 );
not ( n36757 , n36552 );
xor ( n36758 , n36420 , n36421 );
xor ( n36759 , n36758 , n36495 );
buf ( n36760 , n36759 );
buf ( n36761 , n36760 );
and ( n36762 , n36757 , n36761 );
not ( n36763 , n36761 );
and ( n36764 , n36746 , n36747 );
xor ( n36765 , n36763 , n36764 );
and ( n36766 , n36765 , n36552 );
or ( n36767 , n36762 , n36766 );
buf ( n36768 , n36767 );
not ( n36769 , n36768 );
buf ( n36770 , n36769 );
buf ( n36771 , n36770 );
not ( n36772 , n36771 );
or ( n36773 , n36756 , n36772 );
not ( n36774 , n36552 );
xor ( n36775 , n36417 , n36418 );
xor ( n36776 , n36775 , n36498 );
buf ( n36777 , n36776 );
buf ( n36778 , n36777 );
and ( n36779 , n36774 , n36778 );
not ( n36780 , n36778 );
and ( n36781 , n36763 , n36764 );
xor ( n36782 , n36780 , n36781 );
and ( n36783 , n36782 , n36552 );
or ( n36784 , n36779 , n36783 );
buf ( n36785 , n36784 );
not ( n36786 , n36785 );
buf ( n36787 , n36786 );
buf ( n36788 , n36787 );
not ( n36789 , n36788 );
or ( n36790 , n36773 , n36789 );
not ( n36791 , n36552 );
xor ( n36792 , n36414 , n36415 );
xor ( n36793 , n36792 , n36501 );
buf ( n36794 , n36793 );
buf ( n36795 , n36794 );
and ( n36796 , n36791 , n36795 );
not ( n36797 , n36795 );
and ( n36798 , n36780 , n36781 );
xor ( n36799 , n36797 , n36798 );
and ( n36800 , n36799 , n36552 );
or ( n36801 , n36796 , n36800 );
buf ( n36802 , n36801 );
not ( n36803 , n36802 );
buf ( n36804 , n36803 );
buf ( n36805 , n36804 );
not ( n36806 , n36805 );
or ( n36807 , n36790 , n36806 );
not ( n36808 , n36552 );
xor ( n36809 , n36411 , n36412 );
xor ( n36810 , n36809 , n36504 );
buf ( n36811 , n36810 );
buf ( n36812 , n36811 );
and ( n36813 , n36808 , n36812 );
not ( n36814 , n36812 );
and ( n36815 , n36797 , n36798 );
xor ( n36816 , n36814 , n36815 );
and ( n36817 , n36816 , n36552 );
or ( n36818 , n36813 , n36817 );
buf ( n36819 , n36818 );
not ( n36820 , n36819 );
buf ( n36821 , n36820 );
buf ( n36822 , n36821 );
not ( n36823 , n36822 );
or ( n36824 , n36807 , n36823 );
not ( n36825 , n36552 );
xor ( n36826 , n36408 , n36409 );
xor ( n36827 , n36826 , n36507 );
buf ( n36828 , n36827 );
buf ( n36829 , n36828 );
and ( n36830 , n36825 , n36829 );
not ( n36831 , n36829 );
and ( n36832 , n36814 , n36815 );
xor ( n36833 , n36831 , n36832 );
and ( n36834 , n36833 , n36552 );
or ( n36835 , n36830 , n36834 );
buf ( n36836 , n36835 );
not ( n36837 , n36836 );
buf ( n36838 , n36837 );
buf ( n36839 , n36838 );
not ( n36840 , n36839 );
or ( n36841 , n36824 , n36840 );
not ( n36842 , n36552 );
xor ( n36843 , n36405 , n36406 );
xor ( n36844 , n36843 , n36510 );
buf ( n36845 , n36844 );
buf ( n36846 , n36845 );
and ( n36847 , n36842 , n36846 );
not ( n36848 , n36846 );
and ( n36849 , n36831 , n36832 );
xor ( n36850 , n36848 , n36849 );
and ( n36851 , n36850 , n36552 );
or ( n36852 , n36847 , n36851 );
buf ( n36853 , n36852 );
not ( n36854 , n36853 );
buf ( n36855 , n36854 );
buf ( n36856 , n36855 );
not ( n36857 , n36856 );
or ( n36858 , n36841 , n36857 );
not ( n36859 , n36552 );
xor ( n36860 , n36402 , n36403 );
xor ( n36861 , n36860 , n36513 );
buf ( n36862 , n36861 );
buf ( n36863 , n36862 );
and ( n36864 , n36859 , n36863 );
not ( n36865 , n36863 );
and ( n36866 , n36848 , n36849 );
xor ( n36867 , n36865 , n36866 );
and ( n36868 , n36867 , n36552 );
or ( n36869 , n36864 , n36868 );
buf ( n36870 , n36869 );
not ( n36871 , n36870 );
buf ( n36872 , n36871 );
buf ( n36873 , n36872 );
not ( n36874 , n36873 );
or ( n36875 , n36858 , n36874 );
not ( n36876 , n36552 );
xor ( n36877 , n36399 , n36400 );
xor ( n36878 , n36877 , n36516 );
buf ( n36879 , n36878 );
buf ( n36880 , n36879 );
and ( n36881 , n36876 , n36880 );
not ( n36882 , n36880 );
and ( n36883 , n36865 , n36866 );
xor ( n36884 , n36882 , n36883 );
and ( n36885 , n36884 , n36552 );
or ( n36886 , n36881 , n36885 );
buf ( n36887 , n36886 );
not ( n36888 , n36887 );
buf ( n36889 , n36888 );
buf ( n36890 , n36889 );
not ( n36891 , n36890 );
or ( n36892 , n36875 , n36891 );
not ( n36893 , n36552 );
xor ( n36894 , n36396 , n36397 );
xor ( n36895 , n36894 , n36519 );
buf ( n36896 , n36895 );
buf ( n36897 , n36896 );
and ( n36898 , n36893 , n36897 );
not ( n36899 , n36897 );
and ( n36900 , n36882 , n36883 );
xor ( n36901 , n36899 , n36900 );
and ( n36902 , n36901 , n36552 );
or ( n36903 , n36898 , n36902 );
buf ( n36904 , n36903 );
not ( n36905 , n36904 );
buf ( n36906 , n36905 );
buf ( n36907 , n36906 );
not ( n36908 , n36907 );
or ( n36909 , n36892 , n36908 );
not ( n36910 , n36552 );
xor ( n36911 , n36393 , n36394 );
xor ( n36912 , n36911 , n36522 );
buf ( n36913 , n36912 );
buf ( n36914 , n36913 );
and ( n36915 , n36910 , n36914 );
not ( n36916 , n36914 );
and ( n36917 , n36899 , n36900 );
xor ( n36918 , n36916 , n36917 );
and ( n36919 , n36918 , n36552 );
or ( n36920 , n36915 , n36919 );
buf ( n36921 , n36920 );
not ( n36922 , n36921 );
buf ( n36923 , n36922 );
buf ( n36924 , n36923 );
not ( n36925 , n36924 );
or ( n36926 , n36909 , n36925 );
not ( n36927 , n36552 );
xor ( n36928 , n36390 , n36391 );
xor ( n36929 , n36928 , n36525 );
buf ( n36930 , n36929 );
buf ( n36931 , n36930 );
and ( n36932 , n36927 , n36931 );
not ( n36933 , n36931 );
and ( n36934 , n36916 , n36917 );
xor ( n36935 , n36933 , n36934 );
and ( n36936 , n36935 , n36552 );
or ( n36937 , n36932 , n36936 );
buf ( n36938 , n36937 );
not ( n36939 , n36938 );
buf ( n36940 , n36939 );
buf ( n36941 , n36940 );
not ( n36942 , n36941 );
or ( n36943 , n36926 , n36942 );
not ( n36944 , n36552 );
xor ( n36945 , n36387 , n36388 );
xor ( n36946 , n36945 , n36528 );
buf ( n36947 , n36946 );
buf ( n36948 , n36947 );
and ( n36949 , n36944 , n36948 );
not ( n36950 , n36948 );
and ( n36951 , n36933 , n36934 );
xor ( n36952 , n36950 , n36951 );
and ( n36953 , n36952 , n36552 );
or ( n36954 , n36949 , n36953 );
buf ( n36955 , n36954 );
not ( n36956 , n36955 );
buf ( n36957 , n36956 );
buf ( n36958 , n36957 );
not ( n36959 , n36958 );
or ( n36960 , n36943 , n36959 );
not ( n36961 , n36552 );
xor ( n36962 , n36384 , n36385 );
xor ( n36963 , n36962 , n36531 );
buf ( n36964 , n36963 );
buf ( n36965 , n36964 );
and ( n36966 , n36961 , n36965 );
not ( n36967 , n36965 );
and ( n36968 , n36950 , n36951 );
xor ( n36969 , n36967 , n36968 );
and ( n36970 , n36969 , n36552 );
or ( n36971 , n36966 , n36970 );
buf ( n36972 , n36971 );
not ( n36973 , n36972 );
buf ( n36974 , n36973 );
buf ( n36975 , n36974 );
not ( n36976 , n36975 );
or ( n36977 , n36960 , n36976 );
not ( n36978 , n36552 );
xor ( n36979 , n36381 , n36382 );
xor ( n36980 , n36979 , n36534 );
buf ( n36981 , n36980 );
buf ( n36982 , n36981 );
and ( n36983 , n36978 , n36982 );
not ( n36984 , n36982 );
and ( n36985 , n36967 , n36968 );
xor ( n36986 , n36984 , n36985 );
and ( n36987 , n36986 , n36552 );
or ( n36988 , n36983 , n36987 );
buf ( n36989 , n36988 );
not ( n36990 , n36989 );
buf ( n36991 , n36990 );
buf ( n36992 , n36991 );
not ( n36993 , n36992 );
or ( n36994 , n36977 , n36993 );
not ( n36995 , n36552 );
xor ( n36996 , n36378 , n36379 );
xor ( n36997 , n36996 , n36537 );
buf ( n36998 , n36997 );
buf ( n36999 , n36998 );
and ( n37000 , n36995 , n36999 );
not ( n37001 , n36999 );
and ( n37002 , n36984 , n36985 );
xor ( n37003 , n37001 , n37002 );
and ( n37004 , n37003 , n36552 );
or ( n37005 , n37000 , n37004 );
buf ( n37006 , n37005 );
not ( n37007 , n37006 );
buf ( n37008 , n37007 );
buf ( n37009 , n37008 );
not ( n37010 , n37009 );
or ( n37011 , n36994 , n37010 );
not ( n37012 , n36552 );
xor ( n37013 , n36375 , n36376 );
xor ( n37014 , n37013 , n36540 );
buf ( n37015 , n37014 );
buf ( n37016 , n37015 );
and ( n37017 , n37012 , n37016 );
not ( n37018 , n37016 );
and ( n37019 , n37001 , n37002 );
xor ( n37020 , n37018 , n37019 );
and ( n37021 , n37020 , n36552 );
or ( n37022 , n37017 , n37021 );
buf ( n37023 , n37022 );
not ( n37024 , n37023 );
buf ( n37025 , n37024 );
buf ( n37026 , n37025 );
not ( n37027 , n37026 );
or ( n37028 , n37011 , n37027 );
not ( n37029 , n36552 );
xor ( n37030 , n36372 , n36373 );
xor ( n37031 , n37030 , n36543 );
buf ( n37032 , n37031 );
buf ( n37033 , n37032 );
and ( n37034 , n37029 , n37033 );
not ( n37035 , n37033 );
and ( n37036 , n37018 , n37019 );
xor ( n37037 , n37035 , n37036 );
and ( n37038 , n37037 , n36552 );
or ( n37039 , n37034 , n37038 );
buf ( n37040 , n37039 );
not ( n37041 , n37040 );
buf ( n37042 , n37041 );
buf ( n37043 , n37042 );
not ( n37044 , n37043 );
or ( n37045 , n37028 , n37044 );
or ( n37046 , n37045 , C0 );
buf ( n37047 , n37046 );
and ( n37048 , n37047 , n36552 );
not ( n37049 , n37048 );
and ( n37050 , n37049 , n36670 );
xor ( n37051 , n36670 , n36552 );
xor ( n37052 , n36653 , n36552 );
xor ( n37053 , n36636 , n36552 );
xor ( n37054 , n36619 , n36552 );
xor ( n37055 , n36602 , n36552 );
xor ( n37056 , n36585 , n36552 );
xor ( n37057 , n36568 , n36552 );
xor ( n37058 , n36365 , n36552 );
and ( n37059 , n37058 , n36552 );
and ( n37060 , n37057 , n37059 );
and ( n37061 , n37056 , n37060 );
and ( n37062 , n37055 , n37061 );
and ( n37063 , n37054 , n37062 );
and ( n37064 , n37053 , n37063 );
and ( n37065 , n37052 , n37064 );
xor ( n37066 , n37051 , n37065 );
and ( n37067 , n37066 , n37048 );
or ( n37068 , n37050 , n37067 );
buf ( n37069 , n37068 );
and ( n37070 , n37069 , n36345 );
or ( n37071 , n36348 , n36347 );
or ( n37072 , n37071 , n36350 );
or ( n37073 , n37072 , C0 );
and ( n37074 , n13413 , n37073 );
or ( n37075 , n37070 , n37074 );
and ( n37076 , n37075 , n14586 );
buf ( n37077 , n13514 );
buf ( n37078 , n15866 );
xor ( n37079 , n37077 , n37078 );
buf ( n37080 , n37079 );
buf ( n37081 , n37080 );
buf ( n37082 , n37081 );
not ( n37083 , n37082 );
buf ( n37084 , n37083 );
buf ( n37085 , n37084 );
not ( n37086 , n37085 );
buf ( n37087 , n13150 );
buf ( n37088 , n14934 );
not ( n37089 , n37088 );
xor ( n37090 , n37087 , n37089 );
buf ( n37091 , n14611 );
buf ( n37092 , n14952 );
not ( n37093 , n37092 );
and ( n37094 , n37091 , n37093 );
buf ( n37095 , n14964 );
buf ( n37096 , n14977 );
not ( n37097 , n37096 );
and ( n37098 , n37095 , n37097 );
buf ( n37099 , n13162 );
buf ( n37100 , n14992 );
not ( n37101 , n37100 );
and ( n37102 , n37099 , n37101 );
buf ( n37103 , n13175 );
buf ( n37104 , n15007 );
not ( n37105 , n37104 );
and ( n37106 , n37103 , n37105 );
buf ( n37107 , n13187 );
buf ( n37108 , n15022 );
not ( n37109 , n37108 );
and ( n37110 , n37107 , n37109 );
buf ( n37111 , n13199 );
buf ( n37112 , n15037 );
not ( n37113 , n37112 );
and ( n37114 , n37111 , n37113 );
buf ( n37115 , n13211 );
buf ( n37116 , n15052 );
not ( n37117 , n37116 );
and ( n37118 , n37115 , n37117 );
buf ( n37119 , n13223 );
buf ( n37120 , n15067 );
not ( n37121 , n37120 );
and ( n37122 , n37119 , n37121 );
buf ( n37123 , n13235 );
buf ( n37124 , n15082 );
not ( n37125 , n37124 );
and ( n37126 , n37123 , n37125 );
buf ( n37127 , n13247 );
buf ( n37128 , n15097 );
not ( n37129 , n37128 );
and ( n37130 , n37127 , n37129 );
buf ( n37131 , n13259 );
buf ( n37132 , n15112 );
not ( n37133 , n37132 );
and ( n37134 , n37131 , n37133 );
buf ( n37135 , n13271 );
buf ( n37136 , n15449 );
not ( n37137 , n37136 );
and ( n37138 , n37135 , n37137 );
buf ( n37139 , n13283 );
buf ( n37140 , n15471 );
not ( n37141 , n37140 );
and ( n37142 , n37139 , n37141 );
buf ( n37143 , n13295 );
buf ( n37144 , n15493 );
not ( n37145 , n37144 );
and ( n37146 , n37143 , n37145 );
buf ( n37147 , n13307 );
buf ( n37148 , n15515 );
not ( n37149 , n37148 );
and ( n37150 , n37147 , n37149 );
buf ( n37151 , n13319 );
buf ( n37152 , n15537 );
not ( n37153 , n37152 );
and ( n37154 , n37151 , n37153 );
buf ( n37155 , n13331 );
buf ( n37156 , n15559 );
not ( n37157 , n37156 );
and ( n37158 , n37155 , n37157 );
buf ( n37159 , n13343 );
buf ( n37160 , n15581 );
not ( n37161 , n37160 );
and ( n37162 , n37159 , n37161 );
buf ( n37163 , n13355 );
buf ( n37164 , n15603 );
not ( n37165 , n37164 );
and ( n37166 , n37163 , n37165 );
buf ( n37167 , n13367 );
buf ( n37168 , n15625 );
not ( n37169 , n37168 );
and ( n37170 , n37167 , n37169 );
buf ( n37171 , n13379 );
buf ( n37172 , n15647 );
not ( n37173 , n37172 );
and ( n37174 , n37171 , n37173 );
buf ( n37175 , n13391 );
buf ( n37176 , n15669 );
not ( n37177 , n37176 );
and ( n37178 , n37175 , n37177 );
buf ( n37179 , n13403 );
buf ( n37180 , n15691 );
not ( n37181 , n37180 );
and ( n37182 , n37179 , n37181 );
buf ( n37183 , n13415 );
buf ( n37184 , n15713 );
not ( n37185 , n37184 );
and ( n37186 , n37183 , n37185 );
buf ( n37187 , n13427 );
buf ( n37188 , n15735 );
not ( n37189 , n37188 );
and ( n37190 , n37187 , n37189 );
buf ( n37191 , n13439 );
buf ( n37192 , n15757 );
not ( n37193 , n37192 );
and ( n37194 , n37191 , n37193 );
buf ( n37195 , n13451 );
buf ( n37196 , n15779 );
not ( n37197 , n37196 );
and ( n37198 , n37195 , n37197 );
buf ( n37199 , n13463 );
buf ( n37200 , n15801 );
not ( n37201 , n37200 );
and ( n37202 , n37199 , n37201 );
buf ( n37203 , n13480 );
buf ( n37204 , n15823 );
not ( n37205 , n37204 );
and ( n37206 , n37203 , n37205 );
buf ( n37207 , n13497 );
buf ( n37208 , n15845 );
not ( n37209 , n37208 );
and ( n37210 , n37207 , n37209 );
not ( n37211 , n37078 );
or ( n37212 , n37077 , n37211 );
and ( n37213 , n37209 , n37212 );
and ( n37214 , n37207 , n37212 );
or ( n37215 , n37210 , n37213 , n37214 );
and ( n37216 , n37205 , n37215 );
and ( n37217 , n37203 , n37215 );
or ( n37218 , n37206 , n37216 , n37217 );
and ( n37219 , n37201 , n37218 );
and ( n37220 , n37199 , n37218 );
or ( n37221 , n37202 , n37219 , n37220 );
and ( n37222 , n37197 , n37221 );
and ( n37223 , n37195 , n37221 );
or ( n37224 , n37198 , n37222 , n37223 );
and ( n37225 , n37193 , n37224 );
and ( n37226 , n37191 , n37224 );
or ( n37227 , n37194 , n37225 , n37226 );
and ( n37228 , n37189 , n37227 );
and ( n37229 , n37187 , n37227 );
or ( n37230 , n37190 , n37228 , n37229 );
and ( n37231 , n37185 , n37230 );
and ( n37232 , n37183 , n37230 );
or ( n37233 , n37186 , n37231 , n37232 );
and ( n37234 , n37181 , n37233 );
and ( n37235 , n37179 , n37233 );
or ( n37236 , n37182 , n37234 , n37235 );
and ( n37237 , n37177 , n37236 );
and ( n37238 , n37175 , n37236 );
or ( n37239 , n37178 , n37237 , n37238 );
and ( n37240 , n37173 , n37239 );
and ( n37241 , n37171 , n37239 );
or ( n37242 , n37174 , n37240 , n37241 );
and ( n37243 , n37169 , n37242 );
and ( n37244 , n37167 , n37242 );
or ( n37245 , n37170 , n37243 , n37244 );
and ( n37246 , n37165 , n37245 );
and ( n37247 , n37163 , n37245 );
or ( n37248 , n37166 , n37246 , n37247 );
and ( n37249 , n37161 , n37248 );
and ( n37250 , n37159 , n37248 );
or ( n37251 , n37162 , n37249 , n37250 );
and ( n37252 , n37157 , n37251 );
and ( n37253 , n37155 , n37251 );
or ( n37254 , n37158 , n37252 , n37253 );
and ( n37255 , n37153 , n37254 );
and ( n37256 , n37151 , n37254 );
or ( n37257 , n37154 , n37255 , n37256 );
and ( n37258 , n37149 , n37257 );
and ( n37259 , n37147 , n37257 );
or ( n37260 , n37150 , n37258 , n37259 );
and ( n37261 , n37145 , n37260 );
and ( n37262 , n37143 , n37260 );
or ( n37263 , n37146 , n37261 , n37262 );
and ( n37264 , n37141 , n37263 );
and ( n37265 , n37139 , n37263 );
or ( n37266 , n37142 , n37264 , n37265 );
and ( n37267 , n37137 , n37266 );
and ( n37268 , n37135 , n37266 );
or ( n37269 , n37138 , n37267 , n37268 );
and ( n37270 , n37133 , n37269 );
and ( n37271 , n37131 , n37269 );
or ( n37272 , n37134 , n37270 , n37271 );
and ( n37273 , n37129 , n37272 );
and ( n37274 , n37127 , n37272 );
or ( n37275 , n37130 , n37273 , n37274 );
and ( n37276 , n37125 , n37275 );
and ( n37277 , n37123 , n37275 );
or ( n37278 , n37126 , n37276 , n37277 );
and ( n37279 , n37121 , n37278 );
and ( n37280 , n37119 , n37278 );
or ( n37281 , n37122 , n37279 , n37280 );
and ( n37282 , n37117 , n37281 );
and ( n37283 , n37115 , n37281 );
or ( n37284 , n37118 , n37282 , n37283 );
and ( n37285 , n37113 , n37284 );
and ( n37286 , n37111 , n37284 );
or ( n37287 , n37114 , n37285 , n37286 );
and ( n37288 , n37109 , n37287 );
and ( n37289 , n37107 , n37287 );
or ( n37290 , n37110 , n37288 , n37289 );
and ( n37291 , n37105 , n37290 );
and ( n37292 , n37103 , n37290 );
or ( n37293 , n37106 , n37291 , n37292 );
and ( n37294 , n37101 , n37293 );
and ( n37295 , n37099 , n37293 );
or ( n37296 , n37102 , n37294 , n37295 );
and ( n37297 , n37097 , n37296 );
and ( n37298 , n37095 , n37296 );
or ( n37299 , n37098 , n37297 , n37298 );
and ( n37300 , n37093 , n37299 );
and ( n37301 , n37091 , n37299 );
or ( n37302 , n37094 , n37300 , n37301 );
xor ( n37303 , n37090 , n37302 );
buf ( n37304 , n37303 );
buf ( n37305 , n37304 );
not ( n37306 , n37305 );
xor ( n37307 , n37207 , n37209 );
xor ( n37308 , n37307 , n37212 );
buf ( n37309 , n37308 );
buf ( n37310 , n37309 );
and ( n37311 , n37306 , n37310 );
not ( n37312 , n37310 );
not ( n37313 , n37081 );
xor ( n37314 , n37312 , n37313 );
and ( n37315 , n37314 , n37305 );
or ( n37316 , n37311 , n37315 );
buf ( n37317 , n37316 );
not ( n37318 , n37317 );
buf ( n37319 , n37318 );
buf ( n37320 , n37319 );
not ( n37321 , n37320 );
or ( n37322 , n37086 , n37321 );
not ( n37323 , n37305 );
xor ( n37324 , n37203 , n37205 );
xor ( n37325 , n37324 , n37215 );
buf ( n37326 , n37325 );
buf ( n37327 , n37326 );
and ( n37328 , n37323 , n37327 );
not ( n37329 , n37327 );
and ( n37330 , n37312 , n37313 );
xor ( n37331 , n37329 , n37330 );
and ( n37332 , n37331 , n37305 );
or ( n37333 , n37328 , n37332 );
buf ( n37334 , n37333 );
not ( n37335 , n37334 );
buf ( n37336 , n37335 );
buf ( n37337 , n37336 );
not ( n37338 , n37337 );
or ( n37339 , n37322 , n37338 );
not ( n37340 , n37305 );
xor ( n37341 , n37199 , n37201 );
xor ( n37342 , n37341 , n37218 );
buf ( n37343 , n37342 );
buf ( n37344 , n37343 );
and ( n37345 , n37340 , n37344 );
not ( n37346 , n37344 );
and ( n37347 , n37329 , n37330 );
xor ( n37348 , n37346 , n37347 );
and ( n37349 , n37348 , n37305 );
or ( n37350 , n37345 , n37349 );
buf ( n37351 , n37350 );
not ( n37352 , n37351 );
buf ( n37353 , n37352 );
buf ( n37354 , n37353 );
not ( n37355 , n37354 );
or ( n37356 , n37339 , n37355 );
not ( n37357 , n37305 );
xor ( n37358 , n37195 , n37197 );
xor ( n37359 , n37358 , n37221 );
buf ( n37360 , n37359 );
buf ( n37361 , n37360 );
and ( n37362 , n37357 , n37361 );
not ( n37363 , n37361 );
and ( n37364 , n37346 , n37347 );
xor ( n37365 , n37363 , n37364 );
and ( n37366 , n37365 , n37305 );
or ( n37367 , n37362 , n37366 );
buf ( n37368 , n37367 );
not ( n37369 , n37368 );
buf ( n37370 , n37369 );
buf ( n37371 , n37370 );
not ( n37372 , n37371 );
or ( n37373 , n37356 , n37372 );
not ( n37374 , n37305 );
xor ( n37375 , n37191 , n37193 );
xor ( n37376 , n37375 , n37224 );
buf ( n37377 , n37376 );
buf ( n37378 , n37377 );
and ( n37379 , n37374 , n37378 );
not ( n37380 , n37378 );
and ( n37381 , n37363 , n37364 );
xor ( n37382 , n37380 , n37381 );
and ( n37383 , n37382 , n37305 );
or ( n37384 , n37379 , n37383 );
buf ( n37385 , n37384 );
not ( n37386 , n37385 );
buf ( n37387 , n37386 );
buf ( n37388 , n37387 );
not ( n37389 , n37388 );
or ( n37390 , n37373 , n37389 );
not ( n37391 , n37305 );
xor ( n37392 , n37187 , n37189 );
xor ( n37393 , n37392 , n37227 );
buf ( n37394 , n37393 );
buf ( n37395 , n37394 );
and ( n37396 , n37391 , n37395 );
not ( n37397 , n37395 );
and ( n37398 , n37380 , n37381 );
xor ( n37399 , n37397 , n37398 );
and ( n37400 , n37399 , n37305 );
or ( n37401 , n37396 , n37400 );
buf ( n37402 , n37401 );
not ( n37403 , n37402 );
buf ( n37404 , n37403 );
buf ( n37405 , n37404 );
not ( n37406 , n37405 );
or ( n37407 , n37390 , n37406 );
not ( n37408 , n37305 );
xor ( n37409 , n37183 , n37185 );
xor ( n37410 , n37409 , n37230 );
buf ( n37411 , n37410 );
buf ( n37412 , n37411 );
and ( n37413 , n37408 , n37412 );
not ( n37414 , n37412 );
and ( n37415 , n37397 , n37398 );
xor ( n37416 , n37414 , n37415 );
and ( n37417 , n37416 , n37305 );
or ( n37418 , n37413 , n37417 );
buf ( n37419 , n37418 );
not ( n37420 , n37419 );
buf ( n37421 , n37420 );
buf ( n37422 , n37421 );
not ( n37423 , n37422 );
or ( n37424 , n37407 , n37423 );
not ( n37425 , n37305 );
xor ( n37426 , n37179 , n37181 );
xor ( n37427 , n37426 , n37233 );
buf ( n37428 , n37427 );
buf ( n37429 , n37428 );
and ( n37430 , n37425 , n37429 );
not ( n37431 , n37429 );
and ( n37432 , n37414 , n37415 );
xor ( n37433 , n37431 , n37432 );
and ( n37434 , n37433 , n37305 );
or ( n37435 , n37430 , n37434 );
buf ( n37436 , n37435 );
not ( n37437 , n37436 );
buf ( n37438 , n37437 );
buf ( n37439 , n37438 );
not ( n37440 , n37439 );
or ( n37441 , n37424 , n37440 );
not ( n37442 , n37305 );
xor ( n37443 , n37175 , n37177 );
xor ( n37444 , n37443 , n37236 );
buf ( n37445 , n37444 );
buf ( n37446 , n37445 );
and ( n37447 , n37442 , n37446 );
not ( n37448 , n37446 );
and ( n37449 , n37431 , n37432 );
xor ( n37450 , n37448 , n37449 );
and ( n37451 , n37450 , n37305 );
or ( n37452 , n37447 , n37451 );
buf ( n37453 , n37452 );
not ( n37454 , n37453 );
buf ( n37455 , n37454 );
buf ( n37456 , n37455 );
not ( n37457 , n37456 );
or ( n37458 , n37441 , n37457 );
not ( n37459 , n37305 );
xor ( n37460 , n37171 , n37173 );
xor ( n37461 , n37460 , n37239 );
buf ( n37462 , n37461 );
buf ( n37463 , n37462 );
and ( n37464 , n37459 , n37463 );
not ( n37465 , n37463 );
and ( n37466 , n37448 , n37449 );
xor ( n37467 , n37465 , n37466 );
and ( n37468 , n37467 , n37305 );
or ( n37469 , n37464 , n37468 );
buf ( n37470 , n37469 );
not ( n37471 , n37470 );
buf ( n37472 , n37471 );
buf ( n37473 , n37472 );
not ( n37474 , n37473 );
or ( n37475 , n37458 , n37474 );
not ( n37476 , n37305 );
xor ( n37477 , n37167 , n37169 );
xor ( n37478 , n37477 , n37242 );
buf ( n37479 , n37478 );
buf ( n37480 , n37479 );
and ( n37481 , n37476 , n37480 );
not ( n37482 , n37480 );
and ( n37483 , n37465 , n37466 );
xor ( n37484 , n37482 , n37483 );
and ( n37485 , n37484 , n37305 );
or ( n37486 , n37481 , n37485 );
buf ( n37487 , n37486 );
not ( n37488 , n37487 );
buf ( n37489 , n37488 );
buf ( n37490 , n37489 );
not ( n37491 , n37490 );
or ( n37492 , n37475 , n37491 );
not ( n37493 , n37305 );
xor ( n37494 , n37163 , n37165 );
xor ( n37495 , n37494 , n37245 );
buf ( n37496 , n37495 );
buf ( n37497 , n37496 );
and ( n37498 , n37493 , n37497 );
not ( n37499 , n37497 );
and ( n37500 , n37482 , n37483 );
xor ( n37501 , n37499 , n37500 );
and ( n37502 , n37501 , n37305 );
or ( n37503 , n37498 , n37502 );
buf ( n37504 , n37503 );
not ( n37505 , n37504 );
buf ( n37506 , n37505 );
buf ( n37507 , n37506 );
not ( n37508 , n37507 );
or ( n37509 , n37492 , n37508 );
not ( n37510 , n37305 );
xor ( n37511 , n37159 , n37161 );
xor ( n37512 , n37511 , n37248 );
buf ( n37513 , n37512 );
buf ( n37514 , n37513 );
and ( n37515 , n37510 , n37514 );
not ( n37516 , n37514 );
and ( n37517 , n37499 , n37500 );
xor ( n37518 , n37516 , n37517 );
and ( n37519 , n37518 , n37305 );
or ( n37520 , n37515 , n37519 );
buf ( n37521 , n37520 );
not ( n37522 , n37521 );
buf ( n37523 , n37522 );
buf ( n37524 , n37523 );
not ( n37525 , n37524 );
or ( n37526 , n37509 , n37525 );
not ( n37527 , n37305 );
xor ( n37528 , n37155 , n37157 );
xor ( n37529 , n37528 , n37251 );
buf ( n37530 , n37529 );
buf ( n37531 , n37530 );
and ( n37532 , n37527 , n37531 );
not ( n37533 , n37531 );
and ( n37534 , n37516 , n37517 );
xor ( n37535 , n37533 , n37534 );
and ( n37536 , n37535 , n37305 );
or ( n37537 , n37532 , n37536 );
buf ( n37538 , n37537 );
not ( n37539 , n37538 );
buf ( n37540 , n37539 );
buf ( n37541 , n37540 );
not ( n37542 , n37541 );
or ( n37543 , n37526 , n37542 );
not ( n37544 , n37305 );
xor ( n37545 , n37151 , n37153 );
xor ( n37546 , n37545 , n37254 );
buf ( n37547 , n37546 );
buf ( n37548 , n37547 );
and ( n37549 , n37544 , n37548 );
not ( n37550 , n37548 );
and ( n37551 , n37533 , n37534 );
xor ( n37552 , n37550 , n37551 );
and ( n37553 , n37552 , n37305 );
or ( n37554 , n37549 , n37553 );
buf ( n37555 , n37554 );
not ( n37556 , n37555 );
buf ( n37557 , n37556 );
buf ( n37558 , n37557 );
not ( n37559 , n37558 );
or ( n37560 , n37543 , n37559 );
not ( n37561 , n37305 );
xor ( n37562 , n37147 , n37149 );
xor ( n37563 , n37562 , n37257 );
buf ( n37564 , n37563 );
buf ( n37565 , n37564 );
and ( n37566 , n37561 , n37565 );
not ( n37567 , n37565 );
and ( n37568 , n37550 , n37551 );
xor ( n37569 , n37567 , n37568 );
and ( n37570 , n37569 , n37305 );
or ( n37571 , n37566 , n37570 );
buf ( n37572 , n37571 );
not ( n37573 , n37572 );
buf ( n37574 , n37573 );
buf ( n37575 , n37574 );
not ( n37576 , n37575 );
or ( n37577 , n37560 , n37576 );
not ( n37578 , n37305 );
xor ( n37579 , n37143 , n37145 );
xor ( n37580 , n37579 , n37260 );
buf ( n37581 , n37580 );
buf ( n37582 , n37581 );
and ( n37583 , n37578 , n37582 );
not ( n37584 , n37582 );
and ( n37585 , n37567 , n37568 );
xor ( n37586 , n37584 , n37585 );
and ( n37587 , n37586 , n37305 );
or ( n37588 , n37583 , n37587 );
buf ( n37589 , n37588 );
not ( n37590 , n37589 );
buf ( n37591 , n37590 );
buf ( n37592 , n37591 );
not ( n37593 , n37592 );
or ( n37594 , n37577 , n37593 );
not ( n37595 , n37305 );
xor ( n37596 , n37139 , n37141 );
xor ( n37597 , n37596 , n37263 );
buf ( n37598 , n37597 );
buf ( n37599 , n37598 );
and ( n37600 , n37595 , n37599 );
not ( n37601 , n37599 );
and ( n37602 , n37584 , n37585 );
xor ( n37603 , n37601 , n37602 );
and ( n37604 , n37603 , n37305 );
or ( n37605 , n37600 , n37604 );
buf ( n37606 , n37605 );
not ( n37607 , n37606 );
buf ( n37608 , n37607 );
buf ( n37609 , n37608 );
not ( n37610 , n37609 );
or ( n37611 , n37594 , n37610 );
not ( n37612 , n37305 );
xor ( n37613 , n37135 , n37137 );
xor ( n37614 , n37613 , n37266 );
buf ( n37615 , n37614 );
buf ( n37616 , n37615 );
and ( n37617 , n37612 , n37616 );
not ( n37618 , n37616 );
and ( n37619 , n37601 , n37602 );
xor ( n37620 , n37618 , n37619 );
and ( n37621 , n37620 , n37305 );
or ( n37622 , n37617 , n37621 );
buf ( n37623 , n37622 );
not ( n37624 , n37623 );
buf ( n37625 , n37624 );
buf ( n37626 , n37625 );
not ( n37627 , n37626 );
or ( n37628 , n37611 , n37627 );
not ( n37629 , n37305 );
xor ( n37630 , n37131 , n37133 );
xor ( n37631 , n37630 , n37269 );
buf ( n37632 , n37631 );
buf ( n37633 , n37632 );
and ( n37634 , n37629 , n37633 );
not ( n37635 , n37633 );
and ( n37636 , n37618 , n37619 );
xor ( n37637 , n37635 , n37636 );
and ( n37638 , n37637 , n37305 );
or ( n37639 , n37634 , n37638 );
buf ( n37640 , n37639 );
not ( n37641 , n37640 );
buf ( n37642 , n37641 );
buf ( n37643 , n37642 );
not ( n37644 , n37643 );
or ( n37645 , n37628 , n37644 );
not ( n37646 , n37305 );
xor ( n37647 , n37127 , n37129 );
xor ( n37648 , n37647 , n37272 );
buf ( n37649 , n37648 );
buf ( n37650 , n37649 );
and ( n37651 , n37646 , n37650 );
not ( n37652 , n37650 );
and ( n37653 , n37635 , n37636 );
xor ( n37654 , n37652 , n37653 );
and ( n37655 , n37654 , n37305 );
or ( n37656 , n37651 , n37655 );
buf ( n37657 , n37656 );
not ( n37658 , n37657 );
buf ( n37659 , n37658 );
buf ( n37660 , n37659 );
not ( n37661 , n37660 );
or ( n37662 , n37645 , n37661 );
not ( n37663 , n37305 );
xor ( n37664 , n37123 , n37125 );
xor ( n37665 , n37664 , n37275 );
buf ( n37666 , n37665 );
buf ( n37667 , n37666 );
and ( n37668 , n37663 , n37667 );
not ( n37669 , n37667 );
and ( n37670 , n37652 , n37653 );
xor ( n37671 , n37669 , n37670 );
and ( n37672 , n37671 , n37305 );
or ( n37673 , n37668 , n37672 );
buf ( n37674 , n37673 );
not ( n37675 , n37674 );
buf ( n37676 , n37675 );
buf ( n37677 , n37676 );
not ( n37678 , n37677 );
or ( n37679 , n37662 , n37678 );
not ( n37680 , n37305 );
xor ( n37681 , n37119 , n37121 );
xor ( n37682 , n37681 , n37278 );
buf ( n37683 , n37682 );
buf ( n37684 , n37683 );
and ( n37685 , n37680 , n37684 );
not ( n37686 , n37684 );
and ( n37687 , n37669 , n37670 );
xor ( n37688 , n37686 , n37687 );
and ( n37689 , n37688 , n37305 );
or ( n37690 , n37685 , n37689 );
buf ( n37691 , n37690 );
not ( n37692 , n37691 );
buf ( n37693 , n37692 );
buf ( n37694 , n37693 );
not ( n37695 , n37694 );
or ( n37696 , n37679 , n37695 );
not ( n37697 , n37305 );
xor ( n37698 , n37115 , n37117 );
xor ( n37699 , n37698 , n37281 );
buf ( n37700 , n37699 );
buf ( n37701 , n37700 );
and ( n37702 , n37697 , n37701 );
not ( n37703 , n37701 );
and ( n37704 , n37686 , n37687 );
xor ( n37705 , n37703 , n37704 );
and ( n37706 , n37705 , n37305 );
or ( n37707 , n37702 , n37706 );
buf ( n37708 , n37707 );
not ( n37709 , n37708 );
buf ( n37710 , n37709 );
buf ( n37711 , n37710 );
not ( n37712 , n37711 );
or ( n37713 , n37696 , n37712 );
not ( n37714 , n37305 );
xor ( n37715 , n37111 , n37113 );
xor ( n37716 , n37715 , n37284 );
buf ( n37717 , n37716 );
buf ( n37718 , n37717 );
and ( n37719 , n37714 , n37718 );
not ( n37720 , n37718 );
and ( n37721 , n37703 , n37704 );
xor ( n37722 , n37720 , n37721 );
and ( n37723 , n37722 , n37305 );
or ( n37724 , n37719 , n37723 );
buf ( n37725 , n37724 );
not ( n37726 , n37725 );
buf ( n37727 , n37726 );
buf ( n37728 , n37727 );
not ( n37729 , n37728 );
or ( n37730 , n37713 , n37729 );
not ( n37731 , n37305 );
xor ( n37732 , n37107 , n37109 );
xor ( n37733 , n37732 , n37287 );
buf ( n37734 , n37733 );
buf ( n37735 , n37734 );
and ( n37736 , n37731 , n37735 );
not ( n37737 , n37735 );
and ( n37738 , n37720 , n37721 );
xor ( n37739 , n37737 , n37738 );
and ( n37740 , n37739 , n37305 );
or ( n37741 , n37736 , n37740 );
buf ( n37742 , n37741 );
not ( n37743 , n37742 );
buf ( n37744 , n37743 );
buf ( n37745 , n37744 );
not ( n37746 , n37745 );
or ( n37747 , n37730 , n37746 );
not ( n37748 , n37305 );
xor ( n37749 , n37103 , n37105 );
xor ( n37750 , n37749 , n37290 );
buf ( n37751 , n37750 );
buf ( n37752 , n37751 );
and ( n37753 , n37748 , n37752 );
not ( n37754 , n37752 );
and ( n37755 , n37737 , n37738 );
xor ( n37756 , n37754 , n37755 );
and ( n37757 , n37756 , n37305 );
or ( n37758 , n37753 , n37757 );
buf ( n37759 , n37758 );
not ( n37760 , n37759 );
buf ( n37761 , n37760 );
buf ( n37762 , n37761 );
not ( n37763 , n37762 );
or ( n37764 , n37747 , n37763 );
not ( n37765 , n37305 );
xor ( n37766 , n37099 , n37101 );
xor ( n37767 , n37766 , n37293 );
buf ( n37768 , n37767 );
buf ( n37769 , n37768 );
and ( n37770 , n37765 , n37769 );
not ( n37771 , n37769 );
and ( n37772 , n37754 , n37755 );
xor ( n37773 , n37771 , n37772 );
and ( n37774 , n37773 , n37305 );
or ( n37775 , n37770 , n37774 );
buf ( n37776 , n37775 );
not ( n37777 , n37776 );
buf ( n37778 , n37777 );
buf ( n37779 , n37778 );
not ( n37780 , n37779 );
or ( n37781 , n37764 , n37780 );
not ( n37782 , n37305 );
xor ( n37783 , n37095 , n37097 );
xor ( n37784 , n37783 , n37296 );
buf ( n37785 , n37784 );
buf ( n37786 , n37785 );
and ( n37787 , n37782 , n37786 );
not ( n37788 , n37786 );
and ( n37789 , n37771 , n37772 );
xor ( n37790 , n37788 , n37789 );
and ( n37791 , n37790 , n37305 );
or ( n37792 , n37787 , n37791 );
buf ( n37793 , n37792 );
not ( n37794 , n37793 );
buf ( n37795 , n37794 );
buf ( n37796 , n37795 );
not ( n37797 , n37796 );
or ( n37798 , n37781 , n37797 );
or ( n37799 , n37798 , C0 );
buf ( n37800 , n37799 );
and ( n37801 , n37800 , n37305 );
not ( n37802 , n37801 );
and ( n37803 , n37802 , n37423 );
xor ( n37804 , n37423 , n37305 );
xor ( n37805 , n37406 , n37305 );
xor ( n37806 , n37389 , n37305 );
xor ( n37807 , n37372 , n37305 );
xor ( n37808 , n37355 , n37305 );
xor ( n37809 , n37338 , n37305 );
xor ( n37810 , n37321 , n37305 );
xor ( n37811 , n37086 , n37305 );
and ( n37812 , n37811 , n37305 );
and ( n37813 , n37810 , n37812 );
and ( n37814 , n37809 , n37813 );
and ( n37815 , n37808 , n37814 );
and ( n37816 , n37807 , n37815 );
and ( n37817 , n37806 , n37816 );
and ( n37818 , n37805 , n37817 );
xor ( n37819 , n37804 , n37818 );
and ( n37820 , n37819 , n37801 );
or ( n37821 , n37803 , n37820 );
buf ( n37822 , n37821 );
and ( n37823 , n37822 , n36350 );
or ( n37824 , n36349 , n36345 );
or ( n37825 , n37824 , C0 );
and ( n37826 , n13413 , n37825 );
or ( n37827 , n37823 , n37826 );
and ( n37828 , n37827 , n14584 );
and ( n37829 , n37069 , n36350 );
or ( n37830 , n37071 , n36345 );
or ( n37831 , n37830 , C0 );
and ( n37832 , n13413 , n37831 );
or ( n37833 , n37829 , n37832 );
or ( n37834 , n14576 , n14578 );
or ( n37835 , n37834 , n14582 );
and ( n37836 , n37833 , n37835 );
and ( n37837 , n37822 , n36350 );
and ( n37838 , n13413 , n37831 );
or ( n37839 , n37837 , n37838 );
or ( n37840 , n14572 , n14574 );
or ( n37841 , n37840 , n14580 );
and ( n37842 , n37839 , n37841 );
and ( n37843 , n15713 , n36350 );
and ( n37844 , n13413 , n37831 );
or ( n37845 , n37843 , n37844 );
or ( n37846 , n14565 , n14567 );
or ( n37847 , n37846 , n14569 );
and ( n37848 , n37845 , n37847 );
or ( n37849 , n14564 , n14592 );
and ( n37850 , n13413 , n37849 );
or ( n37851 , n36355 , n37076 , n37828 , n37836 , n37842 , n37848 , n37850 );
and ( n37852 , n34822 , n37851 );
and ( n37853 , n13413 , n34821 );
or ( n37854 , n37852 , n37853 );
and ( n37855 , n37854 , n16574 );
and ( n37856 , n13413 , n16576 );
or ( n37857 , n37855 , n37856 );
buf ( n37858 , n37857 );
buf ( n37859 , n37858 );
buf ( n37860 , n10615 );
and ( n37861 , n16984 , n23924 );
and ( n37862 , n21865 , n23926 );
or ( n37863 , n37861 , n37862 );
buf ( n37864 , n37863 );
buf ( n37865 , n37864 );
buf ( n37866 , n10615 );
and ( n37867 , n24325 , n31008 );
and ( n37868 , n29105 , n10618 );
or ( n37869 , n37867 , n37868 );
buf ( n37870 , n37869 );
buf ( n37871 , n37870 );
buf ( n37872 , n10615 );
buf ( n37873 , n10615 );
not ( n37874 , n24800 );
not ( n37875 , n26823 );
and ( n37876 , n37875 , n26071 );
xor ( n37877 , n31021 , n31032 );
and ( n37878 , n37877 , n26823 );
or ( n37879 , n37876 , n37878 );
buf ( n37880 , n37879 );
and ( n37881 , n37880 , n27046 );
and ( n37882 , n37880 , n27049 );
not ( n37883 , n27051 );
and ( n37884 , n37883 , n28016 );
not ( n37885 , n28494 );
and ( n37886 , n37885 , n28028 );
xor ( n37887 , n31049 , n31060 );
and ( n37888 , n37887 , n28494 );
or ( n37889 , n37886 , n37888 );
buf ( n37890 , n37889 );
and ( n37891 , n37890 , n27051 );
or ( n37892 , n37884 , n37891 );
and ( n37893 , n37892 , n28506 );
and ( n37894 , n28016 , n28508 );
or ( n37895 , n37881 , n37882 , n37893 , n37894 );
and ( n37896 , n37895 , n28586 );
and ( n37897 , n26089 , n34573 );
or ( n37898 , n37896 , n37897 );
and ( n37899 , n37898 , n28594 );
not ( n37900 , n30249 );
and ( n37901 , n37900 , n29871 );
xor ( n37902 , n31084 , n31095 );
and ( n37903 , n37902 , n30249 );
or ( n37904 , n37901 , n37903 );
buf ( n37905 , n37904 );
and ( n37906 , n37905 , n28586 );
and ( n37907 , n26089 , n34573 );
or ( n37908 , n37906 , n37907 );
and ( n37909 , n37908 , n30269 );
not ( n37910 , n30963 );
and ( n37911 , n37910 , n30585 );
xor ( n37912 , n31112 , n31123 );
and ( n37913 , n37912 , n30963 );
or ( n37914 , n37911 , n37913 );
buf ( n37915 , n37914 );
and ( n37916 , n37915 , n28586 );
and ( n37917 , n26089 , n34573 );
or ( n37918 , n37916 , n37917 );
and ( n37919 , n37918 , n30982 );
and ( n37920 , n29535 , n28586 );
and ( n37921 , n26089 , n34573 );
or ( n37922 , n37920 , n37921 );
and ( n37923 , n37922 , n30989 );
xor ( n37924 , n31147 , n31163 );
buf ( n37925 , n37924 );
and ( n37926 , n37925 , n28586 );
and ( n37927 , n26089 , n34573 );
or ( n37928 , n37926 , n37927 );
and ( n37929 , n37928 , n31002 );
and ( n37930 , n26089 , n34607 );
or ( n37931 , n37899 , n37909 , n37919 , n37923 , n37929 , n37930 );
and ( n37932 , n37874 , n37931 );
and ( n37933 , n26089 , n24800 );
or ( n37934 , n37932 , n37933 );
and ( n37935 , n37934 , n31008 );
and ( n37936 , n26089 , n10618 );
or ( n37937 , n37935 , n37936 );
buf ( n37938 , n37937 );
buf ( n37939 , n37938 );
buf ( n37940 , n10613 );
buf ( n37941 , n10615 );
buf ( n37942 , n10615 );
buf ( n37943 , n10613 );
buf ( n37944 , n10613 );
not ( n37945 , n17162 );
not ( n37946 , n17450 );
or ( n37947 , n21341 , n17873 );
and ( n37948 , n10673 , n37947 );
buf ( n37949 , n21637 );
buf ( n37950 , n18504 );
xor ( n37951 , n37949 , n37950 );
buf ( n37952 , n37951 );
buf ( n37953 , n37952 );
buf ( n37954 , n37953 );
not ( n37955 , n37954 );
buf ( n37956 , n37955 );
buf ( n37957 , n37956 );
not ( n37958 , n37957 );
buf ( n37959 , n18521 );
buf ( n37960 , n20478 );
buf ( n37961 , n20490 );
buf ( n37962 , n19452 );
buf ( n37963 , n19418 );
buf ( n37964 , n19384 );
buf ( n37965 , n17453 );
buf ( n37966 , n19317 );
buf ( n37967 , n19283 );
buf ( n37968 , n19249 );
buf ( n37969 , n19215 );
buf ( n37970 , n19181 );
buf ( n37971 , n22040 );
buf ( n37972 , n19147 );
and ( n37973 , n37971 , n37972 );
buf ( n37974 , n22060 );
buf ( n37975 , n19113 );
and ( n37976 , n37974 , n37975 );
buf ( n37977 , n22080 );
buf ( n37978 , n19079 );
and ( n37979 , n37977 , n37978 );
buf ( n37980 , n22100 );
buf ( n37981 , n19045 );
and ( n37982 , n37980 , n37981 );
buf ( n37983 , n22120 );
buf ( n37984 , n19011 );
and ( n37985 , n37983 , n37984 );
buf ( n37986 , n22140 );
buf ( n37987 , n18977 );
and ( n37988 , n37986 , n37987 );
buf ( n37989 , n22160 );
buf ( n37990 , n18943 );
and ( n37991 , n37989 , n37990 );
buf ( n37992 , n22180 );
buf ( n37993 , n18909 );
and ( n37994 , n37992 , n37993 );
buf ( n37995 , n22200 );
buf ( n37996 , n18875 );
and ( n37997 , n37995 , n37996 );
buf ( n37998 , n22220 );
buf ( n37999 , n18841 );
and ( n38000 , n37998 , n37999 );
buf ( n38001 , n22240 );
buf ( n38002 , n18807 );
and ( n38003 , n38001 , n38002 );
buf ( n38004 , n22260 );
buf ( n38005 , n18773 );
and ( n38006 , n38004 , n38005 );
buf ( n38007 , n22280 );
buf ( n38008 , n18739 );
and ( n38009 , n38007 , n38008 );
buf ( n38010 , n22300 );
buf ( n38011 , n18705 );
and ( n38012 , n38010 , n38011 );
buf ( n38013 , n22320 );
buf ( n38014 , n18671 );
and ( n38015 , n38013 , n38014 );
buf ( n38016 , n22340 );
buf ( n38017 , n18637 );
and ( n38018 , n38016 , n38017 );
buf ( n38019 , n22360 );
buf ( n38020 , n18604 );
and ( n38021 , n38019 , n38020 );
buf ( n38022 , n22380 );
buf ( n38023 , n18571 );
and ( n38024 , n38022 , n38023 );
buf ( n38025 , n22400 );
buf ( n38026 , n18540 );
and ( n38027 , n38025 , n38026 );
and ( n38028 , n37949 , n37950 );
and ( n38029 , n38026 , n38028 );
and ( n38030 , n38025 , n38028 );
or ( n38031 , n38027 , n38029 , n38030 );
and ( n38032 , n38023 , n38031 );
and ( n38033 , n38022 , n38031 );
or ( n38034 , n38024 , n38032 , n38033 );
and ( n38035 , n38020 , n38034 );
and ( n38036 , n38019 , n38034 );
or ( n38037 , n38021 , n38035 , n38036 );
and ( n38038 , n38017 , n38037 );
and ( n38039 , n38016 , n38037 );
or ( n38040 , n38018 , n38038 , n38039 );
and ( n38041 , n38014 , n38040 );
and ( n38042 , n38013 , n38040 );
or ( n38043 , n38015 , n38041 , n38042 );
and ( n38044 , n38011 , n38043 );
and ( n38045 , n38010 , n38043 );
or ( n38046 , n38012 , n38044 , n38045 );
and ( n38047 , n38008 , n38046 );
and ( n38048 , n38007 , n38046 );
or ( n38049 , n38009 , n38047 , n38048 );
and ( n38050 , n38005 , n38049 );
and ( n38051 , n38004 , n38049 );
or ( n38052 , n38006 , n38050 , n38051 );
and ( n38053 , n38002 , n38052 );
and ( n38054 , n38001 , n38052 );
or ( n38055 , n38003 , n38053 , n38054 );
and ( n38056 , n37999 , n38055 );
and ( n38057 , n37998 , n38055 );
or ( n38058 , n38000 , n38056 , n38057 );
and ( n38059 , n37996 , n38058 );
and ( n38060 , n37995 , n38058 );
or ( n38061 , n37997 , n38059 , n38060 );
and ( n38062 , n37993 , n38061 );
and ( n38063 , n37992 , n38061 );
or ( n38064 , n37994 , n38062 , n38063 );
and ( n38065 , n37990 , n38064 );
and ( n38066 , n37989 , n38064 );
or ( n38067 , n37991 , n38065 , n38066 );
and ( n38068 , n37987 , n38067 );
and ( n38069 , n37986 , n38067 );
or ( n38070 , n37988 , n38068 , n38069 );
and ( n38071 , n37984 , n38070 );
and ( n38072 , n37983 , n38070 );
or ( n38073 , n37985 , n38071 , n38072 );
and ( n38074 , n37981 , n38073 );
and ( n38075 , n37980 , n38073 );
or ( n38076 , n37982 , n38074 , n38075 );
and ( n38077 , n37978 , n38076 );
and ( n38078 , n37977 , n38076 );
or ( n38079 , n37979 , n38077 , n38078 );
and ( n38080 , n37975 , n38079 );
and ( n38081 , n37974 , n38079 );
or ( n38082 , n37976 , n38080 , n38081 );
and ( n38083 , n37972 , n38082 );
and ( n38084 , n37971 , n38082 );
or ( n38085 , n37973 , n38083 , n38084 );
and ( n38086 , n37970 , n38085 );
and ( n38087 , n37969 , n38086 );
and ( n38088 , n37968 , n38087 );
and ( n38089 , n37967 , n38088 );
and ( n38090 , n37966 , n38089 );
and ( n38091 , n37965 , n38090 );
and ( n38092 , n37964 , n38091 );
and ( n38093 , n37963 , n38092 );
and ( n38094 , n37962 , n38093 );
and ( n38095 , n37961 , n38094 );
and ( n38096 , n37960 , n38095 );
xor ( n38097 , n37959 , n38096 );
buf ( n38098 , n38097 );
buf ( n38099 , n38098 );
not ( n38100 , n38099 );
xor ( n38101 , n38025 , n38026 );
xor ( n38102 , n38101 , n38028 );
buf ( n38103 , n38102 );
buf ( n38104 , n38103 );
and ( n38105 , n38100 , n38104 );
not ( n38106 , n38104 );
not ( n38107 , n37953 );
xor ( n38108 , n38106 , n38107 );
and ( n38109 , n38108 , n38099 );
or ( n38110 , n38105 , n38109 );
buf ( n38111 , n38110 );
not ( n38112 , n38111 );
buf ( n38113 , n38112 );
buf ( n38114 , n38113 );
not ( n38115 , n38114 );
or ( n38116 , n37958 , n38115 );
not ( n38117 , n38099 );
xor ( n38118 , n38022 , n38023 );
xor ( n38119 , n38118 , n38031 );
buf ( n38120 , n38119 );
buf ( n38121 , n38120 );
and ( n38122 , n38117 , n38121 );
not ( n38123 , n38121 );
and ( n38124 , n38106 , n38107 );
xor ( n38125 , n38123 , n38124 );
and ( n38126 , n38125 , n38099 );
or ( n38127 , n38122 , n38126 );
buf ( n38128 , n38127 );
not ( n38129 , n38128 );
buf ( n38130 , n38129 );
buf ( n38131 , n38130 );
not ( n38132 , n38131 );
or ( n38133 , n38116 , n38132 );
not ( n38134 , n38099 );
xor ( n38135 , n38019 , n38020 );
xor ( n38136 , n38135 , n38034 );
buf ( n38137 , n38136 );
buf ( n38138 , n38137 );
and ( n38139 , n38134 , n38138 );
not ( n38140 , n38138 );
and ( n38141 , n38123 , n38124 );
xor ( n38142 , n38140 , n38141 );
and ( n38143 , n38142 , n38099 );
or ( n38144 , n38139 , n38143 );
buf ( n38145 , n38144 );
not ( n38146 , n38145 );
buf ( n38147 , n38146 );
buf ( n38148 , n38147 );
not ( n38149 , n38148 );
or ( n38150 , n38133 , n38149 );
not ( n38151 , n38099 );
xor ( n38152 , n38016 , n38017 );
xor ( n38153 , n38152 , n38037 );
buf ( n38154 , n38153 );
buf ( n38155 , n38154 );
and ( n38156 , n38151 , n38155 );
not ( n38157 , n38155 );
and ( n38158 , n38140 , n38141 );
xor ( n38159 , n38157 , n38158 );
and ( n38160 , n38159 , n38099 );
or ( n38161 , n38156 , n38160 );
buf ( n38162 , n38161 );
not ( n38163 , n38162 );
buf ( n38164 , n38163 );
buf ( n38165 , n38164 );
not ( n38166 , n38165 );
or ( n38167 , n38150 , n38166 );
not ( n38168 , n38099 );
xor ( n38169 , n38013 , n38014 );
xor ( n38170 , n38169 , n38040 );
buf ( n38171 , n38170 );
buf ( n38172 , n38171 );
and ( n38173 , n38168 , n38172 );
not ( n38174 , n38172 );
and ( n38175 , n38157 , n38158 );
xor ( n38176 , n38174 , n38175 );
and ( n38177 , n38176 , n38099 );
or ( n38178 , n38173 , n38177 );
buf ( n38179 , n38178 );
not ( n38180 , n38179 );
buf ( n38181 , n38180 );
buf ( n38182 , n38181 );
not ( n38183 , n38182 );
or ( n38184 , n38167 , n38183 );
not ( n38185 , n38099 );
xor ( n38186 , n38010 , n38011 );
xor ( n38187 , n38186 , n38043 );
buf ( n38188 , n38187 );
buf ( n38189 , n38188 );
and ( n38190 , n38185 , n38189 );
not ( n38191 , n38189 );
and ( n38192 , n38174 , n38175 );
xor ( n38193 , n38191 , n38192 );
and ( n38194 , n38193 , n38099 );
or ( n38195 , n38190 , n38194 );
buf ( n38196 , n38195 );
not ( n38197 , n38196 );
buf ( n38198 , n38197 );
buf ( n38199 , n38198 );
not ( n38200 , n38199 );
or ( n38201 , n38184 , n38200 );
not ( n38202 , n38099 );
xor ( n38203 , n38007 , n38008 );
xor ( n38204 , n38203 , n38046 );
buf ( n38205 , n38204 );
buf ( n38206 , n38205 );
and ( n38207 , n38202 , n38206 );
not ( n38208 , n38206 );
and ( n38209 , n38191 , n38192 );
xor ( n38210 , n38208 , n38209 );
and ( n38211 , n38210 , n38099 );
or ( n38212 , n38207 , n38211 );
buf ( n38213 , n38212 );
not ( n38214 , n38213 );
buf ( n38215 , n38214 );
buf ( n38216 , n38215 );
not ( n38217 , n38216 );
or ( n38218 , n38201 , n38217 );
not ( n38219 , n38099 );
xor ( n38220 , n38004 , n38005 );
xor ( n38221 , n38220 , n38049 );
buf ( n38222 , n38221 );
buf ( n38223 , n38222 );
and ( n38224 , n38219 , n38223 );
not ( n38225 , n38223 );
and ( n38226 , n38208 , n38209 );
xor ( n38227 , n38225 , n38226 );
and ( n38228 , n38227 , n38099 );
or ( n38229 , n38224 , n38228 );
buf ( n38230 , n38229 );
not ( n38231 , n38230 );
buf ( n38232 , n38231 );
buf ( n38233 , n38232 );
not ( n38234 , n38233 );
or ( n38235 , n38218 , n38234 );
not ( n38236 , n38099 );
xor ( n38237 , n38001 , n38002 );
xor ( n38238 , n38237 , n38052 );
buf ( n38239 , n38238 );
buf ( n38240 , n38239 );
and ( n38241 , n38236 , n38240 );
not ( n38242 , n38240 );
and ( n38243 , n38225 , n38226 );
xor ( n38244 , n38242 , n38243 );
and ( n38245 , n38244 , n38099 );
or ( n38246 , n38241 , n38245 );
buf ( n38247 , n38246 );
not ( n38248 , n38247 );
buf ( n38249 , n38248 );
buf ( n38250 , n38249 );
not ( n38251 , n38250 );
or ( n38252 , n38235 , n38251 );
not ( n38253 , n38099 );
xor ( n38254 , n37998 , n37999 );
xor ( n38255 , n38254 , n38055 );
buf ( n38256 , n38255 );
buf ( n38257 , n38256 );
and ( n38258 , n38253 , n38257 );
not ( n38259 , n38257 );
and ( n38260 , n38242 , n38243 );
xor ( n38261 , n38259 , n38260 );
and ( n38262 , n38261 , n38099 );
or ( n38263 , n38258 , n38262 );
buf ( n38264 , n38263 );
not ( n38265 , n38264 );
buf ( n38266 , n38265 );
buf ( n38267 , n38266 );
not ( n38268 , n38267 );
or ( n38269 , n38252 , n38268 );
not ( n38270 , n38099 );
xor ( n38271 , n37995 , n37996 );
xor ( n38272 , n38271 , n38058 );
buf ( n38273 , n38272 );
buf ( n38274 , n38273 );
and ( n38275 , n38270 , n38274 );
not ( n38276 , n38274 );
and ( n38277 , n38259 , n38260 );
xor ( n38278 , n38276 , n38277 );
and ( n38279 , n38278 , n38099 );
or ( n38280 , n38275 , n38279 );
buf ( n38281 , n38280 );
not ( n38282 , n38281 );
buf ( n38283 , n38282 );
buf ( n38284 , n38283 );
not ( n38285 , n38284 );
or ( n38286 , n38269 , n38285 );
not ( n38287 , n38099 );
xor ( n38288 , n37992 , n37993 );
xor ( n38289 , n38288 , n38061 );
buf ( n38290 , n38289 );
buf ( n38291 , n38290 );
and ( n38292 , n38287 , n38291 );
not ( n38293 , n38291 );
and ( n38294 , n38276 , n38277 );
xor ( n38295 , n38293 , n38294 );
and ( n38296 , n38295 , n38099 );
or ( n38297 , n38292 , n38296 );
buf ( n38298 , n38297 );
not ( n38299 , n38298 );
buf ( n38300 , n38299 );
buf ( n38301 , n38300 );
not ( n38302 , n38301 );
or ( n38303 , n38286 , n38302 );
not ( n38304 , n38099 );
xor ( n38305 , n37989 , n37990 );
xor ( n38306 , n38305 , n38064 );
buf ( n38307 , n38306 );
buf ( n38308 , n38307 );
and ( n38309 , n38304 , n38308 );
not ( n38310 , n38308 );
and ( n38311 , n38293 , n38294 );
xor ( n38312 , n38310 , n38311 );
and ( n38313 , n38312 , n38099 );
or ( n38314 , n38309 , n38313 );
buf ( n38315 , n38314 );
not ( n38316 , n38315 );
buf ( n38317 , n38316 );
buf ( n38318 , n38317 );
not ( n38319 , n38318 );
or ( n38320 , n38303 , n38319 );
not ( n38321 , n38099 );
xor ( n38322 , n37986 , n37987 );
xor ( n38323 , n38322 , n38067 );
buf ( n38324 , n38323 );
buf ( n38325 , n38324 );
and ( n38326 , n38321 , n38325 );
not ( n38327 , n38325 );
and ( n38328 , n38310 , n38311 );
xor ( n38329 , n38327 , n38328 );
and ( n38330 , n38329 , n38099 );
or ( n38331 , n38326 , n38330 );
buf ( n38332 , n38331 );
not ( n38333 , n38332 );
buf ( n38334 , n38333 );
buf ( n38335 , n38334 );
not ( n38336 , n38335 );
or ( n38337 , n38320 , n38336 );
not ( n38338 , n38099 );
xor ( n38339 , n37983 , n37984 );
xor ( n38340 , n38339 , n38070 );
buf ( n38341 , n38340 );
buf ( n38342 , n38341 );
and ( n38343 , n38338 , n38342 );
not ( n38344 , n38342 );
and ( n38345 , n38327 , n38328 );
xor ( n38346 , n38344 , n38345 );
and ( n38347 , n38346 , n38099 );
or ( n38348 , n38343 , n38347 );
buf ( n38349 , n38348 );
not ( n38350 , n38349 );
buf ( n38351 , n38350 );
buf ( n38352 , n38351 );
not ( n38353 , n38352 );
or ( n38354 , n38337 , n38353 );
not ( n38355 , n38099 );
xor ( n38356 , n37980 , n37981 );
xor ( n38357 , n38356 , n38073 );
buf ( n38358 , n38357 );
buf ( n38359 , n38358 );
and ( n38360 , n38355 , n38359 );
not ( n38361 , n38359 );
and ( n38362 , n38344 , n38345 );
xor ( n38363 , n38361 , n38362 );
and ( n38364 , n38363 , n38099 );
or ( n38365 , n38360 , n38364 );
buf ( n38366 , n38365 );
not ( n38367 , n38366 );
buf ( n38368 , n38367 );
buf ( n38369 , n38368 );
not ( n38370 , n38369 );
or ( n38371 , n38354 , n38370 );
not ( n38372 , n38099 );
xor ( n38373 , n37977 , n37978 );
xor ( n38374 , n38373 , n38076 );
buf ( n38375 , n38374 );
buf ( n38376 , n38375 );
and ( n38377 , n38372 , n38376 );
not ( n38378 , n38376 );
and ( n38379 , n38361 , n38362 );
xor ( n38380 , n38378 , n38379 );
and ( n38381 , n38380 , n38099 );
or ( n38382 , n38377 , n38381 );
buf ( n38383 , n38382 );
not ( n38384 , n38383 );
buf ( n38385 , n38384 );
buf ( n38386 , n38385 );
not ( n38387 , n38386 );
or ( n38388 , n38371 , n38387 );
not ( n38389 , n38099 );
xor ( n38390 , n37974 , n37975 );
xor ( n38391 , n38390 , n38079 );
buf ( n38392 , n38391 );
buf ( n38393 , n38392 );
and ( n38394 , n38389 , n38393 );
not ( n38395 , n38393 );
and ( n38396 , n38378 , n38379 );
xor ( n38397 , n38395 , n38396 );
and ( n38398 , n38397 , n38099 );
or ( n38399 , n38394 , n38398 );
buf ( n38400 , n38399 );
not ( n38401 , n38400 );
buf ( n38402 , n38401 );
buf ( n38403 , n38402 );
not ( n38404 , n38403 );
or ( n38405 , n38388 , n38404 );
not ( n38406 , n38099 );
xor ( n38407 , n37971 , n37972 );
xor ( n38408 , n38407 , n38082 );
buf ( n38409 , n38408 );
buf ( n38410 , n38409 );
and ( n38411 , n38406 , n38410 );
not ( n38412 , n38410 );
and ( n38413 , n38395 , n38396 );
xor ( n38414 , n38412 , n38413 );
and ( n38415 , n38414 , n38099 );
or ( n38416 , n38411 , n38415 );
buf ( n38417 , n38416 );
not ( n38418 , n38417 );
buf ( n38419 , n38418 );
buf ( n38420 , n38419 );
not ( n38421 , n38420 );
or ( n38422 , n38405 , n38421 );
buf ( n38423 , n38422 );
buf ( n38424 , n38423 );
and ( n38425 , n38424 , n38099 );
not ( n38426 , n38425 );
and ( n38427 , n38426 , n38302 );
xor ( n38428 , n38302 , n38099 );
xor ( n38429 , n38285 , n38099 );
xor ( n38430 , n38268 , n38099 );
xor ( n38431 , n38251 , n38099 );
xor ( n38432 , n38234 , n38099 );
xor ( n38433 , n38217 , n38099 );
xor ( n38434 , n38200 , n38099 );
xor ( n38435 , n38183 , n38099 );
xor ( n38436 , n38166 , n38099 );
xor ( n38437 , n38149 , n38099 );
xor ( n38438 , n38132 , n38099 );
xor ( n38439 , n38115 , n38099 );
xor ( n38440 , n37958 , n38099 );
and ( n38441 , n38440 , n38099 );
and ( n38442 , n38439 , n38441 );
and ( n38443 , n38438 , n38442 );
and ( n38444 , n38437 , n38443 );
and ( n38445 , n38436 , n38444 );
and ( n38446 , n38435 , n38445 );
and ( n38447 , n38434 , n38446 );
and ( n38448 , n38433 , n38447 );
and ( n38449 , n38432 , n38448 );
and ( n38450 , n38431 , n38449 );
and ( n38451 , n38430 , n38450 );
and ( n38452 , n38429 , n38451 );
xor ( n38453 , n38428 , n38452 );
and ( n38454 , n38453 , n38425 );
or ( n38455 , n38427 , n38454 );
buf ( n38456 , n38455 );
and ( n38457 , n38456 , n19745 );
buf ( n38458 , n21637 );
buf ( n38459 , n18508 );
xor ( n38460 , n38458 , n38459 );
buf ( n38461 , n38460 );
buf ( n38462 , n38461 );
buf ( n38463 , n38462 );
not ( n38464 , n38463 );
buf ( n38465 , n38464 );
buf ( n38466 , n38465 );
not ( n38467 , n38466 );
buf ( n38468 , n18523 );
buf ( n38469 , n20480 );
buf ( n38470 , n20492 );
buf ( n38471 , n19454 );
buf ( n38472 , n19420 );
buf ( n38473 , n19386 );
buf ( n38474 , n19352 );
buf ( n38475 , n19319 );
buf ( n38476 , n19285 );
buf ( n38477 , n19251 );
buf ( n38478 , n19217 );
buf ( n38479 , n19183 );
buf ( n38480 , n22040 );
buf ( n38481 , n19149 );
and ( n38482 , n38480 , n38481 );
buf ( n38483 , n22060 );
buf ( n38484 , n19115 );
and ( n38485 , n38483 , n38484 );
buf ( n38486 , n22080 );
buf ( n38487 , n19081 );
and ( n38488 , n38486 , n38487 );
buf ( n38489 , n22100 );
buf ( n38490 , n19047 );
and ( n38491 , n38489 , n38490 );
buf ( n38492 , n22120 );
buf ( n38493 , n19013 );
and ( n38494 , n38492 , n38493 );
buf ( n38495 , n22140 );
buf ( n38496 , n18979 );
and ( n38497 , n38495 , n38496 );
buf ( n38498 , n22160 );
buf ( n38499 , n18945 );
and ( n38500 , n38498 , n38499 );
buf ( n38501 , n22180 );
buf ( n38502 , n18911 );
and ( n38503 , n38501 , n38502 );
buf ( n38504 , n22200 );
buf ( n38505 , n18877 );
and ( n38506 , n38504 , n38505 );
buf ( n38507 , n22220 );
buf ( n38508 , n18843 );
and ( n38509 , n38507 , n38508 );
buf ( n38510 , n22240 );
buf ( n38511 , n18809 );
and ( n38512 , n38510 , n38511 );
buf ( n38513 , n22260 );
buf ( n38514 , n18775 );
and ( n38515 , n38513 , n38514 );
buf ( n38516 , n22280 );
buf ( n38517 , n18741 );
and ( n38518 , n38516 , n38517 );
buf ( n38519 , n22300 );
buf ( n38520 , n18707 );
and ( n38521 , n38519 , n38520 );
buf ( n38522 , n22320 );
buf ( n38523 , n18673 );
and ( n38524 , n38522 , n38523 );
buf ( n38525 , n22340 );
buf ( n38526 , n18639 );
and ( n38527 , n38525 , n38526 );
buf ( n38528 , n22360 );
buf ( n38529 , n18606 );
and ( n38530 , n38528 , n38529 );
buf ( n38531 , n22380 );
buf ( n38532 , n18573 );
and ( n38533 , n38531 , n38532 );
buf ( n38534 , n22400 );
buf ( n38535 , n18542 );
and ( n38536 , n38534 , n38535 );
and ( n38537 , n38458 , n38459 );
and ( n38538 , n38535 , n38537 );
and ( n38539 , n38534 , n38537 );
or ( n38540 , n38536 , n38538 , n38539 );
and ( n38541 , n38532 , n38540 );
and ( n38542 , n38531 , n38540 );
or ( n38543 , n38533 , n38541 , n38542 );
and ( n38544 , n38529 , n38543 );
and ( n38545 , n38528 , n38543 );
or ( n38546 , n38530 , n38544 , n38545 );
and ( n38547 , n38526 , n38546 );
and ( n38548 , n38525 , n38546 );
or ( n38549 , n38527 , n38547 , n38548 );
and ( n38550 , n38523 , n38549 );
and ( n38551 , n38522 , n38549 );
or ( n38552 , n38524 , n38550 , n38551 );
and ( n38553 , n38520 , n38552 );
and ( n38554 , n38519 , n38552 );
or ( n38555 , n38521 , n38553 , n38554 );
and ( n38556 , n38517 , n38555 );
and ( n38557 , n38516 , n38555 );
or ( n38558 , n38518 , n38556 , n38557 );
and ( n38559 , n38514 , n38558 );
and ( n38560 , n38513 , n38558 );
or ( n38561 , n38515 , n38559 , n38560 );
and ( n38562 , n38511 , n38561 );
and ( n38563 , n38510 , n38561 );
or ( n38564 , n38512 , n38562 , n38563 );
and ( n38565 , n38508 , n38564 );
and ( n38566 , n38507 , n38564 );
or ( n38567 , n38509 , n38565 , n38566 );
and ( n38568 , n38505 , n38567 );
and ( n38569 , n38504 , n38567 );
or ( n38570 , n38506 , n38568 , n38569 );
and ( n38571 , n38502 , n38570 );
and ( n38572 , n38501 , n38570 );
or ( n38573 , n38503 , n38571 , n38572 );
and ( n38574 , n38499 , n38573 );
and ( n38575 , n38498 , n38573 );
or ( n38576 , n38500 , n38574 , n38575 );
and ( n38577 , n38496 , n38576 );
and ( n38578 , n38495 , n38576 );
or ( n38579 , n38497 , n38577 , n38578 );
and ( n38580 , n38493 , n38579 );
and ( n38581 , n38492 , n38579 );
or ( n38582 , n38494 , n38580 , n38581 );
and ( n38583 , n38490 , n38582 );
and ( n38584 , n38489 , n38582 );
or ( n38585 , n38491 , n38583 , n38584 );
and ( n38586 , n38487 , n38585 );
and ( n38587 , n38486 , n38585 );
or ( n38588 , n38488 , n38586 , n38587 );
and ( n38589 , n38484 , n38588 );
and ( n38590 , n38483 , n38588 );
or ( n38591 , n38485 , n38589 , n38590 );
and ( n38592 , n38481 , n38591 );
and ( n38593 , n38480 , n38591 );
or ( n38594 , n38482 , n38592 , n38593 );
and ( n38595 , n38479 , n38594 );
and ( n38596 , n38478 , n38595 );
and ( n38597 , n38477 , n38596 );
and ( n38598 , n38476 , n38597 );
and ( n38599 , n38475 , n38598 );
and ( n38600 , n38474 , n38599 );
and ( n38601 , n38473 , n38600 );
and ( n38602 , n38472 , n38601 );
and ( n38603 , n38471 , n38602 );
and ( n38604 , n38470 , n38603 );
and ( n38605 , n38469 , n38604 );
xor ( n38606 , n38468 , n38605 );
buf ( n38607 , n38606 );
buf ( n38608 , n38607 );
not ( n38609 , n38608 );
xor ( n38610 , n38534 , n38535 );
xor ( n38611 , n38610 , n38537 );
buf ( n38612 , n38611 );
buf ( n38613 , n38612 );
and ( n38614 , n38609 , n38613 );
not ( n38615 , n38613 );
not ( n38616 , n38462 );
xor ( n38617 , n38615 , n38616 );
and ( n38618 , n38617 , n38608 );
or ( n38619 , n38614 , n38618 );
buf ( n38620 , n38619 );
not ( n38621 , n38620 );
buf ( n38622 , n38621 );
buf ( n38623 , n38622 );
not ( n38624 , n38623 );
or ( n38625 , n38467 , n38624 );
not ( n38626 , n38608 );
xor ( n38627 , n38531 , n38532 );
xor ( n38628 , n38627 , n38540 );
buf ( n38629 , n38628 );
buf ( n38630 , n38629 );
and ( n38631 , n38626 , n38630 );
not ( n38632 , n38630 );
and ( n38633 , n38615 , n38616 );
xor ( n38634 , n38632 , n38633 );
and ( n38635 , n38634 , n38608 );
or ( n38636 , n38631 , n38635 );
buf ( n38637 , n38636 );
not ( n38638 , n38637 );
buf ( n38639 , n38638 );
buf ( n38640 , n38639 );
not ( n38641 , n38640 );
or ( n38642 , n38625 , n38641 );
not ( n38643 , n38608 );
xor ( n38644 , n38528 , n38529 );
xor ( n38645 , n38644 , n38543 );
buf ( n38646 , n38645 );
buf ( n38647 , n38646 );
and ( n38648 , n38643 , n38647 );
not ( n38649 , n38647 );
and ( n38650 , n38632 , n38633 );
xor ( n38651 , n38649 , n38650 );
and ( n38652 , n38651 , n38608 );
or ( n38653 , n38648 , n38652 );
buf ( n38654 , n38653 );
not ( n38655 , n38654 );
buf ( n38656 , n38655 );
buf ( n38657 , n38656 );
not ( n38658 , n38657 );
or ( n38659 , n38642 , n38658 );
not ( n38660 , n38608 );
xor ( n38661 , n38525 , n38526 );
xor ( n38662 , n38661 , n38546 );
buf ( n38663 , n38662 );
buf ( n38664 , n38663 );
and ( n38665 , n38660 , n38664 );
not ( n38666 , n38664 );
and ( n38667 , n38649 , n38650 );
xor ( n38668 , n38666 , n38667 );
and ( n38669 , n38668 , n38608 );
or ( n38670 , n38665 , n38669 );
buf ( n38671 , n38670 );
not ( n38672 , n38671 );
buf ( n38673 , n38672 );
buf ( n38674 , n38673 );
not ( n38675 , n38674 );
or ( n38676 , n38659 , n38675 );
not ( n38677 , n38608 );
xor ( n38678 , n38522 , n38523 );
xor ( n38679 , n38678 , n38549 );
buf ( n38680 , n38679 );
buf ( n38681 , n38680 );
and ( n38682 , n38677 , n38681 );
not ( n38683 , n38681 );
and ( n38684 , n38666 , n38667 );
xor ( n38685 , n38683 , n38684 );
and ( n38686 , n38685 , n38608 );
or ( n38687 , n38682 , n38686 );
buf ( n38688 , n38687 );
not ( n38689 , n38688 );
buf ( n38690 , n38689 );
buf ( n38691 , n38690 );
not ( n38692 , n38691 );
or ( n38693 , n38676 , n38692 );
not ( n38694 , n38608 );
xor ( n38695 , n38519 , n38520 );
xor ( n38696 , n38695 , n38552 );
buf ( n38697 , n38696 );
buf ( n38698 , n38697 );
and ( n38699 , n38694 , n38698 );
not ( n38700 , n38698 );
and ( n38701 , n38683 , n38684 );
xor ( n38702 , n38700 , n38701 );
and ( n38703 , n38702 , n38608 );
or ( n38704 , n38699 , n38703 );
buf ( n38705 , n38704 );
not ( n38706 , n38705 );
buf ( n38707 , n38706 );
buf ( n38708 , n38707 );
not ( n38709 , n38708 );
or ( n38710 , n38693 , n38709 );
not ( n38711 , n38608 );
xor ( n38712 , n38516 , n38517 );
xor ( n38713 , n38712 , n38555 );
buf ( n38714 , n38713 );
buf ( n38715 , n38714 );
and ( n38716 , n38711 , n38715 );
not ( n38717 , n38715 );
and ( n38718 , n38700 , n38701 );
xor ( n38719 , n38717 , n38718 );
and ( n38720 , n38719 , n38608 );
or ( n38721 , n38716 , n38720 );
buf ( n38722 , n38721 );
not ( n38723 , n38722 );
buf ( n38724 , n38723 );
buf ( n38725 , n38724 );
not ( n38726 , n38725 );
or ( n38727 , n38710 , n38726 );
not ( n38728 , n38608 );
xor ( n38729 , n38513 , n38514 );
xor ( n38730 , n38729 , n38558 );
buf ( n38731 , n38730 );
buf ( n38732 , n38731 );
and ( n38733 , n38728 , n38732 );
not ( n38734 , n38732 );
and ( n38735 , n38717 , n38718 );
xor ( n38736 , n38734 , n38735 );
and ( n38737 , n38736 , n38608 );
or ( n38738 , n38733 , n38737 );
buf ( n38739 , n38738 );
not ( n38740 , n38739 );
buf ( n38741 , n38740 );
buf ( n38742 , n38741 );
not ( n38743 , n38742 );
or ( n38744 , n38727 , n38743 );
not ( n38745 , n38608 );
xor ( n38746 , n38510 , n38511 );
xor ( n38747 , n38746 , n38561 );
buf ( n38748 , n38747 );
buf ( n38749 , n38748 );
and ( n38750 , n38745 , n38749 );
not ( n38751 , n38749 );
and ( n38752 , n38734 , n38735 );
xor ( n38753 , n38751 , n38752 );
and ( n38754 , n38753 , n38608 );
or ( n38755 , n38750 , n38754 );
buf ( n38756 , n38755 );
not ( n38757 , n38756 );
buf ( n38758 , n38757 );
buf ( n38759 , n38758 );
not ( n38760 , n38759 );
or ( n38761 , n38744 , n38760 );
not ( n38762 , n38608 );
xor ( n38763 , n38507 , n38508 );
xor ( n38764 , n38763 , n38564 );
buf ( n38765 , n38764 );
buf ( n38766 , n38765 );
and ( n38767 , n38762 , n38766 );
not ( n38768 , n38766 );
and ( n38769 , n38751 , n38752 );
xor ( n38770 , n38768 , n38769 );
and ( n38771 , n38770 , n38608 );
or ( n38772 , n38767 , n38771 );
buf ( n38773 , n38772 );
not ( n38774 , n38773 );
buf ( n38775 , n38774 );
buf ( n38776 , n38775 );
not ( n38777 , n38776 );
or ( n38778 , n38761 , n38777 );
not ( n38779 , n38608 );
xor ( n38780 , n38504 , n38505 );
xor ( n38781 , n38780 , n38567 );
buf ( n38782 , n38781 );
buf ( n38783 , n38782 );
and ( n38784 , n38779 , n38783 );
not ( n38785 , n38783 );
and ( n38786 , n38768 , n38769 );
xor ( n38787 , n38785 , n38786 );
and ( n38788 , n38787 , n38608 );
or ( n38789 , n38784 , n38788 );
buf ( n38790 , n38789 );
not ( n38791 , n38790 );
buf ( n38792 , n38791 );
buf ( n38793 , n38792 );
not ( n38794 , n38793 );
or ( n38795 , n38778 , n38794 );
not ( n38796 , n38608 );
xor ( n38797 , n38501 , n38502 );
xor ( n38798 , n38797 , n38570 );
buf ( n38799 , n38798 );
buf ( n38800 , n38799 );
and ( n38801 , n38796 , n38800 );
not ( n38802 , n38800 );
and ( n38803 , n38785 , n38786 );
xor ( n38804 , n38802 , n38803 );
and ( n38805 , n38804 , n38608 );
or ( n38806 , n38801 , n38805 );
buf ( n38807 , n38806 );
not ( n38808 , n38807 );
buf ( n38809 , n38808 );
buf ( n38810 , n38809 );
not ( n38811 , n38810 );
or ( n38812 , n38795 , n38811 );
not ( n38813 , n38608 );
xor ( n38814 , n38498 , n38499 );
xor ( n38815 , n38814 , n38573 );
buf ( n38816 , n38815 );
buf ( n38817 , n38816 );
and ( n38818 , n38813 , n38817 );
not ( n38819 , n38817 );
and ( n38820 , n38802 , n38803 );
xor ( n38821 , n38819 , n38820 );
and ( n38822 , n38821 , n38608 );
or ( n38823 , n38818 , n38822 );
buf ( n38824 , n38823 );
not ( n38825 , n38824 );
buf ( n38826 , n38825 );
buf ( n38827 , n38826 );
not ( n38828 , n38827 );
or ( n38829 , n38812 , n38828 );
not ( n38830 , n38608 );
xor ( n38831 , n38495 , n38496 );
xor ( n38832 , n38831 , n38576 );
buf ( n38833 , n38832 );
buf ( n38834 , n38833 );
and ( n38835 , n38830 , n38834 );
not ( n38836 , n38834 );
and ( n38837 , n38819 , n38820 );
xor ( n38838 , n38836 , n38837 );
and ( n38839 , n38838 , n38608 );
or ( n38840 , n38835 , n38839 );
buf ( n38841 , n38840 );
not ( n38842 , n38841 );
buf ( n38843 , n38842 );
buf ( n38844 , n38843 );
not ( n38845 , n38844 );
or ( n38846 , n38829 , n38845 );
not ( n38847 , n38608 );
xor ( n38848 , n38492 , n38493 );
xor ( n38849 , n38848 , n38579 );
buf ( n38850 , n38849 );
buf ( n38851 , n38850 );
and ( n38852 , n38847 , n38851 );
not ( n38853 , n38851 );
and ( n38854 , n38836 , n38837 );
xor ( n38855 , n38853 , n38854 );
and ( n38856 , n38855 , n38608 );
or ( n38857 , n38852 , n38856 );
buf ( n38858 , n38857 );
not ( n38859 , n38858 );
buf ( n38860 , n38859 );
buf ( n38861 , n38860 );
not ( n38862 , n38861 );
or ( n38863 , n38846 , n38862 );
not ( n38864 , n38608 );
xor ( n38865 , n38489 , n38490 );
xor ( n38866 , n38865 , n38582 );
buf ( n38867 , n38866 );
buf ( n38868 , n38867 );
and ( n38869 , n38864 , n38868 );
not ( n38870 , n38868 );
and ( n38871 , n38853 , n38854 );
xor ( n38872 , n38870 , n38871 );
and ( n38873 , n38872 , n38608 );
or ( n38874 , n38869 , n38873 );
buf ( n38875 , n38874 );
not ( n38876 , n38875 );
buf ( n38877 , n38876 );
buf ( n38878 , n38877 );
not ( n38879 , n38878 );
or ( n38880 , n38863 , n38879 );
not ( n38881 , n38608 );
xor ( n38882 , n38486 , n38487 );
xor ( n38883 , n38882 , n38585 );
buf ( n38884 , n38883 );
buf ( n38885 , n38884 );
and ( n38886 , n38881 , n38885 );
not ( n38887 , n38885 );
and ( n38888 , n38870 , n38871 );
xor ( n38889 , n38887 , n38888 );
and ( n38890 , n38889 , n38608 );
or ( n38891 , n38886 , n38890 );
buf ( n38892 , n38891 );
not ( n38893 , n38892 );
buf ( n38894 , n38893 );
buf ( n38895 , n38894 );
not ( n38896 , n38895 );
or ( n38897 , n38880 , n38896 );
not ( n38898 , n38608 );
xor ( n38899 , n38483 , n38484 );
xor ( n38900 , n38899 , n38588 );
buf ( n38901 , n38900 );
buf ( n38902 , n38901 );
and ( n38903 , n38898 , n38902 );
not ( n38904 , n38902 );
and ( n38905 , n38887 , n38888 );
xor ( n38906 , n38904 , n38905 );
and ( n38907 , n38906 , n38608 );
or ( n38908 , n38903 , n38907 );
buf ( n38909 , n38908 );
not ( n38910 , n38909 );
buf ( n38911 , n38910 );
buf ( n38912 , n38911 );
not ( n38913 , n38912 );
or ( n38914 , n38897 , n38913 );
not ( n38915 , n38608 );
xor ( n38916 , n38480 , n38481 );
xor ( n38917 , n38916 , n38591 );
buf ( n38918 , n38917 );
buf ( n38919 , n38918 );
and ( n38920 , n38915 , n38919 );
not ( n38921 , n38919 );
and ( n38922 , n38904 , n38905 );
xor ( n38923 , n38921 , n38922 );
and ( n38924 , n38923 , n38608 );
or ( n38925 , n38920 , n38924 );
buf ( n38926 , n38925 );
not ( n38927 , n38926 );
buf ( n38928 , n38927 );
buf ( n38929 , n38928 );
not ( n38930 , n38929 );
or ( n38931 , n38914 , n38930 );
buf ( n38932 , n38931 );
buf ( n38933 , n38932 );
and ( n38934 , n38933 , n38608 );
not ( n38935 , n38934 );
and ( n38936 , n38935 , n38811 );
xor ( n38937 , n38811 , n38608 );
xor ( n38938 , n38794 , n38608 );
xor ( n38939 , n38777 , n38608 );
xor ( n38940 , n38760 , n38608 );
xor ( n38941 , n38743 , n38608 );
xor ( n38942 , n38726 , n38608 );
xor ( n38943 , n38709 , n38608 );
xor ( n38944 , n38692 , n38608 );
xor ( n38945 , n38675 , n38608 );
xor ( n38946 , n38658 , n38608 );
xor ( n38947 , n38641 , n38608 );
xor ( n38948 , n38624 , n38608 );
xor ( n38949 , n38467 , n38608 );
and ( n38950 , n38949 , n38608 );
and ( n38951 , n38948 , n38950 );
and ( n38952 , n38947 , n38951 );
and ( n38953 , n38946 , n38952 );
and ( n38954 , n38945 , n38953 );
and ( n38955 , n38944 , n38954 );
and ( n38956 , n38943 , n38955 );
and ( n38957 , n38942 , n38956 );
and ( n38958 , n38941 , n38957 );
and ( n38959 , n38940 , n38958 );
and ( n38960 , n38939 , n38959 );
and ( n38961 , n38938 , n38960 );
xor ( n38962 , n38937 , n38961 );
and ( n38963 , n38962 , n38934 );
or ( n38964 , n38936 , n38963 );
buf ( n38965 , n38964 );
and ( n38966 , n38965 , n19748 );
and ( n38967 , n22180 , n21253 );
and ( n38968 , n10673 , n21255 );
or ( n38969 , n38457 , n38966 , n38967 , n38968 );
or ( n38970 , n23917 , n23834 );
or ( n38971 , n38970 , n23830 );
or ( n38972 , n38971 , n23831 );
or ( n38973 , n38972 , n23819 );
or ( n38974 , n38973 , n23820 );
or ( n38975 , n38974 , n23058 );
or ( n38976 , n38975 , n23059 );
or ( n38977 , n38976 , n23822 );
or ( n38978 , n38977 , n23061 );
or ( n38979 , n38978 , n23824 );
or ( n38980 , n38979 , n23063 );
and ( n38981 , n38969 , n38980 );
or ( n38982 , n37948 , n38981 );
and ( n38983 , n37946 , n38982 );
or ( n38984 , n38983 , C0 );
and ( n38985 , n37945 , n38984 );
and ( n38986 , n38969 , n17162 );
or ( n38987 , n38985 , n38986 );
and ( n38988 , n38987 , n23924 );
buf ( n38989 , n17875 );
buf ( n38990 , n38989 );
not ( n38991 , n38990 );
buf ( n38992 , n38991 );
buf ( n38993 , n38992 );
not ( n38994 , n38993 );
buf ( n38995 , n17882 );
not ( n38996 , n38995 );
buf ( n38997 , n17885 );
and ( n38998 , n38996 , n38997 );
not ( n38999 , n38997 );
not ( n39000 , n38989 );
xor ( n39001 , n38999 , n39000 );
and ( n39002 , n39001 , n38995 );
or ( n39003 , n38998 , n39002 );
buf ( n39004 , n39003 );
not ( n39005 , n39004 );
buf ( n39006 , n39005 );
buf ( n39007 , n39006 );
not ( n39008 , n39007 );
or ( n39009 , n38994 , n39008 );
not ( n39010 , n38995 );
buf ( n39011 , n17900 );
and ( n39012 , n39010 , n39011 );
not ( n39013 , n39011 );
and ( n39014 , n38999 , n39000 );
xor ( n39015 , n39013 , n39014 );
and ( n39016 , n39015 , n38995 );
or ( n39017 , n39012 , n39016 );
buf ( n39018 , n39017 );
not ( n39019 , n39018 );
buf ( n39020 , n39019 );
buf ( n39021 , n39020 );
not ( n39022 , n39021 );
or ( n39023 , n39009 , n39022 );
not ( n39024 , n38995 );
buf ( n39025 , n17915 );
and ( n39026 , n39024 , n39025 );
not ( n39027 , n39025 );
and ( n39028 , n39013 , n39014 );
xor ( n39029 , n39027 , n39028 );
and ( n39030 , n39029 , n38995 );
or ( n39031 , n39026 , n39030 );
buf ( n39032 , n39031 );
not ( n39033 , n39032 );
buf ( n39034 , n39033 );
buf ( n39035 , n39034 );
not ( n39036 , n39035 );
or ( n39037 , n39023 , n39036 );
not ( n39038 , n38995 );
buf ( n39039 , n17930 );
and ( n39040 , n39038 , n39039 );
not ( n39041 , n39039 );
and ( n39042 , n39027 , n39028 );
xor ( n39043 , n39041 , n39042 );
and ( n39044 , n39043 , n38995 );
or ( n39045 , n39040 , n39044 );
buf ( n39046 , n39045 );
not ( n39047 , n39046 );
buf ( n39048 , n39047 );
buf ( n39049 , n39048 );
not ( n39050 , n39049 );
or ( n39051 , n39037 , n39050 );
not ( n39052 , n38995 );
buf ( n39053 , n17945 );
and ( n39054 , n39052 , n39053 );
not ( n39055 , n39053 );
and ( n39056 , n39041 , n39042 );
xor ( n39057 , n39055 , n39056 );
and ( n39058 , n39057 , n38995 );
or ( n39059 , n39054 , n39058 );
buf ( n39060 , n39059 );
not ( n39061 , n39060 );
buf ( n39062 , n39061 );
buf ( n39063 , n39062 );
not ( n39064 , n39063 );
or ( n39065 , n39051 , n39064 );
not ( n39066 , n38995 );
buf ( n39067 , n17960 );
and ( n39068 , n39066 , n39067 );
not ( n39069 , n39067 );
and ( n39070 , n39055 , n39056 );
xor ( n39071 , n39069 , n39070 );
and ( n39072 , n39071 , n38995 );
or ( n39073 , n39068 , n39072 );
buf ( n39074 , n39073 );
not ( n39075 , n39074 );
buf ( n39076 , n39075 );
buf ( n39077 , n39076 );
not ( n39078 , n39077 );
or ( n39079 , n39065 , n39078 );
not ( n39080 , n38995 );
buf ( n39081 , n17975 );
and ( n39082 , n39080 , n39081 );
not ( n39083 , n39081 );
and ( n39084 , n39069 , n39070 );
xor ( n39085 , n39083 , n39084 );
and ( n39086 , n39085 , n38995 );
or ( n39087 , n39082 , n39086 );
buf ( n39088 , n39087 );
not ( n39089 , n39088 );
buf ( n39090 , n39089 );
buf ( n39091 , n39090 );
not ( n39092 , n39091 );
or ( n39093 , n39079 , n39092 );
not ( n39094 , n38995 );
buf ( n39095 , n17990 );
and ( n39096 , n39094 , n39095 );
not ( n39097 , n39095 );
and ( n39098 , n39083 , n39084 );
xor ( n39099 , n39097 , n39098 );
and ( n39100 , n39099 , n38995 );
or ( n39101 , n39096 , n39100 );
buf ( n39102 , n39101 );
not ( n39103 , n39102 );
buf ( n39104 , n39103 );
buf ( n39105 , n39104 );
not ( n39106 , n39105 );
or ( n39107 , n39093 , n39106 );
not ( n39108 , n38995 );
buf ( n39109 , n18005 );
and ( n39110 , n39108 , n39109 );
not ( n39111 , n39109 );
and ( n39112 , n39097 , n39098 );
xor ( n39113 , n39111 , n39112 );
and ( n39114 , n39113 , n38995 );
or ( n39115 , n39110 , n39114 );
buf ( n39116 , n39115 );
not ( n39117 , n39116 );
buf ( n39118 , n39117 );
buf ( n39119 , n39118 );
not ( n39120 , n39119 );
or ( n39121 , n39107 , n39120 );
not ( n39122 , n38995 );
buf ( n39123 , n18020 );
and ( n39124 , n39122 , n39123 );
not ( n39125 , n39123 );
and ( n39126 , n39111 , n39112 );
xor ( n39127 , n39125 , n39126 );
and ( n39128 , n39127 , n38995 );
or ( n39129 , n39124 , n39128 );
buf ( n39130 , n39129 );
not ( n39131 , n39130 );
buf ( n39132 , n39131 );
buf ( n39133 , n39132 );
not ( n39134 , n39133 );
or ( n39135 , n39121 , n39134 );
not ( n39136 , n38995 );
buf ( n39137 , n18035 );
and ( n39138 , n39136 , n39137 );
not ( n39139 , n39137 );
and ( n39140 , n39125 , n39126 );
xor ( n39141 , n39139 , n39140 );
and ( n39142 , n39141 , n38995 );
or ( n39143 , n39138 , n39142 );
buf ( n39144 , n39143 );
not ( n39145 , n39144 );
buf ( n39146 , n39145 );
buf ( n39147 , n39146 );
not ( n39148 , n39147 );
or ( n39149 , n39135 , n39148 );
not ( n39150 , n38995 );
buf ( n39151 , n18050 );
and ( n39152 , n39150 , n39151 );
not ( n39153 , n39151 );
and ( n39154 , n39139 , n39140 );
xor ( n39155 , n39153 , n39154 );
and ( n39156 , n39155 , n38995 );
or ( n39157 , n39152 , n39156 );
buf ( n39158 , n39157 );
not ( n39159 , n39158 );
buf ( n39160 , n39159 );
buf ( n39161 , n39160 );
not ( n39162 , n39161 );
or ( n39163 , n39149 , n39162 );
not ( n39164 , n38995 );
buf ( n39165 , n18065 );
and ( n39166 , n39164 , n39165 );
not ( n39167 , n39165 );
and ( n39168 , n39153 , n39154 );
xor ( n39169 , n39167 , n39168 );
and ( n39170 , n39169 , n38995 );
or ( n39171 , n39166 , n39170 );
buf ( n39172 , n39171 );
not ( n39173 , n39172 );
buf ( n39174 , n39173 );
buf ( n39175 , n39174 );
not ( n39176 , n39175 );
or ( n39177 , n39163 , n39176 );
not ( n39178 , n38995 );
buf ( n39179 , n18080 );
and ( n39180 , n39178 , n39179 );
not ( n39181 , n39179 );
and ( n39182 , n39167 , n39168 );
xor ( n39183 , n39181 , n39182 );
and ( n39184 , n39183 , n38995 );
or ( n39185 , n39180 , n39184 );
buf ( n39186 , n39185 );
not ( n39187 , n39186 );
buf ( n39188 , n39187 );
buf ( n39189 , n39188 );
not ( n39190 , n39189 );
or ( n39191 , n39177 , n39190 );
not ( n39192 , n38995 );
buf ( n39193 , n18095 );
and ( n39194 , n39192 , n39193 );
not ( n39195 , n39193 );
and ( n39196 , n39181 , n39182 );
xor ( n39197 , n39195 , n39196 );
and ( n39198 , n39197 , n38995 );
or ( n39199 , n39194 , n39198 );
buf ( n39200 , n39199 );
not ( n39201 , n39200 );
buf ( n39202 , n39201 );
buf ( n39203 , n39202 );
not ( n39204 , n39203 );
or ( n39205 , n39191 , n39204 );
not ( n39206 , n38995 );
buf ( n39207 , n18110 );
and ( n39208 , n39206 , n39207 );
not ( n39209 , n39207 );
and ( n39210 , n39195 , n39196 );
xor ( n39211 , n39209 , n39210 );
and ( n39212 , n39211 , n38995 );
or ( n39213 , n39208 , n39212 );
buf ( n39214 , n39213 );
not ( n39215 , n39214 );
buf ( n39216 , n39215 );
buf ( n39217 , n39216 );
not ( n39218 , n39217 );
or ( n39219 , n39205 , n39218 );
not ( n39220 , n38995 );
buf ( n39221 , n18125 );
and ( n39222 , n39220 , n39221 );
not ( n39223 , n39221 );
and ( n39224 , n39209 , n39210 );
xor ( n39225 , n39223 , n39224 );
and ( n39226 , n39225 , n38995 );
or ( n39227 , n39222 , n39226 );
buf ( n39228 , n39227 );
not ( n39229 , n39228 );
buf ( n39230 , n39229 );
buf ( n39231 , n39230 );
not ( n39232 , n39231 );
or ( n39233 , n39219 , n39232 );
not ( n39234 , n38995 );
buf ( n39235 , n18140 );
and ( n39236 , n39234 , n39235 );
not ( n39237 , n39235 );
and ( n39238 , n39223 , n39224 );
xor ( n39239 , n39237 , n39238 );
and ( n39240 , n39239 , n38995 );
or ( n39241 , n39236 , n39240 );
buf ( n39242 , n39241 );
not ( n39243 , n39242 );
buf ( n39244 , n39243 );
buf ( n39245 , n39244 );
not ( n39246 , n39245 );
or ( n39247 , n39233 , n39246 );
not ( n39248 , n38995 );
buf ( n39249 , n18155 );
and ( n39250 , n39248 , n39249 );
not ( n39251 , n39249 );
and ( n39252 , n39237 , n39238 );
xor ( n39253 , n39251 , n39252 );
and ( n39254 , n39253 , n38995 );
or ( n39255 , n39250 , n39254 );
buf ( n39256 , n39255 );
not ( n39257 , n39256 );
buf ( n39258 , n39257 );
buf ( n39259 , n39258 );
not ( n39260 , n39259 );
or ( n39261 , n39247 , n39260 );
buf ( n39262 , n39261 );
buf ( n39263 , n39262 );
and ( n39264 , n39263 , n38995 );
not ( n39265 , n39264 );
and ( n39266 , n39265 , n39162 );
xor ( n39267 , n39162 , n38995 );
xor ( n39268 , n39148 , n38995 );
xor ( n39269 , n39134 , n38995 );
xor ( n39270 , n39120 , n38995 );
xor ( n39271 , n39106 , n38995 );
xor ( n39272 , n39092 , n38995 );
xor ( n39273 , n39078 , n38995 );
xor ( n39274 , n39064 , n38995 );
xor ( n39275 , n39050 , n38995 );
xor ( n39276 , n39036 , n38995 );
xor ( n39277 , n39022 , n38995 );
xor ( n39278 , n39008 , n38995 );
xor ( n39279 , n38994 , n38995 );
and ( n39280 , n39279 , n38995 );
and ( n39281 , n39278 , n39280 );
and ( n39282 , n39277 , n39281 );
and ( n39283 , n39276 , n39282 );
and ( n39284 , n39275 , n39283 );
and ( n39285 , n39274 , n39284 );
and ( n39286 , n39273 , n39285 );
and ( n39287 , n39272 , n39286 );
and ( n39288 , n39271 , n39287 );
and ( n39289 , n39270 , n39288 );
and ( n39290 , n39269 , n39289 );
and ( n39291 , n39268 , n39290 );
xor ( n39292 , n39267 , n39291 );
and ( n39293 , n39292 , n39264 );
or ( n39294 , n39266 , n39293 );
buf ( n39295 , n39294 );
and ( n39296 , n39295 , n23926 );
or ( n39297 , n38988 , n39296 );
buf ( n39298 , n39297 );
buf ( n39299 , n39298 );
and ( n39300 , n11553 , n16574 );
and ( n39301 , n15462 , n16576 );
or ( n39302 , n39300 , n39301 );
buf ( n39303 , n39302 );
buf ( n39304 , n39303 );
not ( n39305 , n17451 );
not ( n39306 , n19474 );
and ( n39307 , n39306 , n19063 );
xor ( n39308 , n19485 , n19517 );
and ( n39309 , n39308 , n19474 );
or ( n39310 , n39307 , n39309 );
buf ( n39311 , n39310 );
and ( n39312 , n39311 , n19745 );
and ( n39313 , n39311 , n19748 );
not ( n39314 , n19750 );
and ( n39315 , n39314 , n20943 );
not ( n39316 , n21193 );
and ( n39317 , n39316 , n20955 );
xor ( n39318 , n21204 , n21238 );
and ( n39319 , n39318 , n21193 );
or ( n39320 , n39317 , n39319 );
buf ( n39321 , n39320 );
and ( n39322 , n39321 , n19750 );
or ( n39323 , n39315 , n39322 );
and ( n39324 , n39323 , n21253 );
and ( n39325 , n20943 , n21255 );
or ( n39326 , n39312 , n39313 , n39324 , n39325 );
and ( n39327 , n39326 , n21334 );
and ( n39328 , n19083 , n34492 );
or ( n39329 , n39327 , n39328 );
and ( n39330 , n39329 , n21341 );
not ( n39331 , n22996 );
and ( n39332 , n39331 , n22788 );
xor ( n39333 , n23007 , n23041 );
and ( n39334 , n39333 , n22996 );
or ( n39335 , n39332 , n39334 );
buf ( n39336 , n39335 );
and ( n39337 , n39336 , n21334 );
and ( n39338 , n19083 , n34492 );
or ( n39339 , n39337 , n39338 );
and ( n39340 , n39339 , n23064 );
not ( n39341 , n23758 );
and ( n39342 , n39341 , n23550 );
xor ( n39343 , n23769 , n23803 );
and ( n39344 , n39343 , n23758 );
or ( n39345 , n39342 , n39344 );
buf ( n39346 , n39345 );
and ( n39347 , n39346 , n21334 );
and ( n39348 , n19083 , n34492 );
or ( n39349 , n39347 , n39348 );
and ( n39350 , n39349 , n23825 );
and ( n39351 , n22082 , n21334 );
and ( n39352 , n19083 , n34492 );
or ( n39353 , n39351 , n39352 );
and ( n39354 , n39353 , n23832 );
xor ( n39355 , n23853 , n23903 );
buf ( n39356 , n39355 );
and ( n39357 , n39356 , n21334 );
and ( n39358 , n19083 , n34492 );
or ( n39359 , n39357 , n39358 );
and ( n39360 , n39359 , n23917 );
and ( n39361 , n19083 , n34526 );
or ( n39362 , n39330 , n39340 , n39350 , n39354 , n39360 , n39361 );
and ( n39363 , n39305 , n39362 );
and ( n39364 , n19083 , n17451 );
or ( n39365 , n39363 , n39364 );
and ( n39366 , n39365 , n23924 );
and ( n39367 , n19083 , n23926 );
or ( n39368 , n39366 , n39367 );
buf ( n39369 , n39368 );
buf ( n39370 , n39369 );
buf ( n39371 , n10615 );
and ( n39372 , n11816 , n16574 );
and ( n39373 , n15050 , n16576 );
or ( n39374 , n39372 , n39373 );
buf ( n39375 , n39374 );
buf ( n39376 , n39375 );
not ( n39377 , n34821 );
not ( n39378 , n13916 );
and ( n39379 , n39378 , n13760 );
xor ( n39380 , n13761 , n13864 );
and ( n39381 , n39380 , n13916 );
or ( n39382 , n39379 , n39381 );
buf ( n39383 , n39382 );
and ( n39384 , n39383 , n14137 );
and ( n39385 , n39383 , n14143 );
not ( n39386 , n14139 );
and ( n39387 , n39386 , n35833 );
not ( n39388 , n36245 );
and ( n39389 , n39388 , n35845 );
xor ( n39390 , n35845 , n35634 );
xor ( n39391 , n35823 , n35634 );
xor ( n39392 , n35801 , n35634 );
and ( n39393 , n36248 , n36262 );
and ( n39394 , n39392 , n39393 );
and ( n39395 , n39391 , n39394 );
xor ( n39396 , n39390 , n39395 );
and ( n39397 , n39396 , n36245 );
or ( n39398 , n39389 , n39397 );
buf ( n39399 , n39398 );
and ( n39400 , n39399 , n14139 );
or ( n39401 , n39387 , n39400 );
and ( n39402 , n39401 , n14140 );
and ( n39403 , n35833 , n14141 );
or ( n39404 , n39384 , n39385 , n39402 , n39403 );
and ( n39405 , n39404 , n36347 );
or ( n39406 , n36345 , n36348 );
or ( n39407 , n39406 , n36350 );
or ( n39408 , n39407 , C0 );
and ( n39409 , n13375 , n39408 );
or ( n39410 , n39405 , n39409 );
and ( n39411 , n39410 , n14562 );
not ( n39412 , n37048 );
and ( n39413 , n39412 , n36721 );
xor ( n39414 , n36721 , n36552 );
xor ( n39415 , n36704 , n36552 );
xor ( n39416 , n36687 , n36552 );
and ( n39417 , n37051 , n37065 );
and ( n39418 , n39416 , n39417 );
and ( n39419 , n39415 , n39418 );
xor ( n39420 , n39414 , n39419 );
and ( n39421 , n39420 , n37048 );
or ( n39422 , n39413 , n39421 );
buf ( n39423 , n39422 );
and ( n39424 , n39423 , n36348 );
or ( n39425 , n36345 , n36347 );
or ( n39426 , n39425 , n36350 );
or ( n39427 , n39426 , C0 );
and ( n39428 , n13375 , n39427 );
or ( n39429 , n39424 , n39428 );
and ( n39430 , n39429 , n14586 );
not ( n39431 , n37801 );
and ( n39432 , n39431 , n37474 );
xor ( n39433 , n37474 , n37305 );
xor ( n39434 , n37457 , n37305 );
xor ( n39435 , n37440 , n37305 );
and ( n39436 , n37804 , n37818 );
and ( n39437 , n39435 , n39436 );
and ( n39438 , n39434 , n39437 );
xor ( n39439 , n39433 , n39438 );
and ( n39440 , n39439 , n37801 );
or ( n39441 , n39432 , n39440 );
buf ( n39442 , n39441 );
and ( n39443 , n39442 , n36347 );
or ( n39444 , n36350 , n36348 );
or ( n39445 , n39444 , n36345 );
or ( n39446 , n39445 , C0 );
and ( n39447 , n13375 , n39446 );
or ( n39448 , n39443 , n39447 );
and ( n39449 , n39448 , n14584 );
and ( n39450 , n39423 , n36348 );
or ( n39451 , n36350 , n36347 );
or ( n39452 , n39451 , n36345 );
or ( n39453 , n39452 , C0 );
and ( n39454 , n13375 , n39453 );
or ( n39455 , n39450 , n39454 );
and ( n39456 , n39455 , n37835 );
and ( n39457 , n39442 , n36348 );
and ( n39458 , n13375 , n39453 );
or ( n39459 , n39457 , n39458 );
and ( n39460 , n39459 , n37841 );
and ( n39461 , n15647 , n36348 );
and ( n39462 , n13375 , n39453 );
or ( n39463 , n39461 , n39462 );
and ( n39464 , n39463 , n37847 );
and ( n39465 , n13375 , n37849 );
or ( n39466 , n39411 , n39430 , n39449 , n39456 , n39460 , n39464 , n39465 );
and ( n39467 , n39377 , n39466 );
and ( n39468 , n13375 , n34821 );
or ( n39469 , n39467 , n39468 );
and ( n39470 , n39469 , n16574 );
and ( n39471 , n13375 , n16576 );
or ( n39472 , n39470 , n39471 );
buf ( n39473 , n39472 );
buf ( n39474 , n39473 );
buf ( n39475 , n10615 );
buf ( n39476 , n10615 );
buf ( n39477 , n10615 );
not ( n39478 , n17451 );
not ( n39479 , n19474 );
and ( n39480 , n39479 , n19097 );
xor ( n39481 , n19484 , n19518 );
and ( n39482 , n39481 , n19474 );
or ( n39483 , n39480 , n39482 );
buf ( n39484 , n39483 );
and ( n39485 , n39484 , n19745 );
and ( n39486 , n39484 , n19748 );
not ( n39487 , n19750 );
and ( n39488 , n39487 , n20965 );
not ( n39489 , n21193 );
and ( n39490 , n39489 , n20977 );
xor ( n39491 , n21203 , n21239 );
and ( n39492 , n39491 , n21193 );
or ( n39493 , n39490 , n39492 );
buf ( n39494 , n39493 );
and ( n39495 , n39494 , n19750 );
or ( n39496 , n39488 , n39495 );
and ( n39497 , n39496 , n21253 );
and ( n39498 , n20965 , n21255 );
or ( n39499 , n39485 , n39486 , n39497 , n39498 );
and ( n39500 , n39499 , n21333 );
and ( n39501 , n19115 , n34758 );
or ( n39502 , n39500 , n39501 );
and ( n39503 , n39502 , n21341 );
not ( n39504 , n22996 );
and ( n39505 , n39504 , n22805 );
xor ( n39506 , n23006 , n23042 );
and ( n39507 , n39506 , n22996 );
or ( n39508 , n39505 , n39507 );
buf ( n39509 , n39508 );
and ( n39510 , n39509 , n21333 );
and ( n39511 , n19115 , n34758 );
or ( n39512 , n39510 , n39511 );
and ( n39513 , n39512 , n23064 );
not ( n39514 , n23758 );
and ( n39515 , n39514 , n23567 );
xor ( n39516 , n23768 , n23804 );
and ( n39517 , n39516 , n23758 );
or ( n39518 , n39515 , n39517 );
buf ( n39519 , n39518 );
and ( n39520 , n39519 , n21333 );
and ( n39521 , n19115 , n34758 );
or ( n39522 , n39520 , n39521 );
and ( n39523 , n39522 , n23825 );
and ( n39524 , n22062 , n21333 );
and ( n39525 , n19115 , n34758 );
or ( n39526 , n39524 , n39525 );
and ( n39527 , n39526 , n23832 );
xor ( n39528 , n23851 , n23904 );
buf ( n39529 , n39528 );
and ( n39530 , n39529 , n21333 );
and ( n39531 , n19115 , n34758 );
or ( n39532 , n39530 , n39531 );
and ( n39533 , n39532 , n23917 );
and ( n39534 , n19115 , n34526 );
or ( n39535 , n39503 , n39513 , n39523 , n39527 , n39533 , n39534 );
and ( n39536 , n39478 , n39535 );
and ( n39537 , n19115 , n17451 );
or ( n39538 , n39536 , n39537 );
and ( n39539 , n39538 , n23924 );
and ( n39540 , n19115 , n23926 );
or ( n39541 , n39539 , n39540 );
buf ( n39542 , n39541 );
buf ( n39543 , n39542 );
buf ( n39544 , n10613 );
buf ( n39545 , n10613 );
and ( n39546 , n16785 , n23924 );
and ( n39547 , n22113 , n23926 );
or ( n39548 , n39546 , n39547 );
buf ( n39549 , n39548 );
buf ( n39550 , n39549 );
buf ( n39551 , n10613 );
buf ( n39552 , n10615 );
buf ( n39553 , n10613 );
buf ( n39554 , n10613 );
not ( n39555 , n17451 );
not ( n39556 , n19474 );
and ( n39557 , n39556 , n19301 );
xor ( n39558 , n19478 , n19524 );
and ( n39559 , n39558 , n19474 );
or ( n39560 , n39557 , n39559 );
buf ( n39561 , n39560 );
and ( n39562 , n39561 , n19745 );
and ( n39563 , n39561 , n19748 );
not ( n39564 , n19750 );
and ( n39565 , n39564 , n21097 );
not ( n39566 , n21193 );
and ( n39567 , n39566 , n21109 );
xor ( n39568 , n21197 , n21245 );
and ( n39569 , n39568 , n21193 );
or ( n39570 , n39567 , n39569 );
buf ( n39571 , n39570 );
and ( n39572 , n39571 , n19750 );
or ( n39573 , n39565 , n39572 );
and ( n39574 , n39573 , n21253 );
and ( n39575 , n21097 , n21255 );
or ( n39576 , n39562 , n39563 , n39574 , n39575 );
and ( n39577 , n39576 , n21334 );
and ( n39578 , n19321 , n34492 );
or ( n39579 , n39577 , n39578 );
and ( n39580 , n39579 , n21341 );
not ( n39581 , n22996 );
and ( n39582 , n39581 , n22907 );
xor ( n39583 , n23000 , n23048 );
and ( n39584 , n39583 , n22996 );
or ( n39585 , n39582 , n39584 );
buf ( n39586 , n39585 );
and ( n39587 , n39586 , n21334 );
and ( n39588 , n19321 , n34492 );
or ( n39589 , n39587 , n39588 );
and ( n39590 , n39589 , n23064 );
not ( n39591 , n23758 );
and ( n39592 , n39591 , n23669 );
xor ( n39593 , n23762 , n23810 );
and ( n39594 , n39593 , n23758 );
or ( n39595 , n39592 , n39594 );
buf ( n39596 , n39595 );
and ( n39597 , n39596 , n21334 );
and ( n39598 , n19321 , n34492 );
or ( n39599 , n39597 , n39598 );
and ( n39600 , n39599 , n23825 );
and ( n39601 , n21932 , n21334 );
and ( n39602 , n19321 , n34492 );
or ( n39603 , n39601 , n39602 );
and ( n39604 , n39603 , n23832 );
xor ( n39605 , n23839 , n23910 );
buf ( n39606 , n39605 );
and ( n39607 , n39606 , n21334 );
and ( n39608 , n19321 , n34492 );
or ( n39609 , n39607 , n39608 );
and ( n39610 , n39609 , n23917 );
and ( n39611 , n19321 , n34526 );
or ( n39612 , n39580 , n39590 , n39600 , n39604 , n39610 , n39611 );
and ( n39613 , n39555 , n39612 );
and ( n39614 , n19321 , n17451 );
or ( n39615 , n39613 , n39614 );
and ( n39616 , n39615 , n23924 );
and ( n39617 , n19321 , n23926 );
or ( n39618 , n39616 , n39617 );
buf ( n39619 , n39618 );
buf ( n39620 , n39619 );
and ( n39621 , n24249 , n31008 );
and ( n39622 , n28604 , n10618 );
or ( n39623 , n39621 , n39622 );
buf ( n39624 , n39623 );
buf ( n39625 , n39624 );
buf ( n39626 , n10613 );
buf ( n39627 , n10613 );
buf ( n39628 , n10615 );
not ( n39629 , n24800 );
not ( n39630 , n26823 );
and ( n39631 , n39630 , n26411 );
xor ( n39632 , n26411 , n25877 );
xor ( n39633 , n26377 , n25877 );
xor ( n39634 , n26343 , n25877 );
and ( n39635 , n34622 , n34629 );
and ( n39636 , n39634 , n39635 );
and ( n39637 , n39633 , n39636 );
xor ( n39638 , n39632 , n39637 );
and ( n39639 , n39638 , n26823 );
or ( n39640 , n39631 , n39639 );
buf ( n39641 , n39640 );
and ( n39642 , n39641 , n27046 );
and ( n39643 , n39641 , n27049 );
not ( n39644 , n27051 );
and ( n39645 , n39644 , n28236 );
not ( n39646 , n28494 );
and ( n39647 , n39646 , n28248 );
xor ( n39648 , n28248 , n27883 );
xor ( n39649 , n28226 , n27883 );
xor ( n39650 , n28204 , n27883 );
and ( n39651 , n34640 , n34647 );
and ( n39652 , n39650 , n39651 );
and ( n39653 , n39649 , n39652 );
xor ( n39654 , n39648 , n39653 );
and ( n39655 , n39654 , n28494 );
or ( n39656 , n39647 , n39655 );
buf ( n39657 , n39656 );
and ( n39658 , n39657 , n27051 );
or ( n39659 , n39645 , n39658 );
and ( n39660 , n39659 , n28506 );
and ( n39661 , n28236 , n28508 );
or ( n39662 , n39642 , n39643 , n39660 , n39661 );
and ( n39663 , n39662 , n28586 );
and ( n39664 , n26429 , n34573 );
or ( n39665 , n39663 , n39664 );
and ( n39666 , n39665 , n28594 );
not ( n39667 , n30249 );
and ( n39668 , n39667 , n30041 );
xor ( n39669 , n30041 , n29753 );
xor ( n39670 , n30024 , n29753 );
xor ( n39671 , n30007 , n29753 );
and ( n39672 , n34663 , n34670 );
and ( n39673 , n39671 , n39672 );
and ( n39674 , n39670 , n39673 );
xor ( n39675 , n39669 , n39674 );
and ( n39676 , n39675 , n30249 );
or ( n39677 , n39668 , n39676 );
buf ( n39678 , n39677 );
and ( n39679 , n39678 , n28586 );
and ( n39680 , n26429 , n34573 );
or ( n39681 , n39679 , n39680 );
and ( n39682 , n39681 , n30269 );
not ( n39683 , n30963 );
and ( n39684 , n39683 , n30755 );
xor ( n39685 , n30755 , n30467 );
xor ( n39686 , n30738 , n30467 );
xor ( n39687 , n30721 , n30467 );
and ( n39688 , n34681 , n34688 );
and ( n39689 , n39687 , n39688 );
and ( n39690 , n39686 , n39689 );
xor ( n39691 , n39685 , n39690 );
and ( n39692 , n39691 , n30963 );
or ( n39693 , n39684 , n39692 );
buf ( n39694 , n39693 );
and ( n39695 , n39694 , n28586 );
and ( n39696 , n26429 , n34573 );
or ( n39697 , n39695 , n39696 );
and ( n39698 , n39697 , n30982 );
and ( n39699 , n29335 , n28586 );
and ( n39700 , n26429 , n34573 );
or ( n39701 , n39699 , n39700 );
and ( n39702 , n39701 , n30989 );
buf ( n39703 , n29335 );
not ( n39704 , n39703 );
buf ( n39705 , n29355 );
not ( n39706 , n39705 );
buf ( n39707 , n29375 );
not ( n39708 , n39707 );
and ( n39709 , n34702 , n34712 );
and ( n39710 , n39708 , n39709 );
and ( n39711 , n39706 , n39710 );
xor ( n39712 , n39704 , n39711 );
buf ( n39713 , n39712 );
and ( n39714 , n39713 , n28586 );
and ( n39715 , n26429 , n34573 );
or ( n39716 , n39714 , n39715 );
and ( n39717 , n39716 , n31002 );
and ( n39718 , n26429 , n34607 );
or ( n39719 , n39666 , n39682 , n39698 , n39702 , n39717 , n39718 );
and ( n39720 , n39629 , n39719 );
and ( n39721 , n26429 , n24800 );
or ( n39722 , n39720 , n39721 );
and ( n39723 , n39722 , n31008 );
and ( n39724 , n26429 , n10618 );
or ( n39725 , n39723 , n39724 );
buf ( n39726 , n39725 );
buf ( n39727 , n39726 );
buf ( n39728 , n10615 );
not ( n39729 , n11333 );
and ( n39730 , n39729 , n11040 );
xor ( n39731 , n11349 , n11353 );
and ( n39732 , n39731 , n11333 );
or ( n39733 , n39730 , n39732 );
buf ( n39734 , n39733 );
buf ( n39735 , n39734 );
not ( n39736 , n11333 );
and ( n39737 , n39736 , n11159 );
xor ( n39738 , n11342 , n11360 );
and ( n39739 , n39738 , n11333 );
or ( n39740 , n39737 , n39739 );
buf ( n39741 , n39740 );
buf ( n39742 , n39741 );
not ( n39743 , n17451 );
and ( n39744 , n18841 , n17873 );
and ( n39745 , n34488 , n21330 );
and ( n39746 , n18841 , n21338 );
or ( n39747 , n39745 , n39746 );
and ( n39748 , n39747 , n21341 );
and ( n39749 , n34501 , n21330 );
and ( n39750 , n18841 , n21338 );
or ( n39751 , n39749 , n39750 );
and ( n39752 , n39751 , n23064 );
and ( n39753 , n34511 , n21330 );
and ( n39754 , n18841 , n21338 );
or ( n39755 , n39753 , n39754 );
and ( n39756 , n39755 , n23825 );
and ( n39757 , n22222 , n21330 );
and ( n39758 , n18841 , n21338 );
or ( n39759 , n39757 , n39758 );
and ( n39760 , n39759 , n23832 );
and ( n39761 , n18839 , n23834 );
and ( n39762 , n34521 , n21330 );
and ( n39763 , n18841 , n21338 );
or ( n39764 , n39762 , n39763 );
and ( n39765 , n39764 , n23917 );
or ( n39766 , n39744 , n39748 , n39752 , n39756 , n39760 , n39761 , n39765 );
and ( n39767 , n39743 , n39766 );
and ( n39768 , n18841 , n17451 );
or ( n39769 , n39767 , n39768 );
and ( n39770 , n39769 , n23924 );
and ( n39771 , n18841 , n23926 );
or ( n39772 , n39770 , n39771 );
buf ( n39773 , n39772 );
buf ( n39774 , n39773 );
buf ( n39775 , n10613 );
buf ( n39776 , n10615 );
buf ( n39777 , n10613 );
buf ( n39778 , n10615 );
buf ( n39779 , n10615 );
buf ( n39780 , n10615 );
buf ( n39781 , n10613 );
not ( n39782 , n24800 );
not ( n39783 , n26823 );
and ( n39784 , n39783 , n26003 );
xor ( n39785 , n31023 , n31030 );
and ( n39786 , n39785 , n26823 );
or ( n39787 , n39784 , n39786 );
buf ( n39788 , n39787 );
and ( n39789 , n39788 , n27046 );
and ( n39790 , n39788 , n27049 );
not ( n39791 , n27051 );
and ( n39792 , n39791 , n27972 );
not ( n39793 , n28494 );
and ( n39794 , n39793 , n27984 );
xor ( n39795 , n31051 , n31058 );
and ( n39796 , n39795 , n28494 );
or ( n39797 , n39794 , n39796 );
buf ( n39798 , n39797 );
and ( n39799 , n39798 , n27051 );
or ( n39800 , n39792 , n39799 );
and ( n39801 , n39800 , n28506 );
and ( n39802 , n27972 , n28508 );
or ( n39803 , n39789 , n39790 , n39801 , n39802 );
and ( n39804 , n39803 , n28587 );
or ( n39805 , n28586 , n28583 );
or ( n39806 , n39805 , n28589 );
or ( n39807 , n39806 , C0 );
and ( n39808 , n26023 , n39807 );
or ( n39809 , n39804 , n39808 );
and ( n39810 , n39809 , n28594 );
not ( n39811 , n30249 );
and ( n39812 , n39811 , n29837 );
xor ( n39813 , n31086 , n31093 );
and ( n39814 , n39813 , n30249 );
or ( n39815 , n39812 , n39814 );
buf ( n39816 , n39815 );
and ( n39817 , n39816 , n28587 );
and ( n39818 , n26023 , n39807 );
or ( n39819 , n39817 , n39818 );
and ( n39820 , n39819 , n30269 );
not ( n39821 , n30963 );
and ( n39822 , n39821 , n30551 );
xor ( n39823 , n31114 , n31121 );
and ( n39824 , n39823 , n30963 );
or ( n39825 , n39822 , n39824 );
buf ( n39826 , n39825 );
and ( n39827 , n39826 , n28587 );
and ( n39828 , n26023 , n39807 );
or ( n39829 , n39827 , n39828 );
and ( n39830 , n39829 , n30982 );
and ( n39831 , n29575 , n28587 );
and ( n39832 , n26023 , n39807 );
or ( n39833 , n39831 , n39832 );
and ( n39834 , n39833 , n30989 );
xor ( n39835 , n31151 , n31161 );
buf ( n39836 , n39835 );
and ( n39837 , n39836 , n28587 );
and ( n39838 , n26023 , n39807 );
or ( n39839 , n39837 , n39838 );
and ( n39840 , n39839 , n31002 );
and ( n39841 , n26023 , n34607 );
or ( n39842 , n39810 , n39820 , n39830 , n39834 , n39840 , n39841 );
and ( n39843 , n39782 , n39842 );
and ( n39844 , n26023 , n24800 );
or ( n39845 , n39843 , n39844 );
and ( n39846 , n39845 , n31008 );
and ( n39847 , n26023 , n10618 );
or ( n39848 , n39846 , n39847 );
buf ( n39849 , n39848 );
buf ( n39850 , n39849 );
not ( n39851 , n17451 );
not ( n39852 , n19474 );
and ( n39853 , n39852 , n19368 );
xor ( n39854 , n19368 , n18528 );
and ( n39855 , n19477 , n19525 );
xor ( n39856 , n39854 , n39855 );
and ( n39857 , n39856 , n19474 );
or ( n39858 , n39853 , n39857 );
buf ( n39859 , n39858 );
and ( n39860 , n39859 , n19745 );
and ( n39861 , n39859 , n19748 );
not ( n39862 , n19750 );
and ( n39863 , n39862 , n21133 );
not ( n39864 , n21193 );
and ( n39865 , n39864 , n21145 );
xor ( n39866 , n21145 , n20582 );
and ( n39867 , n21196 , n21246 );
xor ( n39868 , n39866 , n39867 );
and ( n39869 , n39868 , n21193 );
or ( n39870 , n39865 , n39869 );
buf ( n39871 , n39870 );
and ( n39872 , n39871 , n19750 );
or ( n39873 , n39863 , n39872 );
and ( n39874 , n39873 , n21253 );
and ( n39875 , n21133 , n21255 );
or ( n39876 , n39860 , n39861 , n39874 , n39875 );
and ( n39877 , n39876 , n21334 );
and ( n39878 , n19388 , n34492 );
or ( n39879 , n39877 , n39878 );
and ( n39880 , n39879 , n21341 );
not ( n39881 , n22996 );
and ( n39882 , n39881 , n22941 );
xor ( n39883 , n22941 , n22500 );
and ( n39884 , n22999 , n23049 );
xor ( n39885 , n39883 , n39884 );
and ( n39886 , n39885 , n22996 );
or ( n39887 , n39882 , n39886 );
buf ( n39888 , n39887 );
and ( n39889 , n39888 , n21334 );
and ( n39890 , n19388 , n34492 );
or ( n39891 , n39889 , n39890 );
and ( n39892 , n39891 , n23064 );
not ( n39893 , n23758 );
and ( n39894 , n39893 , n23703 );
xor ( n39895 , n23703 , n23262 );
and ( n39896 , n23761 , n23811 );
xor ( n39897 , n39895 , n39896 );
and ( n39898 , n39897 , n23758 );
or ( n39899 , n39894 , n39898 );
buf ( n39900 , n39899 );
and ( n39901 , n39900 , n21334 );
and ( n39902 , n19388 , n34492 );
or ( n39903 , n39901 , n39902 );
and ( n39904 , n39903 , n23825 );
and ( n39905 , n21906 , n21334 );
and ( n39906 , n19388 , n34492 );
or ( n39907 , n39905 , n39906 );
and ( n39908 , n39907 , n23832 );
buf ( n39909 , n21906 );
not ( n39910 , n39909 );
and ( n39911 , n23837 , n23911 );
xor ( n39912 , n39910 , n39911 );
buf ( n39913 , n39912 );
and ( n39914 , n39913 , n21334 );
and ( n39915 , n19388 , n34492 );
or ( n39916 , n39914 , n39915 );
and ( n39917 , n39916 , n23917 );
and ( n39918 , n19388 , n34526 );
or ( n39919 , n39880 , n39892 , n39904 , n39908 , n39917 , n39918 );
and ( n39920 , n39851 , n39919 );
and ( n39921 , n19388 , n17451 );
or ( n39922 , n39920 , n39921 );
and ( n39923 , n39922 , n23924 );
and ( n39924 , n19388 , n23926 );
or ( n39925 , n39923 , n39924 );
buf ( n39926 , n39925 );
buf ( n39927 , n39926 );
buf ( n39928 , n10615 );
buf ( n39929 , n10615 );
not ( n39930 , n24800 );
and ( n39931 , n25853 , n25222 );
not ( n39932 , n27051 );
and ( n39933 , n39932 , n27156 );
not ( n39934 , n28494 );
and ( n39935 , n39934 , n27162 );
xor ( n39936 , n28498 , n27883 );
and ( n39937 , n39936 , n28494 );
or ( n39938 , n39935 , n39937 );
buf ( n39939 , n39938 );
and ( n39940 , n39939 , n27051 );
or ( n39941 , n39933 , n39940 );
and ( n39942 , n39941 , n28506 );
and ( n39943 , n27156 , n28508 );
or ( n39944 , C0 , C0 , n39942 , n39943 );
and ( n39945 , n39944 , n28583 );
and ( n39946 , n25853 , n28591 );
or ( n39947 , n39945 , n39946 );
and ( n39948 , n39947 , n28594 );
not ( n39949 , n30249 );
and ( n39950 , n39949 , n28901 );
xor ( n39951 , n30253 , n29753 );
and ( n39952 , n39951 , n30249 );
or ( n39953 , n39950 , n39952 );
buf ( n39954 , n39953 );
and ( n39955 , n39954 , n28583 );
and ( n39956 , n25853 , n28591 );
or ( n39957 , n39955 , n39956 );
and ( n39958 , n39957 , n30269 );
not ( n39959 , n30963 );
and ( n39960 , n39959 , n30280 );
xor ( n39961 , n30967 , n30467 );
and ( n39962 , n39961 , n30963 );
or ( n39963 , n39960 , n39962 );
buf ( n39964 , n39963 );
and ( n39965 , n39964 , n28583 );
and ( n39966 , n25853 , n28591 );
or ( n39967 , n39965 , n39966 );
and ( n39968 , n39967 , n30982 );
and ( n39969 , n28892 , n28583 );
and ( n39970 , n25853 , n28591 );
or ( n39971 , n39969 , n39970 );
and ( n39972 , n39971 , n30989 );
and ( n39973 , n25663 , n30991 );
buf ( n39974 , n30995 );
and ( n39975 , n39974 , n28583 );
and ( n39976 , n25853 , n28591 );
or ( n39977 , n39975 , n39976 );
and ( n39978 , n39977 , n31002 );
or ( n39979 , n39931 , n39948 , n39958 , n39968 , n39972 , n39973 , n39978 );
and ( n39980 , n39930 , n39979 );
and ( n39981 , n25853 , n24800 );
or ( n39982 , n39980 , n39981 );
and ( n39983 , n39982 , n31008 );
and ( n39984 , n25853 , n10618 );
or ( n39985 , n39983 , n39984 );
buf ( n39986 , n39985 );
buf ( n39987 , n39986 );
buf ( n39988 , n10615 );
buf ( n39989 , n10615 );
not ( n39990 , n17451 );
not ( n39991 , n19474 );
and ( n39992 , n39991 , n18689 );
xor ( n39993 , n19496 , n19506 );
and ( n39994 , n39993 , n19474 );
or ( n39995 , n39992 , n39994 );
buf ( n39996 , n39995 );
and ( n39997 , n39996 , n19745 );
and ( n39998 , n39996 , n19748 );
not ( n39999 , n19750 );
and ( n40000 , n39999 , n20701 );
not ( n40001 , n21193 );
and ( n40002 , n40001 , n20713 );
xor ( n40003 , n21215 , n21227 );
and ( n40004 , n40003 , n21193 );
or ( n40005 , n40002 , n40004 );
buf ( n40006 , n40005 );
and ( n40007 , n40006 , n19750 );
or ( n40008 , n40000 , n40007 );
and ( n40009 , n40008 , n21253 );
and ( n40010 , n20701 , n21255 );
or ( n40011 , n39997 , n39998 , n40009 , n40010 );
and ( n40012 , n40011 , n21333 );
and ( n40013 , n18707 , n34758 );
or ( n40014 , n40012 , n40013 );
and ( n40015 , n40014 , n21341 );
not ( n40016 , n22996 );
and ( n40017 , n40016 , n22601 );
xor ( n40018 , n23018 , n23030 );
and ( n40019 , n40018 , n22996 );
or ( n40020 , n40017 , n40019 );
buf ( n40021 , n40020 );
and ( n40022 , n40021 , n21333 );
and ( n40023 , n18707 , n34758 );
or ( n40024 , n40022 , n40023 );
and ( n40025 , n40024 , n23064 );
not ( n40026 , n23758 );
and ( n40027 , n40026 , n23363 );
xor ( n40028 , n23780 , n23792 );
and ( n40029 , n40028 , n23758 );
or ( n40030 , n40027 , n40029 );
buf ( n40031 , n40030 );
and ( n40032 , n40031 , n21333 );
and ( n40033 , n18707 , n34758 );
or ( n40034 , n40032 , n40033 );
and ( n40035 , n40034 , n23825 );
and ( n40036 , n22302 , n21333 );
and ( n40037 , n18707 , n34758 );
or ( n40038 , n40036 , n40037 );
and ( n40039 , n40038 , n23832 );
xor ( n40040 , n23875 , n23892 );
buf ( n40041 , n40040 );
and ( n40042 , n40041 , n21333 );
and ( n40043 , n18707 , n34758 );
or ( n40044 , n40042 , n40043 );
and ( n40045 , n40044 , n23917 );
and ( n40046 , n18707 , n34526 );
or ( n40047 , n40015 , n40025 , n40035 , n40039 , n40045 , n40046 );
and ( n40048 , n39990 , n40047 );
and ( n40049 , n18707 , n17451 );
or ( n40050 , n40048 , n40049 );
and ( n40051 , n40050 , n23924 );
and ( n40052 , n18707 , n23926 );
or ( n40053 , n40051 , n40052 );
buf ( n40054 , n40053 );
buf ( n40055 , n40054 );
not ( n40056 , n17451 );
and ( n40057 , n20478 , n17873 );
xor ( n40058 , n19470 , n18528 );
xor ( n40059 , n19436 , n18528 );
xor ( n40060 , n19402 , n18528 );
and ( n40061 , n39854 , n39855 );
and ( n40062 , n40060 , n40061 );
and ( n40063 , n40059 , n40062 );
and ( n40064 , n40058 , n40063 );
buf ( n40065 , n40064 );
and ( n40066 , n40065 , n19474 );
or ( n40067 , C0 , n40066 );
buf ( n40068 , n40067 );
and ( n40069 , n40068 , n19745 );
and ( n40070 , n40068 , n19748 );
not ( n40071 , n19750 );
xor ( n40072 , n20518 , n20575 );
buf ( n40073 , n40072 );
and ( n40074 , n40073 , n19753 );
or ( n40075 , C0 , n40074 );
buf ( n40076 , n40075 );
and ( n40077 , n40071 , n40076 );
or ( n40078 , n40077 , C0 );
and ( n40079 , n40078 , n21253 );
and ( n40080 , n40076 , n21255 );
or ( n40081 , n40069 , n40070 , n40079 , n40080 );
and ( n40082 , n40081 , n21330 );
and ( n40083 , n20478 , n21338 );
or ( n40084 , n40082 , n40083 );
and ( n40085 , n40084 , n21341 );
xor ( n40086 , n22992 , n22500 );
xor ( n40087 , n22975 , n22500 );
xor ( n40088 , n22958 , n22500 );
and ( n40089 , n39883 , n39884 );
and ( n40090 , n40088 , n40089 );
and ( n40091 , n40087 , n40090 );
and ( n40092 , n40086 , n40091 );
buf ( n40093 , n40092 );
and ( n40094 , n40093 , n22996 );
or ( n40095 , C0 , n40094 );
buf ( n40096 , n40095 );
and ( n40097 , n40096 , n21330 );
and ( n40098 , n20478 , n21338 );
or ( n40099 , n40097 , n40098 );
and ( n40100 , n40099 , n23064 );
xor ( n40101 , n23754 , n23262 );
xor ( n40102 , n23737 , n23262 );
xor ( n40103 , n23720 , n23262 );
and ( n40104 , n39895 , n39896 );
and ( n40105 , n40103 , n40104 );
and ( n40106 , n40102 , n40105 );
and ( n40107 , n40101 , n40106 );
buf ( n40108 , n40107 );
and ( n40109 , n40108 , n23758 );
or ( n40110 , C0 , n40109 );
buf ( n40111 , n40110 );
and ( n40112 , n40111 , n21330 );
and ( n40113 , n20478 , n21338 );
or ( n40114 , n40112 , n40113 );
and ( n40115 , n40114 , n23825 );
and ( n40116 , n21854 , n21330 );
and ( n40117 , n20478 , n21338 );
or ( n40118 , n40116 , n40117 );
and ( n40119 , n40118 , n23832 );
and ( n40120 , n20476 , n23834 );
buf ( n40121 , n21854 );
not ( n40122 , n40121 );
buf ( n40123 , n21867 );
not ( n40124 , n40123 );
buf ( n40125 , n21880 );
not ( n40126 , n40125 );
buf ( n40127 , n21893 );
not ( n40128 , n40127 );
and ( n40129 , n39910 , n39911 );
and ( n40130 , n40128 , n40129 );
and ( n40131 , n40126 , n40130 );
and ( n40132 , n40124 , n40131 );
xor ( n40133 , n40122 , n40132 );
buf ( n40134 , n40133 );
and ( n40135 , n40134 , n21330 );
and ( n40136 , n20478 , n21338 );
or ( n40137 , n40135 , n40136 );
and ( n40138 , n40137 , n23917 );
or ( n40139 , n40057 , n40085 , n40100 , n40115 , n40119 , n40120 , n40138 );
and ( n40140 , n40056 , n40139 );
and ( n40141 , n20478 , n17451 );
or ( n40142 , n40140 , n40141 );
and ( n40143 , n40142 , n23924 );
and ( n40144 , n20478 , n23926 );
or ( n40145 , n40143 , n40144 );
buf ( n40146 , n40145 );
buf ( n40147 , n40146 );
buf ( n40148 , n10615 );
buf ( n40149 , n10613 );
buf ( n40150 , n10613 );
buf ( n40151 , n10615 );
not ( n40152 , n24511 );
not ( n40153 , n24799 );
or ( n40154 , n28594 , n25222 );
and ( n40155 , n10660 , n40154 );
buf ( n40156 , n28890 );
buf ( n40157 , n25853 );
xor ( n40158 , n40156 , n40157 );
buf ( n40159 , n40158 );
buf ( n40160 , n40159 );
buf ( n40161 , n40160 );
not ( n40162 , n40161 );
buf ( n40163 , n40162 );
buf ( n40164 , n40163 );
not ( n40165 , n40164 );
buf ( n40166 , n25870 );
buf ( n40167 , n27175 );
buf ( n40168 , n27187 );
buf ( n40169 , n26801 );
buf ( n40170 , n26767 );
buf ( n40171 , n26733 );
buf ( n40172 , n26699 );
buf ( n40173 , n26665 );
buf ( n40174 , n26631 );
buf ( n40175 , n26597 );
buf ( n40176 , n26563 );
buf ( n40177 , n26529 );
buf ( n40178 , n29293 );
buf ( n40179 , n26495 );
and ( n40180 , n40178 , n40179 );
buf ( n40181 , n29313 );
buf ( n40182 , n26461 );
and ( n40183 , n40181 , n40182 );
buf ( n40184 , n29333 );
buf ( n40185 , n26427 );
and ( n40186 , n40184 , n40185 );
buf ( n40187 , n29353 );
buf ( n40188 , n26393 );
and ( n40189 , n40187 , n40188 );
buf ( n40190 , n29373 );
buf ( n40191 , n26359 );
and ( n40192 , n40190 , n40191 );
buf ( n40193 , n29393 );
buf ( n40194 , n26325 );
and ( n40195 , n40193 , n40194 );
buf ( n40196 , n29413 );
buf ( n40197 , n26291 );
and ( n40198 , n40196 , n40197 );
buf ( n40199 , n29433 );
buf ( n40200 , n26257 );
and ( n40201 , n40199 , n40200 );
buf ( n40202 , n29453 );
buf ( n40203 , n26223 );
and ( n40204 , n40202 , n40203 );
buf ( n40205 , n29473 );
buf ( n40206 , n26189 );
and ( n40207 , n40205 , n40206 );
buf ( n40208 , n29493 );
buf ( n40209 , n26155 );
and ( n40210 , n40208 , n40209 );
buf ( n40211 , n29513 );
buf ( n40212 , n26121 );
and ( n40213 , n40211 , n40212 );
buf ( n40214 , n29533 );
buf ( n40215 , n26087 );
and ( n40216 , n40214 , n40215 );
buf ( n40217 , n29553 );
buf ( n40218 , n26053 );
and ( n40219 , n40217 , n40218 );
buf ( n40220 , n29573 );
buf ( n40221 , n26019 );
and ( n40222 , n40220 , n40221 );
buf ( n40223 , n29593 );
buf ( n40224 , n25985 );
and ( n40225 , n40223 , n40224 );
buf ( n40226 , n29613 );
buf ( n40227 , n25952 );
and ( n40228 , n40226 , n40227 );
buf ( n40229 , n29633 );
buf ( n40230 , n25919 );
and ( n40231 , n40229 , n40230 );
buf ( n40232 , n29653 );
buf ( n40233 , n24802 );
and ( n40234 , n40232 , n40233 );
and ( n40235 , n40156 , n40157 );
and ( n40236 , n40233 , n40235 );
and ( n40237 , n40232 , n40235 );
or ( n40238 , n40234 , n40236 , n40237 );
and ( n40239 , n40230 , n40238 );
and ( n40240 , n40229 , n40238 );
or ( n40241 , n40231 , n40239 , n40240 );
and ( n40242 , n40227 , n40241 );
and ( n40243 , n40226 , n40241 );
or ( n40244 , n40228 , n40242 , n40243 );
and ( n40245 , n40224 , n40244 );
and ( n40246 , n40223 , n40244 );
or ( n40247 , n40225 , n40245 , n40246 );
and ( n40248 , n40221 , n40247 );
and ( n40249 , n40220 , n40247 );
or ( n40250 , n40222 , n40248 , n40249 );
and ( n40251 , n40218 , n40250 );
and ( n40252 , n40217 , n40250 );
or ( n40253 , n40219 , n40251 , n40252 );
and ( n40254 , n40215 , n40253 );
and ( n40255 , n40214 , n40253 );
or ( n40256 , n40216 , n40254 , n40255 );
and ( n40257 , n40212 , n40256 );
and ( n40258 , n40211 , n40256 );
or ( n40259 , n40213 , n40257 , n40258 );
and ( n40260 , n40209 , n40259 );
and ( n40261 , n40208 , n40259 );
or ( n40262 , n40210 , n40260 , n40261 );
and ( n40263 , n40206 , n40262 );
and ( n40264 , n40205 , n40262 );
or ( n40265 , n40207 , n40263 , n40264 );
and ( n40266 , n40203 , n40265 );
and ( n40267 , n40202 , n40265 );
or ( n40268 , n40204 , n40266 , n40267 );
and ( n40269 , n40200 , n40268 );
and ( n40270 , n40199 , n40268 );
or ( n40271 , n40201 , n40269 , n40270 );
and ( n40272 , n40197 , n40271 );
and ( n40273 , n40196 , n40271 );
or ( n40274 , n40198 , n40272 , n40273 );
and ( n40275 , n40194 , n40274 );
and ( n40276 , n40193 , n40274 );
or ( n40277 , n40195 , n40275 , n40276 );
and ( n40278 , n40191 , n40277 );
and ( n40279 , n40190 , n40277 );
or ( n40280 , n40192 , n40278 , n40279 );
and ( n40281 , n40188 , n40280 );
and ( n40282 , n40187 , n40280 );
or ( n40283 , n40189 , n40281 , n40282 );
and ( n40284 , n40185 , n40283 );
and ( n40285 , n40184 , n40283 );
or ( n40286 , n40186 , n40284 , n40285 );
and ( n40287 , n40182 , n40286 );
and ( n40288 , n40181 , n40286 );
or ( n40289 , n40183 , n40287 , n40288 );
and ( n40290 , n40179 , n40289 );
and ( n40291 , n40178 , n40289 );
or ( n40292 , n40180 , n40290 , n40291 );
and ( n40293 , n40177 , n40292 );
and ( n40294 , n40176 , n40293 );
and ( n40295 , n40175 , n40294 );
and ( n40296 , n40174 , n40295 );
and ( n40297 , n40173 , n40296 );
and ( n40298 , n40172 , n40297 );
and ( n40299 , n40171 , n40298 );
and ( n40300 , n40170 , n40299 );
and ( n40301 , n40169 , n40300 );
and ( n40302 , n40168 , n40301 );
and ( n40303 , n40167 , n40302 );
xor ( n40304 , n40166 , n40303 );
buf ( n40305 , n40304 );
buf ( n40306 , n40305 );
not ( n40307 , n40306 );
xor ( n40308 , n40232 , n40233 );
xor ( n40309 , n40308 , n40235 );
buf ( n40310 , n40309 );
buf ( n40311 , n40310 );
and ( n40312 , n40307 , n40311 );
not ( n40313 , n40311 );
not ( n40314 , n40160 );
xor ( n40315 , n40313 , n40314 );
and ( n40316 , n40315 , n40306 );
or ( n40317 , n40312 , n40316 );
buf ( n40318 , n40317 );
not ( n40319 , n40318 );
buf ( n40320 , n40319 );
buf ( n40321 , n40320 );
not ( n40322 , n40321 );
or ( n40323 , n40165 , n40322 );
not ( n40324 , n40306 );
xor ( n40325 , n40229 , n40230 );
xor ( n40326 , n40325 , n40238 );
buf ( n40327 , n40326 );
buf ( n40328 , n40327 );
and ( n40329 , n40324 , n40328 );
not ( n40330 , n40328 );
and ( n40331 , n40313 , n40314 );
xor ( n40332 , n40330 , n40331 );
and ( n40333 , n40332 , n40306 );
or ( n40334 , n40329 , n40333 );
buf ( n40335 , n40334 );
not ( n40336 , n40335 );
buf ( n40337 , n40336 );
buf ( n40338 , n40337 );
not ( n40339 , n40338 );
or ( n40340 , n40323 , n40339 );
not ( n40341 , n40306 );
xor ( n40342 , n40226 , n40227 );
xor ( n40343 , n40342 , n40241 );
buf ( n40344 , n40343 );
buf ( n40345 , n40344 );
and ( n40346 , n40341 , n40345 );
not ( n40347 , n40345 );
and ( n40348 , n40330 , n40331 );
xor ( n40349 , n40347 , n40348 );
and ( n40350 , n40349 , n40306 );
or ( n40351 , n40346 , n40350 );
buf ( n40352 , n40351 );
not ( n40353 , n40352 );
buf ( n40354 , n40353 );
buf ( n40355 , n40354 );
not ( n40356 , n40355 );
or ( n40357 , n40340 , n40356 );
not ( n40358 , n40306 );
xor ( n40359 , n40223 , n40224 );
xor ( n40360 , n40359 , n40244 );
buf ( n40361 , n40360 );
buf ( n40362 , n40361 );
and ( n40363 , n40358 , n40362 );
not ( n40364 , n40362 );
and ( n40365 , n40347 , n40348 );
xor ( n40366 , n40364 , n40365 );
and ( n40367 , n40366 , n40306 );
or ( n40368 , n40363 , n40367 );
buf ( n40369 , n40368 );
not ( n40370 , n40369 );
buf ( n40371 , n40370 );
buf ( n40372 , n40371 );
not ( n40373 , n40372 );
or ( n40374 , n40357 , n40373 );
not ( n40375 , n40306 );
xor ( n40376 , n40220 , n40221 );
xor ( n40377 , n40376 , n40247 );
buf ( n40378 , n40377 );
buf ( n40379 , n40378 );
and ( n40380 , n40375 , n40379 );
not ( n40381 , n40379 );
and ( n40382 , n40364 , n40365 );
xor ( n40383 , n40381 , n40382 );
and ( n40384 , n40383 , n40306 );
or ( n40385 , n40380 , n40384 );
buf ( n40386 , n40385 );
not ( n40387 , n40386 );
buf ( n40388 , n40387 );
buf ( n40389 , n40388 );
not ( n40390 , n40389 );
or ( n40391 , n40374 , n40390 );
not ( n40392 , n40306 );
xor ( n40393 , n40217 , n40218 );
xor ( n40394 , n40393 , n40250 );
buf ( n40395 , n40394 );
buf ( n40396 , n40395 );
and ( n40397 , n40392 , n40396 );
not ( n40398 , n40396 );
and ( n40399 , n40381 , n40382 );
xor ( n40400 , n40398 , n40399 );
and ( n40401 , n40400 , n40306 );
or ( n40402 , n40397 , n40401 );
buf ( n40403 , n40402 );
not ( n40404 , n40403 );
buf ( n40405 , n40404 );
buf ( n40406 , n40405 );
not ( n40407 , n40406 );
or ( n40408 , n40391 , n40407 );
not ( n40409 , n40306 );
xor ( n40410 , n40214 , n40215 );
xor ( n40411 , n40410 , n40253 );
buf ( n40412 , n40411 );
buf ( n40413 , n40412 );
and ( n40414 , n40409 , n40413 );
not ( n40415 , n40413 );
and ( n40416 , n40398 , n40399 );
xor ( n40417 , n40415 , n40416 );
and ( n40418 , n40417 , n40306 );
or ( n40419 , n40414 , n40418 );
buf ( n40420 , n40419 );
not ( n40421 , n40420 );
buf ( n40422 , n40421 );
buf ( n40423 , n40422 );
not ( n40424 , n40423 );
or ( n40425 , n40408 , n40424 );
not ( n40426 , n40306 );
xor ( n40427 , n40211 , n40212 );
xor ( n40428 , n40427 , n40256 );
buf ( n40429 , n40428 );
buf ( n40430 , n40429 );
and ( n40431 , n40426 , n40430 );
not ( n40432 , n40430 );
and ( n40433 , n40415 , n40416 );
xor ( n40434 , n40432 , n40433 );
and ( n40435 , n40434 , n40306 );
or ( n40436 , n40431 , n40435 );
buf ( n40437 , n40436 );
not ( n40438 , n40437 );
buf ( n40439 , n40438 );
buf ( n40440 , n40439 );
not ( n40441 , n40440 );
or ( n40442 , n40425 , n40441 );
not ( n40443 , n40306 );
xor ( n40444 , n40208 , n40209 );
xor ( n40445 , n40444 , n40259 );
buf ( n40446 , n40445 );
buf ( n40447 , n40446 );
and ( n40448 , n40443 , n40447 );
not ( n40449 , n40447 );
and ( n40450 , n40432 , n40433 );
xor ( n40451 , n40449 , n40450 );
and ( n40452 , n40451 , n40306 );
or ( n40453 , n40448 , n40452 );
buf ( n40454 , n40453 );
not ( n40455 , n40454 );
buf ( n40456 , n40455 );
buf ( n40457 , n40456 );
not ( n40458 , n40457 );
or ( n40459 , n40442 , n40458 );
not ( n40460 , n40306 );
xor ( n40461 , n40205 , n40206 );
xor ( n40462 , n40461 , n40262 );
buf ( n40463 , n40462 );
buf ( n40464 , n40463 );
and ( n40465 , n40460 , n40464 );
not ( n40466 , n40464 );
and ( n40467 , n40449 , n40450 );
xor ( n40468 , n40466 , n40467 );
and ( n40469 , n40468 , n40306 );
or ( n40470 , n40465 , n40469 );
buf ( n40471 , n40470 );
not ( n40472 , n40471 );
buf ( n40473 , n40472 );
buf ( n40474 , n40473 );
not ( n40475 , n40474 );
or ( n40476 , n40459 , n40475 );
not ( n40477 , n40306 );
xor ( n40478 , n40202 , n40203 );
xor ( n40479 , n40478 , n40265 );
buf ( n40480 , n40479 );
buf ( n40481 , n40480 );
and ( n40482 , n40477 , n40481 );
not ( n40483 , n40481 );
and ( n40484 , n40466 , n40467 );
xor ( n40485 , n40483 , n40484 );
and ( n40486 , n40485 , n40306 );
or ( n40487 , n40482 , n40486 );
buf ( n40488 , n40487 );
not ( n40489 , n40488 );
buf ( n40490 , n40489 );
buf ( n40491 , n40490 );
not ( n40492 , n40491 );
or ( n40493 , n40476 , n40492 );
not ( n40494 , n40306 );
xor ( n40495 , n40199 , n40200 );
xor ( n40496 , n40495 , n40268 );
buf ( n40497 , n40496 );
buf ( n40498 , n40497 );
and ( n40499 , n40494 , n40498 );
not ( n40500 , n40498 );
and ( n40501 , n40483 , n40484 );
xor ( n40502 , n40500 , n40501 );
and ( n40503 , n40502 , n40306 );
or ( n40504 , n40499 , n40503 );
buf ( n40505 , n40504 );
not ( n40506 , n40505 );
buf ( n40507 , n40506 );
buf ( n40508 , n40507 );
not ( n40509 , n40508 );
or ( n40510 , n40493 , n40509 );
not ( n40511 , n40306 );
xor ( n40512 , n40196 , n40197 );
xor ( n40513 , n40512 , n40271 );
buf ( n40514 , n40513 );
buf ( n40515 , n40514 );
and ( n40516 , n40511 , n40515 );
not ( n40517 , n40515 );
and ( n40518 , n40500 , n40501 );
xor ( n40519 , n40517 , n40518 );
and ( n40520 , n40519 , n40306 );
or ( n40521 , n40516 , n40520 );
buf ( n40522 , n40521 );
not ( n40523 , n40522 );
buf ( n40524 , n40523 );
buf ( n40525 , n40524 );
not ( n40526 , n40525 );
or ( n40527 , n40510 , n40526 );
not ( n40528 , n40306 );
xor ( n40529 , n40193 , n40194 );
xor ( n40530 , n40529 , n40274 );
buf ( n40531 , n40530 );
buf ( n40532 , n40531 );
and ( n40533 , n40528 , n40532 );
not ( n40534 , n40532 );
and ( n40535 , n40517 , n40518 );
xor ( n40536 , n40534 , n40535 );
and ( n40537 , n40536 , n40306 );
or ( n40538 , n40533 , n40537 );
buf ( n40539 , n40538 );
not ( n40540 , n40539 );
buf ( n40541 , n40540 );
buf ( n40542 , n40541 );
not ( n40543 , n40542 );
or ( n40544 , n40527 , n40543 );
not ( n40545 , n40306 );
xor ( n40546 , n40190 , n40191 );
xor ( n40547 , n40546 , n40277 );
buf ( n40548 , n40547 );
buf ( n40549 , n40548 );
and ( n40550 , n40545 , n40549 );
not ( n40551 , n40549 );
and ( n40552 , n40534 , n40535 );
xor ( n40553 , n40551 , n40552 );
and ( n40554 , n40553 , n40306 );
or ( n40555 , n40550 , n40554 );
buf ( n40556 , n40555 );
not ( n40557 , n40556 );
buf ( n40558 , n40557 );
buf ( n40559 , n40558 );
not ( n40560 , n40559 );
or ( n40561 , n40544 , n40560 );
not ( n40562 , n40306 );
xor ( n40563 , n40187 , n40188 );
xor ( n40564 , n40563 , n40280 );
buf ( n40565 , n40564 );
buf ( n40566 , n40565 );
and ( n40567 , n40562 , n40566 );
not ( n40568 , n40566 );
and ( n40569 , n40551 , n40552 );
xor ( n40570 , n40568 , n40569 );
and ( n40571 , n40570 , n40306 );
or ( n40572 , n40567 , n40571 );
buf ( n40573 , n40572 );
not ( n40574 , n40573 );
buf ( n40575 , n40574 );
buf ( n40576 , n40575 );
not ( n40577 , n40576 );
or ( n40578 , n40561 , n40577 );
not ( n40579 , n40306 );
xor ( n40580 , n40184 , n40185 );
xor ( n40581 , n40580 , n40283 );
buf ( n40582 , n40581 );
buf ( n40583 , n40582 );
and ( n40584 , n40579 , n40583 );
not ( n40585 , n40583 );
and ( n40586 , n40568 , n40569 );
xor ( n40587 , n40585 , n40586 );
and ( n40588 , n40587 , n40306 );
or ( n40589 , n40584 , n40588 );
buf ( n40590 , n40589 );
not ( n40591 , n40590 );
buf ( n40592 , n40591 );
buf ( n40593 , n40592 );
not ( n40594 , n40593 );
or ( n40595 , n40578 , n40594 );
not ( n40596 , n40306 );
xor ( n40597 , n40181 , n40182 );
xor ( n40598 , n40597 , n40286 );
buf ( n40599 , n40598 );
buf ( n40600 , n40599 );
and ( n40601 , n40596 , n40600 );
not ( n40602 , n40600 );
and ( n40603 , n40585 , n40586 );
xor ( n40604 , n40602 , n40603 );
and ( n40605 , n40604 , n40306 );
or ( n40606 , n40601 , n40605 );
buf ( n40607 , n40606 );
not ( n40608 , n40607 );
buf ( n40609 , n40608 );
buf ( n40610 , n40609 );
not ( n40611 , n40610 );
or ( n40612 , n40595 , n40611 );
not ( n40613 , n40306 );
xor ( n40614 , n40178 , n40179 );
xor ( n40615 , n40614 , n40289 );
buf ( n40616 , n40615 );
buf ( n40617 , n40616 );
and ( n40618 , n40613 , n40617 );
not ( n40619 , n40617 );
and ( n40620 , n40602 , n40603 );
xor ( n40621 , n40619 , n40620 );
and ( n40622 , n40621 , n40306 );
or ( n40623 , n40618 , n40622 );
buf ( n40624 , n40623 );
not ( n40625 , n40624 );
buf ( n40626 , n40625 );
buf ( n40627 , n40626 );
not ( n40628 , n40627 );
or ( n40629 , n40612 , n40628 );
buf ( n40630 , n40629 );
buf ( n40631 , n40630 );
and ( n40632 , n40631 , n40306 );
not ( n40633 , n40632 );
and ( n40634 , n40633 , n40560 );
xor ( n40635 , n40560 , n40306 );
xor ( n40636 , n40543 , n40306 );
xor ( n40637 , n40526 , n40306 );
xor ( n40638 , n40509 , n40306 );
xor ( n40639 , n40492 , n40306 );
xor ( n40640 , n40475 , n40306 );
xor ( n40641 , n40458 , n40306 );
xor ( n40642 , n40441 , n40306 );
xor ( n40643 , n40424 , n40306 );
xor ( n40644 , n40407 , n40306 );
xor ( n40645 , n40390 , n40306 );
xor ( n40646 , n40373 , n40306 );
xor ( n40647 , n40356 , n40306 );
xor ( n40648 , n40339 , n40306 );
xor ( n40649 , n40322 , n40306 );
xor ( n40650 , n40165 , n40306 );
and ( n40651 , n40650 , n40306 );
and ( n40652 , n40649 , n40651 );
and ( n40653 , n40648 , n40652 );
and ( n40654 , n40647 , n40653 );
and ( n40655 , n40646 , n40654 );
and ( n40656 , n40645 , n40655 );
and ( n40657 , n40644 , n40656 );
and ( n40658 , n40643 , n40657 );
and ( n40659 , n40642 , n40658 );
and ( n40660 , n40641 , n40659 );
and ( n40661 , n40640 , n40660 );
and ( n40662 , n40639 , n40661 );
and ( n40663 , n40638 , n40662 );
and ( n40664 , n40637 , n40663 );
and ( n40665 , n40636 , n40664 );
xor ( n40666 , n40635 , n40665 );
and ( n40667 , n40666 , n40632 );
or ( n40668 , n40634 , n40667 );
buf ( n40669 , n40668 );
and ( n40670 , n40669 , n27046 );
buf ( n40671 , n28890 );
buf ( n40672 , n25857 );
xor ( n40673 , n40671 , n40672 );
buf ( n40674 , n40673 );
buf ( n40675 , n40674 );
buf ( n40676 , n40675 );
not ( n40677 , n40676 );
buf ( n40678 , n40677 );
buf ( n40679 , n40678 );
not ( n40680 , n40679 );
buf ( n40681 , n25872 );
buf ( n40682 , n27177 );
buf ( n40683 , n27189 );
buf ( n40684 , n26803 );
buf ( n40685 , n26769 );
buf ( n40686 , n26735 );
buf ( n40687 , n26701 );
buf ( n40688 , n26667 );
buf ( n40689 , n26633 );
buf ( n40690 , n26599 );
buf ( n40691 , n26565 );
buf ( n40692 , n26531 );
buf ( n40693 , n29293 );
buf ( n40694 , n26497 );
and ( n40695 , n40693 , n40694 );
buf ( n40696 , n29313 );
buf ( n40697 , n26463 );
and ( n40698 , n40696 , n40697 );
buf ( n40699 , n29333 );
buf ( n40700 , n26429 );
and ( n40701 , n40699 , n40700 );
buf ( n40702 , n29353 );
buf ( n40703 , n26395 );
and ( n40704 , n40702 , n40703 );
buf ( n40705 , n29373 );
buf ( n40706 , n26361 );
and ( n40707 , n40705 , n40706 );
buf ( n40708 , n29393 );
buf ( n40709 , n26327 );
and ( n40710 , n40708 , n40709 );
buf ( n40711 , n29413 );
buf ( n40712 , n26293 );
and ( n40713 , n40711 , n40712 );
buf ( n40714 , n29433 );
buf ( n40715 , n26259 );
and ( n40716 , n40714 , n40715 );
buf ( n40717 , n29453 );
buf ( n40718 , n26225 );
and ( n40719 , n40717 , n40718 );
buf ( n40720 , n29473 );
buf ( n40721 , n26191 );
and ( n40722 , n40720 , n40721 );
buf ( n40723 , n29493 );
buf ( n40724 , n26157 );
and ( n40725 , n40723 , n40724 );
buf ( n40726 , n29513 );
buf ( n40727 , n26123 );
and ( n40728 , n40726 , n40727 );
buf ( n40729 , n29533 );
buf ( n40730 , n26089 );
and ( n40731 , n40729 , n40730 );
buf ( n40732 , n29553 );
buf ( n40733 , n26055 );
and ( n40734 , n40732 , n40733 );
buf ( n40735 , n29573 );
buf ( n40736 , n26021 );
and ( n40737 , n40735 , n40736 );
buf ( n40738 , n29593 );
buf ( n40739 , n25987 );
and ( n40740 , n40738 , n40739 );
buf ( n40741 , n29613 );
buf ( n40742 , n25954 );
and ( n40743 , n40741 , n40742 );
buf ( n40744 , n29633 );
buf ( n40745 , n25921 );
and ( n40746 , n40744 , n40745 );
buf ( n40747 , n29653 );
buf ( n40748 , n25890 );
and ( n40749 , n40747 , n40748 );
and ( n40750 , n40671 , n40672 );
and ( n40751 , n40748 , n40750 );
and ( n40752 , n40747 , n40750 );
or ( n40753 , n40749 , n40751 , n40752 );
and ( n40754 , n40745 , n40753 );
and ( n40755 , n40744 , n40753 );
or ( n40756 , n40746 , n40754 , n40755 );
and ( n40757 , n40742 , n40756 );
and ( n40758 , n40741 , n40756 );
or ( n40759 , n40743 , n40757 , n40758 );
and ( n40760 , n40739 , n40759 );
and ( n40761 , n40738 , n40759 );
or ( n40762 , n40740 , n40760 , n40761 );
and ( n40763 , n40736 , n40762 );
and ( n40764 , n40735 , n40762 );
or ( n40765 , n40737 , n40763 , n40764 );
and ( n40766 , n40733 , n40765 );
and ( n40767 , n40732 , n40765 );
or ( n40768 , n40734 , n40766 , n40767 );
and ( n40769 , n40730 , n40768 );
and ( n40770 , n40729 , n40768 );
or ( n40771 , n40731 , n40769 , n40770 );
and ( n40772 , n40727 , n40771 );
and ( n40773 , n40726 , n40771 );
or ( n40774 , n40728 , n40772 , n40773 );
and ( n40775 , n40724 , n40774 );
and ( n40776 , n40723 , n40774 );
or ( n40777 , n40725 , n40775 , n40776 );
and ( n40778 , n40721 , n40777 );
and ( n40779 , n40720 , n40777 );
or ( n40780 , n40722 , n40778 , n40779 );
and ( n40781 , n40718 , n40780 );
and ( n40782 , n40717 , n40780 );
or ( n40783 , n40719 , n40781 , n40782 );
and ( n40784 , n40715 , n40783 );
and ( n40785 , n40714 , n40783 );
or ( n40786 , n40716 , n40784 , n40785 );
and ( n40787 , n40712 , n40786 );
and ( n40788 , n40711 , n40786 );
or ( n40789 , n40713 , n40787 , n40788 );
and ( n40790 , n40709 , n40789 );
and ( n40791 , n40708 , n40789 );
or ( n40792 , n40710 , n40790 , n40791 );
and ( n40793 , n40706 , n40792 );
and ( n40794 , n40705 , n40792 );
or ( n40795 , n40707 , n40793 , n40794 );
and ( n40796 , n40703 , n40795 );
and ( n40797 , n40702 , n40795 );
or ( n40798 , n40704 , n40796 , n40797 );
and ( n40799 , n40700 , n40798 );
and ( n40800 , n40699 , n40798 );
or ( n40801 , n40701 , n40799 , n40800 );
and ( n40802 , n40697 , n40801 );
and ( n40803 , n40696 , n40801 );
or ( n40804 , n40698 , n40802 , n40803 );
and ( n40805 , n40694 , n40804 );
and ( n40806 , n40693 , n40804 );
or ( n40807 , n40695 , n40805 , n40806 );
and ( n40808 , n40692 , n40807 );
and ( n40809 , n40691 , n40808 );
and ( n40810 , n40690 , n40809 );
and ( n40811 , n40689 , n40810 );
and ( n40812 , n40688 , n40811 );
and ( n40813 , n40687 , n40812 );
and ( n40814 , n40686 , n40813 );
and ( n40815 , n40685 , n40814 );
and ( n40816 , n40684 , n40815 );
and ( n40817 , n40683 , n40816 );
and ( n40818 , n40682 , n40817 );
xor ( n40819 , n40681 , n40818 );
buf ( n40820 , n40819 );
buf ( n40821 , n40820 );
not ( n40822 , n40821 );
xor ( n40823 , n40747 , n40748 );
xor ( n40824 , n40823 , n40750 );
buf ( n40825 , n40824 );
buf ( n40826 , n40825 );
and ( n40827 , n40822 , n40826 );
not ( n40828 , n40826 );
not ( n40829 , n40675 );
xor ( n40830 , n40828 , n40829 );
and ( n40831 , n40830 , n40821 );
or ( n40832 , n40827 , n40831 );
buf ( n40833 , n40832 );
not ( n40834 , n40833 );
buf ( n40835 , n40834 );
buf ( n40836 , n40835 );
not ( n40837 , n40836 );
or ( n40838 , n40680 , n40837 );
not ( n40839 , n40821 );
xor ( n40840 , n40744 , n40745 );
xor ( n40841 , n40840 , n40753 );
buf ( n40842 , n40841 );
buf ( n40843 , n40842 );
and ( n40844 , n40839 , n40843 );
not ( n40845 , n40843 );
and ( n40846 , n40828 , n40829 );
xor ( n40847 , n40845 , n40846 );
and ( n40848 , n40847 , n40821 );
or ( n40849 , n40844 , n40848 );
buf ( n40850 , n40849 );
not ( n40851 , n40850 );
buf ( n40852 , n40851 );
buf ( n40853 , n40852 );
not ( n40854 , n40853 );
or ( n40855 , n40838 , n40854 );
not ( n40856 , n40821 );
xor ( n40857 , n40741 , n40742 );
xor ( n40858 , n40857 , n40756 );
buf ( n40859 , n40858 );
buf ( n40860 , n40859 );
and ( n40861 , n40856 , n40860 );
not ( n40862 , n40860 );
and ( n40863 , n40845 , n40846 );
xor ( n40864 , n40862 , n40863 );
and ( n40865 , n40864 , n40821 );
or ( n40866 , n40861 , n40865 );
buf ( n40867 , n40866 );
not ( n40868 , n40867 );
buf ( n40869 , n40868 );
buf ( n40870 , n40869 );
not ( n40871 , n40870 );
or ( n40872 , n40855 , n40871 );
not ( n40873 , n40821 );
xor ( n40874 , n40738 , n40739 );
xor ( n40875 , n40874 , n40759 );
buf ( n40876 , n40875 );
buf ( n40877 , n40876 );
and ( n40878 , n40873 , n40877 );
not ( n40879 , n40877 );
and ( n40880 , n40862 , n40863 );
xor ( n40881 , n40879 , n40880 );
and ( n40882 , n40881 , n40821 );
or ( n40883 , n40878 , n40882 );
buf ( n40884 , n40883 );
not ( n40885 , n40884 );
buf ( n40886 , n40885 );
buf ( n40887 , n40886 );
not ( n40888 , n40887 );
or ( n40889 , n40872 , n40888 );
not ( n40890 , n40821 );
xor ( n40891 , n40735 , n40736 );
xor ( n40892 , n40891 , n40762 );
buf ( n40893 , n40892 );
buf ( n40894 , n40893 );
and ( n40895 , n40890 , n40894 );
not ( n40896 , n40894 );
and ( n40897 , n40879 , n40880 );
xor ( n40898 , n40896 , n40897 );
and ( n40899 , n40898 , n40821 );
or ( n40900 , n40895 , n40899 );
buf ( n40901 , n40900 );
not ( n40902 , n40901 );
buf ( n40903 , n40902 );
buf ( n40904 , n40903 );
not ( n40905 , n40904 );
or ( n40906 , n40889 , n40905 );
not ( n40907 , n40821 );
xor ( n40908 , n40732 , n40733 );
xor ( n40909 , n40908 , n40765 );
buf ( n40910 , n40909 );
buf ( n40911 , n40910 );
and ( n40912 , n40907 , n40911 );
not ( n40913 , n40911 );
and ( n40914 , n40896 , n40897 );
xor ( n40915 , n40913 , n40914 );
and ( n40916 , n40915 , n40821 );
or ( n40917 , n40912 , n40916 );
buf ( n40918 , n40917 );
not ( n40919 , n40918 );
buf ( n40920 , n40919 );
buf ( n40921 , n40920 );
not ( n40922 , n40921 );
or ( n40923 , n40906 , n40922 );
not ( n40924 , n40821 );
xor ( n40925 , n40729 , n40730 );
xor ( n40926 , n40925 , n40768 );
buf ( n40927 , n40926 );
buf ( n40928 , n40927 );
and ( n40929 , n40924 , n40928 );
not ( n40930 , n40928 );
and ( n40931 , n40913 , n40914 );
xor ( n40932 , n40930 , n40931 );
and ( n40933 , n40932 , n40821 );
or ( n40934 , n40929 , n40933 );
buf ( n40935 , n40934 );
not ( n40936 , n40935 );
buf ( n40937 , n40936 );
buf ( n40938 , n40937 );
not ( n40939 , n40938 );
or ( n40940 , n40923 , n40939 );
not ( n40941 , n40821 );
xor ( n40942 , n40726 , n40727 );
xor ( n40943 , n40942 , n40771 );
buf ( n40944 , n40943 );
buf ( n40945 , n40944 );
and ( n40946 , n40941 , n40945 );
not ( n40947 , n40945 );
and ( n40948 , n40930 , n40931 );
xor ( n40949 , n40947 , n40948 );
and ( n40950 , n40949 , n40821 );
or ( n40951 , n40946 , n40950 );
buf ( n40952 , n40951 );
not ( n40953 , n40952 );
buf ( n40954 , n40953 );
buf ( n40955 , n40954 );
not ( n40956 , n40955 );
or ( n40957 , n40940 , n40956 );
not ( n40958 , n40821 );
xor ( n40959 , n40723 , n40724 );
xor ( n40960 , n40959 , n40774 );
buf ( n40961 , n40960 );
buf ( n40962 , n40961 );
and ( n40963 , n40958 , n40962 );
not ( n40964 , n40962 );
and ( n40965 , n40947 , n40948 );
xor ( n40966 , n40964 , n40965 );
and ( n40967 , n40966 , n40821 );
or ( n40968 , n40963 , n40967 );
buf ( n40969 , n40968 );
not ( n40970 , n40969 );
buf ( n40971 , n40970 );
buf ( n40972 , n40971 );
not ( n40973 , n40972 );
or ( n40974 , n40957 , n40973 );
not ( n40975 , n40821 );
xor ( n40976 , n40720 , n40721 );
xor ( n40977 , n40976 , n40777 );
buf ( n40978 , n40977 );
buf ( n40979 , n40978 );
and ( n40980 , n40975 , n40979 );
not ( n40981 , n40979 );
and ( n40982 , n40964 , n40965 );
xor ( n40983 , n40981 , n40982 );
and ( n40984 , n40983 , n40821 );
or ( n40985 , n40980 , n40984 );
buf ( n40986 , n40985 );
not ( n40987 , n40986 );
buf ( n40988 , n40987 );
buf ( n40989 , n40988 );
not ( n40990 , n40989 );
or ( n40991 , n40974 , n40990 );
not ( n40992 , n40821 );
xor ( n40993 , n40717 , n40718 );
xor ( n40994 , n40993 , n40780 );
buf ( n40995 , n40994 );
buf ( n40996 , n40995 );
and ( n40997 , n40992 , n40996 );
not ( n40998 , n40996 );
and ( n40999 , n40981 , n40982 );
xor ( n41000 , n40998 , n40999 );
and ( n41001 , n41000 , n40821 );
or ( n41002 , n40997 , n41001 );
buf ( n41003 , n41002 );
not ( n41004 , n41003 );
buf ( n41005 , n41004 );
buf ( n41006 , n41005 );
not ( n41007 , n41006 );
or ( n41008 , n40991 , n41007 );
not ( n41009 , n40821 );
xor ( n41010 , n40714 , n40715 );
xor ( n41011 , n41010 , n40783 );
buf ( n41012 , n41011 );
buf ( n41013 , n41012 );
and ( n41014 , n41009 , n41013 );
not ( n41015 , n41013 );
and ( n41016 , n40998 , n40999 );
xor ( n41017 , n41015 , n41016 );
and ( n41018 , n41017 , n40821 );
or ( n41019 , n41014 , n41018 );
buf ( n41020 , n41019 );
not ( n41021 , n41020 );
buf ( n41022 , n41021 );
buf ( n41023 , n41022 );
not ( n41024 , n41023 );
or ( n41025 , n41008 , n41024 );
not ( n41026 , n40821 );
xor ( n41027 , n40711 , n40712 );
xor ( n41028 , n41027 , n40786 );
buf ( n41029 , n41028 );
buf ( n41030 , n41029 );
and ( n41031 , n41026 , n41030 );
not ( n41032 , n41030 );
and ( n41033 , n41015 , n41016 );
xor ( n41034 , n41032 , n41033 );
and ( n41035 , n41034 , n40821 );
or ( n41036 , n41031 , n41035 );
buf ( n41037 , n41036 );
not ( n41038 , n41037 );
buf ( n41039 , n41038 );
buf ( n41040 , n41039 );
not ( n41041 , n41040 );
or ( n41042 , n41025 , n41041 );
not ( n41043 , n40821 );
xor ( n41044 , n40708 , n40709 );
xor ( n41045 , n41044 , n40789 );
buf ( n41046 , n41045 );
buf ( n41047 , n41046 );
and ( n41048 , n41043 , n41047 );
not ( n41049 , n41047 );
and ( n41050 , n41032 , n41033 );
xor ( n41051 , n41049 , n41050 );
and ( n41052 , n41051 , n40821 );
or ( n41053 , n41048 , n41052 );
buf ( n41054 , n41053 );
not ( n41055 , n41054 );
buf ( n41056 , n41055 );
buf ( n41057 , n41056 );
not ( n41058 , n41057 );
or ( n41059 , n41042 , n41058 );
not ( n41060 , n40821 );
xor ( n41061 , n40705 , n40706 );
xor ( n41062 , n41061 , n40792 );
buf ( n41063 , n41062 );
buf ( n41064 , n41063 );
and ( n41065 , n41060 , n41064 );
not ( n41066 , n41064 );
and ( n41067 , n41049 , n41050 );
xor ( n41068 , n41066 , n41067 );
and ( n41069 , n41068 , n40821 );
or ( n41070 , n41065 , n41069 );
buf ( n41071 , n41070 );
not ( n41072 , n41071 );
buf ( n41073 , n41072 );
buf ( n41074 , n41073 );
not ( n41075 , n41074 );
or ( n41076 , n41059 , n41075 );
not ( n41077 , n40821 );
xor ( n41078 , n40702 , n40703 );
xor ( n41079 , n41078 , n40795 );
buf ( n41080 , n41079 );
buf ( n41081 , n41080 );
and ( n41082 , n41077 , n41081 );
not ( n41083 , n41081 );
and ( n41084 , n41066 , n41067 );
xor ( n41085 , n41083 , n41084 );
and ( n41086 , n41085 , n40821 );
or ( n41087 , n41082 , n41086 );
buf ( n41088 , n41087 );
not ( n41089 , n41088 );
buf ( n41090 , n41089 );
buf ( n41091 , n41090 );
not ( n41092 , n41091 );
or ( n41093 , n41076 , n41092 );
not ( n41094 , n40821 );
xor ( n41095 , n40699 , n40700 );
xor ( n41096 , n41095 , n40798 );
buf ( n41097 , n41096 );
buf ( n41098 , n41097 );
and ( n41099 , n41094 , n41098 );
not ( n41100 , n41098 );
and ( n41101 , n41083 , n41084 );
xor ( n41102 , n41100 , n41101 );
and ( n41103 , n41102 , n40821 );
or ( n41104 , n41099 , n41103 );
buf ( n41105 , n41104 );
not ( n41106 , n41105 );
buf ( n41107 , n41106 );
buf ( n41108 , n41107 );
not ( n41109 , n41108 );
or ( n41110 , n41093 , n41109 );
not ( n41111 , n40821 );
xor ( n41112 , n40696 , n40697 );
xor ( n41113 , n41112 , n40801 );
buf ( n41114 , n41113 );
buf ( n41115 , n41114 );
and ( n41116 , n41111 , n41115 );
not ( n41117 , n41115 );
and ( n41118 , n41100 , n41101 );
xor ( n41119 , n41117 , n41118 );
and ( n41120 , n41119 , n40821 );
or ( n41121 , n41116 , n41120 );
buf ( n41122 , n41121 );
not ( n41123 , n41122 );
buf ( n41124 , n41123 );
buf ( n41125 , n41124 );
not ( n41126 , n41125 );
or ( n41127 , n41110 , n41126 );
not ( n41128 , n40821 );
xor ( n41129 , n40693 , n40694 );
xor ( n41130 , n41129 , n40804 );
buf ( n41131 , n41130 );
buf ( n41132 , n41131 );
and ( n41133 , n41128 , n41132 );
not ( n41134 , n41132 );
and ( n41135 , n41117 , n41118 );
xor ( n41136 , n41134 , n41135 );
and ( n41137 , n41136 , n40821 );
or ( n41138 , n41133 , n41137 );
buf ( n41139 , n41138 );
not ( n41140 , n41139 );
buf ( n41141 , n41140 );
buf ( n41142 , n41141 );
not ( n41143 , n41142 );
or ( n41144 , n41127 , n41143 );
buf ( n41145 , n41144 );
buf ( n41146 , n41145 );
and ( n41147 , n41146 , n40821 );
not ( n41148 , n41147 );
and ( n41149 , n41148 , n41075 );
xor ( n41150 , n41075 , n40821 );
xor ( n41151 , n41058 , n40821 );
xor ( n41152 , n41041 , n40821 );
xor ( n41153 , n41024 , n40821 );
xor ( n41154 , n41007 , n40821 );
xor ( n41155 , n40990 , n40821 );
xor ( n41156 , n40973 , n40821 );
xor ( n41157 , n40956 , n40821 );
xor ( n41158 , n40939 , n40821 );
xor ( n41159 , n40922 , n40821 );
xor ( n41160 , n40905 , n40821 );
xor ( n41161 , n40888 , n40821 );
xor ( n41162 , n40871 , n40821 );
xor ( n41163 , n40854 , n40821 );
xor ( n41164 , n40837 , n40821 );
xor ( n41165 , n40680 , n40821 );
and ( n41166 , n41165 , n40821 );
and ( n41167 , n41164 , n41166 );
and ( n41168 , n41163 , n41167 );
and ( n41169 , n41162 , n41168 );
and ( n41170 , n41161 , n41169 );
and ( n41171 , n41160 , n41170 );
and ( n41172 , n41159 , n41171 );
and ( n41173 , n41158 , n41172 );
and ( n41174 , n41157 , n41173 );
and ( n41175 , n41156 , n41174 );
and ( n41176 , n41155 , n41175 );
and ( n41177 , n41154 , n41176 );
and ( n41178 , n41153 , n41177 );
and ( n41179 , n41152 , n41178 );
and ( n41180 , n41151 , n41179 );
xor ( n41181 , n41150 , n41180 );
and ( n41182 , n41181 , n41147 );
or ( n41183 , n41149 , n41182 );
buf ( n41184 , n41183 );
and ( n41185 , n41184 , n27049 );
and ( n41186 , n29373 , n28506 );
and ( n41187 , n10660 , n28508 );
or ( n41188 , n40670 , n41185 , n41186 , n41187 );
or ( n41189 , n31002 , n30991 );
or ( n41190 , n41189 , n30987 );
or ( n41191 , n41190 , n30988 );
or ( n41192 , n41191 , n30976 );
or ( n41193 , n41192 , n30977 );
or ( n41194 , n41193 , n30263 );
or ( n41195 , n41194 , n30264 );
or ( n41196 , n41195 , n30979 );
or ( n41197 , n41196 , n30266 );
or ( n41198 , n41197 , n30981 );
or ( n41199 , n41198 , n30268 );
and ( n41200 , n41188 , n41199 );
or ( n41201 , n40155 , n41200 );
and ( n41202 , n40153 , n41201 );
buf ( n41203 , n25853 );
buf ( n41204 , n41203 );
not ( n41205 , n41204 );
buf ( n41206 , n41205 );
buf ( n41207 , n41206 );
not ( n41208 , n41207 );
buf ( n41209 , n25870 );
not ( n41210 , n41209 );
buf ( n41211 , n24802 );
and ( n41212 , n41210 , n41211 );
not ( n41213 , n41211 );
not ( n41214 , n41203 );
xor ( n41215 , n41213 , n41214 );
and ( n41216 , n41215 , n41209 );
or ( n41217 , n41212 , n41216 );
buf ( n41218 , n41217 );
not ( n41219 , n41218 );
buf ( n41220 , n41219 );
buf ( n41221 , n41220 );
not ( n41222 , n41221 );
or ( n41223 , n41208 , n41222 );
not ( n41224 , n41209 );
buf ( n41225 , n25919 );
and ( n41226 , n41224 , n41225 );
not ( n41227 , n41225 );
and ( n41228 , n41213 , n41214 );
xor ( n41229 , n41227 , n41228 );
and ( n41230 , n41229 , n41209 );
or ( n41231 , n41226 , n41230 );
buf ( n41232 , n41231 );
not ( n41233 , n41232 );
buf ( n41234 , n41233 );
buf ( n41235 , n41234 );
not ( n41236 , n41235 );
or ( n41237 , n41223 , n41236 );
not ( n41238 , n41209 );
buf ( n41239 , n25952 );
and ( n41240 , n41238 , n41239 );
not ( n41241 , n41239 );
and ( n41242 , n41227 , n41228 );
xor ( n41243 , n41241 , n41242 );
and ( n41244 , n41243 , n41209 );
or ( n41245 , n41240 , n41244 );
buf ( n41246 , n41245 );
not ( n41247 , n41246 );
buf ( n41248 , n41247 );
buf ( n41249 , n41248 );
not ( n41250 , n41249 );
or ( n41251 , n41237 , n41250 );
not ( n41252 , n41209 );
buf ( n41253 , n25985 );
and ( n41254 , n41252 , n41253 );
not ( n41255 , n41253 );
and ( n41256 , n41241 , n41242 );
xor ( n41257 , n41255 , n41256 );
and ( n41258 , n41257 , n41209 );
or ( n41259 , n41254 , n41258 );
buf ( n41260 , n41259 );
not ( n41261 , n41260 );
buf ( n41262 , n41261 );
buf ( n41263 , n41262 );
not ( n41264 , n41263 );
or ( n41265 , n41251 , n41264 );
not ( n41266 , n41209 );
buf ( n41267 , n26019 );
and ( n41268 , n41266 , n41267 );
not ( n41269 , n41267 );
and ( n41270 , n41255 , n41256 );
xor ( n41271 , n41269 , n41270 );
and ( n41272 , n41271 , n41209 );
or ( n41273 , n41268 , n41272 );
buf ( n41274 , n41273 );
not ( n41275 , n41274 );
buf ( n41276 , n41275 );
buf ( n41277 , n41276 );
not ( n41278 , n41277 );
or ( n41279 , n41265 , n41278 );
not ( n41280 , n41209 );
buf ( n41281 , n26053 );
and ( n41282 , n41280 , n41281 );
not ( n41283 , n41281 );
and ( n41284 , n41269 , n41270 );
xor ( n41285 , n41283 , n41284 );
and ( n41286 , n41285 , n41209 );
or ( n41287 , n41282 , n41286 );
buf ( n41288 , n41287 );
not ( n41289 , n41288 );
buf ( n41290 , n41289 );
buf ( n41291 , n41290 );
not ( n41292 , n41291 );
or ( n41293 , n41279 , n41292 );
not ( n41294 , n41209 );
buf ( n41295 , n26087 );
and ( n41296 , n41294 , n41295 );
not ( n41297 , n41295 );
and ( n41298 , n41283 , n41284 );
xor ( n41299 , n41297 , n41298 );
and ( n41300 , n41299 , n41209 );
or ( n41301 , n41296 , n41300 );
buf ( n41302 , n41301 );
not ( n41303 , n41302 );
buf ( n41304 , n41303 );
buf ( n41305 , n41304 );
not ( n41306 , n41305 );
or ( n41307 , n41293 , n41306 );
not ( n41308 , n41209 );
buf ( n41309 , n26121 );
and ( n41310 , n41308 , n41309 );
not ( n41311 , n41309 );
and ( n41312 , n41297 , n41298 );
xor ( n41313 , n41311 , n41312 );
and ( n41314 , n41313 , n41209 );
or ( n41315 , n41310 , n41314 );
buf ( n41316 , n41315 );
not ( n41317 , n41316 );
buf ( n41318 , n41317 );
buf ( n41319 , n41318 );
not ( n41320 , n41319 );
or ( n41321 , n41307 , n41320 );
not ( n41322 , n41209 );
buf ( n41323 , n26155 );
and ( n41324 , n41322 , n41323 );
not ( n41325 , n41323 );
and ( n41326 , n41311 , n41312 );
xor ( n41327 , n41325 , n41326 );
and ( n41328 , n41327 , n41209 );
or ( n41329 , n41324 , n41328 );
buf ( n41330 , n41329 );
not ( n41331 , n41330 );
buf ( n41332 , n41331 );
buf ( n41333 , n41332 );
not ( n41334 , n41333 );
or ( n41335 , n41321 , n41334 );
not ( n41336 , n41209 );
buf ( n41337 , n26189 );
and ( n41338 , n41336 , n41337 );
not ( n41339 , n41337 );
and ( n41340 , n41325 , n41326 );
xor ( n41341 , n41339 , n41340 );
and ( n41342 , n41341 , n41209 );
or ( n41343 , n41338 , n41342 );
buf ( n41344 , n41343 );
not ( n41345 , n41344 );
buf ( n41346 , n41345 );
buf ( n41347 , n41346 );
not ( n41348 , n41347 );
or ( n41349 , n41335 , n41348 );
not ( n41350 , n41209 );
buf ( n41351 , n26223 );
and ( n41352 , n41350 , n41351 );
not ( n41353 , n41351 );
and ( n41354 , n41339 , n41340 );
xor ( n41355 , n41353 , n41354 );
and ( n41356 , n41355 , n41209 );
or ( n41357 , n41352 , n41356 );
buf ( n41358 , n41357 );
not ( n41359 , n41358 );
buf ( n41360 , n41359 );
buf ( n41361 , n41360 );
not ( n41362 , n41361 );
or ( n41363 , n41349 , n41362 );
not ( n41364 , n41209 );
buf ( n41365 , n26257 );
and ( n41366 , n41364 , n41365 );
not ( n41367 , n41365 );
and ( n41368 , n41353 , n41354 );
xor ( n41369 , n41367 , n41368 );
and ( n41370 , n41369 , n41209 );
or ( n41371 , n41366 , n41370 );
buf ( n41372 , n41371 );
not ( n41373 , n41372 );
buf ( n41374 , n41373 );
buf ( n41375 , n41374 );
not ( n41376 , n41375 );
or ( n41377 , n41363 , n41376 );
not ( n41378 , n41209 );
buf ( n41379 , n26291 );
and ( n41380 , n41378 , n41379 );
not ( n41381 , n41379 );
and ( n41382 , n41367 , n41368 );
xor ( n41383 , n41381 , n41382 );
and ( n41384 , n41383 , n41209 );
or ( n41385 , n41380 , n41384 );
buf ( n41386 , n41385 );
not ( n41387 , n41386 );
buf ( n41388 , n41387 );
buf ( n41389 , n41388 );
not ( n41390 , n41389 );
or ( n41391 , n41377 , n41390 );
not ( n41392 , n41209 );
buf ( n41393 , n26325 );
and ( n41394 , n41392 , n41393 );
not ( n41395 , n41393 );
and ( n41396 , n41381 , n41382 );
xor ( n41397 , n41395 , n41396 );
and ( n41398 , n41397 , n41209 );
or ( n41399 , n41394 , n41398 );
buf ( n41400 , n41399 );
not ( n41401 , n41400 );
buf ( n41402 , n41401 );
buf ( n41403 , n41402 );
not ( n41404 , n41403 );
or ( n41405 , n41391 , n41404 );
not ( n41406 , n41209 );
buf ( n41407 , n26359 );
and ( n41408 , n41406 , n41407 );
not ( n41409 , n41407 );
and ( n41410 , n41395 , n41396 );
xor ( n41411 , n41409 , n41410 );
and ( n41412 , n41411 , n41209 );
or ( n41413 , n41408 , n41412 );
buf ( n41414 , n41413 );
not ( n41415 , n41414 );
buf ( n41416 , n41415 );
buf ( n41417 , n41416 );
not ( n41418 , n41417 );
or ( n41419 , n41405 , n41418 );
not ( n41420 , n41209 );
buf ( n41421 , n26393 );
and ( n41422 , n41420 , n41421 );
not ( n41423 , n41421 );
and ( n41424 , n41409 , n41410 );
xor ( n41425 , n41423 , n41424 );
and ( n41426 , n41425 , n41209 );
or ( n41427 , n41422 , n41426 );
buf ( n41428 , n41427 );
not ( n41429 , n41428 );
buf ( n41430 , n41429 );
buf ( n41431 , n41430 );
not ( n41432 , n41431 );
or ( n41433 , n41419 , n41432 );
not ( n41434 , n41209 );
buf ( n41435 , n26427 );
and ( n41436 , n41434 , n41435 );
not ( n41437 , n41435 );
and ( n41438 , n41423 , n41424 );
xor ( n41439 , n41437 , n41438 );
and ( n41440 , n41439 , n41209 );
or ( n41441 , n41436 , n41440 );
buf ( n41442 , n41441 );
not ( n41443 , n41442 );
buf ( n41444 , n41443 );
buf ( n41445 , n41444 );
not ( n41446 , n41445 );
or ( n41447 , n41433 , n41446 );
not ( n41448 , n41209 );
buf ( n41449 , n26461 );
and ( n41450 , n41448 , n41449 );
not ( n41451 , n41449 );
and ( n41452 , n41437 , n41438 );
xor ( n41453 , n41451 , n41452 );
and ( n41454 , n41453 , n41209 );
or ( n41455 , n41450 , n41454 );
buf ( n41456 , n41455 );
not ( n41457 , n41456 );
buf ( n41458 , n41457 );
buf ( n41459 , n41458 );
not ( n41460 , n41459 );
or ( n41461 , n41447 , n41460 );
not ( n41462 , n41209 );
buf ( n41463 , n26495 );
and ( n41464 , n41462 , n41463 );
not ( n41465 , n41463 );
and ( n41466 , n41451 , n41452 );
xor ( n41467 , n41465 , n41466 );
and ( n41468 , n41467 , n41209 );
or ( n41469 , n41464 , n41468 );
buf ( n41470 , n41469 );
not ( n41471 , n41470 );
buf ( n41472 , n41471 );
buf ( n41473 , n41472 );
not ( n41474 , n41473 );
or ( n41475 , n41461 , n41474 );
buf ( n41476 , n41475 );
buf ( n41477 , n41476 );
and ( n41478 , n41477 , n41209 );
not ( n41479 , n41478 );
and ( n41480 , n41479 , n41418 );
xor ( n41481 , n41418 , n41209 );
xor ( n41482 , n41404 , n41209 );
xor ( n41483 , n41390 , n41209 );
xor ( n41484 , n41376 , n41209 );
xor ( n41485 , n41362 , n41209 );
xor ( n41486 , n41348 , n41209 );
xor ( n41487 , n41334 , n41209 );
xor ( n41488 , n41320 , n41209 );
xor ( n41489 , n41306 , n41209 );
xor ( n41490 , n41292 , n41209 );
xor ( n41491 , n41278 , n41209 );
xor ( n41492 , n41264 , n41209 );
xor ( n41493 , n41250 , n41209 );
xor ( n41494 , n41236 , n41209 );
xor ( n41495 , n41222 , n41209 );
xor ( n41496 , n41208 , n41209 );
and ( n41497 , n41496 , n41209 );
and ( n41498 , n41495 , n41497 );
and ( n41499 , n41494 , n41498 );
and ( n41500 , n41493 , n41499 );
and ( n41501 , n41492 , n41500 );
and ( n41502 , n41491 , n41501 );
and ( n41503 , n41490 , n41502 );
and ( n41504 , n41489 , n41503 );
and ( n41505 , n41488 , n41504 );
and ( n41506 , n41487 , n41505 );
and ( n41507 , n41486 , n41506 );
and ( n41508 , n41485 , n41507 );
and ( n41509 , n41484 , n41508 );
and ( n41510 , n41483 , n41509 );
and ( n41511 , n41482 , n41510 );
xor ( n41512 , n41481 , n41511 );
and ( n41513 , n41512 , n41478 );
or ( n41514 , n41480 , n41513 );
buf ( n41515 , n41514 );
buf ( n41516 , n41515 );
buf ( n41517 , n29373 );
not ( n41518 , n41517 );
buf ( n41519 , n41518 );
buf ( n41520 , n41519 );
not ( n41521 , n41520 );
buf ( n41522 , n41521 );
buf ( n41523 , n41522 );
buf ( n41524 , n41523 );
xor ( n41525 , n41516 , n41524 );
not ( n41526 , n41478 );
and ( n41527 , n41526 , n41404 );
xor ( n41528 , n41482 , n41510 );
and ( n41529 , n41528 , n41478 );
or ( n41530 , n41527 , n41529 );
buf ( n41531 , n41530 );
buf ( n41532 , n41531 );
buf ( n41533 , n29393 );
not ( n41534 , n41533 );
buf ( n41535 , n41534 );
buf ( n41536 , n41535 );
not ( n41537 , n41536 );
buf ( n41538 , n41537 );
buf ( n41539 , n41538 );
buf ( n41540 , n41539 );
and ( n41541 , n41532 , n41540 );
not ( n41542 , n41478 );
and ( n41543 , n41542 , n41390 );
xor ( n41544 , n41483 , n41509 );
and ( n41545 , n41544 , n41478 );
or ( n41546 , n41543 , n41545 );
buf ( n41547 , n41546 );
buf ( n41548 , n41547 );
buf ( n41549 , n29413 );
not ( n41550 , n41549 );
buf ( n41551 , n41550 );
buf ( n41552 , n41551 );
not ( n41553 , n41552 );
buf ( n41554 , n41553 );
buf ( n41555 , n41554 );
buf ( n41556 , n41555 );
and ( n41557 , n41548 , n41556 );
not ( n41558 , n41478 );
and ( n41559 , n41558 , n41376 );
xor ( n41560 , n41484 , n41508 );
and ( n41561 , n41560 , n41478 );
or ( n41562 , n41559 , n41561 );
buf ( n41563 , n41562 );
buf ( n41564 , n41563 );
buf ( n41565 , n29433 );
not ( n41566 , n41565 );
buf ( n41567 , n41566 );
buf ( n41568 , n41567 );
not ( n41569 , n41568 );
buf ( n41570 , n41569 );
buf ( n41571 , n41570 );
buf ( n41572 , n41571 );
and ( n41573 , n41564 , n41572 );
not ( n41574 , n41478 );
and ( n41575 , n41574 , n41362 );
xor ( n41576 , n41485 , n41507 );
and ( n41577 , n41576 , n41478 );
or ( n41578 , n41575 , n41577 );
buf ( n41579 , n41578 );
buf ( n41580 , n41579 );
buf ( n41581 , n29453 );
not ( n41582 , n41581 );
buf ( n41583 , n41582 );
buf ( n41584 , n41583 );
not ( n41585 , n41584 );
buf ( n41586 , n41585 );
buf ( n41587 , n41586 );
buf ( n41588 , n41587 );
and ( n41589 , n41580 , n41588 );
not ( n41590 , n41478 );
and ( n41591 , n41590 , n41348 );
xor ( n41592 , n41486 , n41506 );
and ( n41593 , n41592 , n41478 );
or ( n41594 , n41591 , n41593 );
buf ( n41595 , n41594 );
buf ( n41596 , n41595 );
buf ( n41597 , n29473 );
not ( n41598 , n41597 );
buf ( n41599 , n41598 );
buf ( n41600 , n41599 );
not ( n41601 , n41600 );
buf ( n41602 , n41601 );
buf ( n41603 , n41602 );
buf ( n41604 , n41603 );
and ( n41605 , n41596 , n41604 );
not ( n41606 , n41478 );
and ( n41607 , n41606 , n41334 );
xor ( n41608 , n41487 , n41505 );
and ( n41609 , n41608 , n41478 );
or ( n41610 , n41607 , n41609 );
buf ( n41611 , n41610 );
buf ( n41612 , n41611 );
buf ( n41613 , n29493 );
not ( n41614 , n41613 );
buf ( n41615 , n41614 );
buf ( n41616 , n41615 );
not ( n41617 , n41616 );
buf ( n41618 , n41617 );
buf ( n41619 , n41618 );
buf ( n41620 , n41619 );
and ( n41621 , n41612 , n41620 );
not ( n41622 , n41478 );
and ( n41623 , n41622 , n41320 );
xor ( n41624 , n41488 , n41504 );
and ( n41625 , n41624 , n41478 );
or ( n41626 , n41623 , n41625 );
buf ( n41627 , n41626 );
buf ( n41628 , n41627 );
buf ( n41629 , n29513 );
not ( n41630 , n41629 );
buf ( n41631 , n41630 );
buf ( n41632 , n41631 );
not ( n41633 , n41632 );
buf ( n41634 , n41633 );
buf ( n41635 , n41634 );
buf ( n41636 , n41635 );
and ( n41637 , n41628 , n41636 );
not ( n41638 , n41478 );
and ( n41639 , n41638 , n41306 );
xor ( n41640 , n41489 , n41503 );
and ( n41641 , n41640 , n41478 );
or ( n41642 , n41639 , n41641 );
buf ( n41643 , n41642 );
buf ( n41644 , n41643 );
buf ( n41645 , n29533 );
not ( n41646 , n41645 );
buf ( n41647 , n41646 );
buf ( n41648 , n41647 );
not ( n41649 , n41648 );
buf ( n41650 , n41649 );
buf ( n41651 , n41650 );
buf ( n41652 , n41651 );
and ( n41653 , n41644 , n41652 );
not ( n41654 , n41478 );
and ( n41655 , n41654 , n41292 );
xor ( n41656 , n41490 , n41502 );
and ( n41657 , n41656 , n41478 );
or ( n41658 , n41655 , n41657 );
buf ( n41659 , n41658 );
buf ( n41660 , n41659 );
buf ( n41661 , n29553 );
not ( n41662 , n41661 );
buf ( n41663 , n41662 );
buf ( n41664 , n41663 );
not ( n41665 , n41664 );
buf ( n41666 , n41665 );
buf ( n41667 , n41666 );
buf ( n41668 , n41667 );
and ( n41669 , n41660 , n41668 );
not ( n41670 , n41478 );
and ( n41671 , n41670 , n41278 );
xor ( n41672 , n41491 , n41501 );
and ( n41673 , n41672 , n41478 );
or ( n41674 , n41671 , n41673 );
buf ( n41675 , n41674 );
buf ( n41676 , n41675 );
buf ( n41677 , n29573 );
not ( n41678 , n41677 );
buf ( n41679 , n41678 );
buf ( n41680 , n41679 );
not ( n41681 , n41680 );
buf ( n41682 , n41681 );
buf ( n41683 , n41682 );
buf ( n41684 , n41683 );
and ( n41685 , n41676 , n41684 );
not ( n41686 , n41478 );
and ( n41687 , n41686 , n41264 );
xor ( n41688 , n41492 , n41500 );
and ( n41689 , n41688 , n41478 );
or ( n41690 , n41687 , n41689 );
buf ( n41691 , n41690 );
buf ( n41692 , n41691 );
buf ( n41693 , n29593 );
not ( n41694 , n41693 );
buf ( n41695 , n41694 );
buf ( n41696 , n41695 );
not ( n41697 , n41696 );
buf ( n41698 , n41697 );
buf ( n41699 , n41698 );
buf ( n41700 , n41699 );
and ( n41701 , n41692 , n41700 );
not ( n41702 , n41478 );
and ( n41703 , n41702 , n41250 );
xor ( n41704 , n41493 , n41499 );
and ( n41705 , n41704 , n41478 );
or ( n41706 , n41703 , n41705 );
buf ( n41707 , n41706 );
buf ( n41708 , n41707 );
buf ( n41709 , n29613 );
not ( n41710 , n41709 );
buf ( n41711 , n41710 );
buf ( n41712 , n41711 );
not ( n41713 , n41712 );
buf ( n41714 , n41713 );
buf ( n41715 , n41714 );
buf ( n41716 , n41715 );
and ( n41717 , n41708 , n41716 );
not ( n41718 , n41478 );
and ( n41719 , n41718 , n41236 );
xor ( n41720 , n41494 , n41498 );
and ( n41721 , n41720 , n41478 );
or ( n41722 , n41719 , n41721 );
buf ( n41723 , n41722 );
buf ( n41724 , n41723 );
buf ( n41725 , n29633 );
not ( n41726 , n41725 );
buf ( n41727 , n41726 );
buf ( n41728 , n41727 );
not ( n41729 , n41728 );
buf ( n41730 , n41729 );
buf ( n41731 , n41730 );
buf ( n41732 , n41731 );
and ( n41733 , n41724 , n41732 );
not ( n41734 , n41478 );
and ( n41735 , n41734 , n41222 );
xor ( n41736 , n41495 , n41497 );
and ( n41737 , n41736 , n41478 );
or ( n41738 , n41735 , n41737 );
buf ( n41739 , n41738 );
buf ( n41740 , n41739 );
buf ( n41741 , n29653 );
not ( n41742 , n41741 );
buf ( n41743 , n41742 );
buf ( n41744 , n41743 );
not ( n41745 , n41744 );
buf ( n41746 , n41745 );
buf ( n41747 , n41746 );
buf ( n41748 , n41747 );
and ( n41749 , n41740 , n41748 );
not ( n41750 , n41478 );
and ( n41751 , n41750 , n41208 );
xor ( n41752 , n41496 , n41209 );
and ( n41753 , n41752 , n41478 );
or ( n41754 , n41751 , n41753 );
buf ( n41755 , n41754 );
buf ( n41756 , n41755 );
buf ( n41757 , n28890 );
not ( n41758 , n41757 );
buf ( n41759 , n41758 );
not ( n41760 , n41759 );
buf ( n41761 , n41760 );
buf ( n41762 , n41761 );
buf ( n41763 , n41762 );
and ( n41764 , n41756 , n41763 );
and ( n41765 , n41748 , n41764 );
and ( n41766 , n41740 , n41764 );
or ( n41767 , n41749 , n41765 , n41766 );
and ( n41768 , n41732 , n41767 );
and ( n41769 , n41724 , n41767 );
or ( n41770 , n41733 , n41768 , n41769 );
and ( n41771 , n41716 , n41770 );
and ( n41772 , n41708 , n41770 );
or ( n41773 , n41717 , n41771 , n41772 );
and ( n41774 , n41700 , n41773 );
and ( n41775 , n41692 , n41773 );
or ( n41776 , n41701 , n41774 , n41775 );
and ( n41777 , n41684 , n41776 );
and ( n41778 , n41676 , n41776 );
or ( n41779 , n41685 , n41777 , n41778 );
and ( n41780 , n41668 , n41779 );
and ( n41781 , n41660 , n41779 );
or ( n41782 , n41669 , n41780 , n41781 );
and ( n41783 , n41652 , n41782 );
and ( n41784 , n41644 , n41782 );
or ( n41785 , n41653 , n41783 , n41784 );
and ( n41786 , n41636 , n41785 );
and ( n41787 , n41628 , n41785 );
or ( n41788 , n41637 , n41786 , n41787 );
and ( n41789 , n41620 , n41788 );
and ( n41790 , n41612 , n41788 );
or ( n41791 , n41621 , n41789 , n41790 );
and ( n41792 , n41604 , n41791 );
and ( n41793 , n41596 , n41791 );
or ( n41794 , n41605 , n41792 , n41793 );
and ( n41795 , n41588 , n41794 );
and ( n41796 , n41580 , n41794 );
or ( n41797 , n41589 , n41795 , n41796 );
and ( n41798 , n41572 , n41797 );
and ( n41799 , n41564 , n41797 );
or ( n41800 , n41573 , n41798 , n41799 );
and ( n41801 , n41556 , n41800 );
and ( n41802 , n41548 , n41800 );
or ( n41803 , n41557 , n41801 , n41802 );
and ( n41804 , n41540 , n41803 );
and ( n41805 , n41532 , n41803 );
or ( n41806 , n41541 , n41804 , n41805 );
xor ( n41807 , n41525 , n41806 );
buf ( n41808 , n41807 );
and ( n41809 , n41808 , n27046 );
buf ( n41810 , n25857 );
buf ( n41811 , n41810 );
not ( n41812 , n41811 );
buf ( n41813 , n41812 );
buf ( n41814 , n41813 );
not ( n41815 , n41814 );
buf ( n41816 , n25872 );
not ( n41817 , n41816 );
buf ( n41818 , n25890 );
and ( n41819 , n41817 , n41818 );
not ( n41820 , n41818 );
not ( n41821 , n41810 );
xor ( n41822 , n41820 , n41821 );
and ( n41823 , n41822 , n41816 );
or ( n41824 , n41819 , n41823 );
buf ( n41825 , n41824 );
not ( n41826 , n41825 );
buf ( n41827 , n41826 );
buf ( n41828 , n41827 );
not ( n41829 , n41828 );
or ( n41830 , n41815 , n41829 );
not ( n41831 , n41816 );
buf ( n41832 , n25921 );
and ( n41833 , n41831 , n41832 );
not ( n41834 , n41832 );
and ( n41835 , n41820 , n41821 );
xor ( n41836 , n41834 , n41835 );
and ( n41837 , n41836 , n41816 );
or ( n41838 , n41833 , n41837 );
buf ( n41839 , n41838 );
not ( n41840 , n41839 );
buf ( n41841 , n41840 );
buf ( n41842 , n41841 );
not ( n41843 , n41842 );
or ( n41844 , n41830 , n41843 );
not ( n41845 , n41816 );
buf ( n41846 , n25954 );
and ( n41847 , n41845 , n41846 );
not ( n41848 , n41846 );
and ( n41849 , n41834 , n41835 );
xor ( n41850 , n41848 , n41849 );
and ( n41851 , n41850 , n41816 );
or ( n41852 , n41847 , n41851 );
buf ( n41853 , n41852 );
not ( n41854 , n41853 );
buf ( n41855 , n41854 );
buf ( n41856 , n41855 );
not ( n41857 , n41856 );
or ( n41858 , n41844 , n41857 );
not ( n41859 , n41816 );
buf ( n41860 , n25987 );
and ( n41861 , n41859 , n41860 );
not ( n41862 , n41860 );
and ( n41863 , n41848 , n41849 );
xor ( n41864 , n41862 , n41863 );
and ( n41865 , n41864 , n41816 );
or ( n41866 , n41861 , n41865 );
buf ( n41867 , n41866 );
not ( n41868 , n41867 );
buf ( n41869 , n41868 );
buf ( n41870 , n41869 );
not ( n41871 , n41870 );
or ( n41872 , n41858 , n41871 );
not ( n41873 , n41816 );
buf ( n41874 , n26021 );
and ( n41875 , n41873 , n41874 );
not ( n41876 , n41874 );
and ( n41877 , n41862 , n41863 );
xor ( n41878 , n41876 , n41877 );
and ( n41879 , n41878 , n41816 );
or ( n41880 , n41875 , n41879 );
buf ( n41881 , n41880 );
not ( n41882 , n41881 );
buf ( n41883 , n41882 );
buf ( n41884 , n41883 );
not ( n41885 , n41884 );
or ( n41886 , n41872 , n41885 );
not ( n41887 , n41816 );
buf ( n41888 , n26055 );
and ( n41889 , n41887 , n41888 );
not ( n41890 , n41888 );
and ( n41891 , n41876 , n41877 );
xor ( n41892 , n41890 , n41891 );
and ( n41893 , n41892 , n41816 );
or ( n41894 , n41889 , n41893 );
buf ( n41895 , n41894 );
not ( n41896 , n41895 );
buf ( n41897 , n41896 );
buf ( n41898 , n41897 );
not ( n41899 , n41898 );
or ( n41900 , n41886 , n41899 );
not ( n41901 , n41816 );
buf ( n41902 , n26089 );
and ( n41903 , n41901 , n41902 );
not ( n41904 , n41902 );
and ( n41905 , n41890 , n41891 );
xor ( n41906 , n41904 , n41905 );
and ( n41907 , n41906 , n41816 );
or ( n41908 , n41903 , n41907 );
buf ( n41909 , n41908 );
not ( n41910 , n41909 );
buf ( n41911 , n41910 );
buf ( n41912 , n41911 );
not ( n41913 , n41912 );
or ( n41914 , n41900 , n41913 );
not ( n41915 , n41816 );
buf ( n41916 , n26123 );
and ( n41917 , n41915 , n41916 );
not ( n41918 , n41916 );
and ( n41919 , n41904 , n41905 );
xor ( n41920 , n41918 , n41919 );
and ( n41921 , n41920 , n41816 );
or ( n41922 , n41917 , n41921 );
buf ( n41923 , n41922 );
not ( n41924 , n41923 );
buf ( n41925 , n41924 );
buf ( n41926 , n41925 );
not ( n41927 , n41926 );
or ( n41928 , n41914 , n41927 );
not ( n41929 , n41816 );
buf ( n41930 , n26157 );
and ( n41931 , n41929 , n41930 );
not ( n41932 , n41930 );
and ( n41933 , n41918 , n41919 );
xor ( n41934 , n41932 , n41933 );
and ( n41935 , n41934 , n41816 );
or ( n41936 , n41931 , n41935 );
buf ( n41937 , n41936 );
not ( n41938 , n41937 );
buf ( n41939 , n41938 );
buf ( n41940 , n41939 );
not ( n41941 , n41940 );
or ( n41942 , n41928 , n41941 );
not ( n41943 , n41816 );
buf ( n41944 , n26191 );
and ( n41945 , n41943 , n41944 );
not ( n41946 , n41944 );
and ( n41947 , n41932 , n41933 );
xor ( n41948 , n41946 , n41947 );
and ( n41949 , n41948 , n41816 );
or ( n41950 , n41945 , n41949 );
buf ( n41951 , n41950 );
not ( n41952 , n41951 );
buf ( n41953 , n41952 );
buf ( n41954 , n41953 );
not ( n41955 , n41954 );
or ( n41956 , n41942 , n41955 );
not ( n41957 , n41816 );
buf ( n41958 , n26225 );
and ( n41959 , n41957 , n41958 );
not ( n41960 , n41958 );
and ( n41961 , n41946 , n41947 );
xor ( n41962 , n41960 , n41961 );
and ( n41963 , n41962 , n41816 );
or ( n41964 , n41959 , n41963 );
buf ( n41965 , n41964 );
not ( n41966 , n41965 );
buf ( n41967 , n41966 );
buf ( n41968 , n41967 );
not ( n41969 , n41968 );
or ( n41970 , n41956 , n41969 );
not ( n41971 , n41816 );
buf ( n41972 , n26259 );
and ( n41973 , n41971 , n41972 );
not ( n41974 , n41972 );
and ( n41975 , n41960 , n41961 );
xor ( n41976 , n41974 , n41975 );
and ( n41977 , n41976 , n41816 );
or ( n41978 , n41973 , n41977 );
buf ( n41979 , n41978 );
not ( n41980 , n41979 );
buf ( n41981 , n41980 );
buf ( n41982 , n41981 );
not ( n41983 , n41982 );
or ( n41984 , n41970 , n41983 );
not ( n41985 , n41816 );
buf ( n41986 , n26293 );
and ( n41987 , n41985 , n41986 );
not ( n41988 , n41986 );
and ( n41989 , n41974 , n41975 );
xor ( n41990 , n41988 , n41989 );
and ( n41991 , n41990 , n41816 );
or ( n41992 , n41987 , n41991 );
buf ( n41993 , n41992 );
not ( n41994 , n41993 );
buf ( n41995 , n41994 );
buf ( n41996 , n41995 );
not ( n41997 , n41996 );
or ( n41998 , n41984 , n41997 );
not ( n41999 , n41816 );
buf ( n42000 , n26327 );
and ( n42001 , n41999 , n42000 );
not ( n42002 , n42000 );
and ( n42003 , n41988 , n41989 );
xor ( n42004 , n42002 , n42003 );
and ( n42005 , n42004 , n41816 );
or ( n42006 , n42001 , n42005 );
buf ( n42007 , n42006 );
not ( n42008 , n42007 );
buf ( n42009 , n42008 );
buf ( n42010 , n42009 );
not ( n42011 , n42010 );
or ( n42012 , n41998 , n42011 );
not ( n42013 , n41816 );
buf ( n42014 , n26361 );
and ( n42015 , n42013 , n42014 );
not ( n42016 , n42014 );
and ( n42017 , n42002 , n42003 );
xor ( n42018 , n42016 , n42017 );
and ( n42019 , n42018 , n41816 );
or ( n42020 , n42015 , n42019 );
buf ( n42021 , n42020 );
not ( n42022 , n42021 );
buf ( n42023 , n42022 );
buf ( n42024 , n42023 );
not ( n42025 , n42024 );
or ( n42026 , n42012 , n42025 );
not ( n42027 , n41816 );
buf ( n42028 , n26395 );
and ( n42029 , n42027 , n42028 );
not ( n42030 , n42028 );
and ( n42031 , n42016 , n42017 );
xor ( n42032 , n42030 , n42031 );
and ( n42033 , n42032 , n41816 );
or ( n42034 , n42029 , n42033 );
buf ( n42035 , n42034 );
not ( n42036 , n42035 );
buf ( n42037 , n42036 );
buf ( n42038 , n42037 );
not ( n42039 , n42038 );
or ( n42040 , n42026 , n42039 );
not ( n42041 , n41816 );
buf ( n42042 , n26429 );
and ( n42043 , n42041 , n42042 );
not ( n42044 , n42042 );
and ( n42045 , n42030 , n42031 );
xor ( n42046 , n42044 , n42045 );
and ( n42047 , n42046 , n41816 );
or ( n42048 , n42043 , n42047 );
buf ( n42049 , n42048 );
not ( n42050 , n42049 );
buf ( n42051 , n42050 );
buf ( n42052 , n42051 );
not ( n42053 , n42052 );
or ( n42054 , n42040 , n42053 );
not ( n42055 , n41816 );
buf ( n42056 , n26463 );
and ( n42057 , n42055 , n42056 );
not ( n42058 , n42056 );
and ( n42059 , n42044 , n42045 );
xor ( n42060 , n42058 , n42059 );
and ( n42061 , n42060 , n41816 );
or ( n42062 , n42057 , n42061 );
buf ( n42063 , n42062 );
not ( n42064 , n42063 );
buf ( n42065 , n42064 );
buf ( n42066 , n42065 );
not ( n42067 , n42066 );
or ( n42068 , n42054 , n42067 );
not ( n42069 , n41816 );
buf ( n42070 , n26497 );
and ( n42071 , n42069 , n42070 );
not ( n42072 , n42070 );
and ( n42073 , n42058 , n42059 );
xor ( n42074 , n42072 , n42073 );
and ( n42075 , n42074 , n41816 );
or ( n42076 , n42071 , n42075 );
buf ( n42077 , n42076 );
not ( n42078 , n42077 );
buf ( n42079 , n42078 );
buf ( n42080 , n42079 );
not ( n42081 , n42080 );
or ( n42082 , n42068 , n42081 );
buf ( n42083 , n42082 );
buf ( n42084 , n42083 );
and ( n42085 , n42084 , n41816 );
not ( n42086 , n42085 );
and ( n42087 , n42086 , n42025 );
xor ( n42088 , n42025 , n41816 );
xor ( n42089 , n42011 , n41816 );
xor ( n42090 , n41997 , n41816 );
xor ( n42091 , n41983 , n41816 );
xor ( n42092 , n41969 , n41816 );
xor ( n42093 , n41955 , n41816 );
xor ( n42094 , n41941 , n41816 );
xor ( n42095 , n41927 , n41816 );
xor ( n42096 , n41913 , n41816 );
xor ( n42097 , n41899 , n41816 );
xor ( n42098 , n41885 , n41816 );
xor ( n42099 , n41871 , n41816 );
xor ( n42100 , n41857 , n41816 );
xor ( n42101 , n41843 , n41816 );
xor ( n42102 , n41829 , n41816 );
xor ( n42103 , n41815 , n41816 );
and ( n42104 , n42103 , n41816 );
and ( n42105 , n42102 , n42104 );
and ( n42106 , n42101 , n42105 );
and ( n42107 , n42100 , n42106 );
and ( n42108 , n42099 , n42107 );
and ( n42109 , n42098 , n42108 );
and ( n42110 , n42097 , n42109 );
and ( n42111 , n42096 , n42110 );
and ( n42112 , n42095 , n42111 );
and ( n42113 , n42094 , n42112 );
and ( n42114 , n42093 , n42113 );
and ( n42115 , n42092 , n42114 );
and ( n42116 , n42091 , n42115 );
and ( n42117 , n42090 , n42116 );
and ( n42118 , n42089 , n42117 );
xor ( n42119 , n42088 , n42118 );
and ( n42120 , n42119 , n42085 );
or ( n42121 , n42087 , n42120 );
buf ( n42122 , n42121 );
buf ( n42123 , n42122 );
buf ( n42124 , n41523 );
xor ( n42125 , n42123 , n42124 );
not ( n42126 , n42085 );
and ( n42127 , n42126 , n42011 );
xor ( n42128 , n42089 , n42117 );
and ( n42129 , n42128 , n42085 );
or ( n42130 , n42127 , n42129 );
buf ( n42131 , n42130 );
buf ( n42132 , n42131 );
buf ( n42133 , n41539 );
and ( n42134 , n42132 , n42133 );
not ( n42135 , n42085 );
and ( n42136 , n42135 , n41997 );
xor ( n42137 , n42090 , n42116 );
and ( n42138 , n42137 , n42085 );
or ( n42139 , n42136 , n42138 );
buf ( n42140 , n42139 );
buf ( n42141 , n42140 );
buf ( n42142 , n41555 );
and ( n42143 , n42141 , n42142 );
not ( n42144 , n42085 );
and ( n42145 , n42144 , n41983 );
xor ( n42146 , n42091 , n42115 );
and ( n42147 , n42146 , n42085 );
or ( n42148 , n42145 , n42147 );
buf ( n42149 , n42148 );
buf ( n42150 , n42149 );
buf ( n42151 , n41571 );
and ( n42152 , n42150 , n42151 );
not ( n42153 , n42085 );
and ( n42154 , n42153 , n41969 );
xor ( n42155 , n42092 , n42114 );
and ( n42156 , n42155 , n42085 );
or ( n42157 , n42154 , n42156 );
buf ( n42158 , n42157 );
buf ( n42159 , n42158 );
buf ( n42160 , n41587 );
and ( n42161 , n42159 , n42160 );
not ( n42162 , n42085 );
and ( n42163 , n42162 , n41955 );
xor ( n42164 , n42093 , n42113 );
and ( n42165 , n42164 , n42085 );
or ( n42166 , n42163 , n42165 );
buf ( n42167 , n42166 );
buf ( n42168 , n42167 );
buf ( n42169 , n41603 );
and ( n42170 , n42168 , n42169 );
not ( n42171 , n42085 );
and ( n42172 , n42171 , n41941 );
xor ( n42173 , n42094 , n42112 );
and ( n42174 , n42173 , n42085 );
or ( n42175 , n42172 , n42174 );
buf ( n42176 , n42175 );
buf ( n42177 , n42176 );
buf ( n42178 , n41619 );
and ( n42179 , n42177 , n42178 );
not ( n42180 , n42085 );
and ( n42181 , n42180 , n41927 );
xor ( n42182 , n42095 , n42111 );
and ( n42183 , n42182 , n42085 );
or ( n42184 , n42181 , n42183 );
buf ( n42185 , n42184 );
buf ( n42186 , n42185 );
buf ( n42187 , n41635 );
and ( n42188 , n42186 , n42187 );
not ( n42189 , n42085 );
and ( n42190 , n42189 , n41913 );
xor ( n42191 , n42096 , n42110 );
and ( n42192 , n42191 , n42085 );
or ( n42193 , n42190 , n42192 );
buf ( n42194 , n42193 );
buf ( n42195 , n42194 );
buf ( n42196 , n41651 );
and ( n42197 , n42195 , n42196 );
not ( n42198 , n42085 );
and ( n42199 , n42198 , n41899 );
xor ( n42200 , n42097 , n42109 );
and ( n42201 , n42200 , n42085 );
or ( n42202 , n42199 , n42201 );
buf ( n42203 , n42202 );
buf ( n42204 , n42203 );
buf ( n42205 , n41667 );
and ( n42206 , n42204 , n42205 );
not ( n42207 , n42085 );
and ( n42208 , n42207 , n41885 );
xor ( n42209 , n42098 , n42108 );
and ( n42210 , n42209 , n42085 );
or ( n42211 , n42208 , n42210 );
buf ( n42212 , n42211 );
buf ( n42213 , n42212 );
buf ( n42214 , n41683 );
and ( n42215 , n42213 , n42214 );
not ( n42216 , n42085 );
and ( n42217 , n42216 , n41871 );
xor ( n42218 , n42099 , n42107 );
and ( n42219 , n42218 , n42085 );
or ( n42220 , n42217 , n42219 );
buf ( n42221 , n42220 );
buf ( n42222 , n42221 );
buf ( n42223 , n41699 );
and ( n42224 , n42222 , n42223 );
not ( n42225 , n42085 );
and ( n42226 , n42225 , n41857 );
xor ( n42227 , n42100 , n42106 );
and ( n42228 , n42227 , n42085 );
or ( n42229 , n42226 , n42228 );
buf ( n42230 , n42229 );
buf ( n42231 , n42230 );
buf ( n42232 , n41715 );
and ( n42233 , n42231 , n42232 );
not ( n42234 , n42085 );
and ( n42235 , n42234 , n41843 );
xor ( n42236 , n42101 , n42105 );
and ( n42237 , n42236 , n42085 );
or ( n42238 , n42235 , n42237 );
buf ( n42239 , n42238 );
buf ( n42240 , n42239 );
buf ( n42241 , n41731 );
and ( n42242 , n42240 , n42241 );
not ( n42243 , n42085 );
and ( n42244 , n42243 , n41829 );
xor ( n42245 , n42102 , n42104 );
and ( n42246 , n42245 , n42085 );
or ( n42247 , n42244 , n42246 );
buf ( n42248 , n42247 );
buf ( n42249 , n42248 );
buf ( n42250 , n41747 );
and ( n42251 , n42249 , n42250 );
not ( n42252 , n42085 );
and ( n42253 , n42252 , n41815 );
xor ( n42254 , n42103 , n41816 );
and ( n42255 , n42254 , n42085 );
or ( n42256 , n42253 , n42255 );
buf ( n42257 , n42256 );
buf ( n42258 , n42257 );
buf ( n42259 , n41762 );
and ( n42260 , n42258 , n42259 );
and ( n42261 , n42250 , n42260 );
and ( n42262 , n42249 , n42260 );
or ( n42263 , n42251 , n42261 , n42262 );
and ( n42264 , n42241 , n42263 );
and ( n42265 , n42240 , n42263 );
or ( n42266 , n42242 , n42264 , n42265 );
and ( n42267 , n42232 , n42266 );
and ( n42268 , n42231 , n42266 );
or ( n42269 , n42233 , n42267 , n42268 );
and ( n42270 , n42223 , n42269 );
and ( n42271 , n42222 , n42269 );
or ( n42272 , n42224 , n42270 , n42271 );
and ( n42273 , n42214 , n42272 );
and ( n42274 , n42213 , n42272 );
or ( n42275 , n42215 , n42273 , n42274 );
and ( n42276 , n42205 , n42275 );
and ( n42277 , n42204 , n42275 );
or ( n42278 , n42206 , n42276 , n42277 );
and ( n42279 , n42196 , n42278 );
and ( n42280 , n42195 , n42278 );
or ( n42281 , n42197 , n42279 , n42280 );
and ( n42282 , n42187 , n42281 );
and ( n42283 , n42186 , n42281 );
or ( n42284 , n42188 , n42282 , n42283 );
and ( n42285 , n42178 , n42284 );
and ( n42286 , n42177 , n42284 );
or ( n42287 , n42179 , n42285 , n42286 );
and ( n42288 , n42169 , n42287 );
and ( n42289 , n42168 , n42287 );
or ( n42290 , n42170 , n42288 , n42289 );
and ( n42291 , n42160 , n42290 );
and ( n42292 , n42159 , n42290 );
or ( n42293 , n42161 , n42291 , n42292 );
and ( n42294 , n42151 , n42293 );
and ( n42295 , n42150 , n42293 );
or ( n42296 , n42152 , n42294 , n42295 );
and ( n42297 , n42142 , n42296 );
and ( n42298 , n42141 , n42296 );
or ( n42299 , n42143 , n42297 , n42298 );
and ( n42300 , n42133 , n42299 );
and ( n42301 , n42132 , n42299 );
or ( n42302 , n42134 , n42300 , n42301 );
xor ( n42303 , n42125 , n42302 );
buf ( n42304 , n42303 );
and ( n42305 , n42304 , n27049 );
or ( n42306 , n28508 , n28506 );
and ( n42307 , n29373 , n42306 );
or ( n42308 , n41809 , n42305 , n42307 );
buf ( n42309 , n42308 );
and ( n42310 , C1 , n42309 );
or ( n42311 , n42310 , C0 );
buf ( n42312 , n42311 );
not ( n42313 , n42312 );
buf ( n42314 , n42313 );
buf ( n42315 , n42314 );
not ( n42316 , n42315 );
and ( n42317 , C1 , n42316 );
or ( n42318 , n42317 , C0 );
buf ( n42319 , n42318 );
and ( n42320 , n42319 , n24799 );
or ( n42321 , n41202 , n42320 );
and ( n42322 , n40152 , n42321 );
and ( n42323 , n41188 , n24511 );
or ( n42324 , n42322 , n42323 );
and ( n42325 , n42324 , n31008 );
buf ( n42326 , n25224 );
buf ( n42327 , n42326 );
not ( n42328 , n42327 );
buf ( n42329 , n42328 );
buf ( n42330 , n42329 );
not ( n42331 , n42330 );
buf ( n42332 , n25231 );
not ( n42333 , n42332 );
buf ( n42334 , n25234 );
and ( n42335 , n42333 , n42334 );
not ( n42336 , n42334 );
not ( n42337 , n42326 );
xor ( n42338 , n42336 , n42337 );
and ( n42339 , n42338 , n42332 );
or ( n42340 , n42335 , n42339 );
buf ( n42341 , n42340 );
not ( n42342 , n42341 );
buf ( n42343 , n42342 );
buf ( n42344 , n42343 );
not ( n42345 , n42344 );
or ( n42346 , n42331 , n42345 );
not ( n42347 , n42332 );
buf ( n42348 , n25249 );
and ( n42349 , n42347 , n42348 );
not ( n42350 , n42348 );
and ( n42351 , n42336 , n42337 );
xor ( n42352 , n42350 , n42351 );
and ( n42353 , n42352 , n42332 );
or ( n42354 , n42349 , n42353 );
buf ( n42355 , n42354 );
not ( n42356 , n42355 );
buf ( n42357 , n42356 );
buf ( n42358 , n42357 );
not ( n42359 , n42358 );
or ( n42360 , n42346 , n42359 );
not ( n42361 , n42332 );
buf ( n42362 , n25264 );
and ( n42363 , n42361 , n42362 );
not ( n42364 , n42362 );
and ( n42365 , n42350 , n42351 );
xor ( n42366 , n42364 , n42365 );
and ( n42367 , n42366 , n42332 );
or ( n42368 , n42363 , n42367 );
buf ( n42369 , n42368 );
not ( n42370 , n42369 );
buf ( n42371 , n42370 );
buf ( n42372 , n42371 );
not ( n42373 , n42372 );
or ( n42374 , n42360 , n42373 );
not ( n42375 , n42332 );
buf ( n42376 , n25279 );
and ( n42377 , n42375 , n42376 );
not ( n42378 , n42376 );
and ( n42379 , n42364 , n42365 );
xor ( n42380 , n42378 , n42379 );
and ( n42381 , n42380 , n42332 );
or ( n42382 , n42377 , n42381 );
buf ( n42383 , n42382 );
not ( n42384 , n42383 );
buf ( n42385 , n42384 );
buf ( n42386 , n42385 );
not ( n42387 , n42386 );
or ( n42388 , n42374 , n42387 );
not ( n42389 , n42332 );
buf ( n42390 , n25294 );
and ( n42391 , n42389 , n42390 );
not ( n42392 , n42390 );
and ( n42393 , n42378 , n42379 );
xor ( n42394 , n42392 , n42393 );
and ( n42395 , n42394 , n42332 );
or ( n42396 , n42391 , n42395 );
buf ( n42397 , n42396 );
not ( n42398 , n42397 );
buf ( n42399 , n42398 );
buf ( n42400 , n42399 );
not ( n42401 , n42400 );
or ( n42402 , n42388 , n42401 );
not ( n42403 , n42332 );
buf ( n42404 , n25309 );
and ( n42405 , n42403 , n42404 );
not ( n42406 , n42404 );
and ( n42407 , n42392 , n42393 );
xor ( n42408 , n42406 , n42407 );
and ( n42409 , n42408 , n42332 );
or ( n42410 , n42405 , n42409 );
buf ( n42411 , n42410 );
not ( n42412 , n42411 );
buf ( n42413 , n42412 );
buf ( n42414 , n42413 );
not ( n42415 , n42414 );
or ( n42416 , n42402 , n42415 );
not ( n42417 , n42332 );
buf ( n42418 , n25324 );
and ( n42419 , n42417 , n42418 );
not ( n42420 , n42418 );
and ( n42421 , n42406 , n42407 );
xor ( n42422 , n42420 , n42421 );
and ( n42423 , n42422 , n42332 );
or ( n42424 , n42419 , n42423 );
buf ( n42425 , n42424 );
not ( n42426 , n42425 );
buf ( n42427 , n42426 );
buf ( n42428 , n42427 );
not ( n42429 , n42428 );
or ( n42430 , n42416 , n42429 );
not ( n42431 , n42332 );
buf ( n42432 , n25339 );
and ( n42433 , n42431 , n42432 );
not ( n42434 , n42432 );
and ( n42435 , n42420 , n42421 );
xor ( n42436 , n42434 , n42435 );
and ( n42437 , n42436 , n42332 );
or ( n42438 , n42433 , n42437 );
buf ( n42439 , n42438 );
not ( n42440 , n42439 );
buf ( n42441 , n42440 );
buf ( n42442 , n42441 );
not ( n42443 , n42442 );
or ( n42444 , n42430 , n42443 );
not ( n42445 , n42332 );
buf ( n42446 , n25354 );
and ( n42447 , n42445 , n42446 );
not ( n42448 , n42446 );
and ( n42449 , n42434 , n42435 );
xor ( n42450 , n42448 , n42449 );
and ( n42451 , n42450 , n42332 );
or ( n42452 , n42447 , n42451 );
buf ( n42453 , n42452 );
not ( n42454 , n42453 );
buf ( n42455 , n42454 );
buf ( n42456 , n42455 );
not ( n42457 , n42456 );
or ( n42458 , n42444 , n42457 );
not ( n42459 , n42332 );
buf ( n42460 , n25369 );
and ( n42461 , n42459 , n42460 );
not ( n42462 , n42460 );
and ( n42463 , n42448 , n42449 );
xor ( n42464 , n42462 , n42463 );
and ( n42465 , n42464 , n42332 );
or ( n42466 , n42461 , n42465 );
buf ( n42467 , n42466 );
not ( n42468 , n42467 );
buf ( n42469 , n42468 );
buf ( n42470 , n42469 );
not ( n42471 , n42470 );
or ( n42472 , n42458 , n42471 );
not ( n42473 , n42332 );
buf ( n42474 , n25384 );
and ( n42475 , n42473 , n42474 );
not ( n42476 , n42474 );
and ( n42477 , n42462 , n42463 );
xor ( n42478 , n42476 , n42477 );
and ( n42479 , n42478 , n42332 );
or ( n42480 , n42475 , n42479 );
buf ( n42481 , n42480 );
not ( n42482 , n42481 );
buf ( n42483 , n42482 );
buf ( n42484 , n42483 );
not ( n42485 , n42484 );
or ( n42486 , n42472 , n42485 );
not ( n42487 , n42332 );
buf ( n42488 , n25399 );
and ( n42489 , n42487 , n42488 );
not ( n42490 , n42488 );
and ( n42491 , n42476 , n42477 );
xor ( n42492 , n42490 , n42491 );
and ( n42493 , n42492 , n42332 );
or ( n42494 , n42489 , n42493 );
buf ( n42495 , n42494 );
not ( n42496 , n42495 );
buf ( n42497 , n42496 );
buf ( n42498 , n42497 );
not ( n42499 , n42498 );
or ( n42500 , n42486 , n42499 );
not ( n42501 , n42332 );
buf ( n42502 , n25414 );
and ( n42503 , n42501 , n42502 );
not ( n42504 , n42502 );
and ( n42505 , n42490 , n42491 );
xor ( n42506 , n42504 , n42505 );
and ( n42507 , n42506 , n42332 );
or ( n42508 , n42503 , n42507 );
buf ( n42509 , n42508 );
not ( n42510 , n42509 );
buf ( n42511 , n42510 );
buf ( n42512 , n42511 );
not ( n42513 , n42512 );
or ( n42514 , n42500 , n42513 );
not ( n42515 , n42332 );
buf ( n42516 , n25429 );
and ( n42517 , n42515 , n42516 );
not ( n42518 , n42516 );
and ( n42519 , n42504 , n42505 );
xor ( n42520 , n42518 , n42519 );
and ( n42521 , n42520 , n42332 );
or ( n42522 , n42517 , n42521 );
buf ( n42523 , n42522 );
not ( n42524 , n42523 );
buf ( n42525 , n42524 );
buf ( n42526 , n42525 );
not ( n42527 , n42526 );
or ( n42528 , n42514 , n42527 );
not ( n42529 , n42332 );
buf ( n42530 , n25444 );
and ( n42531 , n42529 , n42530 );
not ( n42532 , n42530 );
and ( n42533 , n42518 , n42519 );
xor ( n42534 , n42532 , n42533 );
and ( n42535 , n42534 , n42332 );
or ( n42536 , n42531 , n42535 );
buf ( n42537 , n42536 );
not ( n42538 , n42537 );
buf ( n42539 , n42538 );
buf ( n42540 , n42539 );
not ( n42541 , n42540 );
or ( n42542 , n42528 , n42541 );
not ( n42543 , n42332 );
buf ( n42544 , n25459 );
and ( n42545 , n42543 , n42544 );
not ( n42546 , n42544 );
and ( n42547 , n42532 , n42533 );
xor ( n42548 , n42546 , n42547 );
and ( n42549 , n42548 , n42332 );
or ( n42550 , n42545 , n42549 );
buf ( n42551 , n42550 );
not ( n42552 , n42551 );
buf ( n42553 , n42552 );
buf ( n42554 , n42553 );
not ( n42555 , n42554 );
or ( n42556 , n42542 , n42555 );
not ( n42557 , n42332 );
buf ( n42558 , n25474 );
and ( n42559 , n42557 , n42558 );
not ( n42560 , n42558 );
and ( n42561 , n42546 , n42547 );
xor ( n42562 , n42560 , n42561 );
and ( n42563 , n42562 , n42332 );
or ( n42564 , n42559 , n42563 );
buf ( n42565 , n42564 );
not ( n42566 , n42565 );
buf ( n42567 , n42566 );
buf ( n42568 , n42567 );
not ( n42569 , n42568 );
or ( n42570 , n42556 , n42569 );
not ( n42571 , n42332 );
buf ( n42572 , n25489 );
and ( n42573 , n42571 , n42572 );
not ( n42574 , n42572 );
and ( n42575 , n42560 , n42561 );
xor ( n42576 , n42574 , n42575 );
and ( n42577 , n42576 , n42332 );
or ( n42578 , n42573 , n42577 );
buf ( n42579 , n42578 );
not ( n42580 , n42579 );
buf ( n42581 , n42580 );
buf ( n42582 , n42581 );
not ( n42583 , n42582 );
or ( n42584 , n42570 , n42583 );
not ( n42585 , n42332 );
buf ( n42586 , n25504 );
and ( n42587 , n42585 , n42586 );
not ( n42588 , n42586 );
and ( n42589 , n42574 , n42575 );
xor ( n42590 , n42588 , n42589 );
and ( n42591 , n42590 , n42332 );
or ( n42592 , n42587 , n42591 );
buf ( n42593 , n42592 );
not ( n42594 , n42593 );
buf ( n42595 , n42594 );
buf ( n42596 , n42595 );
not ( n42597 , n42596 );
or ( n42598 , n42584 , n42597 );
buf ( n42599 , n42598 );
buf ( n42600 , n42599 );
and ( n42601 , n42600 , n42332 );
not ( n42602 , n42601 );
and ( n42603 , n42602 , n42541 );
xor ( n42604 , n42541 , n42332 );
xor ( n42605 , n42527 , n42332 );
xor ( n42606 , n42513 , n42332 );
xor ( n42607 , n42499 , n42332 );
xor ( n42608 , n42485 , n42332 );
xor ( n42609 , n42471 , n42332 );
xor ( n42610 , n42457 , n42332 );
xor ( n42611 , n42443 , n42332 );
xor ( n42612 , n42429 , n42332 );
xor ( n42613 , n42415 , n42332 );
xor ( n42614 , n42401 , n42332 );
xor ( n42615 , n42387 , n42332 );
xor ( n42616 , n42373 , n42332 );
xor ( n42617 , n42359 , n42332 );
xor ( n42618 , n42345 , n42332 );
xor ( n42619 , n42331 , n42332 );
and ( n42620 , n42619 , n42332 );
and ( n42621 , n42618 , n42620 );
and ( n42622 , n42617 , n42621 );
and ( n42623 , n42616 , n42622 );
and ( n42624 , n42615 , n42623 );
and ( n42625 , n42614 , n42624 );
and ( n42626 , n42613 , n42625 );
and ( n42627 , n42612 , n42626 );
and ( n42628 , n42611 , n42627 );
and ( n42629 , n42610 , n42628 );
and ( n42630 , n42609 , n42629 );
and ( n42631 , n42608 , n42630 );
and ( n42632 , n42607 , n42631 );
and ( n42633 , n42606 , n42632 );
and ( n42634 , n42605 , n42633 );
xor ( n42635 , n42604 , n42634 );
and ( n42636 , n42635 , n42601 );
or ( n42637 , n42603 , n42636 );
buf ( n42638 , n42637 );
and ( n42639 , n42638 , n10618 );
or ( n42640 , n42325 , n42639 );
buf ( n42641 , n42640 );
buf ( n42642 , n42641 );
buf ( n42643 , n10613 );
buf ( n42644 , n10613 );
buf ( n42645 , n10615 );
not ( n42646 , n17451 );
and ( n42647 , n18540 , n17873 );
and ( n42648 , n34754 , n21330 );
and ( n42649 , n18540 , n21338 );
or ( n42650 , n42648 , n42649 );
and ( n42651 , n42650 , n21341 );
and ( n42652 , n34767 , n21330 );
and ( n42653 , n18540 , n21338 );
or ( n42654 , n42652 , n42653 );
and ( n42655 , n42654 , n23064 );
and ( n42656 , n34777 , n21330 );
and ( n42657 , n18540 , n21338 );
or ( n42658 , n42656 , n42657 );
and ( n42659 , n42658 , n23825 );
and ( n42660 , n22402 , n21330 );
and ( n42661 , n18540 , n21338 );
or ( n42662 , n42660 , n42661 );
and ( n42663 , n42662 , n23832 );
and ( n42664 , n18538 , n23834 );
and ( n42665 , n34787 , n21330 );
and ( n42666 , n18540 , n21338 );
or ( n42667 , n42665 , n42666 );
and ( n42668 , n42667 , n23917 );
or ( n42669 , n42647 , n42651 , n42655 , n42659 , n42663 , n42664 , n42668 );
and ( n42670 , n42646 , n42669 );
and ( n42671 , n18540 , n17451 );
or ( n42672 , n42670 , n42671 );
and ( n42673 , n42672 , n23924 );
and ( n42674 , n18540 , n23926 );
or ( n42675 , n42673 , n42674 );
buf ( n42676 , n42675 );
buf ( n42677 , n42676 );
not ( n42678 , n17451 );
and ( n42679 , n19213 , n17873 );
and ( n42680 , n34421 , n21336 );
or ( n42681 , n21335 , n21330 );
or ( n42682 , n42681 , C0 );
and ( n42683 , n19213 , n42682 );
or ( n42684 , n42680 , n42683 );
and ( n42685 , n42684 , n21341 );
and ( n42686 , n34431 , n21336 );
and ( n42687 , n19213 , n42682 );
or ( n42688 , n42686 , n42687 );
and ( n42689 , n42688 , n23064 );
and ( n42690 , n34441 , n21336 );
and ( n42691 , n19213 , n42682 );
or ( n42692 , n42690 , n42691 );
and ( n42693 , n42692 , n23825 );
and ( n42694 , n21971 , n21336 );
and ( n42695 , n19213 , n42682 );
or ( n42696 , n42694 , n42695 );
and ( n42697 , n42696 , n23832 );
and ( n42698 , n21971 , n23834 );
and ( n42699 , n34452 , n21336 );
and ( n42700 , n19213 , n42682 );
or ( n42701 , n42699 , n42700 );
and ( n42702 , n42701 , n23917 );
or ( n42703 , n42679 , n42685 , n42689 , n42693 , n42697 , n42698 , n42702 );
and ( n42704 , n42678 , n42703 );
and ( n42705 , n19213 , n17451 );
or ( n42706 , n42704 , n42705 );
and ( n42707 , n42706 , n23924 );
and ( n42708 , n18185 , n23926 );
or ( n42709 , n42707 , n42708 );
buf ( n42710 , n42709 );
buf ( n42711 , n42710 );
and ( n42712 , n11641 , n16574 );
and ( n42713 , n15704 , n16576 );
or ( n42714 , n42712 , n42713 );
buf ( n42715 , n42714 );
buf ( n42716 , n42715 );
buf ( n42717 , n10615 );
buf ( n42718 , n10615 );
buf ( n42719 , n10615 );
and ( n42720 , n11593 , n16574 );
and ( n42721 , n15572 , n16576 );
or ( n42722 , n42720 , n42721 );
buf ( n42723 , n42722 );
buf ( n42724 , n42723 );
not ( n42725 , n17451 );
not ( n42726 , n19474 );
and ( n42727 , n42726 , n18927 );
xor ( n42728 , n19489 , n19513 );
and ( n42729 , n42728 , n19474 );
or ( n42730 , n42727 , n42729 );
buf ( n42731 , n42730 );
and ( n42732 , n42731 , n19745 );
and ( n42733 , n42731 , n19748 );
not ( n42734 , n19750 );
and ( n42735 , n42734 , n20855 );
not ( n42736 , n21193 );
and ( n42737 , n42736 , n20867 );
xor ( n42738 , n21208 , n21234 );
and ( n42739 , n42738 , n21193 );
or ( n42740 , n42737 , n42739 );
buf ( n42741 , n42740 );
and ( n42742 , n42741 , n19750 );
or ( n42743 , n42735 , n42742 );
and ( n42744 , n42743 , n21253 );
and ( n42745 , n20855 , n21255 );
or ( n42746 , n42732 , n42733 , n42744 , n42745 );
and ( n42747 , n42746 , n21334 );
and ( n42748 , n18947 , n34492 );
or ( n42749 , n42747 , n42748 );
and ( n42750 , n42749 , n21341 );
not ( n42751 , n22996 );
and ( n42752 , n42751 , n22720 );
xor ( n42753 , n23011 , n23037 );
and ( n42754 , n42753 , n22996 );
or ( n42755 , n42752 , n42754 );
buf ( n42756 , n42755 );
and ( n42757 , n42756 , n21334 );
and ( n42758 , n18947 , n34492 );
or ( n42759 , n42757 , n42758 );
and ( n42760 , n42759 , n23064 );
not ( n42761 , n23758 );
and ( n42762 , n42761 , n23482 );
xor ( n42763 , n23773 , n23799 );
and ( n42764 , n42763 , n23758 );
or ( n42765 , n42762 , n42764 );
buf ( n42766 , n42765 );
and ( n42767 , n42766 , n21334 );
and ( n42768 , n18947 , n34492 );
or ( n42769 , n42767 , n42768 );
and ( n42770 , n42769 , n23825 );
and ( n42771 , n22162 , n21334 );
and ( n42772 , n18947 , n34492 );
or ( n42773 , n42771 , n42772 );
and ( n42774 , n42773 , n23832 );
xor ( n42775 , n23861 , n23899 );
buf ( n42776 , n42775 );
and ( n42777 , n42776 , n21334 );
and ( n42778 , n18947 , n34492 );
or ( n42779 , n42777 , n42778 );
and ( n42780 , n42779 , n23917 );
and ( n42781 , n18947 , n34526 );
or ( n42782 , n42750 , n42760 , n42770 , n42774 , n42780 , n42781 );
and ( n42783 , n42725 , n42782 );
and ( n42784 , n18947 , n17451 );
or ( n42785 , n42783 , n42784 );
and ( n42786 , n42785 , n23924 );
and ( n42787 , n18947 , n23926 );
or ( n42788 , n42786 , n42787 );
buf ( n42789 , n42788 );
buf ( n42790 , n42789 );
buf ( n42791 , n10613 );
not ( n42792 , n17451 );
and ( n42793 , n40011 , n21334 );
and ( n42794 , n18709 , n34492 );
or ( n42795 , n42793 , n42794 );
and ( n42796 , n42795 , n21341 );
and ( n42797 , n40021 , n21334 );
and ( n42798 , n18709 , n34492 );
or ( n42799 , n42797 , n42798 );
and ( n42800 , n42799 , n23064 );
and ( n42801 , n40031 , n21334 );
and ( n42802 , n18709 , n34492 );
or ( n42803 , n42801 , n42802 );
and ( n42804 , n42803 , n23825 );
and ( n42805 , n22302 , n21334 );
and ( n42806 , n18709 , n34492 );
or ( n42807 , n42805 , n42806 );
and ( n42808 , n42807 , n23832 );
and ( n42809 , n40041 , n21334 );
and ( n42810 , n18709 , n34492 );
or ( n42811 , n42809 , n42810 );
and ( n42812 , n42811 , n23917 );
and ( n42813 , n18709 , n34526 );
or ( n42814 , n42796 , n42800 , n42804 , n42808 , n42812 , n42813 );
and ( n42815 , n42792 , n42814 );
and ( n42816 , n18709 , n17451 );
or ( n42817 , n42815 , n42816 );
and ( n42818 , n42817 , n23924 );
and ( n42819 , n18709 , n23926 );
or ( n42820 , n42818 , n42819 );
buf ( n42821 , n42820 );
buf ( n42822 , n42821 );
not ( n42823 , n24800 );
not ( n42824 , n26823 );
and ( n42825 , n42824 , n26581 );
xor ( n42826 , n26581 , n25877 );
xor ( n42827 , n26547 , n25877 );
xor ( n42828 , n26513 , n25877 );
xor ( n42829 , n26479 , n25877 );
xor ( n42830 , n26445 , n25877 );
and ( n42831 , n39632 , n39637 );
and ( n42832 , n42830 , n42831 );
and ( n42833 , n42829 , n42832 );
and ( n42834 , n42828 , n42833 );
and ( n42835 , n42827 , n42834 );
xor ( n42836 , n42826 , n42835 );
and ( n42837 , n42836 , n26823 );
or ( n42838 , n42825 , n42837 );
buf ( n42839 , n42838 );
and ( n42840 , n42839 , n27046 );
and ( n42841 , n42839 , n27049 );
not ( n42842 , n27051 );
and ( n42843 , n42842 , n28346 );
not ( n42844 , n28494 );
and ( n42845 , n42844 , n28358 );
xor ( n42846 , n28358 , n27883 );
xor ( n42847 , n28336 , n27883 );
xor ( n42848 , n28314 , n27883 );
xor ( n42849 , n28292 , n27883 );
xor ( n42850 , n28270 , n27883 );
and ( n42851 , n39648 , n39653 );
and ( n42852 , n42850 , n42851 );
and ( n42853 , n42849 , n42852 );
and ( n42854 , n42848 , n42853 );
and ( n42855 , n42847 , n42854 );
xor ( n42856 , n42846 , n42855 );
and ( n42857 , n42856 , n28494 );
or ( n42858 , n42845 , n42857 );
buf ( n42859 , n42858 );
and ( n42860 , n42859 , n27051 );
or ( n42861 , n42843 , n42860 );
and ( n42862 , n42861 , n28506 );
and ( n42863 , n28346 , n28508 );
or ( n42864 , n42840 , n42841 , n42862 , n42863 );
and ( n42865 , n42864 , n28586 );
and ( n42866 , n26599 , n34573 );
or ( n42867 , n42865 , n42866 );
and ( n42868 , n42867 , n28594 );
not ( n42869 , n30249 );
and ( n42870 , n42869 , n30126 );
xor ( n42871 , n30126 , n29753 );
xor ( n42872 , n30109 , n29753 );
xor ( n42873 , n30092 , n29753 );
xor ( n42874 , n30075 , n29753 );
xor ( n42875 , n30058 , n29753 );
and ( n42876 , n39669 , n39674 );
and ( n42877 , n42875 , n42876 );
and ( n42878 , n42874 , n42877 );
and ( n42879 , n42873 , n42878 );
and ( n42880 , n42872 , n42879 );
xor ( n42881 , n42871 , n42880 );
and ( n42882 , n42881 , n30249 );
or ( n42883 , n42870 , n42882 );
buf ( n42884 , n42883 );
and ( n42885 , n42884 , n28586 );
and ( n42886 , n26599 , n34573 );
or ( n42887 , n42885 , n42886 );
and ( n42888 , n42887 , n30269 );
not ( n42889 , n30963 );
and ( n42890 , n42889 , n30840 );
xor ( n42891 , n30840 , n30467 );
xor ( n42892 , n30823 , n30467 );
xor ( n42893 , n30806 , n30467 );
xor ( n42894 , n30789 , n30467 );
xor ( n42895 , n30772 , n30467 );
and ( n42896 , n39685 , n39690 );
and ( n42897 , n42895 , n42896 );
and ( n42898 , n42894 , n42897 );
and ( n42899 , n42893 , n42898 );
and ( n42900 , n42892 , n42899 );
xor ( n42901 , n42891 , n42900 );
and ( n42902 , n42901 , n30963 );
or ( n42903 , n42890 , n42902 );
buf ( n42904 , n42903 );
and ( n42905 , n42904 , n28586 );
and ( n42906 , n26599 , n34573 );
or ( n42907 , n42905 , n42906 );
and ( n42908 , n42907 , n30982 );
and ( n42909 , n29211 , n28586 );
and ( n42910 , n26599 , n34573 );
or ( n42911 , n42909 , n42910 );
and ( n42912 , n42911 , n30989 );
buf ( n42913 , n29211 );
not ( n42914 , n42913 );
buf ( n42915 , n29224 );
not ( n42916 , n42915 );
buf ( n42917 , n29237 );
not ( n42918 , n42917 );
buf ( n42919 , n29295 );
not ( n42920 , n42919 );
buf ( n42921 , n29315 );
not ( n42922 , n42921 );
and ( n42923 , n39704 , n39711 );
and ( n42924 , n42922 , n42923 );
and ( n42925 , n42920 , n42924 );
and ( n42926 , n42918 , n42925 );
and ( n42927 , n42916 , n42926 );
xor ( n42928 , n42914 , n42927 );
buf ( n42929 , n42928 );
and ( n42930 , n42929 , n28586 );
and ( n42931 , n26599 , n34573 );
or ( n42932 , n42930 , n42931 );
and ( n42933 , n42932 , n31002 );
and ( n42934 , n26599 , n34607 );
or ( n42935 , n42868 , n42888 , n42908 , n42912 , n42933 , n42934 );
and ( n42936 , n42823 , n42935 );
and ( n42937 , n26599 , n24800 );
or ( n42938 , n42936 , n42937 );
and ( n42939 , n42938 , n31008 );
and ( n42940 , n26599 , n10618 );
or ( n42941 , n42939 , n42940 );
buf ( n42942 , n42941 );
buf ( n42943 , n42942 );
buf ( n42944 , n10613 );
buf ( n42945 , n10615 );
buf ( n42946 , n10613 );
buf ( n42947 , n10615 );
not ( n42948 , n17451 );
not ( n42949 , n19474 );
and ( n42950 , n42949 , n18859 );
xor ( n42951 , n19491 , n19511 );
and ( n42952 , n42951 , n19474 );
or ( n42953 , n42950 , n42952 );
buf ( n42954 , n42953 );
and ( n42955 , n42954 , n19745 );
and ( n42956 , n42954 , n19748 );
not ( n42957 , n19750 );
and ( n42958 , n42957 , n20811 );
not ( n42959 , n21193 );
and ( n42960 , n42959 , n20823 );
xor ( n42961 , n21210 , n21232 );
and ( n42962 , n42961 , n21193 );
or ( n42963 , n42960 , n42962 );
buf ( n42964 , n42963 );
and ( n42965 , n42964 , n19750 );
or ( n42966 , n42958 , n42965 );
and ( n42967 , n42966 , n21253 );
and ( n42968 , n20811 , n21255 );
or ( n42969 , n42955 , n42956 , n42967 , n42968 );
and ( n42970 , n42969 , n21334 );
and ( n42971 , n18879 , n34492 );
or ( n42972 , n42970 , n42971 );
and ( n42973 , n42972 , n21341 );
not ( n42974 , n22996 );
and ( n42975 , n42974 , n22686 );
xor ( n42976 , n23013 , n23035 );
and ( n42977 , n42976 , n22996 );
or ( n42978 , n42975 , n42977 );
buf ( n42979 , n42978 );
and ( n42980 , n42979 , n21334 );
and ( n42981 , n18879 , n34492 );
or ( n42982 , n42980 , n42981 );
and ( n42983 , n42982 , n23064 );
not ( n42984 , n23758 );
and ( n42985 , n42984 , n23448 );
xor ( n42986 , n23775 , n23797 );
and ( n42987 , n42986 , n23758 );
or ( n42988 , n42985 , n42987 );
buf ( n42989 , n42988 );
and ( n42990 , n42989 , n21334 );
and ( n42991 , n18879 , n34492 );
or ( n42992 , n42990 , n42991 );
and ( n42993 , n42992 , n23825 );
and ( n42994 , n22202 , n21334 );
and ( n42995 , n18879 , n34492 );
or ( n42996 , n42994 , n42995 );
and ( n42997 , n42996 , n23832 );
xor ( n42998 , n23865 , n23897 );
buf ( n42999 , n42998 );
and ( n43000 , n42999 , n21334 );
and ( n43001 , n18879 , n34492 );
or ( n43002 , n43000 , n43001 );
and ( n43003 , n43002 , n23917 );
and ( n43004 , n18879 , n34526 );
or ( n43005 , n42973 , n42983 , n42993 , n42997 , n43003 , n43004 );
and ( n43006 , n42948 , n43005 );
and ( n43007 , n18879 , n17451 );
or ( n43008 , n43006 , n43007 );
and ( n43009 , n43008 , n23924 );
and ( n43010 , n18879 , n23926 );
or ( n43011 , n43009 , n43010 );
buf ( n43012 , n43011 );
buf ( n43013 , n43012 );
buf ( n43014 , n10613 );
buf ( n43015 , n10613 );
not ( n43016 , n34821 );
not ( n43017 , n13916 );
and ( n43018 , n43017 , n13694 );
xor ( n43019 , n13695 , n13870 );
and ( n43020 , n43019 , n13916 );
or ( n43021 , n43018 , n43020 );
buf ( n43022 , n43021 );
and ( n43023 , n43022 , n14137 );
and ( n43024 , n43022 , n14143 );
not ( n43025 , n14139 );
and ( n43026 , n43025 , n35965 );
not ( n43027 , n36245 );
and ( n43028 , n43027 , n35977 );
xor ( n43029 , n35977 , n35634 );
xor ( n43030 , n35955 , n35634 );
xor ( n43031 , n35933 , n35634 );
xor ( n43032 , n35911 , n35634 );
xor ( n43033 , n35889 , n35634 );
xor ( n43034 , n35867 , n35634 );
and ( n43035 , n39390 , n39395 );
and ( n43036 , n43034 , n43035 );
and ( n43037 , n43033 , n43036 );
and ( n43038 , n43032 , n43037 );
and ( n43039 , n43031 , n43038 );
and ( n43040 , n43030 , n43039 );
xor ( n43041 , n43029 , n43040 );
and ( n43042 , n43041 , n36245 );
or ( n43043 , n43028 , n43042 );
buf ( n43044 , n43043 );
and ( n43045 , n43044 , n14139 );
or ( n43046 , n43026 , n43045 );
and ( n43047 , n43046 , n14140 );
and ( n43048 , n35965 , n14141 );
or ( n43049 , n43023 , n43024 , n43047 , n43048 );
and ( n43050 , n43049 , n36347 );
and ( n43051 , n13303 , n39408 );
or ( n43052 , n43050 , n43051 );
and ( n43053 , n43052 , n14562 );
not ( n43054 , n37048 );
and ( n43055 , n43054 , n36823 );
xor ( n43056 , n36823 , n36552 );
xor ( n43057 , n36806 , n36552 );
xor ( n43058 , n36789 , n36552 );
xor ( n43059 , n36772 , n36552 );
xor ( n43060 , n36755 , n36552 );
xor ( n43061 , n36738 , n36552 );
and ( n43062 , n39414 , n39419 );
and ( n43063 , n43061 , n43062 );
and ( n43064 , n43060 , n43063 );
and ( n43065 , n43059 , n43064 );
and ( n43066 , n43058 , n43065 );
and ( n43067 , n43057 , n43066 );
xor ( n43068 , n43056 , n43067 );
and ( n43069 , n43068 , n37048 );
or ( n43070 , n43055 , n43069 );
buf ( n43071 , n43070 );
and ( n43072 , n43071 , n36348 );
and ( n43073 , n13303 , n39427 );
or ( n43074 , n43072 , n43073 );
and ( n43075 , n43074 , n14586 );
not ( n43076 , n37801 );
and ( n43077 , n43076 , n37576 );
xor ( n43078 , n37576 , n37305 );
xor ( n43079 , n37559 , n37305 );
xor ( n43080 , n37542 , n37305 );
xor ( n43081 , n37525 , n37305 );
xor ( n43082 , n37508 , n37305 );
xor ( n43083 , n37491 , n37305 );
and ( n43084 , n39433 , n39438 );
and ( n43085 , n43083 , n43084 );
and ( n43086 , n43082 , n43085 );
and ( n43087 , n43081 , n43086 );
and ( n43088 , n43080 , n43087 );
and ( n43089 , n43079 , n43088 );
xor ( n43090 , n43078 , n43089 );
and ( n43091 , n43090 , n37801 );
or ( n43092 , n43077 , n43091 );
buf ( n43093 , n43092 );
and ( n43094 , n43093 , n36347 );
and ( n43095 , n13303 , n39446 );
or ( n43096 , n43094 , n43095 );
and ( n43097 , n43096 , n14584 );
and ( n43098 , n43071 , n36348 );
and ( n43099 , n13303 , n39453 );
or ( n43100 , n43098 , n43099 );
and ( n43101 , n43100 , n37835 );
and ( n43102 , n43093 , n36348 );
and ( n43103 , n13303 , n39453 );
or ( n43104 , n43102 , n43103 );
and ( n43105 , n43104 , n37841 );
and ( n43106 , n15515 , n36348 );
and ( n43107 , n13303 , n39453 );
or ( n43108 , n43106 , n43107 );
and ( n43109 , n43108 , n37847 );
and ( n43110 , n13303 , n37849 );
or ( n43111 , n43053 , n43075 , n43097 , n43101 , n43105 , n43109 , n43110 );
and ( n43112 , n43016 , n43111 );
and ( n43113 , n13303 , n34821 );
or ( n43114 , n43112 , n43113 );
and ( n43115 , n43114 , n16574 );
and ( n43116 , n13303 , n16576 );
or ( n43117 , n43115 , n43116 );
buf ( n43118 , n43117 );
buf ( n43119 , n43118 );
buf ( n43120 , n10615 );
not ( n43121 , n34821 );
not ( n43122 , n13916 );
and ( n43123 , n43122 , n13826 );
xor ( n43124 , n13827 , n13858 );
and ( n43125 , n43124 , n13916 );
or ( n43126 , n43123 , n43125 );
buf ( n43127 , n43126 );
and ( n43128 , n43127 , n14137 );
and ( n43129 , n43127 , n14143 );
not ( n43130 , n14139 );
and ( n43131 , n43130 , n35709 );
not ( n43132 , n36245 );
and ( n43133 , n43132 , n35721 );
xor ( n43134 , n36251 , n36259 );
and ( n43135 , n43134 , n36245 );
or ( n43136 , n43133 , n43135 );
buf ( n43137 , n43136 );
and ( n43138 , n43137 , n14139 );
or ( n43139 , n43131 , n43138 );
and ( n43140 , n43139 , n14140 );
and ( n43141 , n35709 , n14141 );
or ( n43142 , n43128 , n43129 , n43140 , n43141 );
and ( n43143 , n43142 , n36345 );
and ( n43144 , n13449 , n36352 );
or ( n43145 , n43143 , n43144 );
and ( n43146 , n43145 , n14562 );
not ( n43147 , n37048 );
and ( n43148 , n43147 , n36619 );
xor ( n43149 , n37054 , n37062 );
and ( n43150 , n43149 , n37048 );
or ( n43151 , n43148 , n43150 );
buf ( n43152 , n43151 );
and ( n43153 , n43152 , n36345 );
and ( n43154 , n13449 , n37073 );
or ( n43155 , n43153 , n43154 );
and ( n43156 , n43155 , n14586 );
not ( n43157 , n37801 );
and ( n43158 , n43157 , n37372 );
xor ( n43159 , n37807 , n37815 );
and ( n43160 , n43159 , n37801 );
or ( n43161 , n43158 , n43160 );
buf ( n43162 , n43161 );
and ( n43163 , n43162 , n36350 );
and ( n43164 , n13449 , n37825 );
or ( n43165 , n43163 , n43164 );
and ( n43166 , n43165 , n14584 );
and ( n43167 , n43152 , n36350 );
and ( n43168 , n13449 , n37831 );
or ( n43169 , n43167 , n43168 );
and ( n43170 , n43169 , n37835 );
and ( n43171 , n43162 , n36350 );
and ( n43172 , n13449 , n37831 );
or ( n43173 , n43171 , n43172 );
and ( n43174 , n43173 , n37841 );
and ( n43175 , n15779 , n36350 );
and ( n43176 , n13449 , n37831 );
or ( n43177 , n43175 , n43176 );
and ( n43178 , n43177 , n37847 );
and ( n43179 , n13449 , n37849 );
or ( n43180 , n43146 , n43156 , n43166 , n43170 , n43174 , n43178 , n43179 );
and ( n43181 , n43121 , n43180 );
and ( n43182 , n13449 , n34821 );
or ( n43183 , n43181 , n43182 );
and ( n43184 , n43183 , n16574 );
and ( n43185 , n13449 , n16576 );
or ( n43186 , n43184 , n43185 );
buf ( n43187 , n43186 );
buf ( n43188 , n43187 );
buf ( n43189 , n10615 );
buf ( n43190 , n10615 );
buf ( n43191 , n10615 );
buf ( n43192 , n10613 );
buf ( n43193 , n10615 );
buf ( n43194 , n10613 );
buf ( n43195 , n10613 );
not ( n43196 , n24800 );
and ( n43197 , n31072 , n28586 );
and ( n43198 , n26191 , n34573 );
or ( n43199 , n43197 , n43198 );
and ( n43200 , n43199 , n28594 );
and ( n43201 , n31102 , n28586 );
and ( n43202 , n26191 , n34573 );
or ( n43203 , n43201 , n43202 );
and ( n43204 , n43203 , n30269 );
and ( n43205 , n31130 , n28586 );
and ( n43206 , n26191 , n34573 );
or ( n43207 , n43205 , n43206 );
and ( n43208 , n43207 , n30982 );
and ( n43209 , n29475 , n28586 );
and ( n43210 , n26191 , n34573 );
or ( n43211 , n43209 , n43210 );
and ( n43212 , n43211 , n30989 );
and ( n43213 , n31168 , n28586 );
and ( n43214 , n26191 , n34573 );
or ( n43215 , n43213 , n43214 );
and ( n43216 , n43215 , n31002 );
and ( n43217 , n26191 , n34607 );
or ( n43218 , n43200 , n43204 , n43208 , n43212 , n43216 , n43217 );
and ( n43219 , n43196 , n43218 );
and ( n43220 , n26191 , n24800 );
or ( n43221 , n43219 , n43220 );
and ( n43222 , n43221 , n31008 );
and ( n43223 , n26191 , n10618 );
or ( n43224 , n43222 , n43223 );
buf ( n43225 , n43224 );
buf ( n43226 , n43225 );
buf ( n43227 , n10613 );
buf ( n43228 , n10615 );
buf ( n43229 , n10615 );
buf ( n43230 , n10615 );
buf ( n43231 , n10613 );
not ( n43232 , n34821 );
and ( n43233 , n43142 , n36347 );
and ( n43234 , n13447 , n39408 );
or ( n43235 , n43233 , n43234 );
and ( n43236 , n43235 , n14562 );
and ( n43237 , n43152 , n36348 );
and ( n43238 , n13447 , n39427 );
or ( n43239 , n43237 , n43238 );
and ( n43240 , n43239 , n14586 );
and ( n43241 , n43162 , n36347 );
and ( n43242 , n13447 , n39446 );
or ( n43243 , n43241 , n43242 );
and ( n43244 , n43243 , n14584 );
and ( n43245 , n43152 , n36348 );
and ( n43246 , n13447 , n39453 );
or ( n43247 , n43245 , n43246 );
and ( n43248 , n43247 , n37835 );
and ( n43249 , n43162 , n36348 );
and ( n43250 , n13447 , n39453 );
or ( n43251 , n43249 , n43250 );
and ( n43252 , n43251 , n37841 );
and ( n43253 , n15779 , n36348 );
and ( n43254 , n13447 , n39453 );
or ( n43255 , n43253 , n43254 );
and ( n43256 , n43255 , n37847 );
and ( n43257 , n13447 , n37849 );
or ( n43258 , n43236 , n43240 , n43244 , n43248 , n43252 , n43256 , n43257 );
and ( n43259 , n43232 , n43258 );
and ( n43260 , n13447 , n34821 );
or ( n43261 , n43259 , n43260 );
and ( n43262 , n43261 , n16574 );
and ( n43263 , n13447 , n16576 );
or ( n43264 , n43262 , n43263 );
buf ( n43265 , n43264 );
buf ( n43266 , n43265 );
not ( n43267 , n17451 );
and ( n43268 , n39876 , n21333 );
and ( n43269 , n19386 , n34758 );
or ( n43270 , n43268 , n43269 );
and ( n43271 , n43270 , n21341 );
and ( n43272 , n39888 , n21333 );
and ( n43273 , n19386 , n34758 );
or ( n43274 , n43272 , n43273 );
and ( n43275 , n43274 , n23064 );
and ( n43276 , n39900 , n21333 );
and ( n43277 , n19386 , n34758 );
or ( n43278 , n43276 , n43277 );
and ( n43279 , n43278 , n23825 );
and ( n43280 , n21906 , n21333 );
and ( n43281 , n19386 , n34758 );
or ( n43282 , n43280 , n43281 );
and ( n43283 , n43282 , n23832 );
and ( n43284 , n39913 , n21333 );
and ( n43285 , n19386 , n34758 );
or ( n43286 , n43284 , n43285 );
and ( n43287 , n43286 , n23917 );
and ( n43288 , n19386 , n34526 );
or ( n43289 , n43271 , n43275 , n43279 , n43283 , n43287 , n43288 );
and ( n43290 , n43267 , n43289 );
and ( n43291 , n19386 , n17451 );
or ( n43292 , n43290 , n43291 );
and ( n43293 , n43292 , n23924 );
and ( n43294 , n19386 , n23926 );
or ( n43295 , n43293 , n43294 );
buf ( n43296 , n43295 );
buf ( n43297 , n43296 );
buf ( n43298 , n10613 );
buf ( n43299 , n10613 );
buf ( n43300 , n10613 );
buf ( n43301 , n10615 );
buf ( n43302 , n10615 );
and ( n43303 , n17016 , n23924 );
and ( n43304 , n21917 , n23926 );
or ( n43305 , n43303 , n43304 );
buf ( n43306 , n43305 );
buf ( n43307 , n43306 );
buf ( n43308 , n10613 );
and ( n43309 , n16889 , n23924 );
and ( n43310 , n22373 , n23926 );
or ( n43311 , n43309 , n43310 );
buf ( n43312 , n43311 );
buf ( n43313 , n43312 );
buf ( n43314 , n10615 );
buf ( n43315 , n10615 );
buf ( n43316 , n10615 );
not ( n43317 , n17451 );
not ( n43318 , n19474 );
and ( n43319 , n43318 , n18893 );
xor ( n43320 , n19490 , n19512 );
and ( n43321 , n43320 , n19474 );
or ( n43322 , n43319 , n43321 );
buf ( n43323 , n43322 );
and ( n43324 , n43323 , n19745 );
and ( n43325 , n43323 , n19748 );
not ( n43326 , n19750 );
and ( n43327 , n43326 , n20833 );
not ( n43328 , n21193 );
and ( n43329 , n43328 , n20845 );
xor ( n43330 , n21209 , n21233 );
and ( n43331 , n43330 , n21193 );
or ( n43332 , n43329 , n43331 );
buf ( n43333 , n43332 );
and ( n43334 , n43333 , n19750 );
or ( n43335 , n43327 , n43334 );
and ( n43336 , n43335 , n21253 );
and ( n43337 , n20833 , n21255 );
or ( n43338 , n43324 , n43325 , n43336 , n43337 );
and ( n43339 , n43338 , n21334 );
and ( n43340 , n18913 , n34492 );
or ( n43341 , n43339 , n43340 );
and ( n43342 , n43341 , n21341 );
not ( n43343 , n22996 );
and ( n43344 , n43343 , n22703 );
xor ( n43345 , n23012 , n23036 );
and ( n43346 , n43345 , n22996 );
or ( n43347 , n43344 , n43346 );
buf ( n43348 , n43347 );
and ( n43349 , n43348 , n21334 );
and ( n43350 , n18913 , n34492 );
or ( n43351 , n43349 , n43350 );
and ( n43352 , n43351 , n23064 );
not ( n43353 , n23758 );
and ( n43354 , n43353 , n23465 );
xor ( n43355 , n23774 , n23798 );
and ( n43356 , n43355 , n23758 );
or ( n43357 , n43354 , n43356 );
buf ( n43358 , n43357 );
and ( n43359 , n43358 , n21334 );
and ( n43360 , n18913 , n34492 );
or ( n43361 , n43359 , n43360 );
and ( n43362 , n43361 , n23825 );
and ( n43363 , n22182 , n21334 );
and ( n43364 , n18913 , n34492 );
or ( n43365 , n43363 , n43364 );
and ( n43366 , n43365 , n23832 );
xor ( n43367 , n23863 , n23898 );
buf ( n43368 , n43367 );
and ( n43369 , n43368 , n21334 );
and ( n43370 , n18913 , n34492 );
or ( n43371 , n43369 , n43370 );
and ( n43372 , n43371 , n23917 );
and ( n43373 , n18913 , n34526 );
or ( n43374 , n43342 , n43352 , n43362 , n43366 , n43372 , n43373 );
and ( n43375 , n43317 , n43374 );
and ( n43376 , n18913 , n17451 );
or ( n43377 , n43375 , n43376 );
and ( n43378 , n43377 , n23924 );
and ( n43379 , n18913 , n23926 );
or ( n43380 , n43378 , n43379 );
buf ( n43381 , n43380 );
buf ( n43382 , n43381 );
buf ( n43383 , n10615 );
buf ( n43384 , n10613 );
buf ( n43385 , n10613 );
buf ( n43386 , n10615 );
not ( n43387 , n24800 );
not ( n43388 , n26823 );
and ( n43389 , n43388 , n26683 );
xor ( n43390 , n26683 , n25877 );
xor ( n43391 , n26649 , n25877 );
xor ( n43392 , n26615 , n25877 );
and ( n43393 , n42826 , n42835 );
and ( n43394 , n43392 , n43393 );
and ( n43395 , n43391 , n43394 );
xor ( n43396 , n43390 , n43395 );
and ( n43397 , n43396 , n26823 );
or ( n43398 , n43389 , n43397 );
buf ( n43399 , n43398 );
and ( n43400 , n43399 , n27046 );
and ( n43401 , n43399 , n27049 );
not ( n43402 , n27051 );
and ( n43403 , n43402 , n28412 );
not ( n43404 , n28494 );
and ( n43405 , n43404 , n28424 );
xor ( n43406 , n28424 , n27883 );
xor ( n43407 , n28402 , n27883 );
xor ( n43408 , n28380 , n27883 );
and ( n43409 , n42846 , n42855 );
and ( n43410 , n43408 , n43409 );
and ( n43411 , n43407 , n43410 );
xor ( n43412 , n43406 , n43411 );
and ( n43413 , n43412 , n28494 );
or ( n43414 , n43405 , n43413 );
buf ( n43415 , n43414 );
and ( n43416 , n43415 , n27051 );
or ( n43417 , n43403 , n43416 );
and ( n43418 , n43417 , n28506 );
and ( n43419 , n28412 , n28508 );
or ( n43420 , n43400 , n43401 , n43418 , n43419 );
and ( n43421 , n43420 , n28587 );
and ( n43422 , n26703 , n39807 );
or ( n43423 , n43421 , n43422 );
and ( n43424 , n43423 , n28594 );
not ( n43425 , n30249 );
and ( n43426 , n43425 , n30177 );
xor ( n43427 , n30177 , n29753 );
xor ( n43428 , n30160 , n29753 );
xor ( n43429 , n30143 , n29753 );
and ( n43430 , n42871 , n42880 );
and ( n43431 , n43429 , n43430 );
and ( n43432 , n43428 , n43431 );
xor ( n43433 , n43427 , n43432 );
and ( n43434 , n43433 , n30249 );
or ( n43435 , n43426 , n43434 );
buf ( n43436 , n43435 );
and ( n43437 , n43436 , n28587 );
and ( n43438 , n26703 , n39807 );
or ( n43439 , n43437 , n43438 );
and ( n43440 , n43439 , n30269 );
not ( n43441 , n30963 );
and ( n43442 , n43441 , n30891 );
xor ( n43443 , n30891 , n30467 );
xor ( n43444 , n30874 , n30467 );
xor ( n43445 , n30857 , n30467 );
and ( n43446 , n42891 , n42900 );
and ( n43447 , n43445 , n43446 );
and ( n43448 , n43444 , n43447 );
xor ( n43449 , n43443 , n43448 );
and ( n43450 , n43449 , n30963 );
or ( n43451 , n43442 , n43450 );
buf ( n43452 , n43451 );
and ( n43453 , n43452 , n28587 );
and ( n43454 , n26703 , n39807 );
or ( n43455 , n43453 , n43454 );
and ( n43456 , n43455 , n30982 );
and ( n43457 , n29172 , n28587 );
and ( n43458 , n26703 , n39807 );
or ( n43459 , n43457 , n43458 );
and ( n43460 , n43459 , n30989 );
buf ( n43461 , n29172 );
not ( n43462 , n43461 );
buf ( n43463 , n29185 );
not ( n43464 , n43463 );
buf ( n43465 , n29198 );
not ( n43466 , n43465 );
and ( n43467 , n42914 , n42927 );
and ( n43468 , n43466 , n43467 );
and ( n43469 , n43464 , n43468 );
xor ( n43470 , n43462 , n43469 );
buf ( n43471 , n43470 );
and ( n43472 , n43471 , n28587 );
and ( n43473 , n26703 , n39807 );
or ( n43474 , n43472 , n43473 );
and ( n43475 , n43474 , n31002 );
and ( n43476 , n26703 , n34607 );
or ( n43477 , n43424 , n43440 , n43456 , n43460 , n43475 , n43476 );
and ( n43478 , n43387 , n43477 );
and ( n43479 , n26703 , n24800 );
or ( n43480 , n43478 , n43479 );
and ( n43481 , n43480 , n31008 );
and ( n43482 , n26703 , n10618 );
or ( n43483 , n43481 , n43482 );
buf ( n43484 , n43483 );
buf ( n43485 , n43484 );
buf ( n43486 , n10613 );
not ( n43487 , n34821 );
and ( n43488 , n43487 , n36343 );
and ( n43489 , n36319 , n34821 );
or ( n43490 , n43488 , n43489 );
and ( n43491 , n43490 , n16574 );
and ( n43492 , n36319 , n16576 );
or ( n43493 , n43491 , n43492 );
buf ( n43494 , n43493 );
buf ( n43495 , n43494 );
buf ( n43496 , n10613 );
buf ( n43497 , n10613 );
buf ( n43498 , n10615 );
buf ( n43499 , n10615 );
buf ( n43500 , n10615 );
buf ( n43501 , n10613 );
buf ( n43502 , n10613 );
buf ( n43503 , n10615 );
not ( n43504 , n34821 );
and ( n43505 , n13491 , n14592 );
not ( n43506 , n13916 );
and ( n43507 , n43506 , n13854 );
xor ( n43508 , n13855 , n13151 );
and ( n43509 , n43508 , n13916 );
or ( n43510 , n43507 , n43509 );
buf ( n43511 , n43510 );
and ( n43512 , n43511 , n14137 );
and ( n43513 , n43511 , n14143 );
not ( n43514 , n14139 );
and ( n43515 , n43514 , n35643 );
not ( n43516 , n36245 );
and ( n43517 , n43516 , n35655 );
xor ( n43518 , n36254 , n36256 );
and ( n43519 , n43518 , n36245 );
or ( n43520 , n43517 , n43519 );
buf ( n43521 , n43520 );
and ( n43522 , n43521 , n14139 );
or ( n43523 , n43515 , n43522 );
and ( n43524 , n43523 , n14140 );
and ( n43525 , n35643 , n14141 );
or ( n43526 , n43512 , n43513 , n43524 , n43525 );
and ( n43527 , n43526 , n36348 );
or ( n43528 , n36347 , n36345 );
or ( n43529 , n43528 , n36350 );
or ( n43530 , n43529 , C0 );
and ( n43531 , n13491 , n43530 );
or ( n43532 , n43527 , n43531 );
and ( n43533 , n43532 , n14562 );
not ( n43534 , n37048 );
and ( n43535 , n43534 , n36568 );
xor ( n43536 , n37057 , n37059 );
and ( n43537 , n43536 , n37048 );
or ( n43538 , n43535 , n43537 );
buf ( n43539 , n43538 );
and ( n43540 , n43539 , n36347 );
or ( n43541 , n36348 , n36345 );
or ( n43542 , n43541 , n36350 );
or ( n43543 , n43542 , C0 );
and ( n43544 , n13491 , n43543 );
or ( n43545 , n43540 , n43544 );
and ( n43546 , n43545 , n14586 );
not ( n43547 , n37801 );
and ( n43548 , n43547 , n37321 );
xor ( n43549 , n37810 , n37812 );
and ( n43550 , n43549 , n37801 );
or ( n43551 , n43548 , n43550 );
buf ( n43552 , n43551 );
and ( n43553 , n43552 , n36348 );
or ( n43554 , n36347 , n36350 );
or ( n43555 , n43554 , n36345 );
or ( n43556 , n43555 , C0 );
and ( n43557 , n13491 , n43556 );
or ( n43558 , n43553 , n43557 );
and ( n43559 , n43558 , n14584 );
and ( n43560 , n43539 , n36347 );
or ( n43561 , n36348 , n36350 );
or ( n43562 , n43561 , n36345 );
or ( n43563 , n43562 , C0 );
and ( n43564 , n13491 , n43563 );
or ( n43565 , n43560 , n43564 );
and ( n43566 , n43565 , n37835 );
and ( n43567 , n43552 , n36347 );
and ( n43568 , n13491 , n43563 );
or ( n43569 , n43567 , n43568 );
and ( n43570 , n43569 , n37841 );
and ( n43571 , n13489 , n14564 );
and ( n43572 , n15845 , n36347 );
and ( n43573 , n13491 , n43563 );
or ( n43574 , n43572 , n43573 );
and ( n43575 , n43574 , n37847 );
or ( n43576 , n43505 , n43533 , n43546 , n43559 , n43566 , n43570 , n43571 , n43575 );
and ( n43577 , n43504 , n43576 );
and ( n43578 , n13491 , n34821 );
or ( n43579 , n43577 , n43578 );
and ( n43580 , n43579 , n16574 );
and ( n43581 , n13491 , n16576 );
or ( n43582 , n43580 , n43581 );
buf ( n43583 , n43582 );
buf ( n43584 , n43583 );
not ( n43585 , n34538 );
and ( n43586 , n43585 , n18610 );
and ( n43587 , n14813 , n34538 );
or ( n43588 , n43586 , n43587 );
and ( n43589 , n43588 , n23924 );
and ( n43590 , n14813 , n23926 );
or ( n43591 , n43589 , n43590 );
buf ( n43592 , n43591 );
buf ( n43593 , n43592 );
buf ( n43594 , n10615 );
not ( n43595 , n34821 );
and ( n43596 , n13337 , n14592 );
not ( n43597 , n13916 );
and ( n43598 , n43597 , n13727 );
xor ( n43599 , n13728 , n13867 );
and ( n43600 , n43599 , n13916 );
or ( n43601 , n43598 , n43600 );
buf ( n43602 , n43601 );
and ( n43603 , n43602 , n14137 );
and ( n43604 , n43602 , n14143 );
not ( n43605 , n14139 );
and ( n43606 , n43605 , n35899 );
not ( n43607 , n36245 );
and ( n43608 , n43607 , n35911 );
xor ( n43609 , n43032 , n43037 );
and ( n43610 , n43609 , n36245 );
or ( n43611 , n43608 , n43610 );
buf ( n43612 , n43611 );
and ( n43613 , n43612 , n14139 );
or ( n43614 , n43606 , n43613 );
and ( n43615 , n43614 , n14140 );
and ( n43616 , n35899 , n14141 );
or ( n43617 , n43603 , n43604 , n43615 , n43616 );
and ( n43618 , n43617 , n36348 );
and ( n43619 , n13337 , n43530 );
or ( n43620 , n43618 , n43619 );
and ( n43621 , n43620 , n14562 );
not ( n43622 , n37048 );
and ( n43623 , n43622 , n36772 );
xor ( n43624 , n43059 , n43064 );
and ( n43625 , n43624 , n37048 );
or ( n43626 , n43623 , n43625 );
buf ( n43627 , n43626 );
and ( n43628 , n43627 , n36347 );
and ( n43629 , n13337 , n43543 );
or ( n43630 , n43628 , n43629 );
and ( n43631 , n43630 , n14586 );
not ( n43632 , n37801 );
and ( n43633 , n43632 , n37525 );
xor ( n43634 , n43081 , n43086 );
and ( n43635 , n43634 , n37801 );
or ( n43636 , n43633 , n43635 );
buf ( n43637 , n43636 );
and ( n43638 , n43637 , n36348 );
and ( n43639 , n13337 , n43556 );
or ( n43640 , n43638 , n43639 );
and ( n43641 , n43640 , n14584 );
and ( n43642 , n43627 , n36347 );
and ( n43643 , n13337 , n43563 );
or ( n43644 , n43642 , n43643 );
and ( n43645 , n43644 , n37835 );
and ( n43646 , n43637 , n36347 );
and ( n43647 , n13337 , n43563 );
or ( n43648 , n43646 , n43647 );
and ( n43649 , n43648 , n37841 );
and ( n43650 , n13335 , n14564 );
and ( n43651 , n15581 , n36347 );
and ( n43652 , n13337 , n43563 );
or ( n43653 , n43651 , n43652 );
and ( n43654 , n43653 , n37847 );
or ( n43655 , n43596 , n43621 , n43631 , n43641 , n43645 , n43649 , n43650 , n43654 );
and ( n43656 , n43595 , n43655 );
and ( n43657 , n13337 , n34821 );
or ( n43658 , n43656 , n43657 );
and ( n43659 , n43658 , n16574 );
and ( n43660 , n13337 , n16576 );
or ( n43661 , n43659 , n43660 );
buf ( n43662 , n43661 );
buf ( n43663 , n43662 );
buf ( n43664 , n10615 );
buf ( n43665 , n10615 );
not ( n43666 , n34821 );
and ( n43667 , n13347 , n14592 );
not ( n43668 , n13916 );
and ( n43669 , n43668 , n13738 );
xor ( n43670 , n13739 , n13866 );
and ( n43671 , n43670 , n13916 );
or ( n43672 , n43669 , n43671 );
buf ( n43673 , n43672 );
and ( n43674 , n43673 , n14137 );
and ( n43675 , n43673 , n14143 );
not ( n43676 , n14139 );
and ( n43677 , n43676 , n35877 );
not ( n43678 , n36245 );
and ( n43679 , n43678 , n35889 );
xor ( n43680 , n43033 , n43036 );
and ( n43681 , n43680 , n36245 );
or ( n43682 , n43679 , n43681 );
buf ( n43683 , n43682 );
and ( n43684 , n43683 , n14139 );
or ( n43685 , n43677 , n43684 );
and ( n43686 , n43685 , n14140 );
and ( n43687 , n35877 , n14141 );
or ( n43688 , n43674 , n43675 , n43686 , n43687 );
and ( n43689 , n43688 , n36350 );
or ( n43690 , n43528 , n36348 );
or ( n43691 , n43690 , C0 );
and ( n43692 , n13347 , n43691 );
or ( n43693 , n43689 , n43692 );
and ( n43694 , n43693 , n14562 );
not ( n43695 , n37048 );
and ( n43696 , n43695 , n36755 );
xor ( n43697 , n43060 , n43063 );
and ( n43698 , n43697 , n37048 );
or ( n43699 , n43696 , n43698 );
buf ( n43700 , n43699 );
and ( n43701 , n43700 , n36350 );
or ( n43702 , n43541 , n36347 );
or ( n43703 , n43702 , C0 );
and ( n43704 , n13347 , n43703 );
or ( n43705 , n43701 , n43704 );
and ( n43706 , n43705 , n14586 );
not ( n43707 , n37801 );
and ( n43708 , n43707 , n37508 );
xor ( n43709 , n43082 , n43085 );
and ( n43710 , n43709 , n37801 );
or ( n43711 , n43708 , n43710 );
buf ( n43712 , n43711 );
and ( n43713 , n43712 , n36345 );
or ( n43714 , n43554 , n36348 );
or ( n43715 , n43714 , C0 );
and ( n43716 , n13347 , n43715 );
or ( n43717 , n43713 , n43716 );
and ( n43718 , n43717 , n14584 );
and ( n43719 , n43700 , n36345 );
or ( n43720 , n43561 , n36347 );
or ( n43721 , n43720 , C0 );
and ( n43722 , n13347 , n43721 );
or ( n43723 , n43719 , n43722 );
and ( n43724 , n43723 , n37835 );
and ( n43725 , n43712 , n36345 );
and ( n43726 , n13347 , n43721 );
or ( n43727 , n43725 , n43726 );
and ( n43728 , n43727 , n37841 );
and ( n43729 , n15603 , n14564 );
and ( n43730 , n15603 , n36345 );
and ( n43731 , n13347 , n43721 );
or ( n43732 , n43730 , n43731 );
and ( n43733 , n43732 , n37847 );
or ( n43734 , n43667 , n43694 , n43706 , n43718 , n43724 , n43728 , n43729 , n43733 );
and ( n43735 , n43666 , n43734 );
and ( n43736 , n13347 , n34821 );
or ( n43737 , n43735 , n43736 );
and ( n43738 , n43737 , n16574 );
and ( n43739 , n12297 , n16576 );
or ( n43740 , n43738 , n43739 );
buf ( n43741 , n43740 );
buf ( n43742 , n43741 );
buf ( n43743 , n10613 );
buf ( n43744 , n10615 );
buf ( n43745 , n10613 );
not ( n43746 , n24511 );
not ( n43747 , n24799 );
and ( n43748 , n10640 , n40154 );
not ( n43749 , n40632 );
and ( n43750 , n43749 , n40628 );
xor ( n43751 , n40628 , n40306 );
xor ( n43752 , n40611 , n40306 );
xor ( n43753 , n40594 , n40306 );
xor ( n43754 , n40577 , n40306 );
and ( n43755 , n40635 , n40665 );
and ( n43756 , n43754 , n43755 );
and ( n43757 , n43753 , n43756 );
and ( n43758 , n43752 , n43757 );
xor ( n43759 , n43751 , n43758 );
and ( n43760 , n43759 , n40632 );
or ( n43761 , n43750 , n43760 );
buf ( n43762 , n43761 );
and ( n43763 , n43762 , n27046 );
not ( n43764 , n41147 );
and ( n43765 , n43764 , n41143 );
xor ( n43766 , n41143 , n40821 );
xor ( n43767 , n41126 , n40821 );
xor ( n43768 , n41109 , n40821 );
xor ( n43769 , n41092 , n40821 );
and ( n43770 , n41150 , n41180 );
and ( n43771 , n43769 , n43770 );
and ( n43772 , n43768 , n43771 );
and ( n43773 , n43767 , n43772 );
xor ( n43774 , n43766 , n43773 );
and ( n43775 , n43774 , n41147 );
or ( n43776 , n43765 , n43775 );
buf ( n43777 , n43776 );
and ( n43778 , n43777 , n27049 );
and ( n43779 , n29293 , n28506 );
and ( n43780 , n10640 , n28508 );
or ( n43781 , n43763 , n43778 , n43779 , n43780 );
and ( n43782 , n43781 , n41199 );
or ( n43783 , n43748 , n43782 );
and ( n43784 , n43747 , n43783 );
not ( n43785 , n41478 );
and ( n43786 , n43785 , n41474 );
xor ( n43787 , n41474 , n41209 );
xor ( n43788 , n41460 , n41209 );
xor ( n43789 , n41446 , n41209 );
xor ( n43790 , n41432 , n41209 );
and ( n43791 , n41481 , n41511 );
and ( n43792 , n43790 , n43791 );
and ( n43793 , n43789 , n43792 );
and ( n43794 , n43788 , n43793 );
xor ( n43795 , n43787 , n43794 );
and ( n43796 , n43795 , n41478 );
or ( n43797 , n43786 , n43796 );
buf ( n43798 , n43797 );
buf ( n43799 , n43798 );
buf ( n43800 , n29293 );
not ( n43801 , n43800 );
buf ( n43802 , n43801 );
buf ( n43803 , n43802 );
not ( n43804 , n43803 );
buf ( n43805 , n43804 );
buf ( n43806 , n43805 );
buf ( n43807 , n43806 );
xor ( n43808 , n43799 , n43807 );
not ( n43809 , n41478 );
and ( n43810 , n43809 , n41460 );
xor ( n43811 , n43788 , n43793 );
and ( n43812 , n43811 , n41478 );
or ( n43813 , n43810 , n43812 );
buf ( n43814 , n43813 );
buf ( n43815 , n43814 );
buf ( n43816 , n29313 );
not ( n43817 , n43816 );
buf ( n43818 , n43817 );
buf ( n43819 , n43818 );
not ( n43820 , n43819 );
buf ( n43821 , n43820 );
buf ( n43822 , n43821 );
buf ( n43823 , n43822 );
and ( n43824 , n43815 , n43823 );
not ( n43825 , n41478 );
and ( n43826 , n43825 , n41446 );
xor ( n43827 , n43789 , n43792 );
and ( n43828 , n43827 , n41478 );
or ( n43829 , n43826 , n43828 );
buf ( n43830 , n43829 );
buf ( n43831 , n43830 );
buf ( n43832 , n29333 );
not ( n43833 , n43832 );
buf ( n43834 , n43833 );
buf ( n43835 , n43834 );
not ( n43836 , n43835 );
buf ( n43837 , n43836 );
buf ( n43838 , n43837 );
buf ( n43839 , n43838 );
and ( n43840 , n43831 , n43839 );
not ( n43841 , n41478 );
and ( n43842 , n43841 , n41432 );
xor ( n43843 , n43790 , n43791 );
and ( n43844 , n43843 , n41478 );
or ( n43845 , n43842 , n43844 );
buf ( n43846 , n43845 );
buf ( n43847 , n43846 );
buf ( n43848 , n29353 );
not ( n43849 , n43848 );
buf ( n43850 , n43849 );
buf ( n43851 , n43850 );
not ( n43852 , n43851 );
buf ( n43853 , n43852 );
buf ( n43854 , n43853 );
buf ( n43855 , n43854 );
and ( n43856 , n43847 , n43855 );
and ( n43857 , n41516 , n41524 );
and ( n43858 , n41524 , n41806 );
and ( n43859 , n41516 , n41806 );
or ( n43860 , n43857 , n43858 , n43859 );
and ( n43861 , n43855 , n43860 );
and ( n43862 , n43847 , n43860 );
or ( n43863 , n43856 , n43861 , n43862 );
and ( n43864 , n43839 , n43863 );
and ( n43865 , n43831 , n43863 );
or ( n43866 , n43840 , n43864 , n43865 );
and ( n43867 , n43823 , n43866 );
and ( n43868 , n43815 , n43866 );
or ( n43869 , n43824 , n43867 , n43868 );
xor ( n43870 , n43808 , n43869 );
buf ( n43871 , n43870 );
and ( n43872 , n43871 , n27046 );
not ( n43873 , n42085 );
and ( n43874 , n43873 , n42081 );
xor ( n43875 , n42081 , n41816 );
xor ( n43876 , n42067 , n41816 );
xor ( n43877 , n42053 , n41816 );
xor ( n43878 , n42039 , n41816 );
and ( n43879 , n42088 , n42118 );
and ( n43880 , n43878 , n43879 );
and ( n43881 , n43877 , n43880 );
and ( n43882 , n43876 , n43881 );
xor ( n43883 , n43875 , n43882 );
and ( n43884 , n43883 , n42085 );
or ( n43885 , n43874 , n43884 );
buf ( n43886 , n43885 );
buf ( n43887 , n43886 );
buf ( n43888 , n43806 );
xor ( n43889 , n43887 , n43888 );
not ( n43890 , n42085 );
and ( n43891 , n43890 , n42067 );
xor ( n43892 , n43876 , n43881 );
and ( n43893 , n43892 , n42085 );
or ( n43894 , n43891 , n43893 );
buf ( n43895 , n43894 );
buf ( n43896 , n43895 );
buf ( n43897 , n43822 );
and ( n43898 , n43896 , n43897 );
not ( n43899 , n42085 );
and ( n43900 , n43899 , n42053 );
xor ( n43901 , n43877 , n43880 );
and ( n43902 , n43901 , n42085 );
or ( n43903 , n43900 , n43902 );
buf ( n43904 , n43903 );
buf ( n43905 , n43904 );
buf ( n43906 , n43838 );
and ( n43907 , n43905 , n43906 );
not ( n43908 , n42085 );
and ( n43909 , n43908 , n42039 );
xor ( n43910 , n43878 , n43879 );
and ( n43911 , n43910 , n42085 );
or ( n43912 , n43909 , n43911 );
buf ( n43913 , n43912 );
buf ( n43914 , n43913 );
buf ( n43915 , n43854 );
and ( n43916 , n43914 , n43915 );
and ( n43917 , n42123 , n42124 );
and ( n43918 , n42124 , n42302 );
and ( n43919 , n42123 , n42302 );
or ( n43920 , n43917 , n43918 , n43919 );
and ( n43921 , n43915 , n43920 );
and ( n43922 , n43914 , n43920 );
or ( n43923 , n43916 , n43921 , n43922 );
and ( n43924 , n43906 , n43923 );
and ( n43925 , n43905 , n43923 );
or ( n43926 , n43907 , n43924 , n43925 );
and ( n43927 , n43897 , n43926 );
and ( n43928 , n43896 , n43926 );
or ( n43929 , n43898 , n43927 , n43928 );
xor ( n43930 , n43889 , n43929 );
buf ( n43931 , n43930 );
and ( n43932 , n43931 , n27049 );
and ( n43933 , n29293 , n42306 );
or ( n43934 , n43872 , n43932 , n43933 );
buf ( n43935 , n43934 );
and ( n43936 , C1 , n43935 );
or ( n43937 , n43936 , C0 );
buf ( n43938 , n43937 );
not ( n43939 , n43938 );
buf ( n43940 , n43939 );
buf ( n43941 , n43940 );
not ( n43942 , n43941 );
and ( n43943 , C1 , n43942 );
or ( n43944 , n43943 , C0 );
buf ( n43945 , n43944 );
and ( n43946 , n43945 , n24799 );
or ( n43947 , n43784 , n43946 );
and ( n43948 , n43746 , n43947 );
and ( n43949 , n43781 , n24511 );
or ( n43950 , n43948 , n43949 );
and ( n43951 , n43950 , n31008 );
not ( n43952 , n42601 );
and ( n43953 , n43952 , n42597 );
xor ( n43954 , n42597 , n42332 );
xor ( n43955 , n42583 , n42332 );
xor ( n43956 , n42569 , n42332 );
xor ( n43957 , n42555 , n42332 );
and ( n43958 , n42604 , n42634 );
and ( n43959 , n43957 , n43958 );
and ( n43960 , n43956 , n43959 );
and ( n43961 , n43955 , n43960 );
xor ( n43962 , n43954 , n43961 );
and ( n43963 , n43962 , n42601 );
or ( n43964 , n43953 , n43963 );
buf ( n43965 , n43964 );
and ( n43966 , n43965 , n10618 );
or ( n43967 , n43951 , n43966 );
buf ( n43968 , n43967 );
buf ( n43969 , n43968 );
buf ( n43970 , n10615 );
not ( n43971 , n34538 );
and ( n43972 , n43971 , n19119 );
and ( n43973 , n14723 , n34538 );
or ( n43974 , n43972 , n43973 );
and ( n43975 , n43974 , n23924 );
and ( n43976 , n14723 , n23926 );
or ( n43977 , n43975 , n43976 );
buf ( n43978 , n43977 );
buf ( n43979 , n43978 );
buf ( n43980 , n10613 );
buf ( n43981 , n10613 );
not ( n43982 , n34538 );
and ( n43983 , n43982 , n18983 );
and ( n43984 , n14747 , n34538 );
or ( n43985 , n43983 , n43984 );
and ( n43986 , n43985 , n23924 );
and ( n43987 , n14747 , n23926 );
or ( n43988 , n43986 , n43987 );
buf ( n43989 , n43988 );
buf ( n43990 , n43989 );
buf ( n43991 , n10613 );
not ( n43992 , n24800 );
and ( n43993 , n26189 , n25222 );
and ( n43994 , n31072 , n28583 );
and ( n43995 , n26189 , n28591 );
or ( n43996 , n43994 , n43995 );
and ( n43997 , n43996 , n28594 );
and ( n43998 , n31102 , n28583 );
and ( n43999 , n26189 , n28591 );
or ( n44000 , n43998 , n43999 );
and ( n44001 , n44000 , n30269 );
and ( n44002 , n31130 , n28583 );
and ( n44003 , n26189 , n28591 );
or ( n44004 , n44002 , n44003 );
and ( n44005 , n44004 , n30982 );
and ( n44006 , n29475 , n28583 );
and ( n44007 , n26189 , n28591 );
or ( n44008 , n44006 , n44007 );
and ( n44009 , n44008 , n30989 );
and ( n44010 , n26187 , n30991 );
and ( n44011 , n31168 , n28583 );
and ( n44012 , n26189 , n28591 );
or ( n44013 , n44011 , n44012 );
and ( n44014 , n44013 , n31002 );
or ( n44015 , n43993 , n43997 , n44001 , n44005 , n44009 , n44010 , n44014 );
and ( n44016 , n43992 , n44015 );
and ( n44017 , n26189 , n24800 );
or ( n44018 , n44016 , n44017 );
and ( n44019 , n44018 , n31008 );
and ( n44020 , n26189 , n10618 );
or ( n44021 , n44019 , n44020 );
buf ( n44022 , n44021 );
buf ( n44023 , n44022 );
buf ( n44024 , n10615 );
buf ( n44025 , n10615 );
buf ( n44026 , n10613 );
buf ( n44027 , n10613 );
buf ( n44028 , n10613 );
buf ( n44029 , n10615 );
buf ( n44030 , n10613 );
buf ( n44031 , n10613 );
buf ( n44032 , n10615 );
and ( n44033 , n16809 , n23924 );
and ( n44034 , n22173 , n23926 );
or ( n44035 , n44033 , n44034 );
buf ( n44036 , n44035 );
buf ( n44037 , n44036 );
not ( n44038 , n34804 );
and ( n44039 , n44038 , n26467 );
and ( n44040 , n14725 , n34804 );
or ( n44041 , n44039 , n44040 );
and ( n44042 , n44041 , n31008 );
and ( n44043 , n14725 , n10618 );
or ( n44044 , n44042 , n44043 );
buf ( n44045 , n44044 );
buf ( n44046 , n44045 );
not ( n44047 , n34821 );
not ( n44048 , n13916 );
and ( n44049 , n44048 , n13804 );
xor ( n44050 , n13805 , n13860 );
and ( n44051 , n44050 , n13916 );
or ( n44052 , n44049 , n44051 );
buf ( n44053 , n44052 );
and ( n44054 , n44053 , n14137 );
and ( n44055 , n44053 , n14143 );
not ( n44056 , n14139 );
and ( n44057 , n44056 , n35753 );
not ( n44058 , n36245 );
and ( n44059 , n44058 , n35765 );
xor ( n44060 , n36249 , n36261 );
and ( n44061 , n44060 , n36245 );
or ( n44062 , n44059 , n44061 );
buf ( n44063 , n44062 );
and ( n44064 , n44063 , n14139 );
or ( n44065 , n44057 , n44064 );
and ( n44066 , n44065 , n14140 );
and ( n44067 , n35753 , n14141 );
or ( n44068 , n44054 , n44055 , n44066 , n44067 );
and ( n44069 , n44068 , n36347 );
and ( n44070 , n13423 , n39408 );
or ( n44071 , n44069 , n44070 );
and ( n44072 , n44071 , n14562 );
not ( n44073 , n37048 );
and ( n44074 , n44073 , n36653 );
xor ( n44075 , n37052 , n37064 );
and ( n44076 , n44075 , n37048 );
or ( n44077 , n44074 , n44076 );
buf ( n44078 , n44077 );
and ( n44079 , n44078 , n36348 );
and ( n44080 , n13423 , n39427 );
or ( n44081 , n44079 , n44080 );
and ( n44082 , n44081 , n14586 );
not ( n44083 , n37801 );
and ( n44084 , n44083 , n37406 );
xor ( n44085 , n37805 , n37817 );
and ( n44086 , n44085 , n37801 );
or ( n44087 , n44084 , n44086 );
buf ( n44088 , n44087 );
and ( n44089 , n44088 , n36347 );
and ( n44090 , n13423 , n39446 );
or ( n44091 , n44089 , n44090 );
and ( n44092 , n44091 , n14584 );
and ( n44093 , n44078 , n36348 );
and ( n44094 , n13423 , n39453 );
or ( n44095 , n44093 , n44094 );
and ( n44096 , n44095 , n37835 );
and ( n44097 , n44088 , n36348 );
and ( n44098 , n13423 , n39453 );
or ( n44099 , n44097 , n44098 );
and ( n44100 , n44099 , n37841 );
and ( n44101 , n15735 , n36348 );
and ( n44102 , n13423 , n39453 );
or ( n44103 , n44101 , n44102 );
and ( n44104 , n44103 , n37847 );
and ( n44105 , n13423 , n37849 );
or ( n44106 , n44072 , n44082 , n44092 , n44096 , n44100 , n44104 , n44105 );
and ( n44107 , n44047 , n44106 );
and ( n44108 , n13423 , n34821 );
or ( n44109 , n44107 , n44108 );
and ( n44110 , n44109 , n16574 );
and ( n44111 , n13423 , n16576 );
or ( n44112 , n44110 , n44111 );
buf ( n44113 , n44112 );
buf ( n44114 , n44113 );
not ( n44115 , n34821 );
and ( n44116 , n13443 , n14592 );
and ( n44117 , n43142 , n36350 );
and ( n44118 , n13443 , n43691 );
or ( n44119 , n44117 , n44118 );
and ( n44120 , n44119 , n14562 );
and ( n44121 , n43152 , n36350 );
and ( n44122 , n13443 , n43703 );
or ( n44123 , n44121 , n44122 );
and ( n44124 , n44123 , n14586 );
and ( n44125 , n43162 , n36345 );
and ( n44126 , n13443 , n43715 );
or ( n44127 , n44125 , n44126 );
and ( n44128 , n44127 , n14584 );
and ( n44129 , n43152 , n36345 );
and ( n44130 , n13443 , n43721 );
or ( n44131 , n44129 , n44130 );
and ( n44132 , n44131 , n37835 );
and ( n44133 , n43162 , n36345 );
and ( n44134 , n13443 , n43721 );
or ( n44135 , n44133 , n44134 );
and ( n44136 , n44135 , n37841 );
and ( n44137 , n15779 , n14564 );
and ( n44138 , n15779 , n36345 );
and ( n44139 , n13443 , n43721 );
or ( n44140 , n44138 , n44139 );
and ( n44141 , n44140 , n37847 );
or ( n44142 , n44116 , n44120 , n44124 , n44128 , n44132 , n44136 , n44137 , n44141 );
and ( n44143 , n44115 , n44142 );
and ( n44144 , n13443 , n34821 );
or ( n44145 , n44143 , n44144 );
and ( n44146 , n44145 , n16574 );
and ( n44147 , n12321 , n16576 );
or ( n44148 , n44146 , n44147 );
buf ( n44149 , n44148 );
buf ( n44150 , n44149 );
buf ( n44151 , n10613 );
buf ( n44152 , n10613 );
not ( n44153 , n34821 );
and ( n44154 , n13472 , n14592 );
not ( n44155 , n13916 );
and ( n44156 , n44155 , n13848 );
xor ( n44157 , n13849 , n13856 );
and ( n44158 , n44157 , n13916 );
or ( n44159 , n44156 , n44158 );
buf ( n44160 , n44159 );
and ( n44161 , n44160 , n14137 );
and ( n44162 , n44160 , n14143 );
not ( n44163 , n14139 );
and ( n44164 , n44163 , n35665 );
not ( n44165 , n36245 );
and ( n44166 , n44165 , n35677 );
xor ( n44167 , n36253 , n36257 );
and ( n44168 , n44167 , n36245 );
or ( n44169 , n44166 , n44168 );
buf ( n44170 , n44169 );
and ( n44171 , n44170 , n14139 );
or ( n44172 , n44164 , n44171 );
and ( n44173 , n44172 , n14140 );
and ( n44174 , n35665 , n14141 );
or ( n44175 , n44161 , n44162 , n44173 , n44174 );
and ( n44176 , n44175 , n36350 );
and ( n44177 , n13472 , n43691 );
or ( n44178 , n44176 , n44177 );
and ( n44179 , n44178 , n14562 );
not ( n44180 , n37048 );
and ( n44181 , n44180 , n36585 );
xor ( n44182 , n37056 , n37060 );
and ( n44183 , n44182 , n37048 );
or ( n44184 , n44181 , n44183 );
buf ( n44185 , n44184 );
and ( n44186 , n44185 , n36350 );
and ( n44187 , n13472 , n43703 );
or ( n44188 , n44186 , n44187 );
and ( n44189 , n44188 , n14586 );
not ( n44190 , n37801 );
and ( n44191 , n44190 , n37338 );
xor ( n44192 , n37809 , n37813 );
and ( n44193 , n44192 , n37801 );
or ( n44194 , n44191 , n44193 );
buf ( n44195 , n44194 );
and ( n44196 , n44195 , n36345 );
and ( n44197 , n13472 , n43715 );
or ( n44198 , n44196 , n44197 );
and ( n44199 , n44198 , n14584 );
and ( n44200 , n44185 , n36345 );
and ( n44201 , n13472 , n43721 );
or ( n44202 , n44200 , n44201 );
and ( n44203 , n44202 , n37835 );
and ( n44204 , n44195 , n36345 );
and ( n44205 , n13472 , n43721 );
or ( n44206 , n44204 , n44205 );
and ( n44207 , n44206 , n37841 );
and ( n44208 , n15823 , n14564 );
and ( n44209 , n15823 , n36345 );
and ( n44210 , n13472 , n43721 );
or ( n44211 , n44209 , n44210 );
and ( n44212 , n44211 , n37847 );
or ( n44213 , n44154 , n44179 , n44189 , n44199 , n44203 , n44207 , n44208 , n44212 );
and ( n44214 , n44153 , n44213 );
and ( n44215 , n13472 , n34821 );
or ( n44216 , n44214 , n44215 );
and ( n44217 , n44216 , n16574 );
and ( n44218 , n12327 , n16576 );
or ( n44219 , n44217 , n44218 );
buf ( n44220 , n44219 );
buf ( n44221 , n44220 );
buf ( n44222 , n10615 );
not ( n44223 , n17162 );
not ( n44224 , n17450 );
and ( n44225 , n10723 , n37947 );
not ( n44226 , n38425 );
and ( n44227 , n44226 , n38132 );
xor ( n44228 , n38438 , n38442 );
and ( n44229 , n44228 , n38425 );
or ( n44230 , n44227 , n44229 );
buf ( n44231 , n44230 );
and ( n44232 , n44231 , n19745 );
not ( n44233 , n38934 );
and ( n44234 , n44233 , n38641 );
xor ( n44235 , n38947 , n38951 );
and ( n44236 , n44235 , n38934 );
or ( n44237 , n44234 , n44236 );
buf ( n44238 , n44237 );
and ( n44239 , n44238 , n19748 );
and ( n44240 , n22380 , n21253 );
and ( n44241 , n10723 , n21255 );
or ( n44242 , n44232 , n44239 , n44240 , n44241 );
and ( n44243 , n44242 , n38980 );
or ( n44244 , n44225 , n44243 );
and ( n44245 , n44224 , n44244 );
buf ( n44246 , n18504 );
buf ( n44247 , n44246 );
not ( n44248 , n44247 );
buf ( n44249 , n44248 );
buf ( n44250 , n44249 );
not ( n44251 , n44250 );
buf ( n44252 , n18521 );
not ( n44253 , n44252 );
buf ( n44254 , n18540 );
and ( n44255 , n44253 , n44254 );
not ( n44256 , n44254 );
not ( n44257 , n44246 );
xor ( n44258 , n44256 , n44257 );
and ( n44259 , n44258 , n44252 );
or ( n44260 , n44255 , n44259 );
buf ( n44261 , n44260 );
not ( n44262 , n44261 );
buf ( n44263 , n44262 );
buf ( n44264 , n44263 );
not ( n44265 , n44264 );
or ( n44266 , n44251 , n44265 );
not ( n44267 , n44252 );
buf ( n44268 , n18571 );
and ( n44269 , n44267 , n44268 );
not ( n44270 , n44268 );
and ( n44271 , n44256 , n44257 );
xor ( n44272 , n44270 , n44271 );
and ( n44273 , n44272 , n44252 );
or ( n44274 , n44269 , n44273 );
buf ( n44275 , n44274 );
not ( n44276 , n44275 );
buf ( n44277 , n44276 );
buf ( n44278 , n44277 );
not ( n44279 , n44278 );
or ( n44280 , n44266 , n44279 );
not ( n44281 , n44252 );
buf ( n44282 , n18604 );
and ( n44283 , n44281 , n44282 );
not ( n44284 , n44282 );
and ( n44285 , n44270 , n44271 );
xor ( n44286 , n44284 , n44285 );
and ( n44287 , n44286 , n44252 );
or ( n44288 , n44283 , n44287 );
buf ( n44289 , n44288 );
not ( n44290 , n44289 );
buf ( n44291 , n44290 );
buf ( n44292 , n44291 );
not ( n44293 , n44292 );
or ( n44294 , n44280 , n44293 );
not ( n44295 , n44252 );
buf ( n44296 , n18637 );
and ( n44297 , n44295 , n44296 );
not ( n44298 , n44296 );
and ( n44299 , n44284 , n44285 );
xor ( n44300 , n44298 , n44299 );
and ( n44301 , n44300 , n44252 );
or ( n44302 , n44297 , n44301 );
buf ( n44303 , n44302 );
not ( n44304 , n44303 );
buf ( n44305 , n44304 );
buf ( n44306 , n44305 );
not ( n44307 , n44306 );
or ( n44308 , n44294 , n44307 );
not ( n44309 , n44252 );
buf ( n44310 , n18671 );
and ( n44311 , n44309 , n44310 );
not ( n44312 , n44310 );
and ( n44313 , n44298 , n44299 );
xor ( n44314 , n44312 , n44313 );
and ( n44315 , n44314 , n44252 );
or ( n44316 , n44311 , n44315 );
buf ( n44317 , n44316 );
not ( n44318 , n44317 );
buf ( n44319 , n44318 );
buf ( n44320 , n44319 );
not ( n44321 , n44320 );
or ( n44322 , n44308 , n44321 );
not ( n44323 , n44252 );
buf ( n44324 , n18705 );
and ( n44325 , n44323 , n44324 );
not ( n44326 , n44324 );
and ( n44327 , n44312 , n44313 );
xor ( n44328 , n44326 , n44327 );
and ( n44329 , n44328 , n44252 );
or ( n44330 , n44325 , n44329 );
buf ( n44331 , n44330 );
not ( n44332 , n44331 );
buf ( n44333 , n44332 );
buf ( n44334 , n44333 );
not ( n44335 , n44334 );
or ( n44336 , n44322 , n44335 );
not ( n44337 , n44252 );
buf ( n44338 , n18739 );
and ( n44339 , n44337 , n44338 );
not ( n44340 , n44338 );
and ( n44341 , n44326 , n44327 );
xor ( n44342 , n44340 , n44341 );
and ( n44343 , n44342 , n44252 );
or ( n44344 , n44339 , n44343 );
buf ( n44345 , n44344 );
not ( n44346 , n44345 );
buf ( n44347 , n44346 );
buf ( n44348 , n44347 );
not ( n44349 , n44348 );
or ( n44350 , n44336 , n44349 );
not ( n44351 , n44252 );
buf ( n44352 , n18773 );
and ( n44353 , n44351 , n44352 );
not ( n44354 , n44352 );
and ( n44355 , n44340 , n44341 );
xor ( n44356 , n44354 , n44355 );
and ( n44357 , n44356 , n44252 );
or ( n44358 , n44353 , n44357 );
buf ( n44359 , n44358 );
not ( n44360 , n44359 );
buf ( n44361 , n44360 );
buf ( n44362 , n44361 );
not ( n44363 , n44362 );
or ( n44364 , n44350 , n44363 );
not ( n44365 , n44252 );
buf ( n44366 , n18807 );
and ( n44367 , n44365 , n44366 );
not ( n44368 , n44366 );
and ( n44369 , n44354 , n44355 );
xor ( n44370 , n44368 , n44369 );
and ( n44371 , n44370 , n44252 );
or ( n44372 , n44367 , n44371 );
buf ( n44373 , n44372 );
not ( n44374 , n44373 );
buf ( n44375 , n44374 );
buf ( n44376 , n44375 );
not ( n44377 , n44376 );
or ( n44378 , n44364 , n44377 );
not ( n44379 , n44252 );
buf ( n44380 , n18841 );
and ( n44381 , n44379 , n44380 );
not ( n44382 , n44380 );
and ( n44383 , n44368 , n44369 );
xor ( n44384 , n44382 , n44383 );
and ( n44385 , n44384 , n44252 );
or ( n44386 , n44381 , n44385 );
buf ( n44387 , n44386 );
not ( n44388 , n44387 );
buf ( n44389 , n44388 );
buf ( n44390 , n44389 );
not ( n44391 , n44390 );
or ( n44392 , n44378 , n44391 );
not ( n44393 , n44252 );
buf ( n44394 , n18875 );
and ( n44395 , n44393 , n44394 );
not ( n44396 , n44394 );
and ( n44397 , n44382 , n44383 );
xor ( n44398 , n44396 , n44397 );
and ( n44399 , n44398 , n44252 );
or ( n44400 , n44395 , n44399 );
buf ( n44401 , n44400 );
not ( n44402 , n44401 );
buf ( n44403 , n44402 );
buf ( n44404 , n44403 );
not ( n44405 , n44404 );
or ( n44406 , n44392 , n44405 );
not ( n44407 , n44252 );
buf ( n44408 , n18909 );
and ( n44409 , n44407 , n44408 );
not ( n44410 , n44408 );
and ( n44411 , n44396 , n44397 );
xor ( n44412 , n44410 , n44411 );
and ( n44413 , n44412 , n44252 );
or ( n44414 , n44409 , n44413 );
buf ( n44415 , n44414 );
not ( n44416 , n44415 );
buf ( n44417 , n44416 );
buf ( n44418 , n44417 );
not ( n44419 , n44418 );
or ( n44420 , n44406 , n44419 );
not ( n44421 , n44252 );
buf ( n44422 , n18943 );
and ( n44423 , n44421 , n44422 );
not ( n44424 , n44422 );
and ( n44425 , n44410 , n44411 );
xor ( n44426 , n44424 , n44425 );
and ( n44427 , n44426 , n44252 );
or ( n44428 , n44423 , n44427 );
buf ( n44429 , n44428 );
not ( n44430 , n44429 );
buf ( n44431 , n44430 );
buf ( n44432 , n44431 );
not ( n44433 , n44432 );
or ( n44434 , n44420 , n44433 );
not ( n44435 , n44252 );
buf ( n44436 , n18977 );
and ( n44437 , n44435 , n44436 );
not ( n44438 , n44436 );
and ( n44439 , n44424 , n44425 );
xor ( n44440 , n44438 , n44439 );
and ( n44441 , n44440 , n44252 );
or ( n44442 , n44437 , n44441 );
buf ( n44443 , n44442 );
not ( n44444 , n44443 );
buf ( n44445 , n44444 );
buf ( n44446 , n44445 );
not ( n44447 , n44446 );
or ( n44448 , n44434 , n44447 );
not ( n44449 , n44252 );
buf ( n44450 , n19011 );
and ( n44451 , n44449 , n44450 );
not ( n44452 , n44450 );
and ( n44453 , n44438 , n44439 );
xor ( n44454 , n44452 , n44453 );
and ( n44455 , n44454 , n44252 );
or ( n44456 , n44451 , n44455 );
buf ( n44457 , n44456 );
not ( n44458 , n44457 );
buf ( n44459 , n44458 );
buf ( n44460 , n44459 );
not ( n44461 , n44460 );
or ( n44462 , n44448 , n44461 );
not ( n44463 , n44252 );
buf ( n44464 , n19045 );
and ( n44465 , n44463 , n44464 );
not ( n44466 , n44464 );
and ( n44467 , n44452 , n44453 );
xor ( n44468 , n44466 , n44467 );
and ( n44469 , n44468 , n44252 );
or ( n44470 , n44465 , n44469 );
buf ( n44471 , n44470 );
not ( n44472 , n44471 );
buf ( n44473 , n44472 );
buf ( n44474 , n44473 );
not ( n44475 , n44474 );
or ( n44476 , n44462 , n44475 );
not ( n44477 , n44252 );
buf ( n44478 , n19079 );
and ( n44479 , n44477 , n44478 );
not ( n44480 , n44478 );
and ( n44481 , n44466 , n44467 );
xor ( n44482 , n44480 , n44481 );
and ( n44483 , n44482 , n44252 );
or ( n44484 , n44479 , n44483 );
buf ( n44485 , n44484 );
not ( n44486 , n44485 );
buf ( n44487 , n44486 );
buf ( n44488 , n44487 );
not ( n44489 , n44488 );
or ( n44490 , n44476 , n44489 );
not ( n44491 , n44252 );
buf ( n44492 , n19113 );
and ( n44493 , n44491 , n44492 );
not ( n44494 , n44492 );
and ( n44495 , n44480 , n44481 );
xor ( n44496 , n44494 , n44495 );
and ( n44497 , n44496 , n44252 );
or ( n44498 , n44493 , n44497 );
buf ( n44499 , n44498 );
not ( n44500 , n44499 );
buf ( n44501 , n44500 );
buf ( n44502 , n44501 );
not ( n44503 , n44502 );
or ( n44504 , n44490 , n44503 );
not ( n44505 , n44252 );
buf ( n44506 , n19147 );
and ( n44507 , n44505 , n44506 );
not ( n44508 , n44506 );
and ( n44509 , n44494 , n44495 );
xor ( n44510 , n44508 , n44509 );
and ( n44511 , n44510 , n44252 );
or ( n44512 , n44507 , n44511 );
buf ( n44513 , n44512 );
not ( n44514 , n44513 );
buf ( n44515 , n44514 );
buf ( n44516 , n44515 );
not ( n44517 , n44516 );
or ( n44518 , n44504 , n44517 );
buf ( n44519 , n44518 );
buf ( n44520 , n44519 );
and ( n44521 , n44520 , n44252 );
not ( n44522 , n44521 );
and ( n44523 , n44522 , n44251 );
xor ( n44524 , n44251 , n44252 );
xor ( n44525 , n44524 , n44252 );
and ( n44526 , n44525 , n44521 );
or ( n44527 , n44523 , n44526 );
buf ( n44528 , n44527 );
buf ( n44529 , n44528 );
buf ( n44530 , n21637 );
not ( n44531 , n44530 );
buf ( n44532 , n44531 );
not ( n44533 , n44532 );
buf ( n44534 , n44533 );
buf ( n44535 , n44534 );
buf ( n44536 , n44535 );
xor ( n44537 , n44529 , n44536 );
buf ( n44538 , n44537 );
and ( n44539 , n44538 , n19745 );
buf ( n44540 , n18508 );
buf ( n44541 , n44540 );
not ( n44542 , n44541 );
buf ( n44543 , n44542 );
buf ( n44544 , n44543 );
not ( n44545 , n44544 );
buf ( n44546 , n18523 );
not ( n44547 , n44546 );
buf ( n44548 , n18542 );
and ( n44549 , n44547 , n44548 );
not ( n44550 , n44548 );
not ( n44551 , n44540 );
xor ( n44552 , n44550 , n44551 );
and ( n44553 , n44552 , n44546 );
or ( n44554 , n44549 , n44553 );
buf ( n44555 , n44554 );
not ( n44556 , n44555 );
buf ( n44557 , n44556 );
buf ( n44558 , n44557 );
not ( n44559 , n44558 );
or ( n44560 , n44545 , n44559 );
not ( n44561 , n44546 );
buf ( n44562 , n18573 );
and ( n44563 , n44561 , n44562 );
not ( n44564 , n44562 );
and ( n44565 , n44550 , n44551 );
xor ( n44566 , n44564 , n44565 );
and ( n44567 , n44566 , n44546 );
or ( n44568 , n44563 , n44567 );
buf ( n44569 , n44568 );
not ( n44570 , n44569 );
buf ( n44571 , n44570 );
buf ( n44572 , n44571 );
not ( n44573 , n44572 );
or ( n44574 , n44560 , n44573 );
not ( n44575 , n44546 );
buf ( n44576 , n18606 );
and ( n44577 , n44575 , n44576 );
not ( n44578 , n44576 );
and ( n44579 , n44564 , n44565 );
xor ( n44580 , n44578 , n44579 );
and ( n44581 , n44580 , n44546 );
or ( n44582 , n44577 , n44581 );
buf ( n44583 , n44582 );
not ( n44584 , n44583 );
buf ( n44585 , n44584 );
buf ( n44586 , n44585 );
not ( n44587 , n44586 );
or ( n44588 , n44574 , n44587 );
not ( n44589 , n44546 );
buf ( n44590 , n18639 );
and ( n44591 , n44589 , n44590 );
not ( n44592 , n44590 );
and ( n44593 , n44578 , n44579 );
xor ( n44594 , n44592 , n44593 );
and ( n44595 , n44594 , n44546 );
or ( n44596 , n44591 , n44595 );
buf ( n44597 , n44596 );
not ( n44598 , n44597 );
buf ( n44599 , n44598 );
buf ( n44600 , n44599 );
not ( n44601 , n44600 );
or ( n44602 , n44588 , n44601 );
not ( n44603 , n44546 );
buf ( n44604 , n18673 );
and ( n44605 , n44603 , n44604 );
not ( n44606 , n44604 );
and ( n44607 , n44592 , n44593 );
xor ( n44608 , n44606 , n44607 );
and ( n44609 , n44608 , n44546 );
or ( n44610 , n44605 , n44609 );
buf ( n44611 , n44610 );
not ( n44612 , n44611 );
buf ( n44613 , n44612 );
buf ( n44614 , n44613 );
not ( n44615 , n44614 );
or ( n44616 , n44602 , n44615 );
not ( n44617 , n44546 );
buf ( n44618 , n18707 );
and ( n44619 , n44617 , n44618 );
not ( n44620 , n44618 );
and ( n44621 , n44606 , n44607 );
xor ( n44622 , n44620 , n44621 );
and ( n44623 , n44622 , n44546 );
or ( n44624 , n44619 , n44623 );
buf ( n44625 , n44624 );
not ( n44626 , n44625 );
buf ( n44627 , n44626 );
buf ( n44628 , n44627 );
not ( n44629 , n44628 );
or ( n44630 , n44616 , n44629 );
not ( n44631 , n44546 );
buf ( n44632 , n18741 );
and ( n44633 , n44631 , n44632 );
not ( n44634 , n44632 );
and ( n44635 , n44620 , n44621 );
xor ( n44636 , n44634 , n44635 );
and ( n44637 , n44636 , n44546 );
or ( n44638 , n44633 , n44637 );
buf ( n44639 , n44638 );
not ( n44640 , n44639 );
buf ( n44641 , n44640 );
buf ( n44642 , n44641 );
not ( n44643 , n44642 );
or ( n44644 , n44630 , n44643 );
not ( n44645 , n44546 );
buf ( n44646 , n18775 );
and ( n44647 , n44645 , n44646 );
not ( n44648 , n44646 );
and ( n44649 , n44634 , n44635 );
xor ( n44650 , n44648 , n44649 );
and ( n44651 , n44650 , n44546 );
or ( n44652 , n44647 , n44651 );
buf ( n44653 , n44652 );
not ( n44654 , n44653 );
buf ( n44655 , n44654 );
buf ( n44656 , n44655 );
not ( n44657 , n44656 );
or ( n44658 , n44644 , n44657 );
not ( n44659 , n44546 );
buf ( n44660 , n18809 );
and ( n44661 , n44659 , n44660 );
not ( n44662 , n44660 );
and ( n44663 , n44648 , n44649 );
xor ( n44664 , n44662 , n44663 );
and ( n44665 , n44664 , n44546 );
or ( n44666 , n44661 , n44665 );
buf ( n44667 , n44666 );
not ( n44668 , n44667 );
buf ( n44669 , n44668 );
buf ( n44670 , n44669 );
not ( n44671 , n44670 );
or ( n44672 , n44658 , n44671 );
not ( n44673 , n44546 );
buf ( n44674 , n18843 );
and ( n44675 , n44673 , n44674 );
not ( n44676 , n44674 );
and ( n44677 , n44662 , n44663 );
xor ( n44678 , n44676 , n44677 );
and ( n44679 , n44678 , n44546 );
or ( n44680 , n44675 , n44679 );
buf ( n44681 , n44680 );
not ( n44682 , n44681 );
buf ( n44683 , n44682 );
buf ( n44684 , n44683 );
not ( n44685 , n44684 );
or ( n44686 , n44672 , n44685 );
not ( n44687 , n44546 );
buf ( n44688 , n18877 );
and ( n44689 , n44687 , n44688 );
not ( n44690 , n44688 );
and ( n44691 , n44676 , n44677 );
xor ( n44692 , n44690 , n44691 );
and ( n44693 , n44692 , n44546 );
or ( n44694 , n44689 , n44693 );
buf ( n44695 , n44694 );
not ( n44696 , n44695 );
buf ( n44697 , n44696 );
buf ( n44698 , n44697 );
not ( n44699 , n44698 );
or ( n44700 , n44686 , n44699 );
not ( n44701 , n44546 );
buf ( n44702 , n18911 );
and ( n44703 , n44701 , n44702 );
not ( n44704 , n44702 );
and ( n44705 , n44690 , n44691 );
xor ( n44706 , n44704 , n44705 );
and ( n44707 , n44706 , n44546 );
or ( n44708 , n44703 , n44707 );
buf ( n44709 , n44708 );
not ( n44710 , n44709 );
buf ( n44711 , n44710 );
buf ( n44712 , n44711 );
not ( n44713 , n44712 );
or ( n44714 , n44700 , n44713 );
not ( n44715 , n44546 );
buf ( n44716 , n18945 );
and ( n44717 , n44715 , n44716 );
not ( n44718 , n44716 );
and ( n44719 , n44704 , n44705 );
xor ( n44720 , n44718 , n44719 );
and ( n44721 , n44720 , n44546 );
or ( n44722 , n44717 , n44721 );
buf ( n44723 , n44722 );
not ( n44724 , n44723 );
buf ( n44725 , n44724 );
buf ( n44726 , n44725 );
not ( n44727 , n44726 );
or ( n44728 , n44714 , n44727 );
not ( n44729 , n44546 );
buf ( n44730 , n18979 );
and ( n44731 , n44729 , n44730 );
not ( n44732 , n44730 );
and ( n44733 , n44718 , n44719 );
xor ( n44734 , n44732 , n44733 );
and ( n44735 , n44734 , n44546 );
or ( n44736 , n44731 , n44735 );
buf ( n44737 , n44736 );
not ( n44738 , n44737 );
buf ( n44739 , n44738 );
buf ( n44740 , n44739 );
not ( n44741 , n44740 );
or ( n44742 , n44728 , n44741 );
not ( n44743 , n44546 );
buf ( n44744 , n19013 );
and ( n44745 , n44743 , n44744 );
not ( n44746 , n44744 );
and ( n44747 , n44732 , n44733 );
xor ( n44748 , n44746 , n44747 );
and ( n44749 , n44748 , n44546 );
or ( n44750 , n44745 , n44749 );
buf ( n44751 , n44750 );
not ( n44752 , n44751 );
buf ( n44753 , n44752 );
buf ( n44754 , n44753 );
not ( n44755 , n44754 );
or ( n44756 , n44742 , n44755 );
not ( n44757 , n44546 );
buf ( n44758 , n19047 );
and ( n44759 , n44757 , n44758 );
not ( n44760 , n44758 );
and ( n44761 , n44746 , n44747 );
xor ( n44762 , n44760 , n44761 );
and ( n44763 , n44762 , n44546 );
or ( n44764 , n44759 , n44763 );
buf ( n44765 , n44764 );
not ( n44766 , n44765 );
buf ( n44767 , n44766 );
buf ( n44768 , n44767 );
not ( n44769 , n44768 );
or ( n44770 , n44756 , n44769 );
not ( n44771 , n44546 );
buf ( n44772 , n19081 );
and ( n44773 , n44771 , n44772 );
not ( n44774 , n44772 );
and ( n44775 , n44760 , n44761 );
xor ( n44776 , n44774 , n44775 );
and ( n44777 , n44776 , n44546 );
or ( n44778 , n44773 , n44777 );
buf ( n44779 , n44778 );
not ( n44780 , n44779 );
buf ( n44781 , n44780 );
buf ( n44782 , n44781 );
not ( n44783 , n44782 );
or ( n44784 , n44770 , n44783 );
not ( n44785 , n44546 );
buf ( n44786 , n19115 );
and ( n44787 , n44785 , n44786 );
not ( n44788 , n44786 );
and ( n44789 , n44774 , n44775 );
xor ( n44790 , n44788 , n44789 );
and ( n44791 , n44790 , n44546 );
or ( n44792 , n44787 , n44791 );
buf ( n44793 , n44792 );
not ( n44794 , n44793 );
buf ( n44795 , n44794 );
buf ( n44796 , n44795 );
not ( n44797 , n44796 );
or ( n44798 , n44784 , n44797 );
not ( n44799 , n44546 );
buf ( n44800 , n19149 );
and ( n44801 , n44799 , n44800 );
not ( n44802 , n44800 );
and ( n44803 , n44788 , n44789 );
xor ( n44804 , n44802 , n44803 );
and ( n44805 , n44804 , n44546 );
or ( n44806 , n44801 , n44805 );
buf ( n44807 , n44806 );
not ( n44808 , n44807 );
buf ( n44809 , n44808 );
buf ( n44810 , n44809 );
not ( n44811 , n44810 );
or ( n44812 , n44798 , n44811 );
buf ( n44813 , n44812 );
buf ( n44814 , n44813 );
and ( n44815 , n44814 , n44546 );
not ( n44816 , n44815 );
and ( n44817 , n44816 , n44545 );
xor ( n44818 , n44545 , n44546 );
xor ( n44819 , n44818 , n44546 );
and ( n44820 , n44819 , n44815 );
or ( n44821 , n44817 , n44820 );
buf ( n44822 , n44821 );
buf ( n44823 , n44822 );
buf ( n44824 , n44535 );
xor ( n44825 , n44823 , n44824 );
buf ( n44826 , n44825 );
and ( n44827 , n44826 , n19748 );
or ( n44828 , n21255 , n21253 );
and ( n44829 , n21637 , n44828 );
or ( n44830 , n44539 , n44827 , n44829 );
buf ( n44831 , n44830 );
buf ( n44832 , n44831 );
not ( n44833 , n44832 );
buf ( n44834 , n44833 );
buf ( n44835 , n44834 );
not ( n44836 , n44835 );
and ( n44837 , C1 , n44836 );
or ( n44838 , n44837 , C0 );
buf ( n44839 , n44838 );
buf ( n44840 , n44839 );
buf ( n44841 , n44840 );
and ( n44842 , n44841 , n17450 );
or ( n44843 , n44245 , n44842 );
and ( n44844 , n44223 , n44843 );
and ( n44845 , n44242 , n17162 );
or ( n44846 , n44844 , n44845 );
and ( n44847 , n44846 , n23924 );
not ( n44848 , n39264 );
and ( n44849 , n44848 , n39022 );
xor ( n44850 , n39277 , n39281 );
and ( n44851 , n44850 , n39264 );
or ( n44852 , n44849 , n44851 );
buf ( n44853 , n44852 );
and ( n44854 , n44853 , n23926 );
or ( n44855 , n44847 , n44854 );
buf ( n44856 , n44855 );
buf ( n44857 , n44856 );
buf ( n44858 , n10613 );
buf ( n44859 , n10613 );
buf ( n44860 , n10615 );
buf ( n44861 , n10615 );
buf ( n44862 , n10615 );
not ( n44863 , n17451 );
and ( n44864 , n34754 , n21334 );
and ( n44865 , n18544 , n34492 );
or ( n44866 , n44864 , n44865 );
and ( n44867 , n44866 , n21341 );
and ( n44868 , n34767 , n21334 );
and ( n44869 , n18544 , n34492 );
or ( n44870 , n44868 , n44869 );
and ( n44871 , n44870 , n23064 );
and ( n44872 , n34777 , n21334 );
and ( n44873 , n18544 , n34492 );
or ( n44874 , n44872 , n44873 );
and ( n44875 , n44874 , n23825 );
and ( n44876 , n22402 , n21334 );
and ( n44877 , n18544 , n34492 );
or ( n44878 , n44876 , n44877 );
and ( n44879 , n44878 , n23832 );
and ( n44880 , n34787 , n21334 );
and ( n44881 , n18544 , n34492 );
or ( n44882 , n44880 , n44881 );
and ( n44883 , n44882 , n23917 );
and ( n44884 , n18544 , n34526 );
or ( n44885 , n44867 , n44871 , n44875 , n44879 , n44883 , n44884 );
and ( n44886 , n44863 , n44885 );
and ( n44887 , n18544 , n17451 );
or ( n44888 , n44886 , n44887 );
and ( n44889 , n44888 , n23924 );
and ( n44890 , n18544 , n23926 );
or ( n44891 , n44889 , n44890 );
buf ( n44892 , n44891 );
buf ( n44893 , n44892 );
buf ( n44894 , n10613 );
not ( n44895 , n34821 );
not ( n44896 , n13916 );
and ( n44897 , n44896 , n13771 );
xor ( n44898 , n13772 , n13863 );
and ( n44899 , n44898 , n13916 );
or ( n44900 , n44897 , n44899 );
buf ( n44901 , n44900 );
and ( n44902 , n44901 , n14137 );
and ( n44903 , n44901 , n14143 );
not ( n44904 , n14139 );
and ( n44905 , n44904 , n35811 );
not ( n44906 , n36245 );
and ( n44907 , n44906 , n35823 );
xor ( n44908 , n39391 , n39394 );
and ( n44909 , n44908 , n36245 );
or ( n44910 , n44907 , n44909 );
buf ( n44911 , n44910 );
and ( n44912 , n44911 , n14139 );
or ( n44913 , n44905 , n44912 );
and ( n44914 , n44913 , n14140 );
and ( n44915 , n35811 , n14141 );
or ( n44916 , n44902 , n44903 , n44914 , n44915 );
and ( n44917 , n44916 , n36345 );
and ( n44918 , n13389 , n36352 );
or ( n44919 , n44917 , n44918 );
and ( n44920 , n44919 , n14562 );
not ( n44921 , n37048 );
and ( n44922 , n44921 , n36704 );
xor ( n44923 , n39415 , n39418 );
and ( n44924 , n44923 , n37048 );
or ( n44925 , n44922 , n44924 );
buf ( n44926 , n44925 );
and ( n44927 , n44926 , n36345 );
and ( n44928 , n13389 , n37073 );
or ( n44929 , n44927 , n44928 );
and ( n44930 , n44929 , n14586 );
not ( n44931 , n37801 );
and ( n44932 , n44931 , n37457 );
xor ( n44933 , n39434 , n39437 );
and ( n44934 , n44933 , n37801 );
or ( n44935 , n44932 , n44934 );
buf ( n44936 , n44935 );
and ( n44937 , n44936 , n36350 );
and ( n44938 , n13389 , n37825 );
or ( n44939 , n44937 , n44938 );
and ( n44940 , n44939 , n14584 );
and ( n44941 , n44926 , n36350 );
and ( n44942 , n13389 , n37831 );
or ( n44943 , n44941 , n44942 );
and ( n44944 , n44943 , n37835 );
and ( n44945 , n44936 , n36350 );
and ( n44946 , n13389 , n37831 );
or ( n44947 , n44945 , n44946 );
and ( n44948 , n44947 , n37841 );
and ( n44949 , n15669 , n36350 );
and ( n44950 , n13389 , n37831 );
or ( n44951 , n44949 , n44950 );
and ( n44952 , n44951 , n37847 );
and ( n44953 , n13389 , n37849 );
or ( n44954 , n44920 , n44930 , n44940 , n44944 , n44948 , n44952 , n44953 );
and ( n44955 , n44895 , n44954 );
and ( n44956 , n13389 , n34821 );
or ( n44957 , n44955 , n44956 );
and ( n44958 , n44957 , n16574 );
and ( n44959 , n13389 , n16576 );
or ( n44960 , n44958 , n44959 );
buf ( n44961 , n44960 );
buf ( n44962 , n44961 );
buf ( n44963 , n10615 );
buf ( n44964 , n10615 );
buf ( n44965 , n10615 );
buf ( n44966 , n10613 );
buf ( n44967 , n10613 );
not ( n44968 , n24800 );
not ( n44969 , n26823 );
and ( n44970 , n44969 , n26241 );
xor ( n44971 , n34624 , n34627 );
and ( n44972 , n44971 , n26823 );
or ( n44973 , n44970 , n44972 );
buf ( n44974 , n44973 );
and ( n44975 , n44974 , n27046 );
and ( n44976 , n44974 , n27049 );
not ( n44977 , n27051 );
and ( n44978 , n44977 , n28126 );
not ( n44979 , n28494 );
and ( n44980 , n44979 , n28138 );
xor ( n44981 , n34642 , n34645 );
and ( n44982 , n44981 , n28494 );
or ( n44983 , n44980 , n44982 );
buf ( n44984 , n44983 );
and ( n44985 , n44984 , n27051 );
or ( n44986 , n44978 , n44985 );
and ( n44987 , n44986 , n28506 );
and ( n44988 , n28126 , n28508 );
or ( n44989 , n44975 , n44976 , n44987 , n44988 );
and ( n44990 , n44989 , n28586 );
and ( n44991 , n26259 , n34573 );
or ( n44992 , n44990 , n44991 );
and ( n44993 , n44992 , n28594 );
not ( n44994 , n30249 );
and ( n44995 , n44994 , n29956 );
xor ( n44996 , n34665 , n34668 );
and ( n44997 , n44996 , n30249 );
or ( n44998 , n44995 , n44997 );
buf ( n44999 , n44998 );
and ( n45000 , n44999 , n28586 );
and ( n45001 , n26259 , n34573 );
or ( n45002 , n45000 , n45001 );
and ( n45003 , n45002 , n30269 );
not ( n45004 , n30963 );
and ( n45005 , n45004 , n30670 );
xor ( n45006 , n34683 , n34686 );
and ( n45007 , n45006 , n30963 );
or ( n45008 , n45005 , n45007 );
buf ( n45009 , n45008 );
and ( n45010 , n45009 , n28586 );
and ( n45011 , n26259 , n34573 );
or ( n45012 , n45010 , n45011 );
and ( n45013 , n45012 , n30982 );
and ( n45014 , n29435 , n28586 );
and ( n45015 , n26259 , n34573 );
or ( n45016 , n45014 , n45015 );
and ( n45017 , n45016 , n30989 );
xor ( n45018 , n34706 , n34710 );
buf ( n45019 , n45018 );
and ( n45020 , n45019 , n28586 );
and ( n45021 , n26259 , n34573 );
or ( n45022 , n45020 , n45021 );
and ( n45023 , n45022 , n31002 );
and ( n45024 , n26259 , n34607 );
or ( n45025 , n44993 , n45003 , n45013 , n45017 , n45023 , n45024 );
and ( n45026 , n44968 , n45025 );
and ( n45027 , n26259 , n24800 );
or ( n45028 , n45026 , n45027 );
and ( n45029 , n45028 , n31008 );
and ( n45030 , n26259 , n10618 );
or ( n45031 , n45029 , n45030 );
buf ( n45032 , n45031 );
buf ( n45033 , n45032 );
not ( n45034 , n24800 );
and ( n45035 , n26425 , n25222 );
and ( n45036 , n39662 , n28589 );
and ( n45037 , n26425 , n31075 );
or ( n45038 , n45036 , n45037 );
and ( n45039 , n45038 , n28594 );
and ( n45040 , n39678 , n28589 );
and ( n45041 , n26425 , n31075 );
or ( n45042 , n45040 , n45041 );
and ( n45043 , n45042 , n30269 );
and ( n45044 , n39694 , n28589 );
and ( n45045 , n26425 , n31075 );
or ( n45046 , n45044 , n45045 );
and ( n45047 , n45046 , n30982 );
and ( n45048 , n29335 , n28589 );
and ( n45049 , n26425 , n31075 );
or ( n45050 , n45048 , n45049 );
and ( n45051 , n45050 , n30989 );
and ( n45052 , n29335 , n30991 );
and ( n45053 , n39713 , n28589 );
and ( n45054 , n26425 , n31075 );
or ( n45055 , n45053 , n45054 );
and ( n45056 , n45055 , n31002 );
or ( n45057 , n45035 , n45039 , n45043 , n45047 , n45051 , n45052 , n45056 );
and ( n45058 , n45034 , n45057 );
and ( n45059 , n26425 , n24800 );
or ( n45060 , n45058 , n45059 );
and ( n45061 , n45060 , n31008 );
and ( n45062 , n25474 , n10618 );
or ( n45063 , n45061 , n45062 );
buf ( n45064 , n45063 );
buf ( n45065 , n45064 );
not ( n45066 , n24800 );
and ( n45067 , n26291 , n25222 );
not ( n45068 , n26823 );
and ( n45069 , n45068 , n26275 );
xor ( n45070 , n34623 , n34628 );
and ( n45071 , n45070 , n26823 );
or ( n45072 , n45069 , n45071 );
buf ( n45073 , n45072 );
and ( n45074 , n45073 , n27046 );
and ( n45075 , n45073 , n27049 );
not ( n45076 , n27051 );
and ( n45077 , n45076 , n28148 );
not ( n45078 , n28494 );
and ( n45079 , n45078 , n28160 );
xor ( n45080 , n34641 , n34646 );
and ( n45081 , n45080 , n28494 );
or ( n45082 , n45079 , n45081 );
buf ( n45083 , n45082 );
and ( n45084 , n45083 , n27051 );
or ( n45085 , n45077 , n45084 );
and ( n45086 , n45085 , n28506 );
and ( n45087 , n28148 , n28508 );
or ( n45088 , n45074 , n45075 , n45086 , n45087 );
and ( n45089 , n45088 , n28583 );
and ( n45090 , n26291 , n28591 );
or ( n45091 , n45089 , n45090 );
and ( n45092 , n45091 , n28594 );
not ( n45093 , n30249 );
and ( n45094 , n45093 , n29973 );
xor ( n45095 , n34664 , n34669 );
and ( n45096 , n45095 , n30249 );
or ( n45097 , n45094 , n45096 );
buf ( n45098 , n45097 );
and ( n45099 , n45098 , n28583 );
and ( n45100 , n26291 , n28591 );
or ( n45101 , n45099 , n45100 );
and ( n45102 , n45101 , n30269 );
not ( n45103 , n30963 );
and ( n45104 , n45103 , n30687 );
xor ( n45105 , n34682 , n34687 );
and ( n45106 , n45105 , n30963 );
or ( n45107 , n45104 , n45106 );
buf ( n45108 , n45107 );
and ( n45109 , n45108 , n28583 );
and ( n45110 , n26291 , n28591 );
or ( n45111 , n45109 , n45110 );
and ( n45112 , n45111 , n30982 );
and ( n45113 , n29415 , n28583 );
and ( n45114 , n26291 , n28591 );
or ( n45115 , n45113 , n45114 );
and ( n45116 , n45115 , n30989 );
and ( n45117 , n26289 , n30991 );
xor ( n45118 , n34704 , n34711 );
buf ( n45119 , n45118 );
and ( n45120 , n45119 , n28583 );
and ( n45121 , n26291 , n28591 );
or ( n45122 , n45120 , n45121 );
and ( n45123 , n45122 , n31002 );
or ( n45124 , n45067 , n45092 , n45102 , n45112 , n45116 , n45117 , n45123 );
and ( n45125 , n45066 , n45124 );
and ( n45126 , n26291 , n24800 );
or ( n45127 , n45125 , n45126 );
and ( n45128 , n45127 , n31008 );
and ( n45129 , n26291 , n10618 );
or ( n45130 , n45128 , n45129 );
buf ( n45131 , n45130 );
buf ( n45132 , n45131 );
buf ( n45133 , n10615 );
buf ( n45134 , n10613 );
buf ( n45135 , n10615 );
buf ( n45136 , n10613 );
buf ( n45137 , n10613 );
not ( n45138 , n34821 );
not ( n45139 , n13916 );
and ( n45140 , n45139 , n13661 );
xor ( n45141 , n13662 , n13873 );
and ( n45142 , n45141 , n13916 );
or ( n45143 , n45140 , n45142 );
buf ( n45144 , n45143 );
and ( n45145 , n45144 , n14137 );
and ( n45146 , n45144 , n14143 );
not ( n45147 , n14139 );
and ( n45148 , n45147 , n36031 );
not ( n45149 , n36245 );
and ( n45150 , n45149 , n36043 );
xor ( n45151 , n36043 , n35634 );
xor ( n45152 , n36021 , n35634 );
xor ( n45153 , n35999 , n35634 );
and ( n45154 , n43029 , n43040 );
and ( n45155 , n45153 , n45154 );
and ( n45156 , n45152 , n45155 );
xor ( n45157 , n45151 , n45156 );
and ( n45158 , n45157 , n36245 );
or ( n45159 , n45150 , n45158 );
buf ( n45160 , n45159 );
and ( n45161 , n45160 , n14139 );
or ( n45162 , n45148 , n45161 );
and ( n45163 , n45162 , n14140 );
and ( n45164 , n36031 , n14141 );
or ( n45165 , n45145 , n45146 , n45163 , n45164 );
and ( n45166 , n45165 , n36347 );
and ( n45167 , n13267 , n39408 );
or ( n45168 , n45166 , n45167 );
and ( n45169 , n45168 , n14562 );
not ( n45170 , n37048 );
and ( n45171 , n45170 , n36874 );
xor ( n45172 , n36874 , n36552 );
xor ( n45173 , n36857 , n36552 );
xor ( n45174 , n36840 , n36552 );
and ( n45175 , n43056 , n43067 );
and ( n45176 , n45174 , n45175 );
and ( n45177 , n45173 , n45176 );
xor ( n45178 , n45172 , n45177 );
and ( n45179 , n45178 , n37048 );
or ( n45180 , n45171 , n45179 );
buf ( n45181 , n45180 );
and ( n45182 , n45181 , n36348 );
and ( n45183 , n13267 , n39427 );
or ( n45184 , n45182 , n45183 );
and ( n45185 , n45184 , n14586 );
not ( n45186 , n37801 );
and ( n45187 , n45186 , n37627 );
xor ( n45188 , n37627 , n37305 );
xor ( n45189 , n37610 , n37305 );
xor ( n45190 , n37593 , n37305 );
and ( n45191 , n43078 , n43089 );
and ( n45192 , n45190 , n45191 );
and ( n45193 , n45189 , n45192 );
xor ( n45194 , n45188 , n45193 );
and ( n45195 , n45194 , n37801 );
or ( n45196 , n45187 , n45195 );
buf ( n45197 , n45196 );
and ( n45198 , n45197 , n36347 );
and ( n45199 , n13267 , n39446 );
or ( n45200 , n45198 , n45199 );
and ( n45201 , n45200 , n14584 );
and ( n45202 , n45181 , n36348 );
and ( n45203 , n13267 , n39453 );
or ( n45204 , n45202 , n45203 );
and ( n45205 , n45204 , n37835 );
and ( n45206 , n45197 , n36348 );
and ( n45207 , n13267 , n39453 );
or ( n45208 , n45206 , n45207 );
and ( n45209 , n45208 , n37841 );
and ( n45210 , n15449 , n36348 );
and ( n45211 , n13267 , n39453 );
or ( n45212 , n45210 , n45211 );
and ( n45213 , n45212 , n37847 );
and ( n45214 , n13267 , n37849 );
or ( n45215 , n45169 , n45185 , n45201 , n45205 , n45209 , n45213 , n45214 );
and ( n45216 , n45138 , n45215 );
and ( n45217 , n13267 , n34821 );
or ( n45218 , n45216 , n45217 );
and ( n45219 , n45218 , n16574 );
and ( n45220 , n13267 , n16576 );
or ( n45221 , n45219 , n45220 );
buf ( n45222 , n45221 );
buf ( n45223 , n45222 );
not ( n45224 , n24800 );
and ( n45225 , n26799 , n25222 );
not ( n45226 , n26823 );
and ( n45227 , n45226 , n26785 );
xor ( n45228 , n26785 , n25877 );
xor ( n45229 , n26751 , n25877 );
xor ( n45230 , n26717 , n25877 );
and ( n45231 , n43390 , n43395 );
and ( n45232 , n45230 , n45231 );
and ( n45233 , n45229 , n45232 );
xor ( n45234 , n45228 , n45233 );
and ( n45235 , n45234 , n26823 );
or ( n45236 , n45227 , n45235 );
buf ( n45237 , n45236 );
and ( n45238 , n45237 , n27046 );
and ( n45239 , n45237 , n27049 );
not ( n45240 , n27051 );
and ( n45241 , n45240 , n28478 );
not ( n45242 , n28494 );
and ( n45243 , n45242 , n28490 );
xor ( n45244 , n28490 , n27883 );
xor ( n45245 , n28468 , n27883 );
xor ( n45246 , n28446 , n27883 );
and ( n45247 , n43406 , n43411 );
and ( n45248 , n45246 , n45247 );
and ( n45249 , n45245 , n45248 );
xor ( n45250 , n45244 , n45249 );
and ( n45251 , n45250 , n28494 );
or ( n45252 , n45243 , n45251 );
buf ( n45253 , n45252 );
and ( n45254 , n45253 , n27051 );
or ( n45255 , n45241 , n45254 );
and ( n45256 , n45255 , n28506 );
and ( n45257 , n28478 , n28508 );
or ( n45258 , n45238 , n45239 , n45256 , n45257 );
and ( n45259 , n45258 , n28589 );
and ( n45260 , n26799 , n31075 );
or ( n45261 , n45259 , n45260 );
and ( n45262 , n45261 , n28594 );
not ( n45263 , n30249 );
and ( n45264 , n45263 , n30228 );
xor ( n45265 , n30228 , n29753 );
xor ( n45266 , n30211 , n29753 );
xor ( n45267 , n30194 , n29753 );
and ( n45268 , n43427 , n43432 );
and ( n45269 , n45267 , n45268 );
and ( n45270 , n45266 , n45269 );
xor ( n45271 , n45265 , n45270 );
and ( n45272 , n45271 , n30249 );
or ( n45273 , n45264 , n45272 );
buf ( n45274 , n45273 );
and ( n45275 , n45274 , n28589 );
and ( n45276 , n26799 , n31075 );
or ( n45277 , n45275 , n45276 );
and ( n45278 , n45277 , n30269 );
not ( n45279 , n30963 );
and ( n45280 , n45279 , n30942 );
xor ( n45281 , n30942 , n30467 );
xor ( n45282 , n30925 , n30467 );
xor ( n45283 , n30908 , n30467 );
and ( n45284 , n43443 , n43448 );
and ( n45285 , n45283 , n45284 );
and ( n45286 , n45282 , n45285 );
xor ( n45287 , n45281 , n45286 );
and ( n45288 , n45287 , n30963 );
or ( n45289 , n45280 , n45288 );
buf ( n45290 , n45289 );
and ( n45291 , n45290 , n28589 );
and ( n45292 , n26799 , n31075 );
or ( n45293 , n45291 , n45292 );
and ( n45294 , n45293 , n30982 );
and ( n45295 , n29133 , n28589 );
and ( n45296 , n26799 , n31075 );
or ( n45297 , n45295 , n45296 );
and ( n45298 , n45297 , n30989 );
and ( n45299 , n29133 , n30991 );
buf ( n45300 , n29133 );
not ( n45301 , n45300 );
buf ( n45302 , n29146 );
not ( n45303 , n45302 );
buf ( n45304 , n29159 );
not ( n45305 , n45304 );
and ( n45306 , n43462 , n43469 );
and ( n45307 , n45305 , n45306 );
and ( n45308 , n45303 , n45307 );
xor ( n45309 , n45301 , n45308 );
buf ( n45310 , n45309 );
and ( n45311 , n45310 , n28589 );
and ( n45312 , n26799 , n31075 );
or ( n45313 , n45311 , n45312 );
and ( n45314 , n45313 , n31002 );
or ( n45315 , n45225 , n45262 , n45278 , n45294 , n45298 , n45299 , n45314 );
and ( n45316 , n45224 , n45315 );
and ( n45317 , n26799 , n24800 );
or ( n45318 , n45316 , n45317 );
and ( n45319 , n45318 , n31008 );
and ( n45320 , n25639 , n10618 );
or ( n45321 , n45319 , n45320 );
buf ( n45322 , n45321 );
buf ( n45323 , n45322 );
and ( n45324 , n24333 , n31008 );
and ( n45325 , n29118 , n10618 );
or ( n45326 , n45324 , n45325 );
buf ( n45327 , n45326 );
buf ( n45328 , n45327 );
not ( n45329 , n17451 );
not ( n45330 , n19474 );
and ( n45331 , n45330 , n19436 );
xor ( n45332 , n40059 , n40062 );
and ( n45333 , n45332 , n19474 );
or ( n45334 , n45331 , n45333 );
buf ( n45335 , n45334 );
and ( n45336 , n45335 , n19745 );
and ( n45337 , n45335 , n19748 );
not ( n45338 , n19750 );
and ( n45339 , n45338 , n21177 );
not ( n45340 , n21193 );
and ( n45341 , n45340 , n21189 );
xor ( n45342 , n21189 , n20582 );
xor ( n45343 , n21167 , n20582 );
and ( n45344 , n39866 , n39867 );
and ( n45345 , n45343 , n45344 );
xor ( n45346 , n45342 , n45345 );
and ( n45347 , n45346 , n21193 );
or ( n45348 , n45341 , n45347 );
buf ( n45349 , n45348 );
and ( n45350 , n45349 , n19750 );
or ( n45351 , n45339 , n45350 );
and ( n45352 , n45351 , n21253 );
and ( n45353 , n21177 , n21255 );
or ( n45354 , n45336 , n45337 , n45352 , n45353 );
and ( n45355 , n45354 , n21333 );
and ( n45356 , n19454 , n34758 );
or ( n45357 , n45355 , n45356 );
and ( n45358 , n45357 , n21341 );
not ( n45359 , n22996 );
and ( n45360 , n45359 , n22975 );
xor ( n45361 , n40087 , n40090 );
and ( n45362 , n45361 , n22996 );
or ( n45363 , n45360 , n45362 );
buf ( n45364 , n45363 );
and ( n45365 , n45364 , n21333 );
and ( n45366 , n19454 , n34758 );
or ( n45367 , n45365 , n45366 );
and ( n45368 , n45367 , n23064 );
not ( n45369 , n23758 );
and ( n45370 , n45369 , n23737 );
xor ( n45371 , n40102 , n40105 );
and ( n45372 , n45371 , n23758 );
or ( n45373 , n45370 , n45372 );
buf ( n45374 , n45373 );
and ( n45375 , n45374 , n21333 );
and ( n45376 , n19454 , n34758 );
or ( n45377 , n45375 , n45376 );
and ( n45378 , n45377 , n23825 );
and ( n45379 , n21880 , n21333 );
and ( n45380 , n19454 , n34758 );
or ( n45381 , n45379 , n45380 );
and ( n45382 , n45381 , n23832 );
xor ( n45383 , n40126 , n40130 );
buf ( n45384 , n45383 );
and ( n45385 , n45384 , n21333 );
and ( n45386 , n19454 , n34758 );
or ( n45387 , n45385 , n45386 );
and ( n45388 , n45387 , n23917 );
and ( n45389 , n19454 , n34526 );
or ( n45390 , n45358 , n45368 , n45378 , n45382 , n45388 , n45389 );
and ( n45391 , n45329 , n45390 );
and ( n45392 , n19454 , n17451 );
or ( n45393 , n45391 , n45392 );
and ( n45394 , n45393 , n23924 );
and ( n45395 , n19454 , n23926 );
or ( n45396 , n45394 , n45395 );
buf ( n45397 , n45396 );
buf ( n45398 , n45397 );
buf ( n45399 , n10613 );
buf ( n45400 , n10615 );
buf ( n45401 , n10615 );
buf ( n45402 , n10615 );
buf ( n45403 , n10615 );
not ( n45404 , n34821 );
not ( n45405 , n13916 );
and ( n45406 , n45405 , n13705 );
xor ( n45407 , n13706 , n13869 );
and ( n45408 , n45407 , n13916 );
or ( n45409 , n45406 , n45408 );
buf ( n45410 , n45409 );
and ( n45411 , n45410 , n14137 );
and ( n45412 , n45410 , n14143 );
not ( n45413 , n14139 );
and ( n45414 , n45413 , n35943 );
not ( n45415 , n36245 );
and ( n45416 , n45415 , n35955 );
xor ( n45417 , n43030 , n43039 );
and ( n45418 , n45417 , n36245 );
or ( n45419 , n45416 , n45418 );
buf ( n45420 , n45419 );
and ( n45421 , n45420 , n14139 );
or ( n45422 , n45414 , n45421 );
and ( n45423 , n45422 , n14140 );
and ( n45424 , n35943 , n14141 );
or ( n45425 , n45411 , n45412 , n45423 , n45424 );
and ( n45426 , n45425 , n36347 );
and ( n45427 , n13315 , n39408 );
or ( n45428 , n45426 , n45427 );
and ( n45429 , n45428 , n14562 );
not ( n45430 , n37048 );
and ( n45431 , n45430 , n36806 );
xor ( n45432 , n43057 , n43066 );
and ( n45433 , n45432 , n37048 );
or ( n45434 , n45431 , n45433 );
buf ( n45435 , n45434 );
and ( n45436 , n45435 , n36348 );
and ( n45437 , n13315 , n39427 );
or ( n45438 , n45436 , n45437 );
and ( n45439 , n45438 , n14586 );
not ( n45440 , n37801 );
and ( n45441 , n45440 , n37559 );
xor ( n45442 , n43079 , n43088 );
and ( n45443 , n45442 , n37801 );
or ( n45444 , n45441 , n45443 );
buf ( n45445 , n45444 );
and ( n45446 , n45445 , n36347 );
and ( n45447 , n13315 , n39446 );
or ( n45448 , n45446 , n45447 );
and ( n45449 , n45448 , n14584 );
and ( n45450 , n45435 , n36348 );
and ( n45451 , n13315 , n39453 );
or ( n45452 , n45450 , n45451 );
and ( n45453 , n45452 , n37835 );
and ( n45454 , n45445 , n36348 );
and ( n45455 , n13315 , n39453 );
or ( n45456 , n45454 , n45455 );
and ( n45457 , n45456 , n37841 );
and ( n45458 , n15537 , n36348 );
and ( n45459 , n13315 , n39453 );
or ( n45460 , n45458 , n45459 );
and ( n45461 , n45460 , n37847 );
and ( n45462 , n13315 , n37849 );
or ( n45463 , n45429 , n45439 , n45449 , n45453 , n45457 , n45461 , n45462 );
and ( n45464 , n45404 , n45463 );
and ( n45465 , n13315 , n34821 );
or ( n45466 , n45464 , n45465 );
and ( n45467 , n45466 , n16574 );
and ( n45468 , n13315 , n16576 );
or ( n45469 , n45467 , n45468 );
buf ( n45470 , n45469 );
buf ( n45471 , n45470 );
buf ( n45472 , n10615 );
buf ( n45473 , n10613 );
buf ( n45474 , n10615 );
not ( n45475 , n34804 );
and ( n45476 , n45475 , n26093 );
and ( n45477 , n14791 , n34804 );
or ( n45478 , n45476 , n45477 );
and ( n45479 , n45478 , n31008 );
and ( n45480 , n14791 , n10618 );
or ( n45481 , n45479 , n45480 );
buf ( n45482 , n45481 );
buf ( n45483 , n45482 );
not ( n45484 , n17162 );
not ( n45485 , n17450 );
and ( n45486 , n10693 , n37947 );
not ( n45487 , n38425 );
and ( n45488 , n45487 , n38234 );
xor ( n45489 , n38432 , n38448 );
and ( n45490 , n45489 , n38425 );
or ( n45491 , n45488 , n45490 );
buf ( n45492 , n45491 );
and ( n45493 , n45492 , n19745 );
not ( n45494 , n38934 );
and ( n45495 , n45494 , n38743 );
xor ( n45496 , n38941 , n38957 );
and ( n45497 , n45496 , n38934 );
or ( n45498 , n45495 , n45497 );
buf ( n45499 , n45498 );
and ( n45500 , n45499 , n19748 );
and ( n45501 , n22260 , n21253 );
and ( n45502 , n10693 , n21255 );
or ( n45503 , n45493 , n45500 , n45501 , n45502 );
and ( n45504 , n45503 , n38980 );
or ( n45505 , n45486 , n45504 );
and ( n45506 , n45485 , n45505 );
or ( n45507 , n45506 , C0 );
and ( n45508 , n45484 , n45507 );
and ( n45509 , n45503 , n17162 );
or ( n45510 , n45508 , n45509 );
and ( n45511 , n45510 , n23924 );
not ( n45512 , n39264 );
and ( n45513 , n45512 , n39106 );
xor ( n45514 , n39271 , n39287 );
and ( n45515 , n45514 , n39264 );
or ( n45516 , n45513 , n45515 );
buf ( n45517 , n45516 );
and ( n45518 , n45517 , n23926 );
or ( n45519 , n45511 , n45518 );
buf ( n45520 , n45519 );
buf ( n45521 , n45520 );
buf ( n45522 , n10615 );
buf ( n45523 , n10613 );
buf ( n45524 , n10613 );
buf ( n45525 , n10615 );
buf ( n45526 , n10613 );
not ( n45527 , n24800 );
and ( n45528 , n25983 , n25222 );
not ( n45529 , n26823 );
and ( n45530 , n45529 , n25970 );
xor ( n45531 , n31024 , n31029 );
and ( n45532 , n45531 , n26823 );
or ( n45533 , n45530 , n45532 );
buf ( n45534 , n45533 );
and ( n45535 , n45534 , n27046 );
and ( n45536 , n45534 , n27049 );
not ( n45537 , n27051 );
and ( n45538 , n45537 , n27950 );
not ( n45539 , n28494 );
and ( n45540 , n45539 , n27962 );
xor ( n45541 , n31052 , n31057 );
and ( n45542 , n45541 , n28494 );
or ( n45543 , n45540 , n45542 );
buf ( n45544 , n45543 );
and ( n45545 , n45544 , n27051 );
or ( n45546 , n45538 , n45545 );
and ( n45547 , n45546 , n28506 );
and ( n45548 , n27950 , n28508 );
or ( n45549 , n45535 , n45536 , n45547 , n45548 );
and ( n45550 , n45549 , n28589 );
and ( n45551 , n25983 , n31075 );
or ( n45552 , n45550 , n45551 );
and ( n45553 , n45552 , n28594 );
not ( n45554 , n30249 );
and ( n45555 , n45554 , n29820 );
xor ( n45556 , n31087 , n31092 );
and ( n45557 , n45556 , n30249 );
or ( n45558 , n45555 , n45557 );
buf ( n45559 , n45558 );
and ( n45560 , n45559 , n28589 );
and ( n45561 , n25983 , n31075 );
or ( n45562 , n45560 , n45561 );
and ( n45563 , n45562 , n30269 );
not ( n45564 , n30963 );
and ( n45565 , n45564 , n30534 );
xor ( n45566 , n31115 , n31120 );
and ( n45567 , n45566 , n30963 );
or ( n45568 , n45565 , n45567 );
buf ( n45569 , n45568 );
and ( n45570 , n45569 , n28589 );
and ( n45571 , n25983 , n31075 );
or ( n45572 , n45570 , n45571 );
and ( n45573 , n45572 , n30982 );
and ( n45574 , n29595 , n28589 );
and ( n45575 , n25983 , n31075 );
or ( n45576 , n45574 , n45575 );
and ( n45577 , n45576 , n30989 );
and ( n45578 , n29595 , n30991 );
xor ( n45579 , n31153 , n31160 );
buf ( n45580 , n45579 );
and ( n45581 , n45580 , n28589 );
and ( n45582 , n25983 , n31075 );
or ( n45583 , n45581 , n45582 );
and ( n45584 , n45583 , n31002 );
or ( n45585 , n45528 , n45553 , n45563 , n45573 , n45577 , n45578 , n45584 );
and ( n45586 , n45527 , n45585 );
and ( n45587 , n25983 , n24800 );
or ( n45588 , n45586 , n45587 );
and ( n45589 , n45588 , n31008 );
and ( n45590 , n25279 , n10618 );
or ( n45591 , n45589 , n45590 );
buf ( n45592 , n45591 );
buf ( n45593 , n45592 );
not ( n45594 , n24800 );
and ( n45595 , n45088 , n28587 );
and ( n45596 , n26295 , n39807 );
or ( n45597 , n45595 , n45596 );
and ( n45598 , n45597 , n28594 );
and ( n45599 , n45098 , n28587 );
and ( n45600 , n26295 , n39807 );
or ( n45601 , n45599 , n45600 );
and ( n45602 , n45601 , n30269 );
and ( n45603 , n45108 , n28587 );
and ( n45604 , n26295 , n39807 );
or ( n45605 , n45603 , n45604 );
and ( n45606 , n45605 , n30982 );
and ( n45607 , n29415 , n28587 );
and ( n45608 , n26295 , n39807 );
or ( n45609 , n45607 , n45608 );
and ( n45610 , n45609 , n30989 );
and ( n45611 , n45119 , n28587 );
and ( n45612 , n26295 , n39807 );
or ( n45613 , n45611 , n45612 );
and ( n45614 , n45613 , n31002 );
and ( n45615 , n26295 , n34607 );
or ( n45616 , n45598 , n45602 , n45606 , n45610 , n45614 , n45615 );
and ( n45617 , n45594 , n45616 );
and ( n45618 , n26295 , n24800 );
or ( n45619 , n45617 , n45618 );
and ( n45620 , n45619 , n31008 );
and ( n45621 , n26295 , n10618 );
or ( n45622 , n45620 , n45621 );
buf ( n45623 , n45622 );
buf ( n45624 , n45623 );
buf ( n45625 , n10615 );
not ( n45626 , n34821 );
not ( n45627 , n13916 );
and ( n45628 , n45627 , n13749 );
xor ( n45629 , n13750 , n13865 );
and ( n45630 , n45629 , n13916 );
or ( n45631 , n45628 , n45630 );
buf ( n45632 , n45631 );
and ( n45633 , n45632 , n14137 );
and ( n45634 , n45632 , n14143 );
not ( n45635 , n14139 );
and ( n45636 , n45635 , n35855 );
not ( n45637 , n36245 );
and ( n45638 , n45637 , n35867 );
xor ( n45639 , n43034 , n43035 );
and ( n45640 , n45639 , n36245 );
or ( n45641 , n45638 , n45640 );
buf ( n45642 , n45641 );
and ( n45643 , n45642 , n14139 );
or ( n45644 , n45636 , n45643 );
and ( n45645 , n45644 , n14140 );
and ( n45646 , n35855 , n14141 );
or ( n45647 , n45633 , n45634 , n45645 , n45646 );
and ( n45648 , n45647 , n36347 );
and ( n45649 , n13363 , n39408 );
or ( n45650 , n45648 , n45649 );
and ( n45651 , n45650 , n14562 );
not ( n45652 , n37048 );
and ( n45653 , n45652 , n36738 );
xor ( n45654 , n43061 , n43062 );
and ( n45655 , n45654 , n37048 );
or ( n45656 , n45653 , n45655 );
buf ( n45657 , n45656 );
and ( n45658 , n45657 , n36348 );
and ( n45659 , n13363 , n39427 );
or ( n45660 , n45658 , n45659 );
and ( n45661 , n45660 , n14586 );
not ( n45662 , n37801 );
and ( n45663 , n45662 , n37491 );
xor ( n45664 , n43083 , n43084 );
and ( n45665 , n45664 , n37801 );
or ( n45666 , n45663 , n45665 );
buf ( n45667 , n45666 );
and ( n45668 , n45667 , n36347 );
and ( n45669 , n13363 , n39446 );
or ( n45670 , n45668 , n45669 );
and ( n45671 , n45670 , n14584 );
and ( n45672 , n45657 , n36348 );
and ( n45673 , n13363 , n39453 );
or ( n45674 , n45672 , n45673 );
and ( n45675 , n45674 , n37835 );
and ( n45676 , n45667 , n36348 );
and ( n45677 , n13363 , n39453 );
or ( n45678 , n45676 , n45677 );
and ( n45679 , n45678 , n37841 );
and ( n45680 , n15625 , n36348 );
and ( n45681 , n13363 , n39453 );
or ( n45682 , n45680 , n45681 );
and ( n45683 , n45682 , n37847 );
and ( n45684 , n13363 , n37849 );
or ( n45685 , n45651 , n45661 , n45671 , n45675 , n45679 , n45683 , n45684 );
and ( n45686 , n45626 , n45685 );
and ( n45687 , n13363 , n34821 );
or ( n45688 , n45686 , n45687 );
and ( n45689 , n45688 , n16574 );
and ( n45690 , n13363 , n16576 );
or ( n45691 , n45689 , n45690 );
buf ( n45692 , n45691 );
buf ( n45693 , n45692 );
buf ( n45694 , n10615 );
buf ( n45695 , n10615 );
buf ( n45696 , n10615 );
buf ( n45697 , n10613 );
buf ( n45698 , n10615 );
buf ( n45699 , n10615 );
buf ( n45700 , n10615 );
buf ( n45701 , n10613 );
buf ( n45702 , n10613 );
buf ( n45703 , n10613 );
buf ( n45704 , n10615 );
buf ( n45705 , n10613 );
not ( n45706 , n34538 );
and ( n45707 , n45706 , n19390 );
and ( n45708 , n14675 , n34538 );
or ( n45709 , n45707 , n45708 );
and ( n45710 , n45709 , n23924 );
and ( n45711 , n14675 , n23926 );
or ( n45712 , n45710 , n45711 );
buf ( n45713 , n45712 );
buf ( n45714 , n45713 );
buf ( n45715 , n10613 );
buf ( n45716 , n10615 );
buf ( n45717 , n10615 );
buf ( n45718 , n10613 );
not ( n45719 , n34821 );
not ( n45720 , n13916 );
and ( n45721 , n45720 , n13628 );
xor ( n45722 , n13629 , n13876 );
and ( n45723 , n45722 , n13916 );
or ( n45724 , n45721 , n45723 );
buf ( n45725 , n45724 );
and ( n45726 , n45725 , n14137 );
and ( n45727 , n45725 , n14143 );
not ( n45728 , n14139 );
and ( n45729 , n45728 , n36097 );
not ( n45730 , n36245 );
and ( n45731 , n45730 , n36109 );
xor ( n45732 , n36109 , n35634 );
xor ( n45733 , n36087 , n35634 );
xor ( n45734 , n36065 , n35634 );
and ( n45735 , n45151 , n45156 );
and ( n45736 , n45734 , n45735 );
and ( n45737 , n45733 , n45736 );
xor ( n45738 , n45732 , n45737 );
and ( n45739 , n45738 , n36245 );
or ( n45740 , n45731 , n45739 );
buf ( n45741 , n45740 );
and ( n45742 , n45741 , n14139 );
or ( n45743 , n45729 , n45742 );
and ( n45744 , n45743 , n14140 );
and ( n45745 , n36097 , n14141 );
or ( n45746 , n45726 , n45727 , n45744 , n45745 );
and ( n45747 , n45746 , n36345 );
and ( n45748 , n13233 , n36352 );
or ( n45749 , n45747 , n45748 );
and ( n45750 , n45749 , n14562 );
not ( n45751 , n37048 );
and ( n45752 , n45751 , n36925 );
xor ( n45753 , n36925 , n36552 );
xor ( n45754 , n36908 , n36552 );
xor ( n45755 , n36891 , n36552 );
and ( n45756 , n45172 , n45177 );
and ( n45757 , n45755 , n45756 );
and ( n45758 , n45754 , n45757 );
xor ( n45759 , n45753 , n45758 );
and ( n45760 , n45759 , n37048 );
or ( n45761 , n45752 , n45760 );
buf ( n45762 , n45761 );
and ( n45763 , n45762 , n36345 );
and ( n45764 , n13233 , n37073 );
or ( n45765 , n45763 , n45764 );
and ( n45766 , n45765 , n14586 );
not ( n45767 , n37801 );
and ( n45768 , n45767 , n37678 );
xor ( n45769 , n37678 , n37305 );
xor ( n45770 , n37661 , n37305 );
xor ( n45771 , n37644 , n37305 );
and ( n45772 , n45188 , n45193 );
and ( n45773 , n45771 , n45772 );
and ( n45774 , n45770 , n45773 );
xor ( n45775 , n45769 , n45774 );
and ( n45776 , n45775 , n37801 );
or ( n45777 , n45768 , n45776 );
buf ( n45778 , n45777 );
and ( n45779 , n45778 , n36350 );
and ( n45780 , n13233 , n37825 );
or ( n45781 , n45779 , n45780 );
and ( n45782 , n45781 , n14584 );
and ( n45783 , n45762 , n36350 );
and ( n45784 , n13233 , n37831 );
or ( n45785 , n45783 , n45784 );
and ( n45786 , n45785 , n37835 );
and ( n45787 , n45778 , n36350 );
and ( n45788 , n13233 , n37831 );
or ( n45789 , n45787 , n45788 );
and ( n45790 , n45789 , n37841 );
and ( n45791 , n15082 , n36350 );
and ( n45792 , n13233 , n37831 );
or ( n45793 , n45791 , n45792 );
and ( n45794 , n45793 , n37847 );
and ( n45795 , n13233 , n37849 );
or ( n45796 , n45750 , n45766 , n45782 , n45786 , n45790 , n45794 , n45795 );
and ( n45797 , n45719 , n45796 );
and ( n45798 , n13233 , n34821 );
or ( n45799 , n45797 , n45798 );
and ( n45800 , n45799 , n16574 );
and ( n45801 , n13233 , n16576 );
or ( n45802 , n45800 , n45801 );
buf ( n45803 , n45802 );
buf ( n45804 , n45803 );
buf ( n45805 , n10613 );
not ( n45806 , n34821 );
and ( n45807 , n43526 , n36345 );
and ( n45808 , n13495 , n36352 );
or ( n45809 , n45807 , n45808 );
and ( n45810 , n45809 , n14562 );
and ( n45811 , n43539 , n36345 );
and ( n45812 , n13495 , n37073 );
or ( n45813 , n45811 , n45812 );
and ( n45814 , n45813 , n14586 );
and ( n45815 , n43552 , n36350 );
and ( n45816 , n13495 , n37825 );
or ( n45817 , n45815 , n45816 );
and ( n45818 , n45817 , n14584 );
and ( n45819 , n43539 , n36350 );
and ( n45820 , n13495 , n37831 );
or ( n45821 , n45819 , n45820 );
and ( n45822 , n45821 , n37835 );
and ( n45823 , n43552 , n36350 );
and ( n45824 , n13495 , n37831 );
or ( n45825 , n45823 , n45824 );
and ( n45826 , n45825 , n37841 );
and ( n45827 , n15845 , n36350 );
and ( n45828 , n13495 , n37831 );
or ( n45829 , n45827 , n45828 );
and ( n45830 , n45829 , n37847 );
and ( n45831 , n13495 , n37849 );
or ( n45832 , n45810 , n45814 , n45818 , n45822 , n45826 , n45830 , n45831 );
and ( n45833 , n45806 , n45832 );
and ( n45834 , n13495 , n34821 );
or ( n45835 , n45833 , n45834 );
and ( n45836 , n45835 , n16574 );
and ( n45837 , n13495 , n16576 );
or ( n45838 , n45836 , n45837 );
buf ( n45839 , n45838 );
buf ( n45840 , n45839 );
buf ( n45841 , n10613 );
and ( n45842 , n24206 , n31008 );
and ( n45843 , n29546 , n10618 );
or ( n45844 , n45842 , n45843 );
buf ( n45845 , n45844 );
buf ( n45846 , n45845 );
buf ( n45847 , n10613 );
buf ( n45848 , n10615 );
buf ( n45849 , n10615 );
buf ( n45850 , n10613 );
buf ( n45851 , n10613 );
not ( n45852 , n24800 );
and ( n45853 , n26561 , n25222 );
not ( n45854 , n26823 );
and ( n45855 , n45854 , n26547 );
xor ( n45856 , n42827 , n42834 );
and ( n45857 , n45856 , n26823 );
or ( n45858 , n45855 , n45857 );
buf ( n45859 , n45858 );
and ( n45860 , n45859 , n27046 );
and ( n45861 , n45859 , n27049 );
not ( n45862 , n27051 );
and ( n45863 , n45862 , n28324 );
not ( n45864 , n28494 );
and ( n45865 , n45864 , n28336 );
xor ( n45866 , n42847 , n42854 );
and ( n45867 , n45866 , n28494 );
or ( n45868 , n45865 , n45867 );
buf ( n45869 , n45868 );
and ( n45870 , n45869 , n27051 );
or ( n45871 , n45863 , n45870 );
and ( n45872 , n45871 , n28506 );
and ( n45873 , n28324 , n28508 );
or ( n45874 , n45860 , n45861 , n45872 , n45873 );
and ( n45875 , n45874 , n28589 );
and ( n45876 , n26561 , n31075 );
or ( n45877 , n45875 , n45876 );
and ( n45878 , n45877 , n28594 );
not ( n45879 , n30249 );
and ( n45880 , n45879 , n30109 );
xor ( n45881 , n42872 , n42879 );
and ( n45882 , n45881 , n30249 );
or ( n45883 , n45880 , n45882 );
buf ( n45884 , n45883 );
and ( n45885 , n45884 , n28589 );
and ( n45886 , n26561 , n31075 );
or ( n45887 , n45885 , n45886 );
and ( n45888 , n45887 , n30269 );
not ( n45889 , n30963 );
and ( n45890 , n45889 , n30823 );
xor ( n45891 , n42892 , n42899 );
and ( n45892 , n45891 , n30963 );
or ( n45893 , n45890 , n45892 );
buf ( n45894 , n45893 );
and ( n45895 , n45894 , n28589 );
and ( n45896 , n26561 , n31075 );
or ( n45897 , n45895 , n45896 );
and ( n45898 , n45897 , n30982 );
and ( n45899 , n29224 , n28589 );
and ( n45900 , n26561 , n31075 );
or ( n45901 , n45899 , n45900 );
and ( n45902 , n45901 , n30989 );
and ( n45903 , n29224 , n30991 );
xor ( n45904 , n42916 , n42926 );
buf ( n45905 , n45904 );
and ( n45906 , n45905 , n28589 );
and ( n45907 , n26561 , n31075 );
or ( n45908 , n45906 , n45907 );
and ( n45909 , n45908 , n31002 );
or ( n45910 , n45853 , n45878 , n45888 , n45898 , n45902 , n45903 , n45909 );
and ( n45911 , n45852 , n45910 );
and ( n45912 , n26561 , n24800 );
or ( n45913 , n45911 , n45912 );
and ( n45914 , n45913 , n31008 );
and ( n45915 , n25534 , n10618 );
or ( n45916 , n45914 , n45915 );
buf ( n45917 , n45916 );
buf ( n45918 , n45917 );
buf ( n45919 , n10615 );
buf ( n45920 , n10615 );
not ( n45921 , n17451 );
and ( n45922 , n19043 , n17873 );
not ( n45923 , n19474 );
and ( n45924 , n45923 , n19029 );
xor ( n45925 , n19486 , n19516 );
and ( n45926 , n45925 , n19474 );
or ( n45927 , n45924 , n45926 );
buf ( n45928 , n45927 );
and ( n45929 , n45928 , n19745 );
and ( n45930 , n45928 , n19748 );
not ( n45931 , n19750 );
and ( n45932 , n45931 , n20921 );
not ( n45933 , n21193 );
and ( n45934 , n45933 , n20933 );
xor ( n45935 , n21205 , n21237 );
and ( n45936 , n45935 , n21193 );
or ( n45937 , n45934 , n45936 );
buf ( n45938 , n45937 );
and ( n45939 , n45938 , n19750 );
or ( n45940 , n45932 , n45939 );
and ( n45941 , n45940 , n21253 );
and ( n45942 , n20921 , n21255 );
or ( n45943 , n45929 , n45930 , n45941 , n45942 );
and ( n45944 , n45943 , n21336 );
and ( n45945 , n19043 , n42682 );
or ( n45946 , n45944 , n45945 );
and ( n45947 , n45946 , n21341 );
not ( n45948 , n22996 );
and ( n45949 , n45948 , n22771 );
xor ( n45950 , n23008 , n23040 );
and ( n45951 , n45950 , n22996 );
or ( n45952 , n45949 , n45951 );
buf ( n45953 , n45952 );
and ( n45954 , n45953 , n21336 );
and ( n45955 , n19043 , n42682 );
or ( n45956 , n45954 , n45955 );
and ( n45957 , n45956 , n23064 );
not ( n45958 , n23758 );
and ( n45959 , n45958 , n23533 );
xor ( n45960 , n23770 , n23802 );
and ( n45961 , n45960 , n23758 );
or ( n45962 , n45959 , n45961 );
buf ( n45963 , n45962 );
and ( n45964 , n45963 , n21336 );
and ( n45965 , n19043 , n42682 );
or ( n45966 , n45964 , n45965 );
and ( n45967 , n45966 , n23825 );
and ( n45968 , n22102 , n21336 );
and ( n45969 , n19043 , n42682 );
or ( n45970 , n45968 , n45969 );
and ( n45971 , n45970 , n23832 );
and ( n45972 , n22102 , n23834 );
xor ( n45973 , n23855 , n23902 );
buf ( n45974 , n45973 );
and ( n45975 , n45974 , n21336 );
and ( n45976 , n19043 , n42682 );
or ( n45977 , n45975 , n45976 );
and ( n45978 , n45977 , n23917 );
or ( n45979 , n45922 , n45947 , n45957 , n45967 , n45971 , n45972 , n45978 );
and ( n45980 , n45921 , n45979 );
and ( n45981 , n19043 , n17451 );
or ( n45982 , n45980 , n45981 );
and ( n45983 , n45982 , n23924 );
and ( n45984 , n18110 , n23926 );
or ( n45985 , n45983 , n45984 );
buf ( n45986 , n45985 );
buf ( n45987 , n45986 );
buf ( n45988 , n10615 );
buf ( n45989 , n10613 );
buf ( n45990 , n10613 );
not ( n45991 , n24511 );
not ( n45992 , n24799 );
and ( n45993 , n10715 , n40154 );
not ( n45994 , n40632 );
and ( n45995 , n45994 , n40373 );
xor ( n45996 , n40646 , n40654 );
and ( n45997 , n45996 , n40632 );
or ( n45998 , n45995 , n45997 );
buf ( n45999 , n45998 );
and ( n46000 , n45999 , n27046 );
not ( n46001 , n41147 );
and ( n46002 , n46001 , n40888 );
xor ( n46003 , n41161 , n41169 );
and ( n46004 , n46003 , n41147 );
or ( n46005 , n46002 , n46004 );
buf ( n46006 , n46005 );
and ( n46007 , n46006 , n27049 );
and ( n46008 , n29593 , n28506 );
and ( n46009 , n10715 , n28508 );
or ( n46010 , n46000 , n46007 , n46008 , n46009 );
and ( n46011 , n46010 , n41199 );
or ( n46012 , n45993 , n46011 );
and ( n46013 , n45992 , n46012 );
xor ( n46014 , n41692 , n41700 );
xor ( n46015 , n46014 , n41773 );
buf ( n46016 , n46015 );
and ( n46017 , n46016 , n27046 );
xor ( n46018 , n42222 , n42223 );
xor ( n46019 , n46018 , n42269 );
buf ( n46020 , n46019 );
and ( n46021 , n46020 , n27049 );
and ( n46022 , n29593 , n42306 );
or ( n46023 , n46017 , n46021 , n46022 );
buf ( n46024 , n46023 );
and ( n46025 , C1 , n46024 );
or ( n46026 , n46025 , C0 );
buf ( n46027 , n46026 );
not ( n46028 , n46027 );
buf ( n46029 , n46028 );
buf ( n46030 , n46029 );
not ( n46031 , n46030 );
and ( n46032 , C1 , n46031 );
or ( n46033 , n46032 , C0 );
buf ( n46034 , n46033 );
and ( n46035 , n46034 , n24799 );
or ( n46036 , n46013 , n46035 );
and ( n46037 , n45991 , n46036 );
and ( n46038 , n46010 , n24511 );
or ( n46039 , n46037 , n46038 );
and ( n46040 , n46039 , n31008 );
not ( n46041 , n42601 );
and ( n46042 , n46041 , n42387 );
xor ( n46043 , n42615 , n42623 );
and ( n46044 , n46043 , n42601 );
or ( n46045 , n46042 , n46044 );
buf ( n46046 , n46045 );
and ( n46047 , n46046 , n10618 );
or ( n46048 , n46040 , n46047 );
buf ( n46049 , n46048 );
buf ( n46050 , n46049 );
buf ( n46051 , n10613 );
buf ( n46052 , n10615 );
buf ( n46053 , n10615 );
buf ( n46054 , n10613 );
not ( n46055 , n17451 );
and ( n46056 , n19181 , n17873 );
not ( n46057 , n19474 );
and ( n46058 , n46057 , n19165 );
xor ( n46059 , n19482 , n19520 );
and ( n46060 , n46059 , n19474 );
or ( n46061 , n46058 , n46060 );
buf ( n46062 , n46061 );
and ( n46063 , n46062 , n19745 );
and ( n46064 , n46062 , n19748 );
not ( n46065 , n19750 );
and ( n46066 , n46065 , n21009 );
not ( n46067 , n21193 );
and ( n46068 , n46067 , n21021 );
xor ( n46069 , n21201 , n21241 );
and ( n46070 , n46069 , n21193 );
or ( n46071 , n46068 , n46070 );
buf ( n46072 , n46071 );
and ( n46073 , n46072 , n19750 );
or ( n46074 , n46066 , n46073 );
and ( n46075 , n46074 , n21253 );
and ( n46076 , n21009 , n21255 );
or ( n46077 , n46063 , n46064 , n46075 , n46076 );
and ( n46078 , n46077 , n21330 );
and ( n46079 , n19181 , n21338 );
or ( n46080 , n46078 , n46079 );
and ( n46081 , n46080 , n21341 );
not ( n46082 , n22996 );
and ( n46083 , n46082 , n22839 );
xor ( n46084 , n23004 , n23044 );
and ( n46085 , n46084 , n22996 );
or ( n46086 , n46083 , n46085 );
buf ( n46087 , n46086 );
and ( n46088 , n46087 , n21330 );
and ( n46089 , n19181 , n21338 );
or ( n46090 , n46088 , n46089 );
and ( n46091 , n46090 , n23064 );
not ( n46092 , n23758 );
and ( n46093 , n46092 , n23601 );
xor ( n46094 , n23766 , n23806 );
and ( n46095 , n46094 , n23758 );
or ( n46096 , n46093 , n46095 );
buf ( n46097 , n46096 );
and ( n46098 , n46097 , n21330 );
and ( n46099 , n19181 , n21338 );
or ( n46100 , n46098 , n46099 );
and ( n46101 , n46100 , n23825 );
and ( n46102 , n21984 , n21330 );
and ( n46103 , n19181 , n21338 );
or ( n46104 , n46102 , n46103 );
and ( n46105 , n46104 , n23832 );
and ( n46106 , n19179 , n23834 );
xor ( n46107 , n23847 , n23906 );
buf ( n46108 , n46107 );
and ( n46109 , n46108 , n21330 );
and ( n46110 , n19181 , n21338 );
or ( n46111 , n46109 , n46110 );
and ( n46112 , n46111 , n23917 );
or ( n46113 , n46056 , n46081 , n46091 , n46101 , n46105 , n46106 , n46112 );
and ( n46114 , n46055 , n46113 );
and ( n46115 , n19181 , n17451 );
or ( n46116 , n46114 , n46115 );
and ( n46117 , n46116 , n23924 );
and ( n46118 , n19181 , n23926 );
or ( n46119 , n46117 , n46118 );
buf ( n46120 , n46119 );
buf ( n46121 , n46120 );
buf ( n46122 , n10613 );
buf ( n46123 , n10615 );
buf ( n46124 , n10613 );
buf ( n46125 , n10613 );
buf ( n46126 , n10613 );
buf ( n46127 , n10615 );
buf ( n46128 , n10615 );
buf ( n46129 , n10615 );
buf ( n46130 , n10613 );
buf ( n46131 , n10613 );
buf ( n46132 , n10615 );
buf ( n46133 , n10613 );
buf ( n46134 , n10613 );
buf ( n46135 , n10615 );
not ( n46136 , n34821 );
and ( n46137 , n13277 , n14592 );
not ( n46138 , n13916 );
and ( n46139 , n46138 , n13672 );
xor ( n46140 , n13673 , n13872 );
and ( n46141 , n46140 , n13916 );
or ( n46142 , n46139 , n46141 );
buf ( n46143 , n46142 );
and ( n46144 , n46143 , n14137 );
and ( n46145 , n46143 , n14143 );
not ( n46146 , n14139 );
and ( n46147 , n46146 , n36009 );
not ( n46148 , n36245 );
and ( n46149 , n46148 , n36021 );
xor ( n46150 , n45152 , n45155 );
and ( n46151 , n46150 , n36245 );
or ( n46152 , n46149 , n46151 );
buf ( n46153 , n46152 );
and ( n46154 , n46153 , n14139 );
or ( n46155 , n46147 , n46154 );
and ( n46156 , n46155 , n14140 );
and ( n46157 , n36009 , n14141 );
or ( n46158 , n46144 , n46145 , n46156 , n46157 );
and ( n46159 , n46158 , n36348 );
and ( n46160 , n13277 , n43530 );
or ( n46161 , n46159 , n46160 );
and ( n46162 , n46161 , n14562 );
not ( n46163 , n37048 );
and ( n46164 , n46163 , n36857 );
xor ( n46165 , n45173 , n45176 );
and ( n46166 , n46165 , n37048 );
or ( n46167 , n46164 , n46166 );
buf ( n46168 , n46167 );
and ( n46169 , n46168 , n36347 );
and ( n46170 , n13277 , n43543 );
or ( n46171 , n46169 , n46170 );
and ( n46172 , n46171 , n14586 );
not ( n46173 , n37801 );
and ( n46174 , n46173 , n37610 );
xor ( n46175 , n45189 , n45192 );
and ( n46176 , n46175 , n37801 );
or ( n46177 , n46174 , n46176 );
buf ( n46178 , n46177 );
and ( n46179 , n46178 , n36348 );
and ( n46180 , n13277 , n43556 );
or ( n46181 , n46179 , n46180 );
and ( n46182 , n46181 , n14584 );
and ( n46183 , n46168 , n36347 );
and ( n46184 , n13277 , n43563 );
or ( n46185 , n46183 , n46184 );
and ( n46186 , n46185 , n37835 );
and ( n46187 , n46178 , n36347 );
and ( n46188 , n13277 , n43563 );
or ( n46189 , n46187 , n46188 );
and ( n46190 , n46189 , n37841 );
and ( n46191 , n13275 , n14564 );
and ( n46192 , n15471 , n36347 );
and ( n46193 , n13277 , n43563 );
or ( n46194 , n46192 , n46193 );
and ( n46195 , n46194 , n37847 );
or ( n46196 , n46137 , n46162 , n46172 , n46182 , n46186 , n46190 , n46191 , n46195 );
and ( n46197 , n46136 , n46196 );
and ( n46198 , n13277 , n34821 );
or ( n46199 , n46197 , n46198 );
and ( n46200 , n46199 , n16574 );
and ( n46201 , n13277 , n16576 );
or ( n46202 , n46200 , n46201 );
buf ( n46203 , n46202 );
buf ( n46204 , n46203 );
buf ( n46205 , n10615 );
not ( n46206 , n17162 );
not ( n46207 , n17450 );
and ( n46208 , n10658 , n37947 );
not ( n46209 , n38425 );
and ( n46210 , n46209 , n38353 );
xor ( n46211 , n38353 , n38099 );
xor ( n46212 , n38336 , n38099 );
xor ( n46213 , n38319 , n38099 );
and ( n46214 , n38428 , n38452 );
and ( n46215 , n46213 , n46214 );
and ( n46216 , n46212 , n46215 );
xor ( n46217 , n46211 , n46216 );
and ( n46218 , n46217 , n38425 );
or ( n46219 , n46210 , n46218 );
buf ( n46220 , n46219 );
and ( n46221 , n46220 , n19745 );
not ( n46222 , n38934 );
and ( n46223 , n46222 , n38862 );
xor ( n46224 , n38862 , n38608 );
xor ( n46225 , n38845 , n38608 );
xor ( n46226 , n38828 , n38608 );
and ( n46227 , n38937 , n38961 );
and ( n46228 , n46226 , n46227 );
and ( n46229 , n46225 , n46228 );
xor ( n46230 , n46224 , n46229 );
and ( n46231 , n46230 , n38934 );
or ( n46232 , n46223 , n46231 );
buf ( n46233 , n46232 );
and ( n46234 , n46233 , n19748 );
and ( n46235 , n22120 , n21253 );
and ( n46236 , n10658 , n21255 );
or ( n46237 , n46221 , n46234 , n46235 , n46236 );
and ( n46238 , n46237 , n38980 );
or ( n46239 , n46208 , n46238 );
and ( n46240 , n46207 , n46239 );
or ( n46241 , n46240 , C0 );
and ( n46242 , n46206 , n46241 );
and ( n46243 , n46237 , n17162 );
or ( n46244 , n46242 , n46243 );
and ( n46245 , n46244 , n23924 );
not ( n46246 , n39264 );
and ( n46247 , n46246 , n39204 );
xor ( n46248 , n39204 , n38995 );
xor ( n46249 , n39190 , n38995 );
xor ( n46250 , n39176 , n38995 );
and ( n46251 , n39267 , n39291 );
and ( n46252 , n46250 , n46251 );
and ( n46253 , n46249 , n46252 );
xor ( n46254 , n46248 , n46253 );
and ( n46255 , n46254 , n39264 );
or ( n46256 , n46247 , n46255 );
buf ( n46257 , n46256 );
and ( n46258 , n46257 , n23926 );
or ( n46259 , n46245 , n46258 );
buf ( n46260 , n46259 );
buf ( n46261 , n46260 );
buf ( n46262 , n10615 );
buf ( n46263 , n10613 );
buf ( n46264 , n10615 );
buf ( n46265 , n10613 );
buf ( n46266 , n10613 );
buf ( n46267 , n10615 );
and ( n46268 , n11529 , n16574 );
and ( n46269 , n15095 , n16576 );
or ( n46270 , n46268 , n46269 );
buf ( n46271 , n46270 );
buf ( n46272 , n46271 );
not ( n46273 , n11333 );
and ( n46274 , n46273 , n11278 );
xor ( n46275 , n11278 , n11007 );
and ( n46276 , n11336 , n11366 );
xor ( n46277 , n46275 , n46276 );
and ( n46278 , n46277 , n11333 );
or ( n46279 , n46274 , n46278 );
buf ( n46280 , n46279 );
buf ( n46281 , n46280 );
not ( n46282 , n34821 );
and ( n46283 , n46158 , n36345 );
and ( n46284 , n13281 , n36352 );
or ( n46285 , n46283 , n46284 );
and ( n46286 , n46285 , n14562 );
and ( n46287 , n46168 , n36345 );
and ( n46288 , n13281 , n37073 );
or ( n46289 , n46287 , n46288 );
and ( n46290 , n46289 , n14586 );
and ( n46291 , n46178 , n36350 );
and ( n46292 , n13281 , n37825 );
or ( n46293 , n46291 , n46292 );
and ( n46294 , n46293 , n14584 );
and ( n46295 , n46168 , n36350 );
and ( n46296 , n13281 , n37831 );
or ( n46297 , n46295 , n46296 );
and ( n46298 , n46297 , n37835 );
and ( n46299 , n46178 , n36350 );
and ( n46300 , n13281 , n37831 );
or ( n46301 , n46299 , n46300 );
and ( n46302 , n46301 , n37841 );
and ( n46303 , n15471 , n36350 );
and ( n46304 , n13281 , n37831 );
or ( n46305 , n46303 , n46304 );
and ( n46306 , n46305 , n37847 );
and ( n46307 , n13281 , n37849 );
or ( n46308 , n46286 , n46290 , n46294 , n46298 , n46302 , n46306 , n46307 );
and ( n46309 , n46282 , n46308 );
and ( n46310 , n13281 , n34821 );
or ( n46311 , n46309 , n46310 );
and ( n46312 , n46311 , n16574 );
and ( n46313 , n13281 , n16576 );
or ( n46314 , n46312 , n46313 );
buf ( n46315 , n46314 );
buf ( n46316 , n46315 );
buf ( n46317 , n10615 );
buf ( n46318 , n10615 );
not ( n46319 , n34821 );
and ( n46320 , n13455 , n14592 );
not ( n46321 , n13916 );
and ( n46322 , n46321 , n13837 );
xor ( n46323 , n13838 , n13857 );
and ( n46324 , n46323 , n13916 );
or ( n46325 , n46322 , n46324 );
buf ( n46326 , n46325 );
and ( n46327 , n46326 , n14137 );
and ( n46328 , n46326 , n14143 );
not ( n46329 , n14139 );
and ( n46330 , n46329 , n35687 );
not ( n46331 , n36245 );
and ( n46332 , n46331 , n35699 );
xor ( n46333 , n36252 , n36258 );
and ( n46334 , n46333 , n36245 );
or ( n46335 , n46332 , n46334 );
buf ( n46336 , n46335 );
and ( n46337 , n46336 , n14139 );
or ( n46338 , n46330 , n46337 );
and ( n46339 , n46338 , n14140 );
and ( n46340 , n35687 , n14141 );
or ( n46341 , n46327 , n46328 , n46339 , n46340 );
and ( n46342 , n46341 , n36350 );
and ( n46343 , n13455 , n43691 );
or ( n46344 , n46342 , n46343 );
and ( n46345 , n46344 , n14562 );
not ( n46346 , n37048 );
and ( n46347 , n46346 , n36602 );
xor ( n46348 , n37055 , n37061 );
and ( n46349 , n46348 , n37048 );
or ( n46350 , n46347 , n46349 );
buf ( n46351 , n46350 );
and ( n46352 , n46351 , n36350 );
and ( n46353 , n13455 , n43703 );
or ( n46354 , n46352 , n46353 );
and ( n46355 , n46354 , n14586 );
not ( n46356 , n37801 );
and ( n46357 , n46356 , n37355 );
xor ( n46358 , n37808 , n37814 );
and ( n46359 , n46358 , n37801 );
or ( n46360 , n46357 , n46359 );
buf ( n46361 , n46360 );
and ( n46362 , n46361 , n36345 );
and ( n46363 , n13455 , n43715 );
or ( n46364 , n46362 , n46363 );
and ( n46365 , n46364 , n14584 );
and ( n46366 , n46351 , n36345 );
and ( n46367 , n13455 , n43721 );
or ( n46368 , n46366 , n46367 );
and ( n46369 , n46368 , n37835 );
and ( n46370 , n46361 , n36345 );
and ( n46371 , n13455 , n43721 );
or ( n46372 , n46370 , n46371 );
and ( n46373 , n46372 , n37841 );
and ( n46374 , n15801 , n14564 );
and ( n46375 , n15801 , n36345 );
and ( n46376 , n13455 , n43721 );
or ( n46377 , n46375 , n46376 );
and ( n46378 , n46377 , n37847 );
or ( n46379 , n46320 , n46345 , n46355 , n46365 , n46369 , n46373 , n46374 , n46378 );
and ( n46380 , n46319 , n46379 );
and ( n46381 , n13455 , n34821 );
or ( n46382 , n46380 , n46381 );
and ( n46383 , n46382 , n16574 );
and ( n46384 , n12324 , n16576 );
or ( n46385 , n46383 , n46384 );
buf ( n46386 , n46385 );
buf ( n46387 , n46386 );
not ( n46388 , n34821 );
and ( n46389 , n13181 , n14592 );
not ( n46390 , n13916 );
and ( n46391 , n46390 , n13584 );
xor ( n46392 , n13585 , n13880 );
and ( n46393 , n46392 , n13916 );
or ( n46394 , n46391 , n46393 );
buf ( n46395 , n46394 );
and ( n46396 , n46395 , n14137 );
and ( n46397 , n46395 , n14143 );
not ( n46398 , n14139 );
and ( n46399 , n46398 , n36185 );
not ( n46400 , n36245 );
and ( n46401 , n46400 , n36197 );
xor ( n46402 , n36197 , n35634 );
xor ( n46403 , n36175 , n35634 );
xor ( n46404 , n36153 , n35634 );
xor ( n46405 , n36131 , n35634 );
and ( n46406 , n45732 , n45737 );
and ( n46407 , n46405 , n46406 );
and ( n46408 , n46404 , n46407 );
and ( n46409 , n46403 , n46408 );
xor ( n46410 , n46402 , n46409 );
and ( n46411 , n46410 , n36245 );
or ( n46412 , n46401 , n46411 );
buf ( n46413 , n46412 );
and ( n46414 , n46413 , n14139 );
or ( n46415 , n46399 , n46414 );
and ( n46416 , n46415 , n14140 );
and ( n46417 , n36185 , n14141 );
or ( n46418 , n46396 , n46397 , n46416 , n46417 );
and ( n46419 , n46418 , n36348 );
and ( n46420 , n13181 , n43530 );
or ( n46421 , n46419 , n46420 );
and ( n46422 , n46421 , n14562 );
not ( n46423 , n37048 );
and ( n46424 , n46423 , n36993 );
xor ( n46425 , n36993 , n36552 );
xor ( n46426 , n36976 , n36552 );
xor ( n46427 , n36959 , n36552 );
xor ( n46428 , n36942 , n36552 );
and ( n46429 , n45753 , n45758 );
and ( n46430 , n46428 , n46429 );
and ( n46431 , n46427 , n46430 );
and ( n46432 , n46426 , n46431 );
xor ( n46433 , n46425 , n46432 );
and ( n46434 , n46433 , n37048 );
or ( n46435 , n46424 , n46434 );
buf ( n46436 , n46435 );
and ( n46437 , n46436 , n36347 );
and ( n46438 , n13181 , n43543 );
or ( n46439 , n46437 , n46438 );
and ( n46440 , n46439 , n14586 );
not ( n46441 , n37801 );
and ( n46442 , n46441 , n37746 );
xor ( n46443 , n37746 , n37305 );
xor ( n46444 , n37729 , n37305 );
xor ( n46445 , n37712 , n37305 );
xor ( n46446 , n37695 , n37305 );
and ( n46447 , n45769 , n45774 );
and ( n46448 , n46446 , n46447 );
and ( n46449 , n46445 , n46448 );
and ( n46450 , n46444 , n46449 );
xor ( n46451 , n46443 , n46450 );
and ( n46452 , n46451 , n37801 );
or ( n46453 , n46442 , n46452 );
buf ( n46454 , n46453 );
and ( n46455 , n46454 , n36348 );
and ( n46456 , n13181 , n43556 );
or ( n46457 , n46455 , n46456 );
and ( n46458 , n46457 , n14584 );
and ( n46459 , n46436 , n36347 );
and ( n46460 , n13181 , n43563 );
or ( n46461 , n46459 , n46460 );
and ( n46462 , n46461 , n37835 );
and ( n46463 , n46454 , n36347 );
and ( n46464 , n13181 , n43563 );
or ( n46465 , n46463 , n46464 );
and ( n46466 , n46465 , n37841 );
and ( n46467 , n13179 , n14564 );
and ( n46468 , n15022 , n36347 );
and ( n46469 , n13181 , n43563 );
or ( n46470 , n46468 , n46469 );
and ( n46471 , n46470 , n37847 );
or ( n46472 , n46389 , n46422 , n46440 , n46458 , n46462 , n46466 , n46467 , n46471 );
and ( n46473 , n46388 , n46472 );
and ( n46474 , n13181 , n34821 );
or ( n46475 , n46473 , n46474 );
and ( n46476 , n46475 , n16574 );
and ( n46477 , n13181 , n16576 );
or ( n46478 , n46476 , n46477 );
buf ( n46479 , n46478 );
buf ( n46480 , n46479 );
buf ( n46481 , n10613 );
not ( n46482 , n24800 );
and ( n46483 , n26323 , n25222 );
and ( n46484 , n34656 , n28589 );
and ( n46485 , n26323 , n31075 );
or ( n46486 , n46484 , n46485 );
and ( n46487 , n46486 , n28594 );
and ( n46488 , n34674 , n28589 );
and ( n46489 , n26323 , n31075 );
or ( n46490 , n46488 , n46489 );
and ( n46491 , n46490 , n30269 );
and ( n46492 , n34692 , n28589 );
and ( n46493 , n26323 , n31075 );
or ( n46494 , n46492 , n46493 );
and ( n46495 , n46494 , n30982 );
and ( n46496 , n29395 , n28589 );
and ( n46497 , n26323 , n31075 );
or ( n46498 , n46496 , n46497 );
and ( n46499 , n46498 , n30989 );
and ( n46500 , n29395 , n30991 );
and ( n46501 , n34714 , n28589 );
and ( n46502 , n26323 , n31075 );
or ( n46503 , n46501 , n46502 );
and ( n46504 , n46503 , n31002 );
or ( n46505 , n46483 , n46487 , n46491 , n46495 , n46499 , n46500 , n46504 );
and ( n46506 , n46482 , n46505 );
and ( n46507 , n26323 , n24800 );
or ( n46508 , n46506 , n46507 );
and ( n46509 , n46508 , n31008 );
and ( n46510 , n25429 , n10618 );
or ( n46511 , n46509 , n46510 );
buf ( n46512 , n46511 );
buf ( n46513 , n46512 );
not ( n46514 , n17451 );
and ( n46515 , n39499 , n21334 );
and ( n46516 , n19117 , n34492 );
or ( n46517 , n46515 , n46516 );
and ( n46518 , n46517 , n21341 );
and ( n46519 , n39509 , n21334 );
and ( n46520 , n19117 , n34492 );
or ( n46521 , n46519 , n46520 );
and ( n46522 , n46521 , n23064 );
and ( n46523 , n39519 , n21334 );
and ( n46524 , n19117 , n34492 );
or ( n46525 , n46523 , n46524 );
and ( n46526 , n46525 , n23825 );
and ( n46527 , n22062 , n21334 );
and ( n46528 , n19117 , n34492 );
or ( n46529 , n46527 , n46528 );
and ( n46530 , n46529 , n23832 );
and ( n46531 , n39529 , n21334 );
and ( n46532 , n19117 , n34492 );
or ( n46533 , n46531 , n46532 );
and ( n46534 , n46533 , n23917 );
and ( n46535 , n19117 , n34526 );
or ( n46536 , n46518 , n46522 , n46526 , n46530 , n46534 , n46535 );
and ( n46537 , n46514 , n46536 );
and ( n46538 , n19117 , n17451 );
or ( n46539 , n46537 , n46538 );
and ( n46540 , n46539 , n23924 );
and ( n46541 , n19117 , n23926 );
or ( n46542 , n46540 , n46541 );
buf ( n46543 , n46542 );
buf ( n46544 , n46543 );
buf ( n46545 , n10615 );
buf ( n46546 , n10613 );
buf ( n46547 , n10613 );
buf ( n46548 , n10615 );
not ( n46549 , n34821 );
and ( n46550 , n46418 , n36345 );
and ( n46551 , n13185 , n36352 );
or ( n46552 , n46550 , n46551 );
and ( n46553 , n46552 , n14562 );
and ( n46554 , n46436 , n36345 );
and ( n46555 , n13185 , n37073 );
or ( n46556 , n46554 , n46555 );
and ( n46557 , n46556 , n14586 );
and ( n46558 , n46454 , n36350 );
and ( n46559 , n13185 , n37825 );
or ( n46560 , n46558 , n46559 );
and ( n46561 , n46560 , n14584 );
and ( n46562 , n46436 , n36350 );
and ( n46563 , n13185 , n37831 );
or ( n46564 , n46562 , n46563 );
and ( n46565 , n46564 , n37835 );
and ( n46566 , n46454 , n36350 );
and ( n46567 , n13185 , n37831 );
or ( n46568 , n46566 , n46567 );
and ( n46569 , n46568 , n37841 );
and ( n46570 , n15022 , n36350 );
and ( n46571 , n13185 , n37831 );
or ( n46572 , n46570 , n46571 );
and ( n46573 , n46572 , n37847 );
and ( n46574 , n13185 , n37849 );
or ( n46575 , n46553 , n46557 , n46561 , n46565 , n46569 , n46573 , n46574 );
and ( n46576 , n46549 , n46575 );
and ( n46577 , n13185 , n34821 );
or ( n46578 , n46576 , n46577 );
and ( n46579 , n46578 , n16574 );
and ( n46580 , n13185 , n16576 );
or ( n46581 , n46579 , n46580 );
buf ( n46582 , n46581 );
buf ( n46583 , n46582 );
buf ( n46584 , n10613 );
not ( n46585 , n17451 );
and ( n46586 , n18771 , n17873 );
not ( n46587 , n19474 );
and ( n46588 , n46587 , n18757 );
xor ( n46589 , n19494 , n19508 );
and ( n46590 , n46589 , n19474 );
or ( n46591 , n46588 , n46590 );
buf ( n46592 , n46591 );
and ( n46593 , n46592 , n19745 );
and ( n46594 , n46592 , n19748 );
not ( n46595 , n19750 );
and ( n46596 , n46595 , n20745 );
not ( n46597 , n21193 );
and ( n46598 , n46597 , n20757 );
xor ( n46599 , n21213 , n21229 );
and ( n46600 , n46599 , n21193 );
or ( n46601 , n46598 , n46600 );
buf ( n46602 , n46601 );
and ( n46603 , n46602 , n19750 );
or ( n46604 , n46596 , n46603 );
and ( n46605 , n46604 , n21253 );
and ( n46606 , n20745 , n21255 );
or ( n46607 , n46593 , n46594 , n46605 , n46606 );
and ( n46608 , n46607 , n21336 );
and ( n46609 , n18771 , n42682 );
or ( n46610 , n46608 , n46609 );
and ( n46611 , n46610 , n21341 );
not ( n46612 , n22996 );
and ( n46613 , n46612 , n22635 );
xor ( n46614 , n23016 , n23032 );
and ( n46615 , n46614 , n22996 );
or ( n46616 , n46613 , n46615 );
buf ( n46617 , n46616 );
and ( n46618 , n46617 , n21336 );
and ( n46619 , n18771 , n42682 );
or ( n46620 , n46618 , n46619 );
and ( n46621 , n46620 , n23064 );
not ( n46622 , n23758 );
and ( n46623 , n46622 , n23397 );
xor ( n46624 , n23778 , n23794 );
and ( n46625 , n46624 , n23758 );
or ( n46626 , n46623 , n46625 );
buf ( n46627 , n46626 );
and ( n46628 , n46627 , n21336 );
and ( n46629 , n18771 , n42682 );
or ( n46630 , n46628 , n46629 );
and ( n46631 , n46630 , n23825 );
and ( n46632 , n22262 , n21336 );
and ( n46633 , n18771 , n42682 );
or ( n46634 , n46632 , n46633 );
and ( n46635 , n46634 , n23832 );
and ( n46636 , n22262 , n23834 );
xor ( n46637 , n23871 , n23894 );
buf ( n46638 , n46637 );
and ( n46639 , n46638 , n21336 );
and ( n46640 , n18771 , n42682 );
or ( n46641 , n46639 , n46640 );
and ( n46642 , n46641 , n23917 );
or ( n46643 , n46586 , n46611 , n46621 , n46631 , n46635 , n46636 , n46642 );
and ( n46644 , n46585 , n46643 );
and ( n46645 , n18771 , n17451 );
or ( n46646 , n46644 , n46645 );
and ( n46647 , n46646 , n23924 );
and ( n46648 , n17990 , n23926 );
or ( n46649 , n46647 , n46648 );
buf ( n46650 , n46649 );
buf ( n46651 , n46650 );
and ( n46652 , n16976 , n23924 );
and ( n46653 , n21852 , n23926 );
or ( n46654 , n46652 , n46653 );
buf ( n46655 , n46654 );
buf ( n46656 , n46655 );
not ( n46657 , n11333 );
and ( n46658 , n46657 , n11057 );
xor ( n46659 , n11348 , n11354 );
and ( n46660 , n46659 , n11333 );
or ( n46661 , n46658 , n46660 );
buf ( n46662 , n46661 );
buf ( n46663 , n46662 );
not ( n46664 , n34821 );
and ( n46665 , n46341 , n36347 );
and ( n46666 , n13459 , n39408 );
or ( n46667 , n46665 , n46666 );
and ( n46668 , n46667 , n14562 );
and ( n46669 , n46351 , n36348 );
and ( n46670 , n13459 , n39427 );
or ( n46671 , n46669 , n46670 );
and ( n46672 , n46671 , n14586 );
and ( n46673 , n46361 , n36347 );
and ( n46674 , n13459 , n39446 );
or ( n46675 , n46673 , n46674 );
and ( n46676 , n46675 , n14584 );
and ( n46677 , n46351 , n36348 );
and ( n46678 , n13459 , n39453 );
or ( n46679 , n46677 , n46678 );
and ( n46680 , n46679 , n37835 );
and ( n46681 , n46361 , n36348 );
and ( n46682 , n13459 , n39453 );
or ( n46683 , n46681 , n46682 );
and ( n46684 , n46683 , n37841 );
and ( n46685 , n15801 , n36348 );
and ( n46686 , n13459 , n39453 );
or ( n46687 , n46685 , n46686 );
and ( n46688 , n46687 , n37847 );
and ( n46689 , n13459 , n37849 );
or ( n46690 , n46668 , n46672 , n46676 , n46680 , n46684 , n46688 , n46689 );
and ( n46691 , n46664 , n46690 );
and ( n46692 , n13459 , n34821 );
or ( n46693 , n46691 , n46692 );
and ( n46694 , n46693 , n16574 );
and ( n46695 , n13459 , n16576 );
or ( n46696 , n46694 , n46695 );
buf ( n46697 , n46696 );
buf ( n46698 , n46697 );
not ( n46699 , n24800 );
and ( n46700 , n26019 , n25222 );
and ( n46701 , n39803 , n28583 );
and ( n46702 , n26019 , n28591 );
or ( n46703 , n46701 , n46702 );
and ( n46704 , n46703 , n28594 );
and ( n46705 , n39816 , n28583 );
and ( n46706 , n26019 , n28591 );
or ( n46707 , n46705 , n46706 );
and ( n46708 , n46707 , n30269 );
and ( n46709 , n39826 , n28583 );
and ( n46710 , n26019 , n28591 );
or ( n46711 , n46709 , n46710 );
and ( n46712 , n46711 , n30982 );
and ( n46713 , n29575 , n28583 );
and ( n46714 , n26019 , n28591 );
or ( n46715 , n46713 , n46714 );
and ( n46716 , n46715 , n30989 );
and ( n46717 , n26017 , n30991 );
and ( n46718 , n39836 , n28583 );
and ( n46719 , n26019 , n28591 );
or ( n46720 , n46718 , n46719 );
and ( n46721 , n46720 , n31002 );
or ( n46722 , n46700 , n46704 , n46708 , n46712 , n46716 , n46717 , n46721 );
and ( n46723 , n46699 , n46722 );
and ( n46724 , n26019 , n24800 );
or ( n46725 , n46723 , n46724 );
and ( n46726 , n46725 , n31008 );
and ( n46727 , n26019 , n10618 );
or ( n46728 , n46726 , n46727 );
buf ( n46729 , n46728 );
buf ( n46730 , n46729 );
buf ( n46731 , n10615 );
buf ( n46732 , n10615 );
and ( n46733 , n24246 , n31008 );
and ( n46734 , n29646 , n10618 );
or ( n46735 , n46733 , n46734 );
buf ( n46736 , n46735 );
buf ( n46737 , n46736 );
not ( n46738 , n17451 );
and ( n46739 , n19145 , n17873 );
not ( n46740 , n19474 );
and ( n46741 , n46740 , n19131 );
xor ( n46742 , n19483 , n19519 );
and ( n46743 , n46742 , n19474 );
or ( n46744 , n46741 , n46743 );
buf ( n46745 , n46744 );
and ( n46746 , n46745 , n19745 );
and ( n46747 , n46745 , n19748 );
not ( n46748 , n19750 );
and ( n46749 , n46748 , n20987 );
not ( n46750 , n21193 );
and ( n46751 , n46750 , n20999 );
xor ( n46752 , n21202 , n21240 );
and ( n46753 , n46752 , n21193 );
or ( n46754 , n46751 , n46753 );
buf ( n46755 , n46754 );
and ( n46756 , n46755 , n19750 );
or ( n46757 , n46749 , n46756 );
and ( n46758 , n46757 , n21253 );
and ( n46759 , n20987 , n21255 );
or ( n46760 , n46746 , n46747 , n46758 , n46759 );
and ( n46761 , n46760 , n21336 );
and ( n46762 , n19145 , n42682 );
or ( n46763 , n46761 , n46762 );
and ( n46764 , n46763 , n21341 );
not ( n46765 , n22996 );
and ( n46766 , n46765 , n22822 );
xor ( n46767 , n23005 , n23043 );
and ( n46768 , n46767 , n22996 );
or ( n46769 , n46766 , n46768 );
buf ( n46770 , n46769 );
and ( n46771 , n46770 , n21336 );
and ( n46772 , n19145 , n42682 );
or ( n46773 , n46771 , n46772 );
and ( n46774 , n46773 , n23064 );
not ( n46775 , n23758 );
and ( n46776 , n46775 , n23584 );
xor ( n46777 , n23767 , n23805 );
and ( n46778 , n46777 , n23758 );
or ( n46779 , n46776 , n46778 );
buf ( n46780 , n46779 );
and ( n46781 , n46780 , n21336 );
and ( n46782 , n19145 , n42682 );
or ( n46783 , n46781 , n46782 );
and ( n46784 , n46783 , n23825 );
and ( n46785 , n22042 , n21336 );
and ( n46786 , n19145 , n42682 );
or ( n46787 , n46785 , n46786 );
and ( n46788 , n46787 , n23832 );
and ( n46789 , n22042 , n23834 );
xor ( n46790 , n23849 , n23905 );
buf ( n46791 , n46790 );
and ( n46792 , n46791 , n21336 );
and ( n46793 , n19145 , n42682 );
or ( n46794 , n46792 , n46793 );
and ( n46795 , n46794 , n23917 );
or ( n46796 , n46739 , n46764 , n46774 , n46784 , n46788 , n46789 , n46795 );
and ( n46797 , n46738 , n46796 );
and ( n46798 , n19145 , n17451 );
or ( n46799 , n46797 , n46798 );
and ( n46800 , n46799 , n23924 );
and ( n46801 , n18155 , n23926 );
or ( n46802 , n46800 , n46801 );
buf ( n46803 , n46802 );
buf ( n46804 , n46803 );
not ( n46805 , n17451 );
and ( n46806 , n18773 , n17873 );
and ( n46807 , n46607 , n21330 );
and ( n46808 , n18773 , n21338 );
or ( n46809 , n46807 , n46808 );
and ( n46810 , n46809 , n21341 );
and ( n46811 , n46617 , n21330 );
and ( n46812 , n18773 , n21338 );
or ( n46813 , n46811 , n46812 );
and ( n46814 , n46813 , n23064 );
and ( n46815 , n46627 , n21330 );
and ( n46816 , n18773 , n21338 );
or ( n46817 , n46815 , n46816 );
and ( n46818 , n46817 , n23825 );
and ( n46819 , n22262 , n21330 );
and ( n46820 , n18773 , n21338 );
or ( n46821 , n46819 , n46820 );
and ( n46822 , n46821 , n23832 );
and ( n46823 , n18771 , n23834 );
and ( n46824 , n46638 , n21330 );
and ( n46825 , n18773 , n21338 );
or ( n46826 , n46824 , n46825 );
and ( n46827 , n46826 , n23917 );
or ( n46828 , n46806 , n46810 , n46814 , n46818 , n46822 , n46823 , n46827 );
and ( n46829 , n46805 , n46828 );
and ( n46830 , n18773 , n17451 );
or ( n46831 , n46829 , n46830 );
and ( n46832 , n46831 , n23924 );
and ( n46833 , n18773 , n23926 );
or ( n46834 , n46832 , n46833 );
buf ( n46835 , n46834 );
buf ( n46836 , n46835 );
not ( n46837 , n17451 );
not ( n46838 , n19474 );
and ( n46839 , n46838 , n18791 );
xor ( n46840 , n19493 , n19509 );
and ( n46841 , n46840 , n19474 );
or ( n46842 , n46839 , n46841 );
buf ( n46843 , n46842 );
and ( n46844 , n46843 , n19745 );
and ( n46845 , n46843 , n19748 );
not ( n46846 , n19750 );
and ( n46847 , n46846 , n20767 );
not ( n46848 , n21193 );
and ( n46849 , n46848 , n20779 );
xor ( n46850 , n21212 , n21230 );
and ( n46851 , n46850 , n21193 );
or ( n46852 , n46849 , n46851 );
buf ( n46853 , n46852 );
and ( n46854 , n46853 , n19750 );
or ( n46855 , n46847 , n46854 );
and ( n46856 , n46855 , n21253 );
and ( n46857 , n20767 , n21255 );
or ( n46858 , n46844 , n46845 , n46856 , n46857 );
and ( n46859 , n46858 , n21333 );
and ( n46860 , n18809 , n34758 );
or ( n46861 , n46859 , n46860 );
and ( n46862 , n46861 , n21341 );
not ( n46863 , n22996 );
and ( n46864 , n46863 , n22652 );
xor ( n46865 , n23015 , n23033 );
and ( n46866 , n46865 , n22996 );
or ( n46867 , n46864 , n46866 );
buf ( n46868 , n46867 );
and ( n46869 , n46868 , n21333 );
and ( n46870 , n18809 , n34758 );
or ( n46871 , n46869 , n46870 );
and ( n46872 , n46871 , n23064 );
not ( n46873 , n23758 );
and ( n46874 , n46873 , n23414 );
xor ( n46875 , n23777 , n23795 );
and ( n46876 , n46875 , n23758 );
or ( n46877 , n46874 , n46876 );
buf ( n46878 , n46877 );
and ( n46879 , n46878 , n21333 );
and ( n46880 , n18809 , n34758 );
or ( n46881 , n46879 , n46880 );
and ( n46882 , n46881 , n23825 );
and ( n46883 , n22242 , n21333 );
and ( n46884 , n18809 , n34758 );
or ( n46885 , n46883 , n46884 );
and ( n46886 , n46885 , n23832 );
xor ( n46887 , n23869 , n23895 );
buf ( n46888 , n46887 );
and ( n46889 , n46888 , n21333 );
and ( n46890 , n18809 , n34758 );
or ( n46891 , n46889 , n46890 );
and ( n46892 , n46891 , n23917 );
and ( n46893 , n18809 , n34526 );
or ( n46894 , n46862 , n46872 , n46882 , n46886 , n46892 , n46893 );
and ( n46895 , n46837 , n46894 );
and ( n46896 , n18809 , n17451 );
or ( n46897 , n46895 , n46896 );
and ( n46898 , n46897 , n23924 );
and ( n46899 , n18809 , n23926 );
or ( n46900 , n46898 , n46899 );
buf ( n46901 , n46900 );
buf ( n46902 , n46901 );
buf ( n46903 , n10615 );
not ( n46904 , n24511 );
not ( n46905 , n24799 );
and ( n46906 , n10700 , n40154 );
not ( n46907 , n40632 );
and ( n46908 , n46907 , n40424 );
xor ( n46909 , n40643 , n40657 );
and ( n46910 , n46909 , n40632 );
or ( n46911 , n46908 , n46910 );
buf ( n46912 , n46911 );
and ( n46913 , n46912 , n27046 );
not ( n46914 , n41147 );
and ( n46915 , n46914 , n40939 );
xor ( n46916 , n41158 , n41172 );
and ( n46917 , n46916 , n41147 );
or ( n46918 , n46915 , n46917 );
buf ( n46919 , n46918 );
and ( n46920 , n46919 , n27049 );
and ( n46921 , n29533 , n28506 );
and ( n46922 , n10700 , n28508 );
or ( n46923 , n46913 , n46920 , n46921 , n46922 );
and ( n46924 , n46923 , n41199 );
or ( n46925 , n46906 , n46924 );
and ( n46926 , n46905 , n46925 );
xor ( n46927 , n41644 , n41652 );
xor ( n46928 , n46927 , n41782 );
buf ( n46929 , n46928 );
and ( n46930 , n46929 , n27046 );
xor ( n46931 , n42195 , n42196 );
xor ( n46932 , n46931 , n42278 );
buf ( n46933 , n46932 );
and ( n46934 , n46933 , n27049 );
and ( n46935 , n29533 , n42306 );
or ( n46936 , n46930 , n46934 , n46935 );
buf ( n46937 , n46936 );
and ( n46938 , C1 , n46937 );
or ( n46939 , n46938 , C0 );
buf ( n46940 , n46939 );
not ( n46941 , n46940 );
buf ( n46942 , n46941 );
buf ( n46943 , n46942 );
not ( n46944 , n46943 );
and ( n46945 , C1 , n46944 );
or ( n46946 , n46945 , C0 );
buf ( n46947 , n46946 );
and ( n46948 , n46947 , n24799 );
or ( n46949 , n46926 , n46948 );
and ( n46950 , n46904 , n46949 );
and ( n46951 , n46923 , n24511 );
or ( n46952 , n46950 , n46951 );
and ( n46953 , n46952 , n31008 );
not ( n46954 , n42601 );
and ( n46955 , n46954 , n42429 );
xor ( n46956 , n42612 , n42626 );
and ( n46957 , n46956 , n42601 );
or ( n46958 , n46955 , n46957 );
buf ( n46959 , n46958 );
and ( n46960 , n46959 , n10618 );
or ( n46961 , n46953 , n46960 );
buf ( n46962 , n46961 );
buf ( n46963 , n46962 );
not ( n46964 , n17451 );
and ( n46965 , n46964 , n21328 );
and ( n46966 , n21304 , n17451 );
or ( n46967 , n46965 , n46966 );
and ( n46968 , n46967 , n23924 );
and ( n46969 , n21304 , n23926 );
or ( n46970 , n46968 , n46969 );
buf ( n46971 , n46970 );
buf ( n46972 , n46971 );
buf ( n46973 , n10613 );
buf ( n46974 , n10613 );
buf ( n46975 , n10613 );
buf ( n46976 , n10613 );
buf ( n46977 , n10613 );
buf ( n46978 , n10615 );
not ( n46979 , n34821 );
and ( n46980 , n13385 , n14592 );
and ( n46981 , n44916 , n36348 );
and ( n46982 , n13385 , n43530 );
or ( n46983 , n46981 , n46982 );
and ( n46984 , n46983 , n14562 );
and ( n46985 , n44926 , n36347 );
and ( n46986 , n13385 , n43543 );
or ( n46987 , n46985 , n46986 );
and ( n46988 , n46987 , n14586 );
and ( n46989 , n44936 , n36348 );
and ( n46990 , n13385 , n43556 );
or ( n46991 , n46989 , n46990 );
and ( n46992 , n46991 , n14584 );
and ( n46993 , n44926 , n36347 );
and ( n46994 , n13385 , n43563 );
or ( n46995 , n46993 , n46994 );
and ( n46996 , n46995 , n37835 );
and ( n46997 , n44936 , n36347 );
and ( n46998 , n13385 , n43563 );
or ( n46999 , n46997 , n46998 );
and ( n47000 , n46999 , n37841 );
and ( n47001 , n13383 , n14564 );
and ( n47002 , n15669 , n36347 );
and ( n47003 , n13385 , n43563 );
or ( n47004 , n47002 , n47003 );
and ( n47005 , n47004 , n37847 );
or ( n47006 , n46980 , n46984 , n46988 , n46992 , n46996 , n47000 , n47001 , n47005 );
and ( n47007 , n46979 , n47006 );
and ( n47008 , n13385 , n34821 );
or ( n47009 , n47007 , n47008 );
and ( n47010 , n47009 , n16574 );
and ( n47011 , n13385 , n16576 );
or ( n47012 , n47010 , n47011 );
buf ( n47013 , n47012 );
buf ( n47014 , n47013 );
buf ( n47015 , n10615 );
buf ( n47016 , n10615 );
not ( n47017 , n17451 );
not ( n47018 , n19474 );
and ( n47019 , n47018 , n19267 );
xor ( n47020 , n19479 , n19523 );
and ( n47021 , n47020 , n19474 );
or ( n47022 , n47019 , n47021 );
buf ( n47023 , n47022 );
and ( n47024 , n47023 , n19745 );
and ( n47025 , n47023 , n19748 );
not ( n47026 , n19750 );
and ( n47027 , n47026 , n21075 );
not ( n47028 , n21193 );
and ( n47029 , n47028 , n21087 );
xor ( n47030 , n21198 , n21244 );
and ( n47031 , n47030 , n21193 );
or ( n47032 , n47029 , n47031 );
buf ( n47033 , n47032 );
and ( n47034 , n47033 , n19750 );
or ( n47035 , n47027 , n47034 );
and ( n47036 , n47035 , n21253 );
and ( n47037 , n21075 , n21255 );
or ( n47038 , n47024 , n47025 , n47036 , n47037 );
and ( n47039 , n47038 , n21333 );
and ( n47040 , n19285 , n34758 );
or ( n47041 , n47039 , n47040 );
and ( n47042 , n47041 , n21341 );
not ( n47043 , n22996 );
and ( n47044 , n47043 , n22890 );
xor ( n47045 , n23001 , n23047 );
and ( n47046 , n47045 , n22996 );
or ( n47047 , n47044 , n47046 );
buf ( n47048 , n47047 );
and ( n47049 , n47048 , n21333 );
and ( n47050 , n19285 , n34758 );
or ( n47051 , n47049 , n47050 );
and ( n47052 , n47051 , n23064 );
not ( n47053 , n23758 );
and ( n47054 , n47053 , n23652 );
xor ( n47055 , n23763 , n23809 );
and ( n47056 , n47055 , n23758 );
or ( n47057 , n47054 , n47056 );
buf ( n47058 , n47057 );
and ( n47059 , n47058 , n21333 );
and ( n47060 , n19285 , n34758 );
or ( n47061 , n47059 , n47060 );
and ( n47062 , n47061 , n23825 );
and ( n47063 , n21945 , n21333 );
and ( n47064 , n19285 , n34758 );
or ( n47065 , n47063 , n47064 );
and ( n47066 , n47065 , n23832 );
xor ( n47067 , n23841 , n23909 );
buf ( n47068 , n47067 );
and ( n47069 , n47068 , n21333 );
and ( n47070 , n19285 , n34758 );
or ( n47071 , n47069 , n47070 );
and ( n47072 , n47071 , n23917 );
and ( n47073 , n19285 , n34526 );
or ( n47074 , n47042 , n47052 , n47062 , n47066 , n47072 , n47073 );
and ( n47075 , n47017 , n47074 );
and ( n47076 , n19285 , n17451 );
or ( n47077 , n47075 , n47076 );
and ( n47078 , n47077 , n23924 );
and ( n47079 , n19285 , n23926 );
or ( n47080 , n47078 , n47079 );
buf ( n47081 , n47080 );
buf ( n47082 , n47081 );
buf ( n47083 , n10615 );
buf ( n47084 , n10615 );
buf ( n47085 , n10615 );
and ( n47086 , n24086 , n31008 );
and ( n47087 , n29222 , n10618 );
or ( n47088 , n47086 , n47087 );
buf ( n47089 , n47088 );
buf ( n47090 , n47089 );
buf ( n47091 , n10613 );
buf ( n47092 , n10615 );
buf ( n47093 , n10615 );
not ( n47094 , n34821 );
and ( n47095 , n43688 , n36347 );
and ( n47096 , n13351 , n39408 );
or ( n47097 , n47095 , n47096 );
and ( n47098 , n47097 , n14562 );
and ( n47099 , n43700 , n36348 );
and ( n47100 , n13351 , n39427 );
or ( n47101 , n47099 , n47100 );
and ( n47102 , n47101 , n14586 );
and ( n47103 , n43712 , n36347 );
and ( n47104 , n13351 , n39446 );
or ( n47105 , n47103 , n47104 );
and ( n47106 , n47105 , n14584 );
and ( n47107 , n43700 , n36348 );
and ( n47108 , n13351 , n39453 );
or ( n47109 , n47107 , n47108 );
and ( n47110 , n47109 , n37835 );
and ( n47111 , n43712 , n36348 );
and ( n47112 , n13351 , n39453 );
or ( n47113 , n47111 , n47112 );
and ( n47114 , n47113 , n37841 );
and ( n47115 , n15603 , n36348 );
and ( n47116 , n13351 , n39453 );
or ( n47117 , n47115 , n47116 );
and ( n47118 , n47117 , n37847 );
and ( n47119 , n13351 , n37849 );
or ( n47120 , n47098 , n47102 , n47106 , n47110 , n47114 , n47118 , n47119 );
and ( n47121 , n47094 , n47120 );
and ( n47122 , n13351 , n34821 );
or ( n47123 , n47121 , n47122 );
and ( n47124 , n47123 , n16574 );
and ( n47125 , n13351 , n16576 );
or ( n47126 , n47124 , n47125 );
buf ( n47127 , n47126 );
buf ( n47128 , n47127 );
not ( n47129 , n11333 );
and ( n47130 , n47129 , n11176 );
xor ( n47131 , n11341 , n11361 );
and ( n47132 , n47131 , n11333 );
or ( n47133 , n47130 , n47132 );
buf ( n47134 , n47133 );
buf ( n47135 , n47134 );
buf ( n47136 , n10615 );
buf ( n47137 , n10613 );
buf ( n47138 , n10615 );
not ( n47139 , n34821 );
and ( n47140 , n13335 , n14592 );
and ( n47141 , n43617 , n36350 );
and ( n47142 , n13335 , n43691 );
or ( n47143 , n47141 , n47142 );
and ( n47144 , n47143 , n14562 );
and ( n47145 , n43627 , n36350 );
and ( n47146 , n13335 , n43703 );
or ( n47147 , n47145 , n47146 );
and ( n47148 , n47147 , n14586 );
and ( n47149 , n43637 , n36345 );
and ( n47150 , n13335 , n43715 );
or ( n47151 , n47149 , n47150 );
and ( n47152 , n47151 , n14584 );
and ( n47153 , n43627 , n36345 );
and ( n47154 , n13335 , n43721 );
or ( n47155 , n47153 , n47154 );
and ( n47156 , n47155 , n37835 );
and ( n47157 , n43637 , n36345 );
and ( n47158 , n13335 , n43721 );
or ( n47159 , n47157 , n47158 );
and ( n47160 , n47159 , n37841 );
and ( n47161 , n15581 , n14564 );
and ( n47162 , n15581 , n36345 );
and ( n47163 , n13335 , n43721 );
or ( n47164 , n47162 , n47163 );
and ( n47165 , n47164 , n37847 );
or ( n47166 , n47140 , n47144 , n47148 , n47152 , n47156 , n47160 , n47161 , n47165 );
and ( n47167 , n47139 , n47166 );
and ( n47168 , n13335 , n34821 );
or ( n47169 , n47167 , n47168 );
and ( n47170 , n47169 , n16574 );
and ( n47171 , n12294 , n16576 );
or ( n47172 , n47170 , n47171 );
buf ( n47173 , n47172 );
buf ( n47174 , n47173 );
buf ( n47175 , n10613 );
not ( n47176 , n24800 );
and ( n47177 , n28510 , n28587 );
and ( n47178 , n25892 , n39807 );
or ( n47179 , n47177 , n47178 );
and ( n47180 , n47179 , n28594 );
and ( n47181 , n30258 , n28587 );
and ( n47182 , n25892 , n39807 );
or ( n47183 , n47181 , n47182 );
and ( n47184 , n47183 , n30269 );
and ( n47185 , n30972 , n28587 );
and ( n47186 , n25892 , n39807 );
or ( n47187 , n47185 , n47186 );
and ( n47188 , n47187 , n30982 );
and ( n47189 , n29655 , n28587 );
and ( n47190 , n25892 , n39807 );
or ( n47191 , n47189 , n47190 );
and ( n47192 , n47191 , n30989 );
and ( n47193 , n30998 , n28587 );
and ( n47194 , n25892 , n39807 );
or ( n47195 , n47193 , n47194 );
and ( n47196 , n47195 , n31002 );
and ( n47197 , n25892 , n34607 );
or ( n47198 , n47180 , n47184 , n47188 , n47192 , n47196 , n47197 );
and ( n47199 , n47176 , n47198 );
and ( n47200 , n25892 , n24800 );
or ( n47201 , n47199 , n47200 );
and ( n47202 , n47201 , n31008 );
and ( n47203 , n25892 , n10618 );
or ( n47204 , n47202 , n47203 );
buf ( n47205 , n47204 );
buf ( n47206 , n47205 );
not ( n47207 , n34821 );
not ( n47208 , n14139 );
and ( n47209 , n47208 , n35633 );
or ( n47210 , n47209 , C0 );
and ( n47211 , n47210 , n14140 );
and ( n47212 , n35633 , n14141 );
or ( n47213 , C0 , C0 , n47211 , n47212 );
and ( n47214 , n47213 , n36347 );
and ( n47215 , n13144 , n39408 );
or ( n47216 , n47214 , n47215 );
and ( n47217 , n47216 , n14562 );
and ( n47218 , n13144 , n39427 );
or ( n47219 , C0 , n47218 );
and ( n47220 , n47219 , n14586 );
and ( n47221 , n13144 , n39446 );
or ( n47222 , C0 , n47221 );
and ( n47223 , n47222 , n14584 );
and ( n47224 , n13144 , n39453 );
or ( n47225 , C0 , n47224 );
and ( n47226 , n47225 , n37835 );
and ( n47227 , n13144 , n39453 );
or ( n47228 , C0 , n47227 );
and ( n47229 , n47228 , n37841 );
and ( n47230 , n14934 , n36348 );
and ( n47231 , n13144 , n39453 );
or ( n47232 , n47230 , n47231 );
and ( n47233 , n47232 , n37847 );
and ( n47234 , n13144 , n37849 );
or ( n47235 , n47217 , n47220 , n47223 , n47226 , n47229 , n47233 , n47234 );
and ( n47236 , n47207 , n47235 );
and ( n47237 , n13144 , n34821 );
or ( n47238 , n47236 , n47237 );
and ( n47239 , n47238 , n16574 );
and ( n47240 , n13144 , n16576 );
or ( n47241 , n47239 , n47240 );
buf ( n47242 , n47241 );
buf ( n47243 , n47242 );
not ( n47244 , n34804 );
and ( n47245 , n47244 , n26263 );
and ( n47246 , n14761 , n34804 );
or ( n47247 , n47245 , n47246 );
and ( n47248 , n47247 , n31008 );
and ( n47249 , n14761 , n10618 );
or ( n47250 , n47248 , n47249 );
buf ( n47251 , n47250 );
buf ( n47252 , n47251 );
buf ( n47253 , n10613 );
buf ( n47254 , n10613 );
buf ( n47255 , n10615 );
buf ( n47256 , n10615 );
buf ( n47257 , n10615 );
buf ( n47258 , n10615 );
buf ( n47259 , n10615 );
buf ( n47260 , n10613 );
buf ( n47261 , n10615 );
buf ( n47262 , n10613 );
buf ( n47263 , n10615 );
buf ( n47264 , n10615 );
buf ( n47265 , n10613 );
buf ( n47266 , n10615 );
buf ( n47267 , n10615 );
and ( n47268 , n24110 , n31008 );
and ( n47269 , n29306 , n10618 );
or ( n47270 , n47268 , n47269 );
buf ( n47271 , n47270 );
buf ( n47272 , n47271 );
buf ( n47273 , n10613 );
not ( n47274 , n17451 );
and ( n47275 , n18907 , n17873 );
and ( n47276 , n43338 , n21336 );
and ( n47277 , n18907 , n42682 );
or ( n47278 , n47276 , n47277 );
and ( n47279 , n47278 , n21341 );
and ( n47280 , n43348 , n21336 );
and ( n47281 , n18907 , n42682 );
or ( n47282 , n47280 , n47281 );
and ( n47283 , n47282 , n23064 );
and ( n47284 , n43358 , n21336 );
and ( n47285 , n18907 , n42682 );
or ( n47286 , n47284 , n47285 );
and ( n47287 , n47286 , n23825 );
and ( n47288 , n22182 , n21336 );
and ( n47289 , n18907 , n42682 );
or ( n47290 , n47288 , n47289 );
and ( n47291 , n47290 , n23832 );
and ( n47292 , n22182 , n23834 );
and ( n47293 , n43368 , n21336 );
and ( n47294 , n18907 , n42682 );
or ( n47295 , n47293 , n47294 );
and ( n47296 , n47295 , n23917 );
or ( n47297 , n47275 , n47279 , n47283 , n47287 , n47291 , n47292 , n47296 );
and ( n47298 , n47274 , n47297 );
and ( n47299 , n18907 , n17451 );
or ( n47300 , n47298 , n47299 );
and ( n47301 , n47300 , n23924 );
and ( n47302 , n18050 , n23926 );
or ( n47303 , n47301 , n47302 );
buf ( n47304 , n47303 );
buf ( n47305 , n47304 );
not ( n47306 , n17451 );
and ( n47307 , n34421 , n21334 );
and ( n47308 , n19219 , n34492 );
or ( n47309 , n47307 , n47308 );
and ( n47310 , n47309 , n21341 );
and ( n47311 , n34431 , n21334 );
and ( n47312 , n19219 , n34492 );
or ( n47313 , n47311 , n47312 );
and ( n47314 , n47313 , n23064 );
and ( n47315 , n34441 , n21334 );
and ( n47316 , n19219 , n34492 );
or ( n47317 , n47315 , n47316 );
and ( n47318 , n47317 , n23825 );
and ( n47319 , n21971 , n21334 );
and ( n47320 , n19219 , n34492 );
or ( n47321 , n47319 , n47320 );
and ( n47322 , n47321 , n23832 );
and ( n47323 , n34452 , n21334 );
and ( n47324 , n19219 , n34492 );
or ( n47325 , n47323 , n47324 );
and ( n47326 , n47325 , n23917 );
and ( n47327 , n19219 , n34526 );
or ( n47328 , n47310 , n47314 , n47318 , n47322 , n47326 , n47327 );
and ( n47329 , n47306 , n47328 );
and ( n47330 , n19219 , n17451 );
or ( n47331 , n47329 , n47330 );
and ( n47332 , n47331 , n23924 );
and ( n47333 , n19219 , n23926 );
or ( n47334 , n47332 , n47333 );
buf ( n47335 , n47334 );
buf ( n47336 , n47335 );
buf ( n47337 , n10615 );
buf ( n47338 , n10613 );
buf ( n47339 , n10615 );
buf ( n47340 , n10613 );
not ( n47341 , n17451 );
and ( n47342 , n18635 , n17873 );
not ( n47343 , n19474 );
and ( n47344 , n47343 , n18622 );
xor ( n47345 , n19498 , n19504 );
and ( n47346 , n47345 , n19474 );
or ( n47347 , n47344 , n47346 );
buf ( n47348 , n47347 );
and ( n47349 , n47348 , n19745 );
and ( n47350 , n47348 , n19748 );
not ( n47351 , n19750 );
and ( n47352 , n47351 , n20657 );
not ( n47353 , n21193 );
and ( n47354 , n47353 , n20669 );
xor ( n47355 , n21217 , n21225 );
and ( n47356 , n47355 , n21193 );
or ( n47357 , n47354 , n47356 );
buf ( n47358 , n47357 );
and ( n47359 , n47358 , n19750 );
or ( n47360 , n47352 , n47359 );
and ( n47361 , n47360 , n21253 );
and ( n47362 , n20657 , n21255 );
or ( n47363 , n47349 , n47350 , n47361 , n47362 );
and ( n47364 , n47363 , n21336 );
and ( n47365 , n18635 , n42682 );
or ( n47366 , n47364 , n47365 );
and ( n47367 , n47366 , n21341 );
not ( n47368 , n22996 );
and ( n47369 , n47368 , n22567 );
xor ( n47370 , n23020 , n23028 );
and ( n47371 , n47370 , n22996 );
or ( n47372 , n47369 , n47371 );
buf ( n47373 , n47372 );
and ( n47374 , n47373 , n21336 );
and ( n47375 , n18635 , n42682 );
or ( n47376 , n47374 , n47375 );
and ( n47377 , n47376 , n23064 );
not ( n47378 , n23758 );
and ( n47379 , n47378 , n23329 );
xor ( n47380 , n23782 , n23790 );
and ( n47381 , n47380 , n23758 );
or ( n47382 , n47379 , n47381 );
buf ( n47383 , n47382 );
and ( n47384 , n47383 , n21336 );
and ( n47385 , n18635 , n42682 );
or ( n47386 , n47384 , n47385 );
and ( n47387 , n47386 , n23825 );
and ( n47388 , n22342 , n21336 );
and ( n47389 , n18635 , n42682 );
or ( n47390 , n47388 , n47389 );
and ( n47391 , n47390 , n23832 );
and ( n47392 , n22342 , n23834 );
xor ( n47393 , n23879 , n23890 );
buf ( n47394 , n47393 );
and ( n47395 , n47394 , n21336 );
and ( n47396 , n18635 , n42682 );
or ( n47397 , n47395 , n47396 );
and ( n47398 , n47397 , n23917 );
or ( n47399 , n47342 , n47367 , n47377 , n47387 , n47391 , n47392 , n47398 );
and ( n47400 , n47341 , n47399 );
and ( n47401 , n18635 , n17451 );
or ( n47402 , n47400 , n47401 );
and ( n47403 , n47402 , n23924 );
and ( n47404 , n17930 , n23926 );
or ( n47405 , n47403 , n47404 );
buf ( n47406 , n47405 );
buf ( n47407 , n47406 );
not ( n47408 , n17451 );
and ( n47409 , n19247 , n17873 );
not ( n47410 , n19474 );
and ( n47411 , n47410 , n19233 );
xor ( n47412 , n19480 , n19522 );
and ( n47413 , n47412 , n19474 );
or ( n47414 , n47411 , n47413 );
buf ( n47415 , n47414 );
and ( n47416 , n47415 , n19745 );
and ( n47417 , n47415 , n19748 );
not ( n47418 , n19750 );
and ( n47419 , n47418 , n21053 );
not ( n47420 , n21193 );
and ( n47421 , n47420 , n21065 );
xor ( n47422 , n21199 , n21243 );
and ( n47423 , n47422 , n21193 );
or ( n47424 , n47421 , n47423 );
buf ( n47425 , n47424 );
and ( n47426 , n47425 , n19750 );
or ( n47427 , n47419 , n47426 );
and ( n47428 , n47427 , n21253 );
and ( n47429 , n21053 , n21255 );
or ( n47430 , n47416 , n47417 , n47428 , n47429 );
and ( n47431 , n47430 , n21336 );
and ( n47432 , n19247 , n42682 );
or ( n47433 , n47431 , n47432 );
and ( n47434 , n47433 , n21341 );
not ( n47435 , n22996 );
and ( n47436 , n47435 , n22873 );
xor ( n47437 , n23002 , n23046 );
and ( n47438 , n47437 , n22996 );
or ( n47439 , n47436 , n47438 );
buf ( n47440 , n47439 );
and ( n47441 , n47440 , n21336 );
and ( n47442 , n19247 , n42682 );
or ( n47443 , n47441 , n47442 );
and ( n47444 , n47443 , n23064 );
not ( n47445 , n23758 );
and ( n47446 , n47445 , n23635 );
xor ( n47447 , n23764 , n23808 );
and ( n47448 , n47447 , n23758 );
or ( n47449 , n47446 , n47448 );
buf ( n47450 , n47449 );
and ( n47451 , n47450 , n21336 );
and ( n47452 , n19247 , n42682 );
or ( n47453 , n47451 , n47452 );
and ( n47454 , n47453 , n23825 );
and ( n47455 , n21958 , n21336 );
and ( n47456 , n19247 , n42682 );
or ( n47457 , n47455 , n47456 );
and ( n47458 , n47457 , n23832 );
and ( n47459 , n21958 , n23834 );
xor ( n47460 , n23843 , n23908 );
buf ( n47461 , n47460 );
and ( n47462 , n47461 , n21336 );
and ( n47463 , n19247 , n42682 );
or ( n47464 , n47462 , n47463 );
and ( n47465 , n47464 , n23917 );
or ( n47466 , n47409 , n47434 , n47444 , n47454 , n47458 , n47459 , n47465 );
and ( n47467 , n47408 , n47466 );
and ( n47468 , n19247 , n17451 );
or ( n47469 , n47467 , n47468 );
and ( n47470 , n47469 , n23924 );
and ( n47471 , n18200 , n23926 );
or ( n47472 , n47470 , n47471 );
buf ( n47473 , n47472 );
buf ( n47474 , n47473 );
buf ( n47475 , n10615 );
buf ( n47476 , n10615 );
buf ( n47477 , n10615 );
not ( n47478 , n24800 );
and ( n47479 , n26493 , n25222 );
not ( n47480 , n26823 );
and ( n47481 , n47480 , n26479 );
xor ( n47482 , n42829 , n42832 );
and ( n47483 , n47482 , n26823 );
or ( n47484 , n47481 , n47483 );
buf ( n47485 , n47484 );
and ( n47486 , n47485 , n27046 );
and ( n47487 , n47485 , n27049 );
not ( n47488 , n27051 );
and ( n47489 , n47488 , n28280 );
not ( n47490 , n28494 );
and ( n47491 , n47490 , n28292 );
xor ( n47492 , n42849 , n42852 );
and ( n47493 , n47492 , n28494 );
or ( n47494 , n47491 , n47493 );
buf ( n47495 , n47494 );
and ( n47496 , n47495 , n27051 );
or ( n47497 , n47489 , n47496 );
and ( n47498 , n47497 , n28506 );
and ( n47499 , n28280 , n28508 );
or ( n47500 , n47486 , n47487 , n47498 , n47499 );
and ( n47501 , n47500 , n28589 );
and ( n47502 , n26493 , n31075 );
or ( n47503 , n47501 , n47502 );
and ( n47504 , n47503 , n28594 );
not ( n47505 , n30249 );
and ( n47506 , n47505 , n30075 );
xor ( n47507 , n42874 , n42877 );
and ( n47508 , n47507 , n30249 );
or ( n47509 , n47506 , n47508 );
buf ( n47510 , n47509 );
and ( n47511 , n47510 , n28589 );
and ( n47512 , n26493 , n31075 );
or ( n47513 , n47511 , n47512 );
and ( n47514 , n47513 , n30269 );
not ( n47515 , n30963 );
and ( n47516 , n47515 , n30789 );
xor ( n47517 , n42894 , n42897 );
and ( n47518 , n47517 , n30963 );
or ( n47519 , n47516 , n47518 );
buf ( n47520 , n47519 );
and ( n47521 , n47520 , n28589 );
and ( n47522 , n26493 , n31075 );
or ( n47523 , n47521 , n47522 );
and ( n47524 , n47523 , n30982 );
and ( n47525 , n29295 , n28589 );
and ( n47526 , n26493 , n31075 );
or ( n47527 , n47525 , n47526 );
and ( n47528 , n47527 , n30989 );
and ( n47529 , n29295 , n30991 );
xor ( n47530 , n42920 , n42924 );
buf ( n47531 , n47530 );
and ( n47532 , n47531 , n28589 );
and ( n47533 , n26493 , n31075 );
or ( n47534 , n47532 , n47533 );
and ( n47535 , n47534 , n31002 );
or ( n47536 , n47479 , n47504 , n47514 , n47524 , n47528 , n47529 , n47535 );
and ( n47537 , n47478 , n47536 );
and ( n47538 , n26493 , n24800 );
or ( n47539 , n47537 , n47538 );
and ( n47540 , n47539 , n31008 );
and ( n47541 , n25504 , n10618 );
or ( n47542 , n47540 , n47541 );
buf ( n47543 , n47542 );
buf ( n47544 , n47543 );
buf ( n47545 , n10613 );
buf ( n47546 , n10615 );
buf ( n47547 , n10613 );
not ( n47548 , n24800 );
and ( n47549 , n26801 , n25222 );
and ( n47550 , n45258 , n28583 );
and ( n47551 , n26801 , n28591 );
or ( n47552 , n47550 , n47551 );
and ( n47553 , n47552 , n28594 );
and ( n47554 , n45274 , n28583 );
and ( n47555 , n26801 , n28591 );
or ( n47556 , n47554 , n47555 );
and ( n47557 , n47556 , n30269 );
and ( n47558 , n45290 , n28583 );
and ( n47559 , n26801 , n28591 );
or ( n47560 , n47558 , n47559 );
and ( n47561 , n47560 , n30982 );
and ( n47562 , n29133 , n28583 );
and ( n47563 , n26801 , n28591 );
or ( n47564 , n47562 , n47563 );
and ( n47565 , n47564 , n30989 );
and ( n47566 , n26799 , n30991 );
and ( n47567 , n45310 , n28583 );
and ( n47568 , n26801 , n28591 );
or ( n47569 , n47567 , n47568 );
and ( n47570 , n47569 , n31002 );
or ( n47571 , n47549 , n47553 , n47557 , n47561 , n47565 , n47566 , n47570 );
and ( n47572 , n47548 , n47571 );
and ( n47573 , n26801 , n24800 );
or ( n47574 , n47572 , n47573 );
and ( n47575 , n47574 , n31008 );
and ( n47576 , n26801 , n10618 );
or ( n47577 , n47575 , n47576 );
buf ( n47578 , n47577 );
buf ( n47579 , n47578 );
buf ( n47580 , n10613 );
buf ( n47581 , n10615 );
buf ( n47582 , n10613 );
buf ( n47583 , n10613 );
buf ( n47584 , n10615 );
buf ( n47585 , n10615 );
buf ( n47586 , n10615 );
not ( n47587 , n24800 );
and ( n47588 , n45258 , n28586 );
and ( n47589 , n26803 , n34573 );
or ( n47590 , n47588 , n47589 );
and ( n47591 , n47590 , n28594 );
and ( n47592 , n45274 , n28586 );
and ( n47593 , n26803 , n34573 );
or ( n47594 , n47592 , n47593 );
and ( n47595 , n47594 , n30269 );
and ( n47596 , n45290 , n28586 );
and ( n47597 , n26803 , n34573 );
or ( n47598 , n47596 , n47597 );
and ( n47599 , n47598 , n30982 );
and ( n47600 , n29133 , n28586 );
and ( n47601 , n26803 , n34573 );
or ( n47602 , n47600 , n47601 );
and ( n47603 , n47602 , n30989 );
and ( n47604 , n45310 , n28586 );
and ( n47605 , n26803 , n34573 );
or ( n47606 , n47604 , n47605 );
and ( n47607 , n47606 , n31002 );
and ( n47608 , n26803 , n34607 );
or ( n47609 , n47591 , n47595 , n47599 , n47603 , n47607 , n47608 );
and ( n47610 , n47587 , n47609 );
and ( n47611 , n26803 , n24800 );
or ( n47612 , n47610 , n47611 );
and ( n47613 , n47612 , n31008 );
and ( n47614 , n26803 , n10618 );
or ( n47615 , n47613 , n47614 );
buf ( n47616 , n47615 );
buf ( n47617 , n47616 );
buf ( n47618 , n10615 );
buf ( n47619 , n10613 );
buf ( n47620 , n10613 );
not ( n47621 , n24800 );
not ( n47622 , n26823 );
and ( n47623 , n47622 , n26445 );
xor ( n47624 , n42830 , n42831 );
and ( n47625 , n47624 , n26823 );
or ( n47626 , n47623 , n47625 );
buf ( n47627 , n47626 );
and ( n47628 , n47627 , n27046 );
and ( n47629 , n47627 , n27049 );
not ( n47630 , n27051 );
and ( n47631 , n47630 , n28258 );
not ( n47632 , n28494 );
and ( n47633 , n47632 , n28270 );
xor ( n47634 , n42850 , n42851 );
and ( n47635 , n47634 , n28494 );
or ( n47636 , n47633 , n47635 );
buf ( n47637 , n47636 );
and ( n47638 , n47637 , n27051 );
or ( n47639 , n47631 , n47638 );
and ( n47640 , n47639 , n28506 );
and ( n47641 , n28258 , n28508 );
or ( n47642 , n47628 , n47629 , n47640 , n47641 );
and ( n47643 , n47642 , n28587 );
and ( n47644 , n26465 , n39807 );
or ( n47645 , n47643 , n47644 );
and ( n47646 , n47645 , n28594 );
not ( n47647 , n30249 );
and ( n47648 , n47647 , n30058 );
xor ( n47649 , n42875 , n42876 );
and ( n47650 , n47649 , n30249 );
or ( n47651 , n47648 , n47650 );
buf ( n47652 , n47651 );
and ( n47653 , n47652 , n28587 );
and ( n47654 , n26465 , n39807 );
or ( n47655 , n47653 , n47654 );
and ( n47656 , n47655 , n30269 );
not ( n47657 , n30963 );
and ( n47658 , n47657 , n30772 );
xor ( n47659 , n42895 , n42896 );
and ( n47660 , n47659 , n30963 );
or ( n47661 , n47658 , n47660 );
buf ( n47662 , n47661 );
and ( n47663 , n47662 , n28587 );
and ( n47664 , n26465 , n39807 );
or ( n47665 , n47663 , n47664 );
and ( n47666 , n47665 , n30982 );
and ( n47667 , n29315 , n28587 );
and ( n47668 , n26465 , n39807 );
or ( n47669 , n47667 , n47668 );
and ( n47670 , n47669 , n30989 );
xor ( n47671 , n42922 , n42923 );
buf ( n47672 , n47671 );
and ( n47673 , n47672 , n28587 );
and ( n47674 , n26465 , n39807 );
or ( n47675 , n47673 , n47674 );
and ( n47676 , n47675 , n31002 );
and ( n47677 , n26465 , n34607 );
or ( n47678 , n47646 , n47656 , n47666 , n47670 , n47676 , n47677 );
and ( n47679 , n47621 , n47678 );
and ( n47680 , n26465 , n24800 );
or ( n47681 , n47679 , n47680 );
and ( n47682 , n47681 , n31008 );
and ( n47683 , n26465 , n10618 );
or ( n47684 , n47682 , n47683 );
buf ( n47685 , n47684 );
buf ( n47686 , n47685 );
buf ( n47687 , n10613 );
buf ( n47688 , n10613 );
buf ( n47689 , n10615 );
buf ( n47690 , n10615 );
buf ( n47691 , n10613 );
buf ( n47692 , n10613 );
buf ( n47693 , n10615 );
buf ( n47694 , n10615 );
not ( n47695 , n34804 );
and ( n47696 , n47695 , n26603 );
and ( n47697 , n14701 , n34804 );
or ( n47698 , n47696 , n47697 );
and ( n47699 , n47698 , n31008 );
and ( n47700 , n14701 , n10618 );
or ( n47701 , n47699 , n47700 );
buf ( n47702 , n47701 );
buf ( n47703 , n47702 );
buf ( n47704 , n10615 );
buf ( n47705 , n10613 );
buf ( n47706 , n10613 );
buf ( n47707 , n10613 );
buf ( n47708 , n10613 );
buf ( n47709 , n10613 );
not ( n47710 , n34821 );
and ( n47711 , n14958 , n14592 );
not ( n47712 , n13916 );
and ( n47713 , n47712 , n13551 );
xor ( n47714 , n13552 , n13883 );
and ( n47715 , n47714 , n13916 );
or ( n47716 , n47713 , n47715 );
buf ( n47717 , n47716 );
and ( n47718 , n47717 , n14137 );
and ( n47719 , n47717 , n14143 );
not ( n47720 , n14139 );
not ( n47721 , n34833 );
buf ( n47722 , n35286 );
and ( n47723 , n47721 , n47722 );
xor ( n47724 , n35288 , n35626 );
buf ( n47725 , n47724 );
and ( n47726 , n47725 , n34833 );
or ( n47727 , n47723 , n47726 );
buf ( n47728 , n47727 );
and ( n47729 , n47720 , n47728 );
xor ( n47730 , n36241 , n35634 );
xor ( n47731 , n36219 , n35634 );
and ( n47732 , n46402 , n46409 );
and ( n47733 , n47731 , n47732 );
and ( n47734 , n47730 , n47733 );
buf ( n47735 , n47734 );
and ( n47736 , n47735 , n36245 );
or ( n47737 , C0 , n47736 );
buf ( n47738 , n47737 );
and ( n47739 , n47738 , n14139 );
or ( n47740 , n47729 , n47739 );
and ( n47741 , n47740 , n14140 );
and ( n47742 , n47728 , n14141 );
or ( n47743 , n47718 , n47719 , n47741 , n47742 );
and ( n47744 , n47743 , n36348 );
and ( n47745 , n14958 , n43530 );
or ( n47746 , n47744 , n47745 );
and ( n47747 , n47746 , n14562 );
not ( n47748 , n37048 );
and ( n47749 , n47748 , n37044 );
xor ( n47750 , n37044 , n36552 );
xor ( n47751 , n37027 , n36552 );
xor ( n47752 , n37010 , n36552 );
and ( n47753 , n46425 , n46432 );
and ( n47754 , n47752 , n47753 );
and ( n47755 , n47751 , n47754 );
xor ( n47756 , n47750 , n47755 );
and ( n47757 , n47756 , n37048 );
or ( n47758 , n47749 , n47757 );
buf ( n47759 , n47758 );
and ( n47760 , n47759 , n36347 );
and ( n47761 , n14958 , n43543 );
or ( n47762 , n47760 , n47761 );
and ( n47763 , n47762 , n14586 );
not ( n47764 , n37801 );
and ( n47765 , n47764 , n37797 );
xor ( n47766 , n37797 , n37305 );
xor ( n47767 , n37780 , n37305 );
xor ( n47768 , n37763 , n37305 );
and ( n47769 , n46443 , n46450 );
and ( n47770 , n47768 , n47769 );
and ( n47771 , n47767 , n47770 );
xor ( n47772 , n47766 , n47771 );
and ( n47773 , n47772 , n37801 );
or ( n47774 , n47765 , n47773 );
buf ( n47775 , n47774 );
and ( n47776 , n47775 , n36348 );
and ( n47777 , n14958 , n43556 );
or ( n47778 , n47776 , n47777 );
and ( n47779 , n47778 , n14584 );
and ( n47780 , n47759 , n36347 );
and ( n47781 , n14958 , n43563 );
or ( n47782 , n47780 , n47781 );
and ( n47783 , n47782 , n37835 );
and ( n47784 , n47775 , n36347 );
and ( n47785 , n14958 , n43563 );
or ( n47786 , n47784 , n47785 );
and ( n47787 , n47786 , n37841 );
and ( n47788 , n14956 , n14564 );
and ( n47789 , n14977 , n36347 );
and ( n47790 , n14958 , n43563 );
or ( n47791 , n47789 , n47790 );
and ( n47792 , n47791 , n37847 );
or ( n47793 , n47711 , n47747 , n47763 , n47779 , n47783 , n47787 , n47788 , n47792 );
and ( n47794 , n47710 , n47793 );
and ( n47795 , n14958 , n34821 );
or ( n47796 , n47794 , n47795 );
and ( n47797 , n47796 , n16574 );
and ( n47798 , n14958 , n16576 );
or ( n47799 , n47797 , n47798 );
buf ( n47800 , n47799 );
buf ( n47801 , n47800 );
buf ( n47802 , n10615 );
and ( n47803 , n17024 , n23924 );
and ( n47804 , n21930 , n23926 );
or ( n47805 , n47803 , n47804 );
buf ( n47806 , n47805 );
buf ( n47807 , n47806 );
not ( n47808 , n34821 );
and ( n47809 , n44175 , n36347 );
and ( n47810 , n13476 , n39408 );
or ( n47811 , n47809 , n47810 );
and ( n47812 , n47811 , n14562 );
and ( n47813 , n44185 , n36348 );
and ( n47814 , n13476 , n39427 );
or ( n47815 , n47813 , n47814 );
and ( n47816 , n47815 , n14586 );
and ( n47817 , n44195 , n36347 );
and ( n47818 , n13476 , n39446 );
or ( n47819 , n47817 , n47818 );
and ( n47820 , n47819 , n14584 );
and ( n47821 , n44185 , n36348 );
and ( n47822 , n13476 , n39453 );
or ( n47823 , n47821 , n47822 );
and ( n47824 , n47823 , n37835 );
and ( n47825 , n44195 , n36348 );
and ( n47826 , n13476 , n39453 );
or ( n47827 , n47825 , n47826 );
and ( n47828 , n47827 , n37841 );
and ( n47829 , n15823 , n36348 );
and ( n47830 , n13476 , n39453 );
or ( n47831 , n47829 , n47830 );
and ( n47832 , n47831 , n37847 );
and ( n47833 , n13476 , n37849 );
or ( n47834 , n47812 , n47816 , n47820 , n47824 , n47828 , n47832 , n47833 );
and ( n47835 , n47808 , n47834 );
and ( n47836 , n13476 , n34821 );
or ( n47837 , n47835 , n47836 );
and ( n47838 , n47837 , n16574 );
and ( n47839 , n13476 , n16576 );
or ( n47840 , n47838 , n47839 );
buf ( n47841 , n47840 );
buf ( n47842 , n47841 );
not ( n47843 , n24800 );
and ( n47844 , n39944 , n28587 );
and ( n47845 , n25860 , n39807 );
or ( n47846 , n47844 , n47845 );
and ( n47847 , n47846 , n28594 );
and ( n47848 , n39954 , n28587 );
and ( n47849 , n25860 , n39807 );
or ( n47850 , n47848 , n47849 );
and ( n47851 , n47850 , n30269 );
and ( n47852 , n39964 , n28587 );
and ( n47853 , n25860 , n39807 );
or ( n47854 , n47852 , n47853 );
and ( n47855 , n47854 , n30982 );
and ( n47856 , n28892 , n28587 );
and ( n47857 , n25860 , n39807 );
or ( n47858 , n47856 , n47857 );
and ( n47859 , n47858 , n30989 );
and ( n47860 , n39974 , n28587 );
and ( n47861 , n25860 , n39807 );
or ( n47862 , n47860 , n47861 );
and ( n47863 , n47862 , n31002 );
and ( n47864 , n25860 , n34607 );
or ( n47865 , n47847 , n47851 , n47855 , n47859 , n47863 , n47864 );
and ( n47866 , n47843 , n47865 );
and ( n47867 , n25860 , n24800 );
or ( n47868 , n47866 , n47867 );
and ( n47869 , n47868 , n31008 );
and ( n47870 , n25860 , n10618 );
or ( n47871 , n47869 , n47870 );
buf ( n47872 , n47871 );
buf ( n47873 , n47872 );
buf ( n47874 , n10615 );
buf ( n47875 , n10615 );
buf ( n47876 , n10615 );
buf ( n47877 , n10615 );
buf ( n47878 , n10615 );
not ( n47879 , n24800 );
and ( n47880 , n42864 , n28587 );
and ( n47881 , n26601 , n39807 );
or ( n47882 , n47880 , n47881 );
and ( n47883 , n47882 , n28594 );
and ( n47884 , n42884 , n28587 );
and ( n47885 , n26601 , n39807 );
or ( n47886 , n47884 , n47885 );
and ( n47887 , n47886 , n30269 );
and ( n47888 , n42904 , n28587 );
and ( n47889 , n26601 , n39807 );
or ( n47890 , n47888 , n47889 );
and ( n47891 , n47890 , n30982 );
and ( n47892 , n29211 , n28587 );
and ( n47893 , n26601 , n39807 );
or ( n47894 , n47892 , n47893 );
and ( n47895 , n47894 , n30989 );
and ( n47896 , n42929 , n28587 );
and ( n47897 , n26601 , n39807 );
or ( n47898 , n47896 , n47897 );
and ( n47899 , n47898 , n31002 );
and ( n47900 , n26601 , n34607 );
or ( n47901 , n47883 , n47887 , n47891 , n47895 , n47899 , n47900 );
and ( n47902 , n47879 , n47901 );
and ( n47903 , n26601 , n24800 );
or ( n47904 , n47902 , n47903 );
and ( n47905 , n47904 , n31008 );
and ( n47906 , n26601 , n10618 );
or ( n47907 , n47905 , n47906 );
buf ( n47908 , n47907 );
buf ( n47909 , n47908 );
buf ( n47910 , n10615 );
not ( n47911 , n34821 );
not ( n47912 , n13916 );
and ( n47913 , n47912 , n13606 );
xor ( n47914 , n13607 , n13878 );
and ( n47915 , n47914 , n13916 );
or ( n47916 , n47913 , n47915 );
buf ( n47917 , n47916 );
and ( n47918 , n47917 , n14137 );
and ( n47919 , n47917 , n14143 );
not ( n47920 , n14139 );
and ( n47921 , n47920 , n36141 );
not ( n47922 , n36245 );
and ( n47923 , n47922 , n36153 );
xor ( n47924 , n46404 , n46407 );
and ( n47925 , n47924 , n36245 );
or ( n47926 , n47923 , n47925 );
buf ( n47927 , n47926 );
and ( n47928 , n47927 , n14139 );
or ( n47929 , n47921 , n47928 );
and ( n47930 , n47929 , n14140 );
and ( n47931 , n36141 , n14141 );
or ( n47932 , n47918 , n47919 , n47930 , n47931 );
and ( n47933 , n47932 , n36345 );
and ( n47934 , n13209 , n36352 );
or ( n47935 , n47933 , n47934 );
and ( n47936 , n47935 , n14562 );
not ( n47937 , n37048 );
and ( n47938 , n47937 , n36959 );
xor ( n47939 , n46427 , n46430 );
and ( n47940 , n47939 , n37048 );
or ( n47941 , n47938 , n47940 );
buf ( n47942 , n47941 );
and ( n47943 , n47942 , n36345 );
and ( n47944 , n13209 , n37073 );
or ( n47945 , n47943 , n47944 );
and ( n47946 , n47945 , n14586 );
not ( n47947 , n37801 );
and ( n47948 , n47947 , n37712 );
xor ( n47949 , n46445 , n46448 );
and ( n47950 , n47949 , n37801 );
or ( n47951 , n47948 , n47950 );
buf ( n47952 , n47951 );
and ( n47953 , n47952 , n36350 );
and ( n47954 , n13209 , n37825 );
or ( n47955 , n47953 , n47954 );
and ( n47956 , n47955 , n14584 );
and ( n47957 , n47942 , n36350 );
and ( n47958 , n13209 , n37831 );
or ( n47959 , n47957 , n47958 );
and ( n47960 , n47959 , n37835 );
and ( n47961 , n47952 , n36350 );
and ( n47962 , n13209 , n37831 );
or ( n47963 , n47961 , n47962 );
and ( n47964 , n47963 , n37841 );
and ( n47965 , n15052 , n36350 );
and ( n47966 , n13209 , n37831 );
or ( n47967 , n47965 , n47966 );
and ( n47968 , n47967 , n37847 );
and ( n47969 , n13209 , n37849 );
or ( n47970 , n47936 , n47946 , n47956 , n47960 , n47964 , n47968 , n47969 );
and ( n47971 , n47911 , n47970 );
and ( n47972 , n13209 , n34821 );
or ( n47973 , n47971 , n47972 );
and ( n47974 , n47973 , n16574 );
and ( n47975 , n13209 , n16576 );
or ( n47976 , n47974 , n47975 );
buf ( n47977 , n47976 );
buf ( n47978 , n47977 );
not ( n47979 , n17162 );
not ( n47980 , n17450 );
and ( n47981 , n10678 , n37947 );
not ( n47982 , n38425 );
and ( n47983 , n47982 , n38285 );
xor ( n47984 , n38429 , n38451 );
and ( n47985 , n47984 , n38425 );
or ( n47986 , n47983 , n47985 );
buf ( n47987 , n47986 );
and ( n47988 , n47987 , n19745 );
not ( n47989 , n38934 );
and ( n47990 , n47989 , n38794 );
xor ( n47991 , n38938 , n38960 );
and ( n47992 , n47991 , n38934 );
or ( n47993 , n47990 , n47992 );
buf ( n47994 , n47993 );
and ( n47995 , n47994 , n19748 );
and ( n47996 , n22200 , n21253 );
and ( n47997 , n10678 , n21255 );
or ( n47998 , n47988 , n47995 , n47996 , n47997 );
and ( n47999 , n47998 , n38980 );
or ( n48000 , n47981 , n47999 );
and ( n48001 , n47980 , n48000 );
or ( n48002 , n48001 , C0 );
and ( n48003 , n47979 , n48002 );
and ( n48004 , n47998 , n17162 );
or ( n48005 , n48003 , n48004 );
and ( n48006 , n48005 , n23924 );
not ( n48007 , n39264 );
and ( n48008 , n48007 , n39148 );
xor ( n48009 , n39268 , n39290 );
and ( n48010 , n48009 , n39264 );
or ( n48011 , n48008 , n48010 );
buf ( n48012 , n48011 );
and ( n48013 , n48012 , n23926 );
or ( n48014 , n48006 , n48013 );
buf ( n48015 , n48014 );
buf ( n48016 , n48015 );
and ( n48017 , n11808 , n16574 );
and ( n48018 , n15035 , n16576 );
or ( n48019 , n48017 , n48018 );
buf ( n48020 , n48019 );
buf ( n48021 , n48020 );
not ( n48022 , n24800 );
and ( n48023 , n26663 , n25222 );
not ( n48024 , n26823 );
and ( n48025 , n48024 , n26649 );
xor ( n48026 , n43391 , n43394 );
and ( n48027 , n48026 , n26823 );
or ( n48028 , n48025 , n48027 );
buf ( n48029 , n48028 );
and ( n48030 , n48029 , n27046 );
and ( n48031 , n48029 , n27049 );
not ( n48032 , n27051 );
and ( n48033 , n48032 , n28390 );
not ( n48034 , n28494 );
and ( n48035 , n48034 , n28402 );
xor ( n48036 , n43407 , n43410 );
and ( n48037 , n48036 , n28494 );
or ( n48038 , n48035 , n48037 );
buf ( n48039 , n48038 );
and ( n48040 , n48039 , n27051 );
or ( n48041 , n48033 , n48040 );
and ( n48042 , n48041 , n28506 );
and ( n48043 , n28390 , n28508 );
or ( n48044 , n48030 , n48031 , n48042 , n48043 );
and ( n48045 , n48044 , n28589 );
and ( n48046 , n26663 , n31075 );
or ( n48047 , n48045 , n48046 );
and ( n48048 , n48047 , n28594 );
not ( n48049 , n30249 );
and ( n48050 , n48049 , n30160 );
xor ( n48051 , n43428 , n43431 );
and ( n48052 , n48051 , n30249 );
or ( n48053 , n48050 , n48052 );
buf ( n48054 , n48053 );
and ( n48055 , n48054 , n28589 );
and ( n48056 , n26663 , n31075 );
or ( n48057 , n48055 , n48056 );
and ( n48058 , n48057 , n30269 );
not ( n48059 , n30963 );
and ( n48060 , n48059 , n30874 );
xor ( n48061 , n43444 , n43447 );
and ( n48062 , n48061 , n30963 );
or ( n48063 , n48060 , n48062 );
buf ( n48064 , n48063 );
and ( n48065 , n48064 , n28589 );
and ( n48066 , n26663 , n31075 );
or ( n48067 , n48065 , n48066 );
and ( n48068 , n48067 , n30982 );
and ( n48069 , n29185 , n28589 );
and ( n48070 , n26663 , n31075 );
or ( n48071 , n48069 , n48070 );
and ( n48072 , n48071 , n30989 );
and ( n48073 , n29185 , n30991 );
xor ( n48074 , n43464 , n43468 );
buf ( n48075 , n48074 );
and ( n48076 , n48075 , n28589 );
and ( n48077 , n26663 , n31075 );
or ( n48078 , n48076 , n48077 );
and ( n48079 , n48078 , n31002 );
or ( n48080 , n48023 , n48048 , n48058 , n48068 , n48072 , n48073 , n48079 );
and ( n48081 , n48022 , n48080 );
and ( n48082 , n26663 , n24800 );
or ( n48083 , n48081 , n48082 );
and ( n48084 , n48083 , n31008 );
and ( n48085 , n25579 , n10618 );
or ( n48086 , n48084 , n48085 );
buf ( n48087 , n48086 );
buf ( n48088 , n48087 );
buf ( n48089 , n10613 );
buf ( n48090 , n10613 );
not ( n48091 , n24800 );
and ( n48092 , n26393 , n25222 );
not ( n48093 , n26823 );
and ( n48094 , n48093 , n26377 );
xor ( n48095 , n39633 , n39636 );
and ( n48096 , n48095 , n26823 );
or ( n48097 , n48094 , n48096 );
buf ( n48098 , n48097 );
and ( n48099 , n48098 , n27046 );
and ( n48100 , n48098 , n27049 );
not ( n48101 , n27051 );
and ( n48102 , n48101 , n28214 );
not ( n48103 , n28494 );
and ( n48104 , n48103 , n28226 );
xor ( n48105 , n39649 , n39652 );
and ( n48106 , n48105 , n28494 );
or ( n48107 , n48104 , n48106 );
buf ( n48108 , n48107 );
and ( n48109 , n48108 , n27051 );
or ( n48110 , n48102 , n48109 );
and ( n48111 , n48110 , n28506 );
and ( n48112 , n28214 , n28508 );
or ( n48113 , n48099 , n48100 , n48111 , n48112 );
and ( n48114 , n48113 , n28583 );
and ( n48115 , n26393 , n28591 );
or ( n48116 , n48114 , n48115 );
and ( n48117 , n48116 , n28594 );
not ( n48118 , n30249 );
and ( n48119 , n48118 , n30024 );
xor ( n48120 , n39670 , n39673 );
and ( n48121 , n48120 , n30249 );
or ( n48122 , n48119 , n48121 );
buf ( n48123 , n48122 );
and ( n48124 , n48123 , n28583 );
and ( n48125 , n26393 , n28591 );
or ( n48126 , n48124 , n48125 );
and ( n48127 , n48126 , n30269 );
not ( n48128 , n30963 );
and ( n48129 , n48128 , n30738 );
xor ( n48130 , n39686 , n39689 );
and ( n48131 , n48130 , n30963 );
or ( n48132 , n48129 , n48131 );
buf ( n48133 , n48132 );
and ( n48134 , n48133 , n28583 );
and ( n48135 , n26393 , n28591 );
or ( n48136 , n48134 , n48135 );
and ( n48137 , n48136 , n30982 );
and ( n48138 , n29355 , n28583 );
and ( n48139 , n26393 , n28591 );
or ( n48140 , n48138 , n48139 );
and ( n48141 , n48140 , n30989 );
and ( n48142 , n26391 , n30991 );
xor ( n48143 , n39706 , n39710 );
buf ( n48144 , n48143 );
and ( n48145 , n48144 , n28583 );
and ( n48146 , n26393 , n28591 );
or ( n48147 , n48145 , n48146 );
and ( n48148 , n48147 , n31002 );
or ( n48149 , n48092 , n48117 , n48127 , n48137 , n48141 , n48142 , n48148 );
and ( n48150 , n48091 , n48149 );
and ( n48151 , n26393 , n24800 );
or ( n48152 , n48150 , n48151 );
and ( n48153 , n48152 , n31008 );
and ( n48154 , n26393 , n10618 );
or ( n48155 , n48153 , n48154 );
buf ( n48156 , n48155 );
buf ( n48157 , n48156 );
not ( n48158 , n17451 );
and ( n48159 , n48158 , n21297 );
and ( n48160 , n21272 , n17451 );
or ( n48161 , n48159 , n48160 );
and ( n48162 , n48161 , n23924 );
and ( n48163 , n21272 , n23926 );
or ( n48164 , n48162 , n48163 );
buf ( n48165 , n48164 );
buf ( n48166 , n48165 );
buf ( n48167 , n10613 );
buf ( n48168 , n10613 );
buf ( n48169 , n10613 );
buf ( n48170 , n10615 );
buf ( n48171 , n10615 );
not ( n48172 , n34821 );
and ( n48173 , n13489 , n14592 );
and ( n48174 , n43526 , n36350 );
and ( n48175 , n13489 , n43691 );
or ( n48176 , n48174 , n48175 );
and ( n48177 , n48176 , n14562 );
and ( n48178 , n43539 , n36350 );
and ( n48179 , n13489 , n43703 );
or ( n48180 , n48178 , n48179 );
and ( n48181 , n48180 , n14586 );
and ( n48182 , n43552 , n36345 );
and ( n48183 , n13489 , n43715 );
or ( n48184 , n48182 , n48183 );
and ( n48185 , n48184 , n14584 );
and ( n48186 , n43539 , n36345 );
and ( n48187 , n13489 , n43721 );
or ( n48188 , n48186 , n48187 );
and ( n48189 , n48188 , n37835 );
and ( n48190 , n43552 , n36345 );
and ( n48191 , n13489 , n43721 );
or ( n48192 , n48190 , n48191 );
and ( n48193 , n48192 , n37841 );
and ( n48194 , n15845 , n14564 );
and ( n48195 , n15845 , n36345 );
and ( n48196 , n13489 , n43721 );
or ( n48197 , n48195 , n48196 );
and ( n48198 , n48197 , n37847 );
or ( n48199 , n48173 , n48177 , n48181 , n48185 , n48189 , n48193 , n48194 , n48198 );
and ( n48200 , n48172 , n48199 );
and ( n48201 , n13489 , n34821 );
or ( n48202 , n48200 , n48201 );
and ( n48203 , n48202 , n16574 );
and ( n48204 , n12330 , n16576 );
or ( n48205 , n48203 , n48204 );
buf ( n48206 , n48205 );
buf ( n48207 , n48206 );
not ( n48208 , n34821 );
and ( n48209 , n13373 , n14592 );
and ( n48210 , n39404 , n36348 );
and ( n48211 , n13373 , n43530 );
or ( n48212 , n48210 , n48211 );
and ( n48213 , n48212 , n14562 );
and ( n48214 , n39423 , n36347 );
and ( n48215 , n13373 , n43543 );
or ( n48216 , n48214 , n48215 );
and ( n48217 , n48216 , n14586 );
and ( n48218 , n39442 , n36348 );
and ( n48219 , n13373 , n43556 );
or ( n48220 , n48218 , n48219 );
and ( n48221 , n48220 , n14584 );
and ( n48222 , n39423 , n36347 );
and ( n48223 , n13373 , n43563 );
or ( n48224 , n48222 , n48223 );
and ( n48225 , n48224 , n37835 );
and ( n48226 , n39442 , n36347 );
and ( n48227 , n13373 , n43563 );
or ( n48228 , n48226 , n48227 );
and ( n48229 , n48228 , n37841 );
and ( n48230 , n13371 , n14564 );
and ( n48231 , n15647 , n36347 );
and ( n48232 , n13373 , n43563 );
or ( n48233 , n48231 , n48232 );
and ( n48234 , n48233 , n37847 );
or ( n48235 , n48209 , n48213 , n48217 , n48221 , n48225 , n48229 , n48230 , n48234 );
and ( n48236 , n48208 , n48235 );
and ( n48237 , n13373 , n34821 );
or ( n48238 , n48236 , n48237 );
and ( n48239 , n48238 , n16574 );
and ( n48240 , n13373 , n16576 );
or ( n48241 , n48239 , n48240 );
buf ( n48242 , n48241 );
buf ( n48243 , n48242 );
not ( n48244 , n17451 );
and ( n48245 , n19418 , n17873 );
not ( n48246 , n19474 );
and ( n48247 , n48246 , n19402 );
xor ( n48248 , n40060 , n40061 );
and ( n48249 , n48248 , n19474 );
or ( n48250 , n48247 , n48249 );
buf ( n48251 , n48250 );
and ( n48252 , n48251 , n19745 );
and ( n48253 , n48251 , n19748 );
not ( n48254 , n19750 );
and ( n48255 , n48254 , n21155 );
not ( n48256 , n21193 );
and ( n48257 , n48256 , n21167 );
xor ( n48258 , n45343 , n45344 );
and ( n48259 , n48258 , n21193 );
or ( n48260 , n48257 , n48259 );
buf ( n48261 , n48260 );
and ( n48262 , n48261 , n19750 );
or ( n48263 , n48255 , n48262 );
and ( n48264 , n48263 , n21253 );
and ( n48265 , n21155 , n21255 );
or ( n48266 , n48252 , n48253 , n48264 , n48265 );
and ( n48267 , n48266 , n21330 );
and ( n48268 , n19418 , n21338 );
or ( n48269 , n48267 , n48268 );
and ( n48270 , n48269 , n21341 );
not ( n48271 , n22996 );
and ( n48272 , n48271 , n22958 );
xor ( n48273 , n40088 , n40089 );
and ( n48274 , n48273 , n22996 );
or ( n48275 , n48272 , n48274 );
buf ( n48276 , n48275 );
and ( n48277 , n48276 , n21330 );
and ( n48278 , n19418 , n21338 );
or ( n48279 , n48277 , n48278 );
and ( n48280 , n48279 , n23064 );
not ( n48281 , n23758 );
and ( n48282 , n48281 , n23720 );
xor ( n48283 , n40103 , n40104 );
and ( n48284 , n48283 , n23758 );
or ( n48285 , n48282 , n48284 );
buf ( n48286 , n48285 );
and ( n48287 , n48286 , n21330 );
and ( n48288 , n19418 , n21338 );
or ( n48289 , n48287 , n48288 );
and ( n48290 , n48289 , n23825 );
and ( n48291 , n21893 , n21330 );
and ( n48292 , n19418 , n21338 );
or ( n48293 , n48291 , n48292 );
and ( n48294 , n48293 , n23832 );
and ( n48295 , n19416 , n23834 );
xor ( n48296 , n40128 , n40129 );
buf ( n48297 , n48296 );
and ( n48298 , n48297 , n21330 );
and ( n48299 , n19418 , n21338 );
or ( n48300 , n48298 , n48299 );
and ( n48301 , n48300 , n23917 );
or ( n48302 , n48245 , n48270 , n48280 , n48290 , n48294 , n48295 , n48301 );
and ( n48303 , n48244 , n48302 );
and ( n48304 , n19418 , n17451 );
or ( n48305 , n48303 , n48304 );
and ( n48306 , n48305 , n23924 );
and ( n48307 , n19418 , n23926 );
or ( n48308 , n48306 , n48307 );
buf ( n48309 , n48308 );
buf ( n48310 , n48309 );
buf ( n48311 , n10615 );
buf ( n48312 , n10615 );
not ( n48313 , n24800 );
not ( n48314 , n26823 );
and ( n48315 , n48314 , n25937 );
xor ( n48316 , n31025 , n31028 );
and ( n48317 , n48316 , n26823 );
or ( n48318 , n48315 , n48317 );
buf ( n48319 , n48318 );
and ( n48320 , n48319 , n27046 );
and ( n48321 , n48319 , n27049 );
not ( n48322 , n27051 );
and ( n48323 , n48322 , n27928 );
not ( n48324 , n28494 );
and ( n48325 , n48324 , n27940 );
xor ( n48326 , n31053 , n31056 );
and ( n48327 , n48326 , n28494 );
or ( n48328 , n48325 , n48327 );
buf ( n48329 , n48328 );
and ( n48330 , n48329 , n27051 );
or ( n48331 , n48323 , n48330 );
and ( n48332 , n48331 , n28506 );
and ( n48333 , n27928 , n28508 );
or ( n48334 , n48320 , n48321 , n48332 , n48333 );
and ( n48335 , n48334 , n28587 );
and ( n48336 , n25956 , n39807 );
or ( n48337 , n48335 , n48336 );
and ( n48338 , n48337 , n28594 );
not ( n48339 , n30249 );
and ( n48340 , n48339 , n29803 );
xor ( n48341 , n31088 , n31091 );
and ( n48342 , n48341 , n30249 );
or ( n48343 , n48340 , n48342 );
buf ( n48344 , n48343 );
and ( n48345 , n48344 , n28587 );
and ( n48346 , n25956 , n39807 );
or ( n48347 , n48345 , n48346 );
and ( n48348 , n48347 , n30269 );
not ( n48349 , n30963 );
and ( n48350 , n48349 , n30517 );
xor ( n48351 , n31116 , n31119 );
and ( n48352 , n48351 , n30963 );
or ( n48353 , n48350 , n48352 );
buf ( n48354 , n48353 );
and ( n48355 , n48354 , n28587 );
and ( n48356 , n25956 , n39807 );
or ( n48357 , n48355 , n48356 );
and ( n48358 , n48357 , n30982 );
and ( n48359 , n29615 , n28587 );
and ( n48360 , n25956 , n39807 );
or ( n48361 , n48359 , n48360 );
and ( n48362 , n48361 , n30989 );
xor ( n48363 , n31155 , n31159 );
buf ( n48364 , n48363 );
and ( n48365 , n48364 , n28587 );
and ( n48366 , n25956 , n39807 );
or ( n48367 , n48365 , n48366 );
and ( n48368 , n48367 , n31002 );
and ( n48369 , n25956 , n34607 );
or ( n48370 , n48338 , n48348 , n48358 , n48362 , n48368 , n48369 );
and ( n48371 , n48313 , n48370 );
and ( n48372 , n25956 , n24800 );
or ( n48373 , n48371 , n48372 );
and ( n48374 , n48373 , n31008 );
and ( n48375 , n25956 , n10618 );
or ( n48376 , n48374 , n48375 );
buf ( n48377 , n48376 );
buf ( n48378 , n48377 );
not ( n48379 , n34821 );
and ( n48380 , n13397 , n14592 );
not ( n48381 , n13916 );
and ( n48382 , n48381 , n13782 );
xor ( n48383 , n13783 , n13862 );
and ( n48384 , n48383 , n13916 );
or ( n48385 , n48382 , n48384 );
buf ( n48386 , n48385 );
and ( n48387 , n48386 , n14137 );
and ( n48388 , n48386 , n14143 );
not ( n48389 , n14139 );
and ( n48390 , n48389 , n35789 );
not ( n48391 , n36245 );
and ( n48392 , n48391 , n35801 );
xor ( n48393 , n39392 , n39393 );
and ( n48394 , n48393 , n36245 );
or ( n48395 , n48392 , n48394 );
buf ( n48396 , n48395 );
and ( n48397 , n48396 , n14139 );
or ( n48398 , n48390 , n48397 );
and ( n48399 , n48398 , n14140 );
and ( n48400 , n35789 , n14141 );
or ( n48401 , n48387 , n48388 , n48399 , n48400 );
and ( n48402 , n48401 , n36348 );
and ( n48403 , n13397 , n43530 );
or ( n48404 , n48402 , n48403 );
and ( n48405 , n48404 , n14562 );
not ( n48406 , n37048 );
and ( n48407 , n48406 , n36687 );
xor ( n48408 , n39416 , n39417 );
and ( n48409 , n48408 , n37048 );
or ( n48410 , n48407 , n48409 );
buf ( n48411 , n48410 );
and ( n48412 , n48411 , n36347 );
and ( n48413 , n13397 , n43543 );
or ( n48414 , n48412 , n48413 );
and ( n48415 , n48414 , n14586 );
not ( n48416 , n37801 );
and ( n48417 , n48416 , n37440 );
xor ( n48418 , n39435 , n39436 );
and ( n48419 , n48418 , n37801 );
or ( n48420 , n48417 , n48419 );
buf ( n48421 , n48420 );
and ( n48422 , n48421 , n36348 );
and ( n48423 , n13397 , n43556 );
or ( n48424 , n48422 , n48423 );
and ( n48425 , n48424 , n14584 );
and ( n48426 , n48411 , n36347 );
and ( n48427 , n13397 , n43563 );
or ( n48428 , n48426 , n48427 );
and ( n48429 , n48428 , n37835 );
and ( n48430 , n48421 , n36347 );
and ( n48431 , n13397 , n43563 );
or ( n48432 , n48430 , n48431 );
and ( n48433 , n48432 , n37841 );
and ( n48434 , n13395 , n14564 );
and ( n48435 , n15691 , n36347 );
and ( n48436 , n13397 , n43563 );
or ( n48437 , n48435 , n48436 );
and ( n48438 , n48437 , n37847 );
or ( n48439 , n48380 , n48405 , n48415 , n48425 , n48429 , n48433 , n48434 , n48438 );
and ( n48440 , n48379 , n48439 );
and ( n48441 , n13397 , n34821 );
or ( n48442 , n48440 , n48441 );
and ( n48443 , n48442 , n16574 );
and ( n48444 , n13397 , n16576 );
or ( n48445 , n48443 , n48444 );
buf ( n48446 , n48445 );
buf ( n48447 , n48446 );
buf ( n48448 , n10613 );
buf ( n48449 , n10613 );
buf ( n48450 , n10615 );
not ( n48451 , n34538 );
and ( n48452 , n48451 , n18949 );
and ( n48453 , n14753 , n34538 );
or ( n48454 , n48452 , n48453 );
and ( n48455 , n48454 , n23924 );
and ( n48456 , n14753 , n23926 );
or ( n48457 , n48455 , n48456 );
buf ( n48458 , n48457 );
buf ( n48459 , n48458 );
buf ( n48460 , n10613 );
buf ( n48461 , n10615 );
not ( n48462 , n24800 );
and ( n48463 , n25663 , n25222 );
and ( n48464 , n39944 , n28589 );
and ( n48465 , n25663 , n31075 );
or ( n48466 , n48464 , n48465 );
and ( n48467 , n48466 , n28594 );
and ( n48468 , n39954 , n28589 );
and ( n48469 , n25663 , n31075 );
or ( n48470 , n48468 , n48469 );
and ( n48471 , n48470 , n30269 );
and ( n48472 , n39964 , n28589 );
and ( n48473 , n25663 , n31075 );
or ( n48474 , n48472 , n48473 );
and ( n48475 , n48474 , n30982 );
and ( n48476 , n28892 , n28589 );
and ( n48477 , n25663 , n31075 );
or ( n48478 , n48476 , n48477 );
and ( n48479 , n48478 , n30989 );
and ( n48480 , n28892 , n30991 );
and ( n48481 , n39974 , n28589 );
and ( n48482 , n25663 , n31075 );
or ( n48483 , n48481 , n48482 );
and ( n48484 , n48483 , n31002 );
or ( n48485 , n48463 , n48467 , n48471 , n48475 , n48479 , n48480 , n48484 );
and ( n48486 , n48462 , n48485 );
and ( n48487 , n25663 , n24800 );
or ( n48488 , n48486 , n48487 );
and ( n48489 , n48488 , n31008 );
and ( n48490 , n25224 , n10618 );
or ( n48491 , n48489 , n48490 );
buf ( n48492 , n48491 );
buf ( n48493 , n48492 );
not ( n48494 , n24800 );
not ( n48495 , n27051 );
and ( n48496 , n48495 , n27882 );
or ( n48497 , n48496 , C0 );
and ( n48498 , n48497 , n28506 );
and ( n48499 , n27882 , n28508 );
or ( n48500 , C0 , C0 , n48498 , n48499 );
and ( n48501 , n48500 , n28586 );
and ( n48502 , n25872 , n34573 );
or ( n48503 , n48501 , n48502 );
and ( n48504 , n48503 , n28594 );
and ( n48505 , n25872 , n34573 );
buf ( n48506 , n48505 );
and ( n48507 , n48506 , n30269 );
and ( n48508 , n25872 , n34573 );
buf ( n48509 , n48508 );
and ( n48510 , n48509 , n30982 );
and ( n48511 , n29094 , n28586 );
and ( n48512 , n25872 , n34573 );
or ( n48513 , n48511 , n48512 );
and ( n48514 , n48513 , n30989 );
buf ( n48515 , n29094 );
not ( n48516 , n48515 );
buf ( n48517 , n29107 );
not ( n48518 , n48517 );
buf ( n48519 , n29120 );
not ( n48520 , n48519 );
and ( n48521 , n45301 , n45308 );
and ( n48522 , n48520 , n48521 );
and ( n48523 , n48518 , n48522 );
xor ( n48524 , n48516 , n48523 );
buf ( n48525 , n48524 );
and ( n48526 , n48525 , n28586 );
and ( n48527 , n25872 , n34573 );
or ( n48528 , n48526 , n48527 );
and ( n48529 , n48528 , n31002 );
and ( n48530 , n25872 , n34607 );
or ( n48531 , n48504 , n48507 , n48510 , n48514 , n48529 , n48530 );
and ( n48532 , n48494 , n48531 );
and ( n48533 , n25872 , n24800 );
or ( n48534 , n48532 , n48533 );
and ( n48535 , n48534 , n31008 );
and ( n48536 , n25872 , n10618 );
or ( n48537 , n48535 , n48536 );
buf ( n48538 , n48537 );
buf ( n48539 , n48538 );
buf ( n48540 , n10613 );
not ( n48541 , n24800 );
and ( n48542 , n26085 , n25222 );
and ( n48543 , n37895 , n28589 );
and ( n48544 , n26085 , n31075 );
or ( n48545 , n48543 , n48544 );
and ( n48546 , n48545 , n28594 );
and ( n48547 , n37905 , n28589 );
and ( n48548 , n26085 , n31075 );
or ( n48549 , n48547 , n48548 );
and ( n48550 , n48549 , n30269 );
and ( n48551 , n37915 , n28589 );
and ( n48552 , n26085 , n31075 );
or ( n48553 , n48551 , n48552 );
and ( n48554 , n48553 , n30982 );
and ( n48555 , n29535 , n28589 );
and ( n48556 , n26085 , n31075 );
or ( n48557 , n48555 , n48556 );
and ( n48558 , n48557 , n30989 );
and ( n48559 , n29535 , n30991 );
and ( n48560 , n37925 , n28589 );
and ( n48561 , n26085 , n31075 );
or ( n48562 , n48560 , n48561 );
and ( n48563 , n48562 , n31002 );
or ( n48564 , n48542 , n48546 , n48550 , n48554 , n48558 , n48559 , n48563 );
and ( n48565 , n48541 , n48564 );
and ( n48566 , n26085 , n24800 );
or ( n48567 , n48565 , n48566 );
and ( n48568 , n48567 , n31008 );
and ( n48569 , n25324 , n10618 );
or ( n48570 , n48568 , n48569 );
buf ( n48571 , n48570 );
buf ( n48572 , n48571 );
buf ( n48573 , n10615 );
not ( n48574 , n34821 );
and ( n48575 , n45746 , n36347 );
and ( n48576 , n13231 , n39408 );
or ( n48577 , n48575 , n48576 );
and ( n48578 , n48577 , n14562 );
and ( n48579 , n45762 , n36348 );
and ( n48580 , n13231 , n39427 );
or ( n48581 , n48579 , n48580 );
and ( n48582 , n48581 , n14586 );
and ( n48583 , n45778 , n36347 );
and ( n48584 , n13231 , n39446 );
or ( n48585 , n48583 , n48584 );
and ( n48586 , n48585 , n14584 );
and ( n48587 , n45762 , n36348 );
and ( n48588 , n13231 , n39453 );
or ( n48589 , n48587 , n48588 );
and ( n48590 , n48589 , n37835 );
and ( n48591 , n45778 , n36348 );
and ( n48592 , n13231 , n39453 );
or ( n48593 , n48591 , n48592 );
and ( n48594 , n48593 , n37841 );
and ( n48595 , n15082 , n36348 );
and ( n48596 , n13231 , n39453 );
or ( n48597 , n48595 , n48596 );
and ( n48598 , n48597 , n37847 );
and ( n48599 , n13231 , n37849 );
or ( n48600 , n48578 , n48582 , n48586 , n48590 , n48594 , n48598 , n48599 );
and ( n48601 , n48574 , n48600 );
and ( n48602 , n13231 , n34821 );
or ( n48603 , n48601 , n48602 );
and ( n48604 , n48603 , n16574 );
and ( n48605 , n13231 , n16576 );
or ( n48606 , n48604 , n48605 );
buf ( n48607 , n48606 );
buf ( n48608 , n48607 );
buf ( n48609 , n10613 );
not ( n48610 , n34821 );
and ( n48611 , n13227 , n14592 );
and ( n48612 , n45746 , n36350 );
and ( n48613 , n13227 , n43691 );
or ( n48614 , n48612 , n48613 );
and ( n48615 , n48614 , n14562 );
and ( n48616 , n45762 , n36350 );
and ( n48617 , n13227 , n43703 );
or ( n48618 , n48616 , n48617 );
and ( n48619 , n48618 , n14586 );
and ( n48620 , n45778 , n36345 );
and ( n48621 , n13227 , n43715 );
or ( n48622 , n48620 , n48621 );
and ( n48623 , n48622 , n14584 );
and ( n48624 , n45762 , n36345 );
and ( n48625 , n13227 , n43721 );
or ( n48626 , n48624 , n48625 );
and ( n48627 , n48626 , n37835 );
and ( n48628 , n45778 , n36345 );
and ( n48629 , n13227 , n43721 );
or ( n48630 , n48628 , n48629 );
and ( n48631 , n48630 , n37841 );
and ( n48632 , n15082 , n14564 );
and ( n48633 , n15082 , n36345 );
and ( n48634 , n13227 , n43721 );
or ( n48635 , n48633 , n48634 );
and ( n48636 , n48635 , n37847 );
or ( n48637 , n48611 , n48615 , n48619 , n48623 , n48627 , n48631 , n48632 , n48636 );
and ( n48638 , n48610 , n48637 );
and ( n48639 , n13227 , n34821 );
or ( n48640 , n48638 , n48639 );
and ( n48641 , n48640 , n16574 );
and ( n48642 , n12267 , n16576 );
or ( n48643 , n48641 , n48642 );
buf ( n48644 , n48643 );
buf ( n48645 , n48644 );
buf ( n48646 , n10615 );
not ( n48647 , n34821 );
and ( n48648 , n13323 , n14592 );
not ( n48649 , n13916 );
and ( n48650 , n48649 , n13716 );
xor ( n48651 , n13717 , n13868 );
and ( n48652 , n48651 , n13916 );
or ( n48653 , n48650 , n48652 );
buf ( n48654 , n48653 );
and ( n48655 , n48654 , n14137 );
and ( n48656 , n48654 , n14143 );
not ( n48657 , n14139 );
and ( n48658 , n48657 , n35921 );
not ( n48659 , n36245 );
and ( n48660 , n48659 , n35933 );
xor ( n48661 , n43031 , n43038 );
and ( n48662 , n48661 , n36245 );
or ( n48663 , n48660 , n48662 );
buf ( n48664 , n48663 );
and ( n48665 , n48664 , n14139 );
or ( n48666 , n48658 , n48665 );
and ( n48667 , n48666 , n14140 );
and ( n48668 , n35921 , n14141 );
or ( n48669 , n48655 , n48656 , n48667 , n48668 );
and ( n48670 , n48669 , n36350 );
and ( n48671 , n13323 , n43691 );
or ( n48672 , n48670 , n48671 );
and ( n48673 , n48672 , n14562 );
not ( n48674 , n37048 );
and ( n48675 , n48674 , n36789 );
xor ( n48676 , n43058 , n43065 );
and ( n48677 , n48676 , n37048 );
or ( n48678 , n48675 , n48677 );
buf ( n48679 , n48678 );
and ( n48680 , n48679 , n36350 );
and ( n48681 , n13323 , n43703 );
or ( n48682 , n48680 , n48681 );
and ( n48683 , n48682 , n14586 );
not ( n48684 , n37801 );
and ( n48685 , n48684 , n37542 );
xor ( n48686 , n43080 , n43087 );
and ( n48687 , n48686 , n37801 );
or ( n48688 , n48685 , n48687 );
buf ( n48689 , n48688 );
and ( n48690 , n48689 , n36345 );
and ( n48691 , n13323 , n43715 );
or ( n48692 , n48690 , n48691 );
and ( n48693 , n48692 , n14584 );
and ( n48694 , n48679 , n36345 );
and ( n48695 , n13323 , n43721 );
or ( n48696 , n48694 , n48695 );
and ( n48697 , n48696 , n37835 );
and ( n48698 , n48689 , n36345 );
and ( n48699 , n13323 , n43721 );
or ( n48700 , n48698 , n48699 );
and ( n48701 , n48700 , n37841 );
and ( n48702 , n15559 , n14564 );
and ( n48703 , n15559 , n36345 );
and ( n48704 , n13323 , n43721 );
or ( n48705 , n48703 , n48704 );
and ( n48706 , n48705 , n37847 );
or ( n48707 , n48648 , n48673 , n48683 , n48693 , n48697 , n48701 , n48702 , n48706 );
and ( n48708 , n48647 , n48707 );
and ( n48709 , n13323 , n34821 );
or ( n48710 , n48708 , n48709 );
and ( n48711 , n48710 , n16574 );
and ( n48712 , n12291 , n16576 );
or ( n48713 , n48711 , n48712 );
buf ( n48714 , n48713 );
buf ( n48715 , n48714 );
buf ( n48716 , n10615 );
buf ( n48717 , n10613 );
not ( n48718 , n17451 );
not ( n48719 , n19474 );
and ( n48720 , n48719 , n19470 );
xor ( n48721 , n40058 , n40063 );
and ( n48722 , n48721 , n19474 );
or ( n48723 , n48720 , n48722 );
buf ( n48724 , n48723 );
and ( n48725 , n48724 , n19745 );
and ( n48726 , n48724 , n19748 );
not ( n48727 , n19750 );
not ( n48728 , n19753 );
buf ( n48729 , n20529 );
and ( n48730 , n48728 , n48729 );
xor ( n48731 , n20531 , n20574 );
buf ( n48732 , n48731 );
and ( n48733 , n48732 , n19753 );
or ( n48734 , n48730 , n48733 );
buf ( n48735 , n48734 );
and ( n48736 , n48727 , n48735 );
and ( n48737 , n45342 , n45345 );
buf ( n48738 , n48737 );
and ( n48739 , n48738 , n21193 );
or ( n48740 , C0 , n48739 );
buf ( n48741 , n48740 );
and ( n48742 , n48741 , n19750 );
or ( n48743 , n48736 , n48742 );
and ( n48744 , n48743 , n21253 );
and ( n48745 , n48735 , n21255 );
or ( n48746 , n48725 , n48726 , n48744 , n48745 );
and ( n48747 , n48746 , n21334 );
and ( n48748 , n20494 , n34492 );
or ( n48749 , n48747 , n48748 );
and ( n48750 , n48749 , n21341 );
not ( n48751 , n22996 );
and ( n48752 , n48751 , n22992 );
xor ( n48753 , n40086 , n40091 );
and ( n48754 , n48753 , n22996 );
or ( n48755 , n48752 , n48754 );
buf ( n48756 , n48755 );
and ( n48757 , n48756 , n21334 );
and ( n48758 , n20494 , n34492 );
or ( n48759 , n48757 , n48758 );
and ( n48760 , n48759 , n23064 );
not ( n48761 , n23758 );
and ( n48762 , n48761 , n23754 );
xor ( n48763 , n40101 , n40106 );
and ( n48764 , n48763 , n23758 );
or ( n48765 , n48762 , n48764 );
buf ( n48766 , n48765 );
and ( n48767 , n48766 , n21334 );
and ( n48768 , n20494 , n34492 );
or ( n48769 , n48767 , n48768 );
and ( n48770 , n48769 , n23825 );
and ( n48771 , n21867 , n21334 );
and ( n48772 , n20494 , n34492 );
or ( n48773 , n48771 , n48772 );
and ( n48774 , n48773 , n23832 );
xor ( n48775 , n40124 , n40131 );
buf ( n48776 , n48775 );
and ( n48777 , n48776 , n21334 );
and ( n48778 , n20494 , n34492 );
or ( n48779 , n48777 , n48778 );
and ( n48780 , n48779 , n23917 );
and ( n48781 , n20494 , n34526 );
or ( n48782 , n48750 , n48760 , n48770 , n48774 , n48780 , n48781 );
and ( n48783 , n48718 , n48782 );
and ( n48784 , n20494 , n17451 );
or ( n48785 , n48783 , n48784 );
and ( n48786 , n48785 , n23924 );
and ( n48787 , n20494 , n23926 );
or ( n48788 , n48786 , n48787 );
buf ( n48789 , n48788 );
buf ( n48790 , n48789 );
buf ( n48791 , n10615 );
buf ( n48792 , n10615 );
and ( n48793 , n16777 , n23924 );
and ( n48794 , n22093 , n23926 );
or ( n48795 , n48793 , n48794 );
buf ( n48796 , n48795 );
buf ( n48797 , n48796 );
buf ( n48798 , n10613 );
and ( n48799 , n11504 , n16574 );
and ( n48800 , n14930 , n16576 );
or ( n48801 , n48799 , n48800 );
buf ( n48802 , n48801 );
buf ( n48803 , n48802 );
not ( n48804 , n24511 );
not ( n48805 , n24799 );
and ( n48806 , n10725 , n40154 );
not ( n48807 , n40632 );
and ( n48808 , n48807 , n40339 );
xor ( n48809 , n40648 , n40652 );
and ( n48810 , n48809 , n40632 );
or ( n48811 , n48808 , n48810 );
buf ( n48812 , n48811 );
and ( n48813 , n48812 , n27046 );
not ( n48814 , n41147 );
and ( n48815 , n48814 , n40854 );
xor ( n48816 , n41163 , n41167 );
and ( n48817 , n48816 , n41147 );
or ( n48818 , n48815 , n48817 );
buf ( n48819 , n48818 );
and ( n48820 , n48819 , n27049 );
and ( n48821 , n29633 , n28506 );
and ( n48822 , n10725 , n28508 );
or ( n48823 , n48813 , n48820 , n48821 , n48822 );
and ( n48824 , n48823 , n41199 );
or ( n48825 , n48806 , n48824 );
and ( n48826 , n48805 , n48825 );
xor ( n48827 , n41724 , n41732 );
xor ( n48828 , n48827 , n41767 );
buf ( n48829 , n48828 );
and ( n48830 , n48829 , n27046 );
xor ( n48831 , n42240 , n42241 );
xor ( n48832 , n48831 , n42263 );
buf ( n48833 , n48832 );
and ( n48834 , n48833 , n27049 );
and ( n48835 , n29633 , n42306 );
or ( n48836 , n48830 , n48834 , n48835 );
buf ( n48837 , n48836 );
and ( n48838 , C1 , n48837 );
or ( n48839 , n48838 , C0 );
buf ( n48840 , n48839 );
not ( n48841 , n48840 );
buf ( n48842 , n48841 );
buf ( n48843 , n48842 );
not ( n48844 , n48843 );
and ( n48845 , C1 , n48844 );
or ( n48846 , n48845 , C0 );
buf ( n48847 , n48846 );
and ( n48848 , n48847 , n24799 );
or ( n48849 , n48826 , n48848 );
and ( n48850 , n48804 , n48849 );
and ( n48851 , n48823 , n24511 );
or ( n48852 , n48850 , n48851 );
and ( n48853 , n48852 , n31008 );
not ( n48854 , n42601 );
and ( n48855 , n48854 , n42359 );
xor ( n48856 , n42617 , n42621 );
and ( n48857 , n48856 , n42601 );
or ( n48858 , n48855 , n48857 );
buf ( n48859 , n48858 );
and ( n48860 , n48859 , n10618 );
or ( n48861 , n48853 , n48860 );
buf ( n48862 , n48861 );
buf ( n48863 , n48862 );
buf ( n48864 , n10615 );
not ( n48865 , n17451 );
not ( n48866 , n19474 );
and ( n48867 , n48866 , n18655 );
xor ( n48868 , n19497 , n19505 );
and ( n48869 , n48868 , n19474 );
or ( n48870 , n48867 , n48869 );
buf ( n48871 , n48870 );
and ( n48872 , n48871 , n19745 );
and ( n48873 , n48871 , n19748 );
not ( n48874 , n19750 );
and ( n48875 , n48874 , n20679 );
not ( n48876 , n21193 );
and ( n48877 , n48876 , n20691 );
xor ( n48878 , n21216 , n21226 );
and ( n48879 , n48878 , n21193 );
or ( n48880 , n48877 , n48879 );
buf ( n48881 , n48880 );
and ( n48882 , n48881 , n19750 );
or ( n48883 , n48875 , n48882 );
and ( n48884 , n48883 , n21253 );
and ( n48885 , n20679 , n21255 );
or ( n48886 , n48872 , n48873 , n48884 , n48885 );
and ( n48887 , n48886 , n21333 );
and ( n48888 , n18673 , n34758 );
or ( n48889 , n48887 , n48888 );
and ( n48890 , n48889 , n21341 );
not ( n48891 , n22996 );
and ( n48892 , n48891 , n22584 );
xor ( n48893 , n23019 , n23029 );
and ( n48894 , n48893 , n22996 );
or ( n48895 , n48892 , n48894 );
buf ( n48896 , n48895 );
and ( n48897 , n48896 , n21333 );
and ( n48898 , n18673 , n34758 );
or ( n48899 , n48897 , n48898 );
and ( n48900 , n48899 , n23064 );
not ( n48901 , n23758 );
and ( n48902 , n48901 , n23346 );
xor ( n48903 , n23781 , n23791 );
and ( n48904 , n48903 , n23758 );
or ( n48905 , n48902 , n48904 );
buf ( n48906 , n48905 );
and ( n48907 , n48906 , n21333 );
and ( n48908 , n18673 , n34758 );
or ( n48909 , n48907 , n48908 );
and ( n48910 , n48909 , n23825 );
and ( n48911 , n22322 , n21333 );
and ( n48912 , n18673 , n34758 );
or ( n48913 , n48911 , n48912 );
and ( n48914 , n48913 , n23832 );
xor ( n48915 , n23877 , n23891 );
buf ( n48916 , n48915 );
and ( n48917 , n48916 , n21333 );
and ( n48918 , n18673 , n34758 );
or ( n48919 , n48917 , n48918 );
and ( n48920 , n48919 , n23917 );
and ( n48921 , n18673 , n34526 );
or ( n48922 , n48890 , n48900 , n48910 , n48914 , n48920 , n48921 );
and ( n48923 , n48865 , n48922 );
and ( n48924 , n18673 , n17451 );
or ( n48925 , n48923 , n48924 );
and ( n48926 , n48925 , n23924 );
and ( n48927 , n18673 , n23926 );
or ( n48928 , n48926 , n48927 );
buf ( n48929 , n48928 );
buf ( n48930 , n48929 );
not ( n48931 , n17451 );
not ( n48932 , n19474 );
and ( n48933 , n48932 , n18589 );
xor ( n48934 , n19499 , n19503 );
and ( n48935 , n48934 , n19474 );
or ( n48936 , n48933 , n48935 );
buf ( n48937 , n48936 );
and ( n48938 , n48937 , n19745 );
and ( n48939 , n48937 , n19748 );
not ( n48940 , n19750 );
and ( n48941 , n48940 , n20635 );
not ( n48942 , n21193 );
and ( n48943 , n48942 , n20647 );
xor ( n48944 , n21218 , n21224 );
and ( n48945 , n48944 , n21193 );
or ( n48946 , n48943 , n48945 );
buf ( n48947 , n48946 );
and ( n48948 , n48947 , n19750 );
or ( n48949 , n48941 , n48948 );
and ( n48950 , n48949 , n21253 );
and ( n48951 , n20635 , n21255 );
or ( n48952 , n48938 , n48939 , n48950 , n48951 );
and ( n48953 , n48952 , n21334 );
and ( n48954 , n18608 , n34492 );
or ( n48955 , n48953 , n48954 );
and ( n48956 , n48955 , n21341 );
not ( n48957 , n22996 );
and ( n48958 , n48957 , n22550 );
xor ( n48959 , n23021 , n23027 );
and ( n48960 , n48959 , n22996 );
or ( n48961 , n48958 , n48960 );
buf ( n48962 , n48961 );
and ( n48963 , n48962 , n21334 );
and ( n48964 , n18608 , n34492 );
or ( n48965 , n48963 , n48964 );
and ( n48966 , n48965 , n23064 );
not ( n48967 , n23758 );
and ( n48968 , n48967 , n23312 );
xor ( n48969 , n23783 , n23789 );
and ( n48970 , n48969 , n23758 );
or ( n48971 , n48968 , n48970 );
buf ( n48972 , n48971 );
and ( n48973 , n48972 , n21334 );
and ( n48974 , n18608 , n34492 );
or ( n48975 , n48973 , n48974 );
and ( n48976 , n48975 , n23825 );
and ( n48977 , n22362 , n21334 );
and ( n48978 , n18608 , n34492 );
or ( n48979 , n48977 , n48978 );
and ( n48980 , n48979 , n23832 );
xor ( n48981 , n23881 , n23889 );
buf ( n48982 , n48981 );
and ( n48983 , n48982 , n21334 );
and ( n48984 , n18608 , n34492 );
or ( n48985 , n48983 , n48984 );
and ( n48986 , n48985 , n23917 );
and ( n48987 , n18608 , n34526 );
or ( n48988 , n48956 , n48966 , n48976 , n48980 , n48986 , n48987 );
and ( n48989 , n48931 , n48988 );
and ( n48990 , n18608 , n17451 );
or ( n48991 , n48989 , n48990 );
and ( n48992 , n48991 , n23924 );
and ( n48993 , n18608 , n23926 );
or ( n48994 , n48992 , n48993 );
buf ( n48995 , n48994 );
buf ( n48996 , n48995 );
buf ( n48997 , n10613 );
not ( n48998 , n34821 );
and ( n48999 , n43526 , n36347 );
and ( n49000 , n13493 , n39408 );
or ( n49001 , n48999 , n49000 );
and ( n49002 , n49001 , n14562 );
and ( n49003 , n43539 , n36348 );
and ( n49004 , n13493 , n39427 );
or ( n49005 , n49003 , n49004 );
and ( n49006 , n49005 , n14586 );
and ( n49007 , n43552 , n36347 );
and ( n49008 , n13493 , n39446 );
or ( n49009 , n49007 , n49008 );
and ( n49010 , n49009 , n14584 );
and ( n49011 , n43539 , n36348 );
and ( n49012 , n13493 , n39453 );
or ( n49013 , n49011 , n49012 );
and ( n49014 , n49013 , n37835 );
and ( n49015 , n43552 , n36348 );
and ( n49016 , n13493 , n39453 );
or ( n49017 , n49015 , n49016 );
and ( n49018 , n49017 , n37841 );
and ( n49019 , n15845 , n36348 );
and ( n49020 , n13493 , n39453 );
or ( n49021 , n49019 , n49020 );
and ( n49022 , n49021 , n37847 );
and ( n49023 , n13493 , n37849 );
or ( n49024 , n49002 , n49006 , n49010 , n49014 , n49018 , n49022 , n49023 );
and ( n49025 , n48998 , n49024 );
and ( n49026 , n13493 , n34821 );
or ( n49027 , n49025 , n49026 );
and ( n49028 , n49027 , n16574 );
and ( n49029 , n13493 , n16576 );
or ( n49030 , n49028 , n49029 );
buf ( n49031 , n49030 );
buf ( n49032 , n49031 );
buf ( n49033 , n10613 );
buf ( n49034 , n10615 );
not ( n49035 , n34821 );
and ( n49036 , n13167 , n14592 );
not ( n49037 , n13916 );
and ( n49038 , n49037 , n13573 );
xor ( n49039 , n13574 , n13881 );
and ( n49040 , n49039 , n13916 );
or ( n49041 , n49038 , n49040 );
buf ( n49042 , n49041 );
and ( n49043 , n49042 , n14137 );
and ( n49044 , n49042 , n14143 );
not ( n49045 , n14139 );
and ( n49046 , n49045 , n36207 );
not ( n49047 , n36245 );
and ( n49048 , n49047 , n36219 );
xor ( n49049 , n47731 , n47732 );
and ( n49050 , n49049 , n36245 );
or ( n49051 , n49048 , n49050 );
buf ( n49052 , n49051 );
and ( n49053 , n49052 , n14139 );
or ( n49054 , n49046 , n49053 );
and ( n49055 , n49054 , n14140 );
and ( n49056 , n36207 , n14141 );
or ( n49057 , n49043 , n49044 , n49055 , n49056 );
and ( n49058 , n49057 , n36350 );
and ( n49059 , n13167 , n43691 );
or ( n49060 , n49058 , n49059 );
and ( n49061 , n49060 , n14562 );
not ( n49062 , n37048 );
and ( n49063 , n49062 , n37010 );
xor ( n49064 , n47752 , n47753 );
and ( n49065 , n49064 , n37048 );
or ( n49066 , n49063 , n49065 );
buf ( n49067 , n49066 );
and ( n49068 , n49067 , n36350 );
and ( n49069 , n13167 , n43703 );
or ( n49070 , n49068 , n49069 );
and ( n49071 , n49070 , n14586 );
not ( n49072 , n37801 );
and ( n49073 , n49072 , n37763 );
xor ( n49074 , n47768 , n47769 );
and ( n49075 , n49074 , n37801 );
or ( n49076 , n49073 , n49075 );
buf ( n49077 , n49076 );
and ( n49078 , n49077 , n36345 );
and ( n49079 , n13167 , n43715 );
or ( n49080 , n49078 , n49079 );
and ( n49081 , n49080 , n14584 );
and ( n49082 , n49067 , n36345 );
and ( n49083 , n13167 , n43721 );
or ( n49084 , n49082 , n49083 );
and ( n49085 , n49084 , n37835 );
and ( n49086 , n49077 , n36345 );
and ( n49087 , n13167 , n43721 );
or ( n49088 , n49086 , n49087 );
and ( n49089 , n49088 , n37841 );
and ( n49090 , n15007 , n14564 );
and ( n49091 , n15007 , n36345 );
and ( n49092 , n13167 , n43721 );
or ( n49093 , n49091 , n49092 );
and ( n49094 , n49093 , n37847 );
or ( n49095 , n49036 , n49061 , n49071 , n49081 , n49085 , n49089 , n49090 , n49094 );
and ( n49096 , n49035 , n49095 );
and ( n49097 , n13167 , n34821 );
or ( n49098 , n49096 , n49097 );
and ( n49099 , n49098 , n16574 );
and ( n49100 , n12252 , n16576 );
or ( n49101 , n49099 , n49100 );
buf ( n49102 , n49101 );
buf ( n49103 , n49102 );
not ( n49104 , n17451 );
and ( n49105 , n18975 , n17873 );
not ( n49106 , n19474 );
and ( n49107 , n49106 , n18961 );
xor ( n49108 , n19488 , n19514 );
and ( n49109 , n49108 , n19474 );
or ( n49110 , n49107 , n49109 );
buf ( n49111 , n49110 );
and ( n49112 , n49111 , n19745 );
and ( n49113 , n49111 , n19748 );
not ( n49114 , n19750 );
and ( n49115 , n49114 , n20877 );
not ( n49116 , n21193 );
and ( n49117 , n49116 , n20889 );
xor ( n49118 , n21207 , n21235 );
and ( n49119 , n49118 , n21193 );
or ( n49120 , n49117 , n49119 );
buf ( n49121 , n49120 );
and ( n49122 , n49121 , n19750 );
or ( n49123 , n49115 , n49122 );
and ( n49124 , n49123 , n21253 );
and ( n49125 , n20877 , n21255 );
or ( n49126 , n49112 , n49113 , n49124 , n49125 );
and ( n49127 , n49126 , n21336 );
and ( n49128 , n18975 , n42682 );
or ( n49129 , n49127 , n49128 );
and ( n49130 , n49129 , n21341 );
not ( n49131 , n22996 );
and ( n49132 , n49131 , n22737 );
xor ( n49133 , n23010 , n23038 );
and ( n49134 , n49133 , n22996 );
or ( n49135 , n49132 , n49134 );
buf ( n49136 , n49135 );
and ( n49137 , n49136 , n21336 );
and ( n49138 , n18975 , n42682 );
or ( n49139 , n49137 , n49138 );
and ( n49140 , n49139 , n23064 );
not ( n49141 , n23758 );
and ( n49142 , n49141 , n23499 );
xor ( n49143 , n23772 , n23800 );
and ( n49144 , n49143 , n23758 );
or ( n49145 , n49142 , n49144 );
buf ( n49146 , n49145 );
and ( n49147 , n49146 , n21336 );
and ( n49148 , n18975 , n42682 );
or ( n49149 , n49147 , n49148 );
and ( n49150 , n49149 , n23825 );
and ( n49151 , n22142 , n21336 );
and ( n49152 , n18975 , n42682 );
or ( n49153 , n49151 , n49152 );
and ( n49154 , n49153 , n23832 );
and ( n49155 , n22142 , n23834 );
xor ( n49156 , n23859 , n23900 );
buf ( n49157 , n49156 );
and ( n49158 , n49157 , n21336 );
and ( n49159 , n18975 , n42682 );
or ( n49160 , n49158 , n49159 );
and ( n49161 , n49160 , n23917 );
or ( n49162 , n49105 , n49130 , n49140 , n49150 , n49154 , n49155 , n49161 );
and ( n49163 , n49104 , n49162 );
and ( n49164 , n18975 , n17451 );
or ( n49165 , n49163 , n49164 );
and ( n49166 , n49165 , n23924 );
and ( n49167 , n18080 , n23926 );
or ( n49168 , n49166 , n49167 );
buf ( n49169 , n49168 );
buf ( n49170 , n49169 );
buf ( n49171 , n10613 );
buf ( n49172 , n10615 );
and ( n49173 , n24061 , n31008 );
and ( n49174 , n29092 , n10618 );
or ( n49175 , n49173 , n49174 );
buf ( n49176 , n49175 );
buf ( n49177 , n49176 );
buf ( n49178 , n10613 );
not ( n49179 , n34821 );
not ( n49180 , n13916 );
and ( n49181 , n49180 , n13595 );
xor ( n49182 , n13596 , n13879 );
and ( n49183 , n49182 , n13916 );
or ( n49184 , n49181 , n49183 );
buf ( n49185 , n49184 );
and ( n49186 , n49185 , n14137 );
and ( n49187 , n49185 , n14143 );
not ( n49188 , n14139 );
and ( n49189 , n49188 , n36163 );
not ( n49190 , n36245 );
and ( n49191 , n49190 , n36175 );
xor ( n49192 , n46403 , n46408 );
and ( n49193 , n49192 , n36245 );
or ( n49194 , n49191 , n49193 );
buf ( n49195 , n49194 );
and ( n49196 , n49195 , n14139 );
or ( n49197 , n49189 , n49196 );
and ( n49198 , n49197 , n14140 );
and ( n49199 , n36163 , n14141 );
or ( n49200 , n49186 , n49187 , n49198 , n49199 );
and ( n49201 , n49200 , n36347 );
and ( n49202 , n13195 , n39408 );
or ( n49203 , n49201 , n49202 );
and ( n49204 , n49203 , n14562 );
not ( n49205 , n37048 );
and ( n49206 , n49205 , n36976 );
xor ( n49207 , n46426 , n46431 );
and ( n49208 , n49207 , n37048 );
or ( n49209 , n49206 , n49208 );
buf ( n49210 , n49209 );
and ( n49211 , n49210 , n36348 );
and ( n49212 , n13195 , n39427 );
or ( n49213 , n49211 , n49212 );
and ( n49214 , n49213 , n14586 );
not ( n49215 , n37801 );
and ( n49216 , n49215 , n37729 );
xor ( n49217 , n46444 , n46449 );
and ( n49218 , n49217 , n37801 );
or ( n49219 , n49216 , n49218 );
buf ( n49220 , n49219 );
and ( n49221 , n49220 , n36347 );
and ( n49222 , n13195 , n39446 );
or ( n49223 , n49221 , n49222 );
and ( n49224 , n49223 , n14584 );
and ( n49225 , n49210 , n36348 );
and ( n49226 , n13195 , n39453 );
or ( n49227 , n49225 , n49226 );
and ( n49228 , n49227 , n37835 );
and ( n49229 , n49220 , n36348 );
and ( n49230 , n13195 , n39453 );
or ( n49231 , n49229 , n49230 );
and ( n49232 , n49231 , n37841 );
and ( n49233 , n15037 , n36348 );
and ( n49234 , n13195 , n39453 );
or ( n49235 , n49233 , n49234 );
and ( n49236 , n49235 , n37847 );
and ( n49237 , n13195 , n37849 );
or ( n49238 , n49204 , n49214 , n49224 , n49228 , n49232 , n49236 , n49237 );
and ( n49239 , n49179 , n49238 );
and ( n49240 , n13195 , n34821 );
or ( n49241 , n49239 , n49240 );
and ( n49242 , n49241 , n16574 );
and ( n49243 , n13195 , n16576 );
or ( n49244 , n49242 , n49243 );
buf ( n49245 , n49244 );
buf ( n49246 , n49245 );
not ( n49247 , n34821 );
and ( n49248 , n47743 , n36345 );
and ( n49249 , n14962 , n36352 );
or ( n49250 , n49248 , n49249 );
and ( n49251 , n49250 , n14562 );
and ( n49252 , n47759 , n36345 );
and ( n49253 , n14962 , n37073 );
or ( n49254 , n49252 , n49253 );
and ( n49255 , n49254 , n14586 );
and ( n49256 , n47775 , n36350 );
and ( n49257 , n14962 , n37825 );
or ( n49258 , n49256 , n49257 );
and ( n49259 , n49258 , n14584 );
and ( n49260 , n47759 , n36350 );
and ( n49261 , n14962 , n37831 );
or ( n49262 , n49260 , n49261 );
and ( n49263 , n49262 , n37835 );
and ( n49264 , n47775 , n36350 );
and ( n49265 , n14962 , n37831 );
or ( n49266 , n49264 , n49265 );
and ( n49267 , n49266 , n37841 );
and ( n49268 , n14977 , n36350 );
and ( n49269 , n14962 , n37831 );
or ( n49270 , n49268 , n49269 );
and ( n49271 , n49270 , n37847 );
and ( n49272 , n14962 , n37849 );
or ( n49273 , n49251 , n49255 , n49259 , n49263 , n49267 , n49271 , n49272 );
and ( n49274 , n49247 , n49273 );
and ( n49275 , n14962 , n34821 );
or ( n49276 , n49274 , n49275 );
and ( n49277 , n49276 , n16574 );
and ( n49278 , n14962 , n16576 );
or ( n49279 , n49277 , n49278 );
buf ( n49280 , n49279 );
buf ( n49281 , n49280 );
buf ( n49282 , n10613 );
buf ( n49283 , n10613 );
buf ( n49284 , n10613 );
buf ( n49285 , n10615 );
buf ( n49286 , n10613 );
buf ( n49287 , n10613 );
buf ( n49288 , n10615 );
not ( n49289 , n34821 );
and ( n49290 , n13311 , n14592 );
and ( n49291 , n45425 , n36350 );
and ( n49292 , n13311 , n43691 );
or ( n49293 , n49291 , n49292 );
and ( n49294 , n49293 , n14562 );
and ( n49295 , n45435 , n36350 );
and ( n49296 , n13311 , n43703 );
or ( n49297 , n49295 , n49296 );
and ( n49298 , n49297 , n14586 );
and ( n49299 , n45445 , n36345 );
and ( n49300 , n13311 , n43715 );
or ( n49301 , n49299 , n49300 );
and ( n49302 , n49301 , n14584 );
and ( n49303 , n45435 , n36345 );
and ( n49304 , n13311 , n43721 );
or ( n49305 , n49303 , n49304 );
and ( n49306 , n49305 , n37835 );
and ( n49307 , n45445 , n36345 );
and ( n49308 , n13311 , n43721 );
or ( n49309 , n49307 , n49308 );
and ( n49310 , n49309 , n37841 );
and ( n49311 , n15537 , n14564 );
and ( n49312 , n15537 , n36345 );
and ( n49313 , n13311 , n43721 );
or ( n49314 , n49312 , n49313 );
and ( n49315 , n49314 , n37847 );
or ( n49316 , n49290 , n49294 , n49298 , n49302 , n49306 , n49310 , n49311 , n49315 );
and ( n49317 , n49289 , n49316 );
and ( n49318 , n13311 , n34821 );
or ( n49319 , n49317 , n49318 );
and ( n49320 , n49319 , n16574 );
and ( n49321 , n12288 , n16576 );
or ( n49322 , n49320 , n49321 );
buf ( n49323 , n49322 );
buf ( n49324 , n49323 );
and ( n49325 , n16833 , n23924 );
and ( n49326 , n22233 , n23926 );
or ( n49327 , n49325 , n49326 );
buf ( n49328 , n49327 );
buf ( n49329 , n49328 );
buf ( n49330 , n10613 );
buf ( n49331 , n10613 );
not ( n49332 , n24800 );
and ( n49333 , n26053 , n25222 );
not ( n49334 , n26823 );
and ( n49335 , n49334 , n26037 );
xor ( n49336 , n31022 , n31031 );
and ( n49337 , n49336 , n26823 );
or ( n49338 , n49335 , n49337 );
buf ( n49339 , n49338 );
and ( n49340 , n49339 , n27046 );
and ( n49341 , n49339 , n27049 );
not ( n49342 , n27051 );
and ( n49343 , n49342 , n27994 );
not ( n49344 , n28494 );
and ( n49345 , n49344 , n28006 );
xor ( n49346 , n31050 , n31059 );
and ( n49347 , n49346 , n28494 );
or ( n49348 , n49345 , n49347 );
buf ( n49349 , n49348 );
and ( n49350 , n49349 , n27051 );
or ( n49351 , n49343 , n49350 );
and ( n49352 , n49351 , n28506 );
and ( n49353 , n27994 , n28508 );
or ( n49354 , n49340 , n49341 , n49352 , n49353 );
and ( n49355 , n49354 , n28583 );
and ( n49356 , n26053 , n28591 );
or ( n49357 , n49355 , n49356 );
and ( n49358 , n49357 , n28594 );
not ( n49359 , n30249 );
and ( n49360 , n49359 , n29854 );
xor ( n49361 , n31085 , n31094 );
and ( n49362 , n49361 , n30249 );
or ( n49363 , n49360 , n49362 );
buf ( n49364 , n49363 );
and ( n49365 , n49364 , n28583 );
and ( n49366 , n26053 , n28591 );
or ( n49367 , n49365 , n49366 );
and ( n49368 , n49367 , n30269 );
not ( n49369 , n30963 );
and ( n49370 , n49369 , n30568 );
xor ( n49371 , n31113 , n31122 );
and ( n49372 , n49371 , n30963 );
or ( n49373 , n49370 , n49372 );
buf ( n49374 , n49373 );
and ( n49375 , n49374 , n28583 );
and ( n49376 , n26053 , n28591 );
or ( n49377 , n49375 , n49376 );
and ( n49378 , n49377 , n30982 );
and ( n49379 , n29555 , n28583 );
and ( n49380 , n26053 , n28591 );
or ( n49381 , n49379 , n49380 );
and ( n49382 , n49381 , n30989 );
and ( n49383 , n26051 , n30991 );
xor ( n49384 , n31149 , n31162 );
buf ( n49385 , n49384 );
and ( n49386 , n49385 , n28583 );
and ( n49387 , n26053 , n28591 );
or ( n49388 , n49386 , n49387 );
and ( n49389 , n49388 , n31002 );
or ( n49390 , n49333 , n49358 , n49368 , n49378 , n49382 , n49383 , n49389 );
and ( n49391 , n49332 , n49390 );
and ( n49392 , n26053 , n24800 );
or ( n49393 , n49391 , n49392 );
and ( n49394 , n49393 , n31008 );
and ( n49395 , n26053 , n10618 );
or ( n49396 , n49394 , n49395 );
buf ( n49397 , n49396 );
buf ( n49398 , n49397 );
buf ( n49399 , n10615 );
buf ( n49400 , n10615 );
not ( n49401 , n24800 );
and ( n49402 , n48044 , n28586 );
and ( n49403 , n26667 , n34573 );
or ( n49404 , n49402 , n49403 );
and ( n49405 , n49404 , n28594 );
and ( n49406 , n48054 , n28586 );
and ( n49407 , n26667 , n34573 );
or ( n49408 , n49406 , n49407 );
and ( n49409 , n49408 , n30269 );
and ( n49410 , n48064 , n28586 );
and ( n49411 , n26667 , n34573 );
or ( n49412 , n49410 , n49411 );
and ( n49413 , n49412 , n30982 );
and ( n49414 , n29185 , n28586 );
and ( n49415 , n26667 , n34573 );
or ( n49416 , n49414 , n49415 );
and ( n49417 , n49416 , n30989 );
and ( n49418 , n48075 , n28586 );
and ( n49419 , n26667 , n34573 );
or ( n49420 , n49418 , n49419 );
and ( n49421 , n49420 , n31002 );
and ( n49422 , n26667 , n34607 );
or ( n49423 , n49405 , n49409 , n49413 , n49417 , n49421 , n49422 );
and ( n49424 , n49401 , n49423 );
and ( n49425 , n26667 , n24800 );
or ( n49426 , n49424 , n49425 );
and ( n49427 , n49426 , n31008 );
and ( n49428 , n26667 , n10618 );
or ( n49429 , n49427 , n49428 );
buf ( n49430 , n49429 );
buf ( n49431 , n49430 );
buf ( n49432 , n10613 );
buf ( n49433 , n10615 );
buf ( n49434 , n10615 );
not ( n49435 , n17451 );
and ( n49436 , n18875 , n17873 );
and ( n49437 , n42969 , n21330 );
and ( n49438 , n18875 , n21338 );
or ( n49439 , n49437 , n49438 );
and ( n49440 , n49439 , n21341 );
and ( n49441 , n42979 , n21330 );
and ( n49442 , n18875 , n21338 );
or ( n49443 , n49441 , n49442 );
and ( n49444 , n49443 , n23064 );
and ( n49445 , n42989 , n21330 );
and ( n49446 , n18875 , n21338 );
or ( n49447 , n49445 , n49446 );
and ( n49448 , n49447 , n23825 );
and ( n49449 , n22202 , n21330 );
and ( n49450 , n18875 , n21338 );
or ( n49451 , n49449 , n49450 );
and ( n49452 , n49451 , n23832 );
and ( n49453 , n18873 , n23834 );
and ( n49454 , n42999 , n21330 );
and ( n49455 , n18875 , n21338 );
or ( n49456 , n49454 , n49455 );
and ( n49457 , n49456 , n23917 );
or ( n49458 , n49436 , n49440 , n49444 , n49448 , n49452 , n49453 , n49457 );
and ( n49459 , n49435 , n49458 );
and ( n49460 , n18875 , n17451 );
or ( n49461 , n49459 , n49460 );
and ( n49462 , n49461 , n23924 );
and ( n49463 , n18875 , n23926 );
or ( n49464 , n49462 , n49463 );
buf ( n49465 , n49464 );
buf ( n49466 , n49465 );
buf ( n49467 , n10613 );
buf ( n49468 , n10613 );
buf ( n49469 , n10615 );
buf ( n49470 , n10613 );
buf ( n49471 , n10613 );
not ( n49472 , n24511 );
not ( n49473 , n24799 );
and ( n49474 , n10670 , n40154 );
not ( n49475 , n40632 );
and ( n49476 , n49475 , n40526 );
xor ( n49477 , n40637 , n40663 );
and ( n49478 , n49477 , n40632 );
or ( n49479 , n49476 , n49478 );
buf ( n49480 , n49479 );
and ( n49481 , n49480 , n27046 );
not ( n49482 , n41147 );
and ( n49483 , n49482 , n41041 );
xor ( n49484 , n41152 , n41178 );
and ( n49485 , n49484 , n41147 );
or ( n49486 , n49483 , n49485 );
buf ( n49487 , n49486 );
and ( n49488 , n49487 , n27049 );
and ( n49489 , n29413 , n28506 );
and ( n49490 , n10670 , n28508 );
or ( n49491 , n49481 , n49488 , n49489 , n49490 );
and ( n49492 , n49491 , n41199 );
or ( n49493 , n49474 , n49492 );
and ( n49494 , n49473 , n49493 );
xor ( n49495 , n41548 , n41556 );
xor ( n49496 , n49495 , n41800 );
buf ( n49497 , n49496 );
and ( n49498 , n49497 , n27046 );
xor ( n49499 , n42141 , n42142 );
xor ( n49500 , n49499 , n42296 );
buf ( n49501 , n49500 );
and ( n49502 , n49501 , n27049 );
and ( n49503 , n29413 , n42306 );
or ( n49504 , n49498 , n49502 , n49503 );
buf ( n49505 , n49504 );
and ( n49506 , C1 , n49505 );
or ( n49507 , n49506 , C0 );
buf ( n49508 , n49507 );
not ( n49509 , n49508 );
buf ( n49510 , n49509 );
buf ( n49511 , n49510 );
not ( n49512 , n49511 );
and ( n49513 , C1 , n49512 );
or ( n49514 , n49513 , C0 );
buf ( n49515 , n49514 );
and ( n49516 , n49515 , n24799 );
or ( n49517 , n49494 , n49516 );
and ( n49518 , n49472 , n49517 );
and ( n49519 , n49491 , n24511 );
or ( n49520 , n49518 , n49519 );
and ( n49521 , n49520 , n31008 );
not ( n49522 , n42601 );
and ( n49523 , n49522 , n42513 );
xor ( n49524 , n42606 , n42632 );
and ( n49525 , n49524 , n42601 );
or ( n49526 , n49523 , n49525 );
buf ( n49527 , n49526 );
and ( n49528 , n49527 , n10618 );
or ( n49529 , n49521 , n49528 );
buf ( n49530 , n49529 );
buf ( n49531 , n49530 );
not ( n49532 , n34804 );
and ( n49533 , n49532 , n25991 );
and ( n49534 , n14809 , n34804 );
or ( n49535 , n49533 , n49534 );
and ( n49536 , n49535 , n31008 );
and ( n49537 , n14809 , n10618 );
or ( n49538 , n49536 , n49537 );
buf ( n49539 , n49538 );
buf ( n49540 , n49539 );
not ( n49541 , n24800 );
not ( n49542 , n26823 );
and ( n49543 , n49542 , n26717 );
xor ( n49544 , n45230 , n45231 );
and ( n49545 , n49544 , n26823 );
or ( n49546 , n49543 , n49545 );
buf ( n49547 , n49546 );
and ( n49548 , n49547 , n27046 );
and ( n49549 , n49547 , n27049 );
not ( n49550 , n27051 );
and ( n49551 , n49550 , n28434 );
not ( n49552 , n28494 );
and ( n49553 , n49552 , n28446 );
xor ( n49554 , n45246 , n45247 );
and ( n49555 , n49554 , n28494 );
or ( n49556 , n49553 , n49555 );
buf ( n49557 , n49556 );
and ( n49558 , n49557 , n27051 );
or ( n49559 , n49551 , n49558 );
and ( n49560 , n49559 , n28506 );
and ( n49561 , n28434 , n28508 );
or ( n49562 , n49548 , n49549 , n49560 , n49561 );
and ( n49563 , n49562 , n28587 );
and ( n49564 , n26737 , n39807 );
or ( n49565 , n49563 , n49564 );
and ( n49566 , n49565 , n28594 );
not ( n49567 , n30249 );
and ( n49568 , n49567 , n30194 );
xor ( n49569 , n45267 , n45268 );
and ( n49570 , n49569 , n30249 );
or ( n49571 , n49568 , n49570 );
buf ( n49572 , n49571 );
and ( n49573 , n49572 , n28587 );
and ( n49574 , n26737 , n39807 );
or ( n49575 , n49573 , n49574 );
and ( n49576 , n49575 , n30269 );
not ( n49577 , n30963 );
and ( n49578 , n49577 , n30908 );
xor ( n49579 , n45283 , n45284 );
and ( n49580 , n49579 , n30963 );
or ( n49581 , n49578 , n49580 );
buf ( n49582 , n49581 );
and ( n49583 , n49582 , n28587 );
and ( n49584 , n26737 , n39807 );
or ( n49585 , n49583 , n49584 );
and ( n49586 , n49585 , n30982 );
and ( n49587 , n29159 , n28587 );
and ( n49588 , n26737 , n39807 );
or ( n49589 , n49587 , n49588 );
and ( n49590 , n49589 , n30989 );
xor ( n49591 , n45305 , n45306 );
buf ( n49592 , n49591 );
and ( n49593 , n49592 , n28587 );
and ( n49594 , n26737 , n39807 );
or ( n49595 , n49593 , n49594 );
and ( n49596 , n49595 , n31002 );
and ( n49597 , n26737 , n34607 );
or ( n49598 , n49566 , n49576 , n49586 , n49590 , n49596 , n49597 );
and ( n49599 , n49541 , n49598 );
and ( n49600 , n26737 , n24800 );
or ( n49601 , n49599 , n49600 );
and ( n49602 , n49601 , n31008 );
and ( n49603 , n26737 , n10618 );
or ( n49604 , n49602 , n49603 );
buf ( n49605 , n49604 );
buf ( n49606 , n49605 );
buf ( n49607 , n10613 );
buf ( n49608 , n10615 );
buf ( n49609 , n10613 );
and ( n49610 , n16825 , n23924 );
and ( n49611 , n22213 , n23926 );
or ( n49612 , n49610 , n49611 );
buf ( n49613 , n49612 );
buf ( n49614 , n49613 );
buf ( n49615 , n10615 );
buf ( n49616 , n10613 );
buf ( n49617 , n10613 );
buf ( n49618 , n10613 );
buf ( n49619 , n10613 );
buf ( n49620 , n10613 );
buf ( n49621 , n10613 );
buf ( n49622 , n10615 );
buf ( n49623 , n10613 );
not ( n49624 , n24800 );
and ( n49625 , n47642 , n28586 );
and ( n49626 , n26463 , n34573 );
or ( n49627 , n49625 , n49626 );
and ( n49628 , n49627 , n28594 );
and ( n49629 , n47652 , n28586 );
and ( n49630 , n26463 , n34573 );
or ( n49631 , n49629 , n49630 );
and ( n49632 , n49631 , n30269 );
and ( n49633 , n47662 , n28586 );
and ( n49634 , n26463 , n34573 );
or ( n49635 , n49633 , n49634 );
and ( n49636 , n49635 , n30982 );
and ( n49637 , n29315 , n28586 );
and ( n49638 , n26463 , n34573 );
or ( n49639 , n49637 , n49638 );
and ( n49640 , n49639 , n30989 );
and ( n49641 , n47672 , n28586 );
and ( n49642 , n26463 , n34573 );
or ( n49643 , n49641 , n49642 );
and ( n49644 , n49643 , n31002 );
and ( n49645 , n26463 , n34607 );
or ( n49646 , n49628 , n49632 , n49636 , n49640 , n49644 , n49645 );
and ( n49647 , n49624 , n49646 );
and ( n49648 , n26463 , n24800 );
or ( n49649 , n49647 , n49648 );
and ( n49650 , n49649 , n31008 );
and ( n49651 , n26463 , n10618 );
or ( n49652 , n49650 , n49651 );
buf ( n49653 , n49652 );
buf ( n49654 , n49653 );
buf ( n49655 , n10613 );
not ( n49656 , n34821 );
and ( n49657 , n13325 , n14592 );
and ( n49658 , n48669 , n36348 );
and ( n49659 , n13325 , n43530 );
or ( n49660 , n49658 , n49659 );
and ( n49661 , n49660 , n14562 );
and ( n49662 , n48679 , n36347 );
and ( n49663 , n13325 , n43543 );
or ( n49664 , n49662 , n49663 );
and ( n49665 , n49664 , n14586 );
and ( n49666 , n48689 , n36348 );
and ( n49667 , n13325 , n43556 );
or ( n49668 , n49666 , n49667 );
and ( n49669 , n49668 , n14584 );
and ( n49670 , n48679 , n36347 );
and ( n49671 , n13325 , n43563 );
or ( n49672 , n49670 , n49671 );
and ( n49673 , n49672 , n37835 );
and ( n49674 , n48689 , n36347 );
and ( n49675 , n13325 , n43563 );
or ( n49676 , n49674 , n49675 );
and ( n49677 , n49676 , n37841 );
and ( n49678 , n13323 , n14564 );
and ( n49679 , n15559 , n36347 );
and ( n49680 , n13325 , n43563 );
or ( n49681 , n49679 , n49680 );
and ( n49682 , n49681 , n37847 );
or ( n49683 , n49657 , n49661 , n49665 , n49669 , n49673 , n49677 , n49678 , n49682 );
and ( n49684 , n49656 , n49683 );
and ( n49685 , n13325 , n34821 );
or ( n49686 , n49684 , n49685 );
and ( n49687 , n49686 , n16574 );
and ( n49688 , n13325 , n16576 );
or ( n49689 , n49687 , n49688 );
buf ( n49690 , n49689 );
buf ( n49691 , n49690 );
buf ( n49692 , n10613 );
buf ( n49693 , n10615 );
buf ( n49694 , n10615 );
buf ( n49695 , n10615 );
buf ( n49696 , n10615 );
buf ( n49697 , n10613 );
buf ( n49698 , n10613 );
not ( n49699 , n17162 );
not ( n49700 , n17450 );
and ( n49701 , n10728 , n37947 );
not ( n49702 , n38425 );
and ( n49703 , n49702 , n38115 );
xor ( n49704 , n38439 , n38441 );
and ( n49705 , n49704 , n38425 );
or ( n49706 , n49703 , n49705 );
buf ( n49707 , n49706 );
and ( n49708 , n49707 , n19745 );
not ( n49709 , n38934 );
and ( n49710 , n49709 , n38624 );
xor ( n49711 , n38948 , n38950 );
and ( n49712 , n49711 , n38934 );
or ( n49713 , n49710 , n49712 );
buf ( n49714 , n49713 );
and ( n49715 , n49714 , n19748 );
and ( n49716 , n22400 , n21253 );
and ( n49717 , n10728 , n21255 );
or ( n49718 , n49708 , n49715 , n49716 , n49717 );
and ( n49719 , n49718 , n38980 );
or ( n49720 , n49701 , n49719 );
and ( n49721 , n49700 , n49720 );
or ( n49722 , n49721 , C0 );
and ( n49723 , n49699 , n49722 );
and ( n49724 , n49718 , n17162 );
or ( n49725 , n49723 , n49724 );
and ( n49726 , n49725 , n23924 );
not ( n49727 , n39264 );
and ( n49728 , n49727 , n39008 );
xor ( n49729 , n39278 , n39280 );
and ( n49730 , n49729 , n39264 );
or ( n49731 , n49728 , n49730 );
buf ( n49732 , n49731 );
and ( n49733 , n49732 , n23926 );
or ( n49734 , n49726 , n49733 );
buf ( n49735 , n49734 );
buf ( n49736 , n49735 );
buf ( n49737 , n10613 );
buf ( n49738 , n10615 );
not ( n49739 , n34804 );
and ( n49740 , n49739 , n26399 );
and ( n49741 , n14737 , n34804 );
or ( n49742 , n49740 , n49741 );
and ( n49743 , n49742 , n31008 );
and ( n49744 , n14737 , n10618 );
or ( n49745 , n49743 , n49744 );
buf ( n49746 , n49745 );
buf ( n49747 , n49746 );
buf ( n49748 , n10615 );
buf ( n49749 , n10613 );
buf ( n49750 , n10615 );
not ( n49751 , n17162 );
not ( n49752 , n17450 );
and ( n49753 , n10708 , n37947 );
not ( n49754 , n38425 );
and ( n49755 , n49754 , n38183 );
xor ( n49756 , n38435 , n38445 );
and ( n49757 , n49756 , n38425 );
or ( n49758 , n49755 , n49757 );
buf ( n49759 , n49758 );
and ( n49760 , n49759 , n19745 );
not ( n49761 , n38934 );
and ( n49762 , n49761 , n38692 );
xor ( n49763 , n38944 , n38954 );
and ( n49764 , n49763 , n38934 );
or ( n49765 , n49762 , n49764 );
buf ( n49766 , n49765 );
and ( n49767 , n49766 , n19748 );
and ( n49768 , n22320 , n21253 );
and ( n49769 , n10708 , n21255 );
or ( n49770 , n49760 , n49767 , n49768 , n49769 );
and ( n49771 , n49770 , n38980 );
or ( n49772 , n49753 , n49771 );
and ( n49773 , n49752 , n49772 );
or ( n49774 , n49773 , C0 );
and ( n49775 , n49751 , n49774 );
and ( n49776 , n49770 , n17162 );
or ( n49777 , n49775 , n49776 );
and ( n49778 , n49777 , n23924 );
not ( n49779 , n39264 );
and ( n49780 , n49779 , n39064 );
xor ( n49781 , n39274 , n39284 );
and ( n49782 , n49781 , n39264 );
or ( n49783 , n49780 , n49782 );
buf ( n49784 , n49783 );
and ( n49785 , n49784 , n23926 );
or ( n49786 , n49778 , n49785 );
buf ( n49787 , n49786 );
buf ( n49788 , n49787 );
buf ( n49789 , n10615 );
buf ( n49790 , n10615 );
not ( n49791 , n17451 );
and ( n49792 , n19450 , n17873 );
and ( n49793 , n45354 , n21336 );
and ( n49794 , n19450 , n42682 );
or ( n49795 , n49793 , n49794 );
and ( n49796 , n49795 , n21341 );
and ( n49797 , n45364 , n21336 );
and ( n49798 , n19450 , n42682 );
or ( n49799 , n49797 , n49798 );
and ( n49800 , n49799 , n23064 );
and ( n49801 , n45374 , n21336 );
and ( n49802 , n19450 , n42682 );
or ( n49803 , n49801 , n49802 );
and ( n49804 , n49803 , n23825 );
and ( n49805 , n21880 , n21336 );
and ( n49806 , n19450 , n42682 );
or ( n49807 , n49805 , n49806 );
and ( n49808 , n49807 , n23832 );
and ( n49809 , n21880 , n23834 );
and ( n49810 , n45384 , n21336 );
and ( n49811 , n19450 , n42682 );
or ( n49812 , n49810 , n49811 );
and ( n49813 , n49812 , n23917 );
or ( n49814 , n49792 , n49796 , n49800 , n49804 , n49808 , n49809 , n49813 );
and ( n49815 , n49791 , n49814 );
and ( n49816 , n19450 , n17451 );
or ( n49817 , n49815 , n49816 );
and ( n49818 , n49817 , n23924 );
and ( n49819 , n18290 , n23926 );
or ( n49820 , n49818 , n49819 );
buf ( n49821 , n49820 );
buf ( n49822 , n49821 );
buf ( n49823 , n10613 );
buf ( n49824 , n10615 );
not ( n49825 , n24800 );
not ( n49826 , n26823 );
and ( n49827 , n49826 , n26105 );
xor ( n49828 , n31020 , n31033 );
and ( n49829 , n49828 , n26823 );
or ( n49830 , n49827 , n49829 );
buf ( n49831 , n49830 );
and ( n49832 , n49831 , n27046 );
and ( n49833 , n49831 , n27049 );
not ( n49834 , n27051 );
and ( n49835 , n49834 , n28038 );
not ( n49836 , n28494 );
and ( n49837 , n49836 , n28050 );
xor ( n49838 , n31048 , n31061 );
and ( n49839 , n49838 , n28494 );
or ( n49840 , n49837 , n49839 );
buf ( n49841 , n49840 );
and ( n49842 , n49841 , n27051 );
or ( n49843 , n49835 , n49842 );
and ( n49844 , n49843 , n28506 );
and ( n49845 , n28038 , n28508 );
or ( n49846 , n49832 , n49833 , n49844 , n49845 );
and ( n49847 , n49846 , n28586 );
and ( n49848 , n26123 , n34573 );
or ( n49849 , n49847 , n49848 );
and ( n49850 , n49849 , n28594 );
not ( n49851 , n30249 );
and ( n49852 , n49851 , n29888 );
xor ( n49853 , n31083 , n31096 );
and ( n49854 , n49853 , n30249 );
or ( n49855 , n49852 , n49854 );
buf ( n49856 , n49855 );
and ( n49857 , n49856 , n28586 );
and ( n49858 , n26123 , n34573 );
or ( n49859 , n49857 , n49858 );
and ( n49860 , n49859 , n30269 );
not ( n49861 , n30963 );
and ( n49862 , n49861 , n30602 );
xor ( n49863 , n31111 , n31124 );
and ( n49864 , n49863 , n30963 );
or ( n49865 , n49862 , n49864 );
buf ( n49866 , n49865 );
and ( n49867 , n49866 , n28586 );
and ( n49868 , n26123 , n34573 );
or ( n49869 , n49867 , n49868 );
and ( n49870 , n49869 , n30982 );
and ( n49871 , n29515 , n28586 );
and ( n49872 , n26123 , n34573 );
or ( n49873 , n49871 , n49872 );
and ( n49874 , n49873 , n30989 );
xor ( n49875 , n31145 , n31164 );
buf ( n49876 , n49875 );
and ( n49877 , n49876 , n28586 );
and ( n49878 , n26123 , n34573 );
or ( n49879 , n49877 , n49878 );
and ( n49880 , n49879 , n31002 );
and ( n49881 , n26123 , n34607 );
or ( n49882 , n49850 , n49860 , n49870 , n49874 , n49880 , n49881 );
and ( n49883 , n49825 , n49882 );
and ( n49884 , n26123 , n24800 );
or ( n49885 , n49883 , n49884 );
and ( n49886 , n49885 , n31008 );
and ( n49887 , n26123 , n10618 );
or ( n49888 , n49886 , n49887 );
buf ( n49889 , n49888 );
buf ( n49890 , n49889 );
buf ( n49891 , n10613 );
buf ( n49892 , n10613 );
buf ( n49893 , n23926 );
buf ( n49894 , n49893 );
not ( n49895 , n17451 );
and ( n49896 , n19317 , n17873 );
and ( n49897 , n39576 , n21330 );
and ( n49898 , n19317 , n21338 );
or ( n49899 , n49897 , n49898 );
and ( n49900 , n49899 , n21341 );
and ( n49901 , n39586 , n21330 );
and ( n49902 , n19317 , n21338 );
or ( n49903 , n49901 , n49902 );
and ( n49904 , n49903 , n23064 );
and ( n49905 , n39596 , n21330 );
and ( n49906 , n19317 , n21338 );
or ( n49907 , n49905 , n49906 );
and ( n49908 , n49907 , n23825 );
and ( n49909 , n21932 , n21330 );
and ( n49910 , n19317 , n21338 );
or ( n49911 , n49909 , n49910 );
and ( n49912 , n49911 , n23832 );
and ( n49913 , n19315 , n23834 );
and ( n49914 , n39606 , n21330 );
and ( n49915 , n19317 , n21338 );
or ( n49916 , n49914 , n49915 );
and ( n49917 , n49916 , n23917 );
or ( n49918 , n49896 , n49900 , n49904 , n49908 , n49912 , n49913 , n49917 );
and ( n49919 , n49895 , n49918 );
and ( n49920 , n19317 , n17451 );
or ( n49921 , n49919 , n49920 );
and ( n49922 , n49921 , n23924 );
and ( n49923 , n19317 , n23926 );
or ( n49924 , n49922 , n49923 );
buf ( n49925 , n49924 );
buf ( n49926 , n49925 );
not ( n49927 , n17451 );
and ( n49928 , n18805 , n17873 );
and ( n49929 , n46858 , n21336 );
and ( n49930 , n18805 , n42682 );
or ( n49931 , n49929 , n49930 );
and ( n49932 , n49931 , n21341 );
and ( n49933 , n46868 , n21336 );
and ( n49934 , n18805 , n42682 );
or ( n49935 , n49933 , n49934 );
and ( n49936 , n49935 , n23064 );
and ( n49937 , n46878 , n21336 );
and ( n49938 , n18805 , n42682 );
or ( n49939 , n49937 , n49938 );
and ( n49940 , n49939 , n23825 );
and ( n49941 , n22242 , n21336 );
and ( n49942 , n18805 , n42682 );
or ( n49943 , n49941 , n49942 );
and ( n49944 , n49943 , n23832 );
and ( n49945 , n22242 , n23834 );
and ( n49946 , n46888 , n21336 );
and ( n49947 , n18805 , n42682 );
or ( n49948 , n49946 , n49947 );
and ( n49949 , n49948 , n23917 );
or ( n49950 , n49928 , n49932 , n49936 , n49940 , n49944 , n49945 , n49949 );
and ( n49951 , n49927 , n49950 );
and ( n49952 , n18805 , n17451 );
or ( n49953 , n49951 , n49952 );
and ( n49954 , n49953 , n23924 );
and ( n49955 , n18005 , n23926 );
or ( n49956 , n49954 , n49955 );
buf ( n49957 , n49956 );
buf ( n49958 , n49957 );
not ( n49959 , n11333 );
and ( n49960 , n49959 , n11074 );
xor ( n49961 , n11347 , n11355 );
and ( n49962 , n49961 , n11333 );
or ( n49963 , n49960 , n49962 );
buf ( n49964 , n49963 );
buf ( n49965 , n49964 );
buf ( n49966 , n10615 );
buf ( n49967 , n10615 );
buf ( n49968 , n10613 );
buf ( n49969 , n10615 );
buf ( n49970 , n10613 );
buf ( n49971 , n10613 );
buf ( n49972 , n10613 );
and ( n49973 , n11768 , n16574 );
and ( n49974 , n14950 , n16576 );
or ( n49975 , n49973 , n49974 );
buf ( n49976 , n49975 );
buf ( n49977 , n49976 );
buf ( n49978 , n10613 );
not ( n49979 , n24800 );
and ( n49980 , n26155 , n25222 );
not ( n49981 , n26823 );
and ( n49982 , n49981 , n26139 );
xor ( n49983 , n31019 , n31034 );
and ( n49984 , n49983 , n26823 );
or ( n49985 , n49982 , n49984 );
buf ( n49986 , n49985 );
and ( n49987 , n49986 , n27046 );
and ( n49988 , n49986 , n27049 );
not ( n49989 , n27051 );
and ( n49990 , n49989 , n28060 );
not ( n49991 , n28494 );
and ( n49992 , n49991 , n28072 );
xor ( n49993 , n31047 , n31062 );
and ( n49994 , n49993 , n28494 );
or ( n49995 , n49992 , n49994 );
buf ( n49996 , n49995 );
and ( n49997 , n49996 , n27051 );
or ( n49998 , n49990 , n49997 );
and ( n49999 , n49998 , n28506 );
and ( n50000 , n28060 , n28508 );
or ( n50001 , n49987 , n49988 , n49999 , n50000 );
and ( n50002 , n50001 , n28583 );
and ( n50003 , n26155 , n28591 );
or ( n50004 , n50002 , n50003 );
and ( n50005 , n50004 , n28594 );
not ( n50006 , n30249 );
and ( n50007 , n50006 , n29905 );
xor ( n50008 , n31082 , n31097 );
and ( n50009 , n50008 , n30249 );
or ( n50010 , n50007 , n50009 );
buf ( n50011 , n50010 );
and ( n50012 , n50011 , n28583 );
and ( n50013 , n26155 , n28591 );
or ( n50014 , n50012 , n50013 );
and ( n50015 , n50014 , n30269 );
not ( n50016 , n30963 );
and ( n50017 , n50016 , n30619 );
xor ( n50018 , n31110 , n31125 );
and ( n50019 , n50018 , n30963 );
or ( n50020 , n50017 , n50019 );
buf ( n50021 , n50020 );
and ( n50022 , n50021 , n28583 );
and ( n50023 , n26155 , n28591 );
or ( n50024 , n50022 , n50023 );
and ( n50025 , n50024 , n30982 );
and ( n50026 , n29495 , n28583 );
and ( n50027 , n26155 , n28591 );
or ( n50028 , n50026 , n50027 );
and ( n50029 , n50028 , n30989 );
and ( n50030 , n26153 , n30991 );
xor ( n50031 , n31143 , n31165 );
buf ( n50032 , n50031 );
and ( n50033 , n50032 , n28583 );
and ( n50034 , n26155 , n28591 );
or ( n50035 , n50033 , n50034 );
and ( n50036 , n50035 , n31002 );
or ( n50037 , n49980 , n50005 , n50015 , n50025 , n50029 , n50030 , n50036 );
and ( n50038 , n49979 , n50037 );
and ( n50039 , n26155 , n24800 );
or ( n50040 , n50038 , n50039 );
and ( n50041 , n50040 , n31008 );
and ( n50042 , n26155 , n10618 );
or ( n50043 , n50041 , n50042 );
buf ( n50044 , n50043 );
buf ( n50045 , n50044 );
buf ( n50046 , n10613 );
buf ( n50047 , n10615 );
not ( n50048 , n17451 );
and ( n50049 , n46760 , n21333 );
and ( n50050 , n19149 , n34758 );
or ( n50051 , n50049 , n50050 );
and ( n50052 , n50051 , n21341 );
and ( n50053 , n46770 , n21333 );
and ( n50054 , n19149 , n34758 );
or ( n50055 , n50053 , n50054 );
and ( n50056 , n50055 , n23064 );
and ( n50057 , n46780 , n21333 );
and ( n50058 , n19149 , n34758 );
or ( n50059 , n50057 , n50058 );
and ( n50060 , n50059 , n23825 );
and ( n50061 , n22042 , n21333 );
and ( n50062 , n19149 , n34758 );
or ( n50063 , n50061 , n50062 );
and ( n50064 , n50063 , n23832 );
and ( n50065 , n46791 , n21333 );
and ( n50066 , n19149 , n34758 );
or ( n50067 , n50065 , n50066 );
and ( n50068 , n50067 , n23917 );
and ( n50069 , n19149 , n34526 );
or ( n50070 , n50052 , n50056 , n50060 , n50064 , n50068 , n50069 );
and ( n50071 , n50048 , n50070 );
and ( n50072 , n19149 , n17451 );
or ( n50073 , n50071 , n50072 );
and ( n50074 , n50073 , n23924 );
and ( n50075 , n19149 , n23926 );
or ( n50076 , n50074 , n50075 );
buf ( n50077 , n50076 );
buf ( n50078 , n50077 );
buf ( n50079 , n10613 );
buf ( n50080 , n10613 );
buf ( n50081 , n10615 );
not ( n50082 , n34821 );
and ( n50083 , n13395 , n14592 );
and ( n50084 , n48401 , n36350 );
and ( n50085 , n13395 , n43691 );
or ( n50086 , n50084 , n50085 );
and ( n50087 , n50086 , n14562 );
and ( n50088 , n48411 , n36350 );
and ( n50089 , n13395 , n43703 );
or ( n50090 , n50088 , n50089 );
and ( n50091 , n50090 , n14586 );
and ( n50092 , n48421 , n36345 );
and ( n50093 , n13395 , n43715 );
or ( n50094 , n50092 , n50093 );
and ( n50095 , n50094 , n14584 );
and ( n50096 , n48411 , n36345 );
and ( n50097 , n13395 , n43721 );
or ( n50098 , n50096 , n50097 );
and ( n50099 , n50098 , n37835 );
and ( n50100 , n48421 , n36345 );
and ( n50101 , n13395 , n43721 );
or ( n50102 , n50100 , n50101 );
and ( n50103 , n50102 , n37841 );
and ( n50104 , n15691 , n14564 );
and ( n50105 , n15691 , n36345 );
and ( n50106 , n13395 , n43721 );
or ( n50107 , n50105 , n50106 );
and ( n50108 , n50107 , n37847 );
or ( n50109 , n50083 , n50087 , n50091 , n50095 , n50099 , n50103 , n50104 , n50108 );
and ( n50110 , n50082 , n50109 );
and ( n50111 , n13395 , n34821 );
or ( n50112 , n50110 , n50111 );
and ( n50113 , n50112 , n16574 );
and ( n50114 , n12309 , n16576 );
or ( n50115 , n50113 , n50114 );
buf ( n50116 , n50115 );
buf ( n50117 , n50116 );
not ( n50118 , n34804 );
and ( n50119 , n50118 , n26127 );
and ( n50120 , n14785 , n34804 );
or ( n50121 , n50119 , n50120 );
and ( n50122 , n50121 , n31008 );
and ( n50123 , n14785 , n10618 );
or ( n50124 , n50122 , n50123 );
buf ( n50125 , n50124 );
buf ( n50126 , n50125 );
buf ( n50127 , n10613 );
buf ( n50128 , n10615 );
not ( n50129 , n24800 );
and ( n50130 , n26087 , n25222 );
and ( n50131 , n37895 , n28583 );
and ( n50132 , n26087 , n28591 );
or ( n50133 , n50131 , n50132 );
and ( n50134 , n50133 , n28594 );
and ( n50135 , n37905 , n28583 );
and ( n50136 , n26087 , n28591 );
or ( n50137 , n50135 , n50136 );
and ( n50138 , n50137 , n30269 );
and ( n50139 , n37915 , n28583 );
and ( n50140 , n26087 , n28591 );
or ( n50141 , n50139 , n50140 );
and ( n50142 , n50141 , n30982 );
and ( n50143 , n29535 , n28583 );
and ( n50144 , n26087 , n28591 );
or ( n50145 , n50143 , n50144 );
and ( n50146 , n50145 , n30989 );
and ( n50147 , n26085 , n30991 );
and ( n50148 , n37925 , n28583 );
and ( n50149 , n26087 , n28591 );
or ( n50150 , n50148 , n50149 );
and ( n50151 , n50150 , n31002 );
or ( n50152 , n50130 , n50134 , n50138 , n50142 , n50146 , n50147 , n50151 );
and ( n50153 , n50129 , n50152 );
and ( n50154 , n26087 , n24800 );
or ( n50155 , n50153 , n50154 );
and ( n50156 , n50155 , n31008 );
and ( n50157 , n26087 , n10618 );
or ( n50158 , n50156 , n50157 );
buf ( n50159 , n50158 );
buf ( n50160 , n50159 );
not ( n50161 , n24800 );
and ( n50162 , n49562 , n28586 );
and ( n50163 , n26735 , n34573 );
or ( n50164 , n50162 , n50163 );
and ( n50165 , n50164 , n28594 );
and ( n50166 , n49572 , n28586 );
and ( n50167 , n26735 , n34573 );
or ( n50168 , n50166 , n50167 );
and ( n50169 , n50168 , n30269 );
and ( n50170 , n49582 , n28586 );
and ( n50171 , n26735 , n34573 );
or ( n50172 , n50170 , n50171 );
and ( n50173 , n50172 , n30982 );
and ( n50174 , n29159 , n28586 );
and ( n50175 , n26735 , n34573 );
or ( n50176 , n50174 , n50175 );
and ( n50177 , n50176 , n30989 );
and ( n50178 , n49592 , n28586 );
and ( n50179 , n26735 , n34573 );
or ( n50180 , n50178 , n50179 );
and ( n50181 , n50180 , n31002 );
and ( n50182 , n26735 , n34607 );
or ( n50183 , n50165 , n50169 , n50173 , n50177 , n50181 , n50182 );
and ( n50184 , n50161 , n50183 );
and ( n50185 , n26735 , n24800 );
or ( n50186 , n50184 , n50185 );
and ( n50187 , n50186 , n31008 );
and ( n50188 , n26735 , n10618 );
or ( n50189 , n50187 , n50188 );
buf ( n50190 , n50189 );
buf ( n50191 , n50190 );
not ( n50192 , n24800 );
and ( n50193 , n26257 , n25222 );
and ( n50194 , n44989 , n28583 );
and ( n50195 , n26257 , n28591 );
or ( n50196 , n50194 , n50195 );
and ( n50197 , n50196 , n28594 );
and ( n50198 , n44999 , n28583 );
and ( n50199 , n26257 , n28591 );
or ( n50200 , n50198 , n50199 );
and ( n50201 , n50200 , n30269 );
and ( n50202 , n45009 , n28583 );
and ( n50203 , n26257 , n28591 );
or ( n50204 , n50202 , n50203 );
and ( n50205 , n50204 , n30982 );
and ( n50206 , n29435 , n28583 );
and ( n50207 , n26257 , n28591 );
or ( n50208 , n50206 , n50207 );
and ( n50209 , n50208 , n30989 );
and ( n50210 , n26255 , n30991 );
and ( n50211 , n45019 , n28583 );
and ( n50212 , n26257 , n28591 );
or ( n50213 , n50211 , n50212 );
and ( n50214 , n50213 , n31002 );
or ( n50215 , n50193 , n50197 , n50201 , n50205 , n50209 , n50210 , n50214 );
and ( n50216 , n50192 , n50215 );
and ( n50217 , n26257 , n24800 );
or ( n50218 , n50216 , n50217 );
and ( n50219 , n50218 , n31008 );
and ( n50220 , n26257 , n10618 );
or ( n50221 , n50219 , n50220 );
buf ( n50222 , n50221 );
buf ( n50223 , n50222 );
not ( n50224 , n34804 );
and ( n50225 , n50224 , n26331 );
and ( n50226 , n14749 , n34804 );
or ( n50227 , n50225 , n50226 );
and ( n50228 , n50227 , n31008 );
and ( n50229 , n14749 , n10618 );
or ( n50230 , n50228 , n50229 );
buf ( n50231 , n50230 );
buf ( n50232 , n50231 );
buf ( n50233 , n10613 );
not ( n50234 , n34821 );
and ( n50235 , n46341 , n36345 );
and ( n50236 , n13461 , n36352 );
or ( n50237 , n50235 , n50236 );
and ( n50238 , n50237 , n14562 );
and ( n50239 , n46351 , n36345 );
and ( n50240 , n13461 , n37073 );
or ( n50241 , n50239 , n50240 );
and ( n50242 , n50241 , n14586 );
and ( n50243 , n46361 , n36350 );
and ( n50244 , n13461 , n37825 );
or ( n50245 , n50243 , n50244 );
and ( n50246 , n50245 , n14584 );
and ( n50247 , n46351 , n36350 );
and ( n50248 , n13461 , n37831 );
or ( n50249 , n50247 , n50248 );
and ( n50250 , n50249 , n37835 );
and ( n50251 , n46361 , n36350 );
and ( n50252 , n13461 , n37831 );
or ( n50253 , n50251 , n50252 );
and ( n50254 , n50253 , n37841 );
and ( n50255 , n15801 , n36350 );
and ( n50256 , n13461 , n37831 );
or ( n50257 , n50255 , n50256 );
and ( n50258 , n50257 , n37847 );
and ( n50259 , n13461 , n37849 );
or ( n50260 , n50238 , n50242 , n50246 , n50250 , n50254 , n50258 , n50259 );
and ( n50261 , n50234 , n50260 );
and ( n50262 , n13461 , n34821 );
or ( n50263 , n50261 , n50262 );
and ( n50264 , n50263 , n16574 );
and ( n50265 , n13461 , n16576 );
or ( n50266 , n50264 , n50265 );
buf ( n50267 , n50266 );
buf ( n50268 , n50267 );
not ( n50269 , n17451 );
and ( n50270 , n19281 , n17873 );
and ( n50271 , n47038 , n21336 );
and ( n50272 , n19281 , n42682 );
or ( n50273 , n50271 , n50272 );
and ( n50274 , n50273 , n21341 );
and ( n50275 , n47048 , n21336 );
and ( n50276 , n19281 , n42682 );
or ( n50277 , n50275 , n50276 );
and ( n50278 , n50277 , n23064 );
and ( n50279 , n47058 , n21336 );
and ( n50280 , n19281 , n42682 );
or ( n50281 , n50279 , n50280 );
and ( n50282 , n50281 , n23825 );
and ( n50283 , n21945 , n21336 );
and ( n50284 , n19281 , n42682 );
or ( n50285 , n50283 , n50284 );
and ( n50286 , n50285 , n23832 );
and ( n50287 , n21945 , n23834 );
and ( n50288 , n47068 , n21336 );
and ( n50289 , n19281 , n42682 );
or ( n50290 , n50288 , n50289 );
and ( n50291 , n50290 , n23917 );
or ( n50292 , n50270 , n50274 , n50278 , n50282 , n50286 , n50287 , n50291 );
and ( n50293 , n50269 , n50292 );
and ( n50294 , n19281 , n17451 );
or ( n50295 , n50293 , n50294 );
and ( n50296 , n50295 , n23924 );
and ( n50297 , n18215 , n23926 );
or ( n50298 , n50296 , n50297 );
buf ( n50299 , n50298 );
buf ( n50300 , n50299 );
not ( n50301 , n34821 );
and ( n50302 , n44175 , n36345 );
and ( n50303 , n13478 , n36352 );
or ( n50304 , n50302 , n50303 );
and ( n50305 , n50304 , n14562 );
and ( n50306 , n44185 , n36345 );
and ( n50307 , n13478 , n37073 );
or ( n50308 , n50306 , n50307 );
and ( n50309 , n50308 , n14586 );
and ( n50310 , n44195 , n36350 );
and ( n50311 , n13478 , n37825 );
or ( n50312 , n50310 , n50311 );
and ( n50313 , n50312 , n14584 );
and ( n50314 , n44185 , n36350 );
and ( n50315 , n13478 , n37831 );
or ( n50316 , n50314 , n50315 );
and ( n50317 , n50316 , n37835 );
and ( n50318 , n44195 , n36350 );
and ( n50319 , n13478 , n37831 );
or ( n50320 , n50318 , n50319 );
and ( n50321 , n50320 , n37841 );
and ( n50322 , n15823 , n36350 );
and ( n50323 , n13478 , n37831 );
or ( n50324 , n50322 , n50323 );
and ( n50325 , n50324 , n37847 );
and ( n50326 , n13478 , n37849 );
or ( n50327 , n50305 , n50309 , n50313 , n50317 , n50321 , n50325 , n50326 );
and ( n50328 , n50301 , n50327 );
and ( n50329 , n13478 , n34821 );
or ( n50330 , n50328 , n50329 );
and ( n50331 , n50330 , n16574 );
and ( n50332 , n13478 , n16576 );
or ( n50333 , n50331 , n50332 );
buf ( n50334 , n50333 );
buf ( n50335 , n50334 );
buf ( n50336 , n10615 );
buf ( n50337 , n10615 );
buf ( n50338 , n10613 );
buf ( n50339 , n10615 );
buf ( n50340 , n10615 );
buf ( n50341 , n10615 );
buf ( n50342 , n10613 );
buf ( n50343 , n10613 );
buf ( n50344 , n10615 );
buf ( n50345 , n10615 );
buf ( n50346 , n10615 );
buf ( n50347 , n10615 );
buf ( n50348 , n10613 );
buf ( n50349 , n10615 );
buf ( n50350 , n10615 );
not ( n50351 , n11954 );
not ( n50352 , n12243 );
and ( n50353 , n10869 , n31187 );
not ( n50354 , n31697 );
and ( n50355 , n50354 , n31540 );
xor ( n50356 , n31540 , n31371 );
xor ( n50357 , n31523 , n31371 );
xor ( n50358 , n31506 , n31371 );
xor ( n50359 , n31489 , n31371 );
xor ( n50360 , n31472 , n31371 );
xor ( n50361 , n31455 , n31371 );
xor ( n50362 , n31438 , n31371 );
xor ( n50363 , n31421 , n31371 );
xor ( n50364 , n31404 , n31371 );
xor ( n50365 , n31387 , n31371 );
and ( n50366 , n31700 , n31371 );
and ( n50367 , n50365 , n50366 );
and ( n50368 , n50364 , n50367 );
and ( n50369 , n50363 , n50368 );
and ( n50370 , n50362 , n50369 );
and ( n50371 , n50361 , n50370 );
and ( n50372 , n50360 , n50371 );
and ( n50373 , n50359 , n50372 );
and ( n50374 , n50358 , n50373 );
and ( n50375 , n50357 , n50374 );
xor ( n50376 , n50356 , n50375 );
and ( n50377 , n50376 , n31697 );
or ( n50378 , n50355 , n50377 );
buf ( n50379 , n50378 );
and ( n50380 , n50379 , n14140 );
not ( n50381 , n32214 );
and ( n50382 , n50381 , n32057 );
xor ( n50383 , n32057 , n31888 );
xor ( n50384 , n32040 , n31888 );
xor ( n50385 , n32023 , n31888 );
xor ( n50386 , n32006 , n31888 );
xor ( n50387 , n31989 , n31888 );
xor ( n50388 , n31972 , n31888 );
xor ( n50389 , n31955 , n31888 );
xor ( n50390 , n31938 , n31888 );
xor ( n50391 , n31921 , n31888 );
xor ( n50392 , n31904 , n31888 );
and ( n50393 , n32217 , n31888 );
and ( n50394 , n50392 , n50393 );
and ( n50395 , n50391 , n50394 );
and ( n50396 , n50390 , n50395 );
and ( n50397 , n50389 , n50396 );
and ( n50398 , n50388 , n50397 );
and ( n50399 , n50387 , n50398 );
and ( n50400 , n50386 , n50399 );
and ( n50401 , n50385 , n50400 );
and ( n50402 , n50384 , n50401 );
xor ( n50403 , n50383 , n50402 );
and ( n50404 , n50403 , n32214 );
or ( n50405 , n50382 , n50404 );
buf ( n50406 , n50405 );
and ( n50407 , n50406 , n14137 );
and ( n50408 , n15645 , n14143 );
and ( n50409 , n10869 , n14141 );
or ( n50410 , n50380 , n50407 , n50408 , n50409 );
and ( n50411 , n50410 , n32236 );
or ( n50412 , n50353 , n50411 );
and ( n50413 , n50352 , n50412 );
not ( n50414 , n34038 );
and ( n50415 , n50414 , n33818 );
xor ( n50416 , n33818 , n33579 );
xor ( n50417 , n33794 , n33579 );
xor ( n50418 , n33770 , n33579 );
xor ( n50419 , n33746 , n33579 );
xor ( n50420 , n33722 , n33579 );
xor ( n50421 , n33698 , n33579 );
xor ( n50422 , n33674 , n33579 );
xor ( n50423 , n33650 , n33579 );
xor ( n50424 , n33626 , n33579 );
xor ( n50425 , n33602 , n33579 );
and ( n50426 , n34041 , n33579 );
and ( n50427 , n50425 , n50426 );
and ( n50428 , n50424 , n50427 );
and ( n50429 , n50423 , n50428 );
and ( n50430 , n50422 , n50429 );
and ( n50431 , n50421 , n50430 );
and ( n50432 , n50420 , n50431 );
and ( n50433 , n50419 , n50432 );
and ( n50434 , n50418 , n50433 );
and ( n50435 , n50417 , n50434 );
xor ( n50436 , n50416 , n50435 );
and ( n50437 , n50436 , n34038 );
or ( n50438 , n50415 , n50437 );
buf ( n50439 , n50438 );
and ( n50440 , n50439 , n12243 );
or ( n50441 , n50413 , n50440 );
and ( n50442 , n50351 , n50441 );
and ( n50443 , n50410 , n11954 );
or ( n50444 , n50442 , n50443 );
and ( n50445 , n50444 , n16574 );
not ( n50446 , n34327 );
and ( n50447 , n50446 , n34197 );
xor ( n50448 , n34197 , n34058 );
xor ( n50449 , n34183 , n34058 );
xor ( n50450 , n34169 , n34058 );
xor ( n50451 , n34155 , n34058 );
xor ( n50452 , n34141 , n34058 );
xor ( n50453 , n34127 , n34058 );
xor ( n50454 , n34113 , n34058 );
xor ( n50455 , n34099 , n34058 );
xor ( n50456 , n34085 , n34058 );
xor ( n50457 , n34071 , n34058 );
and ( n50458 , n34330 , n34058 );
and ( n50459 , n50457 , n50458 );
and ( n50460 , n50456 , n50459 );
and ( n50461 , n50455 , n50460 );
and ( n50462 , n50454 , n50461 );
and ( n50463 , n50453 , n50462 );
and ( n50464 , n50452 , n50463 );
and ( n50465 , n50451 , n50464 );
and ( n50466 , n50450 , n50465 );
and ( n50467 , n50449 , n50466 );
xor ( n50468 , n50448 , n50467 );
and ( n50469 , n50468 , n34327 );
or ( n50470 , n50447 , n50469 );
buf ( n50471 , n50470 );
and ( n50472 , n50471 , n16576 );
or ( n50473 , n50445 , n50472 );
buf ( n50474 , n50473 );
buf ( n50475 , n50474 );
and ( n50476 , n11601 , n16574 );
and ( n50477 , n15594 , n16576 );
or ( n50478 , n50476 , n50477 );
buf ( n50479 , n50478 );
buf ( n50480 , n50479 );
not ( n50481 , n11333 );
and ( n50482 , n50481 , n11295 );
xor ( n50483 , n11295 , n11007 );
and ( n50484 , n46275 , n46276 );
xor ( n50485 , n50483 , n50484 );
and ( n50486 , n50485 , n11333 );
or ( n50487 , n50482 , n50486 );
buf ( n50488 , n50487 );
buf ( n50489 , n50488 );
not ( n50490 , n17451 );
and ( n50491 , n20490 , n17873 );
and ( n50492 , n48746 , n21330 );
and ( n50493 , n20490 , n21338 );
or ( n50494 , n50492 , n50493 );
and ( n50495 , n50494 , n21341 );
and ( n50496 , n48756 , n21330 );
and ( n50497 , n20490 , n21338 );
or ( n50498 , n50496 , n50497 );
and ( n50499 , n50498 , n23064 );
and ( n50500 , n48766 , n21330 );
and ( n50501 , n20490 , n21338 );
or ( n50502 , n50500 , n50501 );
and ( n50503 , n50502 , n23825 );
and ( n50504 , n21867 , n21330 );
and ( n50505 , n20490 , n21338 );
or ( n50506 , n50504 , n50505 );
and ( n50507 , n50506 , n23832 );
and ( n50508 , n20488 , n23834 );
and ( n50509 , n48776 , n21330 );
and ( n50510 , n20490 , n21338 );
or ( n50511 , n50509 , n50510 );
and ( n50512 , n50511 , n23917 );
or ( n50513 , n50491 , n50495 , n50499 , n50503 , n50507 , n50508 , n50512 );
and ( n50514 , n50490 , n50513 );
and ( n50515 , n20490 , n17451 );
or ( n50516 , n50514 , n50515 );
and ( n50517 , n50516 , n23924 );
and ( n50518 , n20490 , n23926 );
or ( n50519 , n50517 , n50518 );
buf ( n50520 , n50519 );
buf ( n50521 , n50520 );
not ( n50522 , n34821 );
and ( n50523 , n13265 , n14592 );
and ( n50524 , n45165 , n36348 );
and ( n50525 , n13265 , n43530 );
or ( n50526 , n50524 , n50525 );
and ( n50527 , n50526 , n14562 );
and ( n50528 , n45181 , n36347 );
and ( n50529 , n13265 , n43543 );
or ( n50530 , n50528 , n50529 );
and ( n50531 , n50530 , n14586 );
and ( n50532 , n45197 , n36348 );
and ( n50533 , n13265 , n43556 );
or ( n50534 , n50532 , n50533 );
and ( n50535 , n50534 , n14584 );
and ( n50536 , n45181 , n36347 );
and ( n50537 , n13265 , n43563 );
or ( n50538 , n50536 , n50537 );
and ( n50539 , n50538 , n37835 );
and ( n50540 , n45197 , n36347 );
and ( n50541 , n13265 , n43563 );
or ( n50542 , n50540 , n50541 );
and ( n50543 , n50542 , n37841 );
and ( n50544 , n13263 , n14564 );
and ( n50545 , n15449 , n36347 );
and ( n50546 , n13265 , n43563 );
or ( n50547 , n50545 , n50546 );
and ( n50548 , n50547 , n37847 );
or ( n50549 , n50523 , n50527 , n50531 , n50535 , n50539 , n50543 , n50544 , n50548 );
and ( n50550 , n50522 , n50549 );
and ( n50551 , n13265 , n34821 );
or ( n50552 , n50550 , n50551 );
and ( n50553 , n50552 , n16574 );
and ( n50554 , n13265 , n16576 );
or ( n50555 , n50553 , n50554 );
buf ( n50556 , n50555 );
buf ( n50557 , n50556 );
buf ( n50558 , n10613 );
buf ( n50559 , n10615 );
buf ( n50560 , n10615 );
buf ( n50561 , n10615 );
buf ( n50562 , n10615 );
buf ( n50563 , n10613 );
buf ( n50564 , n10615 );
buf ( n50565 , n10615 );
not ( n50566 , n24800 );
and ( n50567 , n39803 , n28586 );
and ( n50568 , n26021 , n34573 );
or ( n50569 , n50567 , n50568 );
and ( n50570 , n50569 , n28594 );
and ( n50571 , n39816 , n28586 );
and ( n50572 , n26021 , n34573 );
or ( n50573 , n50571 , n50572 );
and ( n50574 , n50573 , n30269 );
and ( n50575 , n39826 , n28586 );
and ( n50576 , n26021 , n34573 );
or ( n50577 , n50575 , n50576 );
and ( n50578 , n50577 , n30982 );
and ( n50579 , n29575 , n28586 );
and ( n50580 , n26021 , n34573 );
or ( n50581 , n50579 , n50580 );
and ( n50582 , n50581 , n30989 );
and ( n50583 , n39836 , n28586 );
and ( n50584 , n26021 , n34573 );
or ( n50585 , n50583 , n50584 );
and ( n50586 , n50585 , n31002 );
and ( n50587 , n26021 , n34607 );
or ( n50588 , n50570 , n50574 , n50578 , n50582 , n50586 , n50587 );
and ( n50589 , n50566 , n50588 );
and ( n50590 , n26021 , n24800 );
or ( n50591 , n50589 , n50590 );
and ( n50592 , n50591 , n31008 );
and ( n50593 , n26021 , n10618 );
or ( n50594 , n50592 , n50593 );
buf ( n50595 , n50594 );
buf ( n50596 , n50595 );
not ( n50597 , n34538 );
and ( n50598 , n50597 , n20484 );
and ( n50599 , n14651 , n34538 );
or ( n50600 , n50598 , n50599 );
and ( n50601 , n50600 , n23924 );
and ( n50602 , n14651 , n23926 );
or ( n50603 , n50601 , n50602 );
buf ( n50604 , n50603 );
buf ( n50605 , n50604 );
buf ( n50606 , n10615 );
buf ( n50607 , n10613 );
and ( n50608 , n11633 , n16574 );
and ( n50609 , n15682 , n16576 );
or ( n50610 , n50608 , n50609 );
buf ( n50611 , n50610 );
buf ( n50612 , n50611 );
buf ( n50613 , n10615 );
and ( n50614 , n16992 , n23924 );
and ( n50615 , n21878 , n23926 );
or ( n50616 , n50614 , n50615 );
buf ( n50617 , n50616 );
buf ( n50618 , n50617 );
not ( n50619 , n24800 );
and ( n50620 , n26121 , n25222 );
and ( n50621 , n49846 , n28583 );
and ( n50622 , n26121 , n28591 );
or ( n50623 , n50621 , n50622 );
and ( n50624 , n50623 , n28594 );
and ( n50625 , n49856 , n28583 );
and ( n50626 , n26121 , n28591 );
or ( n50627 , n50625 , n50626 );
and ( n50628 , n50627 , n30269 );
and ( n50629 , n49866 , n28583 );
and ( n50630 , n26121 , n28591 );
or ( n50631 , n50629 , n50630 );
and ( n50632 , n50631 , n30982 );
and ( n50633 , n29515 , n28583 );
and ( n50634 , n26121 , n28591 );
or ( n50635 , n50633 , n50634 );
and ( n50636 , n50635 , n30989 );
and ( n50637 , n26119 , n30991 );
and ( n50638 , n49876 , n28583 );
and ( n50639 , n26121 , n28591 );
or ( n50640 , n50638 , n50639 );
and ( n50641 , n50640 , n31002 );
or ( n50642 , n50620 , n50624 , n50628 , n50632 , n50636 , n50637 , n50641 );
and ( n50643 , n50619 , n50642 );
and ( n50644 , n26121 , n24800 );
or ( n50645 , n50643 , n50644 );
and ( n50646 , n50645 , n31008 );
and ( n50647 , n26121 , n10618 );
or ( n50648 , n50646 , n50647 );
buf ( n50649 , n50648 );
buf ( n50650 , n50649 );
buf ( n50651 , n10615 );
buf ( n50652 , n10613 );
not ( n50653 , n17451 );
and ( n50654 , n48886 , n21334 );
and ( n50655 , n18675 , n34492 );
or ( n50656 , n50654 , n50655 );
and ( n50657 , n50656 , n21341 );
and ( n50658 , n48896 , n21334 );
and ( n50659 , n18675 , n34492 );
or ( n50660 , n50658 , n50659 );
and ( n50661 , n50660 , n23064 );
and ( n50662 , n48906 , n21334 );
and ( n50663 , n18675 , n34492 );
or ( n50664 , n50662 , n50663 );
and ( n50665 , n50664 , n23825 );
and ( n50666 , n22322 , n21334 );
and ( n50667 , n18675 , n34492 );
or ( n50668 , n50666 , n50667 );
and ( n50669 , n50668 , n23832 );
and ( n50670 , n48916 , n21334 );
and ( n50671 , n18675 , n34492 );
or ( n50672 , n50670 , n50671 );
and ( n50673 , n50672 , n23917 );
and ( n50674 , n18675 , n34526 );
or ( n50675 , n50657 , n50661 , n50665 , n50669 , n50673 , n50674 );
and ( n50676 , n50653 , n50675 );
and ( n50677 , n18675 , n17451 );
or ( n50678 , n50676 , n50677 );
and ( n50679 , n50678 , n23924 );
and ( n50680 , n18675 , n23926 );
or ( n50681 , n50679 , n50680 );
buf ( n50682 , n50681 );
buf ( n50683 , n50682 );
buf ( n50684 , n10613 );
not ( n50685 , n34538 );
and ( n50686 , n50685 , n18677 );
and ( n50687 , n14801 , n34538 );
or ( n50688 , n50686 , n50687 );
and ( n50689 , n50688 , n23924 );
and ( n50690 , n14801 , n23926 );
or ( n50691 , n50689 , n50690 );
buf ( n50692 , n50691 );
buf ( n50693 , n50692 );
not ( n50694 , n17451 );
and ( n50695 , n18571 , n17873 );
not ( n50696 , n19474 );
and ( n50697 , n50696 , n18558 );
xor ( n50698 , n19500 , n19502 );
and ( n50699 , n50698 , n19474 );
or ( n50700 , n50697 , n50699 );
buf ( n50701 , n50700 );
and ( n50702 , n50701 , n19745 );
and ( n50703 , n50701 , n19748 );
not ( n50704 , n19750 );
and ( n50705 , n50704 , n20613 );
not ( n50706 , n21193 );
and ( n50707 , n50706 , n20625 );
xor ( n50708 , n21219 , n21223 );
and ( n50709 , n50708 , n21193 );
or ( n50710 , n50707 , n50709 );
buf ( n50711 , n50710 );
and ( n50712 , n50711 , n19750 );
or ( n50713 , n50705 , n50712 );
and ( n50714 , n50713 , n21253 );
and ( n50715 , n20613 , n21255 );
or ( n50716 , n50702 , n50703 , n50714 , n50715 );
and ( n50717 , n50716 , n21330 );
and ( n50718 , n18571 , n21338 );
or ( n50719 , n50717 , n50718 );
and ( n50720 , n50719 , n21341 );
not ( n50721 , n22996 );
and ( n50722 , n50721 , n22533 );
xor ( n50723 , n23022 , n23026 );
and ( n50724 , n50723 , n22996 );
or ( n50725 , n50722 , n50724 );
buf ( n50726 , n50725 );
and ( n50727 , n50726 , n21330 );
and ( n50728 , n18571 , n21338 );
or ( n50729 , n50727 , n50728 );
and ( n50730 , n50729 , n23064 );
not ( n50731 , n23758 );
and ( n50732 , n50731 , n23295 );
xor ( n50733 , n23784 , n23788 );
and ( n50734 , n50733 , n23758 );
or ( n50735 , n50732 , n50734 );
buf ( n50736 , n50735 );
and ( n50737 , n50736 , n21330 );
and ( n50738 , n18571 , n21338 );
or ( n50739 , n50737 , n50738 );
and ( n50740 , n50739 , n23825 );
and ( n50741 , n22382 , n21330 );
and ( n50742 , n18571 , n21338 );
or ( n50743 , n50741 , n50742 );
and ( n50744 , n50743 , n23832 );
and ( n50745 , n18569 , n23834 );
xor ( n50746 , n23883 , n23888 );
buf ( n50747 , n50746 );
and ( n50748 , n50747 , n21330 );
and ( n50749 , n18571 , n21338 );
or ( n50750 , n50748 , n50749 );
and ( n50751 , n50750 , n23917 );
or ( n50752 , n50695 , n50720 , n50730 , n50740 , n50744 , n50745 , n50751 );
and ( n50753 , n50694 , n50752 );
and ( n50754 , n18571 , n17451 );
or ( n50755 , n50753 , n50754 );
and ( n50756 , n50755 , n23924 );
and ( n50757 , n18571 , n23926 );
or ( n50758 , n50756 , n50757 );
buf ( n50759 , n50758 );
buf ( n50760 , n50759 );
not ( n50761 , n11333 );
and ( n50762 , n50761 , n11193 );
xor ( n50763 , n11340 , n11362 );
and ( n50764 , n50763 , n11333 );
or ( n50765 , n50762 , n50764 );
buf ( n50766 , n50765 );
buf ( n50767 , n50766 );
buf ( n50768 , n10615 );
not ( n50769 , n24800 );
and ( n50770 , n50769 , n28581 );
and ( n50771 , n28557 , n24800 );
or ( n50772 , n50770 , n50771 );
and ( n50773 , n50772 , n31008 );
and ( n50774 , n28557 , n10618 );
or ( n50775 , n50773 , n50774 );
buf ( n50776 , n50775 );
buf ( n50777 , n50776 );
buf ( n50778 , n10613 );
not ( n50779 , n24511 );
not ( n50780 , n24799 );
and ( n50781 , n10680 , n40154 );
not ( n50782 , n40632 );
and ( n50783 , n50782 , n40492 );
xor ( n50784 , n40639 , n40661 );
and ( n50785 , n50784 , n40632 );
or ( n50786 , n50783 , n50785 );
buf ( n50787 , n50786 );
and ( n50788 , n50787 , n27046 );
not ( n50789 , n41147 );
and ( n50790 , n50789 , n41007 );
xor ( n50791 , n41154 , n41176 );
and ( n50792 , n50791 , n41147 );
or ( n50793 , n50790 , n50792 );
buf ( n50794 , n50793 );
and ( n50795 , n50794 , n27049 );
and ( n50796 , n29453 , n28506 );
and ( n50797 , n10680 , n28508 );
or ( n50798 , n50788 , n50795 , n50796 , n50797 );
and ( n50799 , n50798 , n41199 );
or ( n50800 , n50781 , n50799 );
and ( n50801 , n50780 , n50800 );
xor ( n50802 , n41580 , n41588 );
xor ( n50803 , n50802 , n41794 );
buf ( n50804 , n50803 );
and ( n50805 , n50804 , n27046 );
xor ( n50806 , n42159 , n42160 );
xor ( n50807 , n50806 , n42290 );
buf ( n50808 , n50807 );
and ( n50809 , n50808 , n27049 );
and ( n50810 , n29453 , n42306 );
or ( n50811 , n50805 , n50809 , n50810 );
buf ( n50812 , n50811 );
and ( n50813 , C1 , n50812 );
or ( n50814 , n50813 , C0 );
buf ( n50815 , n50814 );
not ( n50816 , n50815 );
buf ( n50817 , n50816 );
buf ( n50818 , n50817 );
not ( n50819 , n50818 );
and ( n50820 , C1 , n50819 );
or ( n50821 , n50820 , C0 );
buf ( n50822 , n50821 );
and ( n50823 , n50822 , n24799 );
or ( n50824 , n50801 , n50823 );
and ( n50825 , n50779 , n50824 );
and ( n50826 , n50798 , n24511 );
or ( n50827 , n50825 , n50826 );
and ( n50828 , n50827 , n31008 );
not ( n50829 , n42601 );
and ( n50830 , n50829 , n42485 );
xor ( n50831 , n42608 , n42630 );
and ( n50832 , n50831 , n42601 );
or ( n50833 , n50830 , n50832 );
buf ( n50834 , n50833 );
and ( n50835 , n50834 , n10618 );
or ( n50836 , n50828 , n50835 );
buf ( n50837 , n50836 );
buf ( n50838 , n50837 );
buf ( n50839 , n10615 );
not ( n50840 , n17451 );
and ( n50841 , n46607 , n21334 );
and ( n50842 , n18777 , n34492 );
or ( n50843 , n50841 , n50842 );
and ( n50844 , n50843 , n21341 );
and ( n50845 , n46617 , n21334 );
and ( n50846 , n18777 , n34492 );
or ( n50847 , n50845 , n50846 );
and ( n50848 , n50847 , n23064 );
and ( n50849 , n46627 , n21334 );
and ( n50850 , n18777 , n34492 );
or ( n50851 , n50849 , n50850 );
and ( n50852 , n50851 , n23825 );
and ( n50853 , n22262 , n21334 );
and ( n50854 , n18777 , n34492 );
or ( n50855 , n50853 , n50854 );
and ( n50856 , n50855 , n23832 );
and ( n50857 , n46638 , n21334 );
and ( n50858 , n18777 , n34492 );
or ( n50859 , n50857 , n50858 );
and ( n50860 , n50859 , n23917 );
and ( n50861 , n18777 , n34526 );
or ( n50862 , n50844 , n50848 , n50852 , n50856 , n50860 , n50861 );
and ( n50863 , n50840 , n50862 );
and ( n50864 , n18777 , n17451 );
or ( n50865 , n50863 , n50864 );
and ( n50866 , n50865 , n23924 );
and ( n50867 , n18777 , n23926 );
or ( n50868 , n50866 , n50867 );
buf ( n50869 , n50868 );
buf ( n50870 , n50869 );
buf ( n50871 , n16576 );
buf ( n50872 , n50871 );
buf ( n50873 , n10613 );
not ( n50874 , n24800 );
and ( n50875 , n39662 , n28587 );
and ( n50876 , n26431 , n39807 );
or ( n50877 , n50875 , n50876 );
and ( n50878 , n50877 , n28594 );
and ( n50879 , n39678 , n28587 );
and ( n50880 , n26431 , n39807 );
or ( n50881 , n50879 , n50880 );
and ( n50882 , n50881 , n30269 );
and ( n50883 , n39694 , n28587 );
and ( n50884 , n26431 , n39807 );
or ( n50885 , n50883 , n50884 );
and ( n50886 , n50885 , n30982 );
and ( n50887 , n29335 , n28587 );
and ( n50888 , n26431 , n39807 );
or ( n50889 , n50887 , n50888 );
and ( n50890 , n50889 , n30989 );
and ( n50891 , n39713 , n28587 );
and ( n50892 , n26431 , n39807 );
or ( n50893 , n50891 , n50892 );
and ( n50894 , n50893 , n31002 );
and ( n50895 , n26431 , n34607 );
or ( n50896 , n50878 , n50882 , n50886 , n50890 , n50894 , n50895 );
and ( n50897 , n50874 , n50896 );
and ( n50898 , n26431 , n24800 );
or ( n50899 , n50897 , n50898 );
and ( n50900 , n50899 , n31008 );
and ( n50901 , n26431 , n10618 );
or ( n50902 , n50900 , n50901 );
buf ( n50903 , n50902 );
buf ( n50904 , n50903 );
and ( n50905 , n11657 , n16574 );
and ( n50906 , n15748 , n16576 );
or ( n50907 , n50905 , n50906 );
buf ( n50908 , n50907 );
buf ( n50909 , n50908 );
not ( n50910 , n34538 );
and ( n50911 , n50910 , n19187 );
and ( n50912 , n14711 , n34538 );
or ( n50913 , n50911 , n50912 );
and ( n50914 , n50913 , n23924 );
and ( n50915 , n14711 , n23926 );
or ( n50916 , n50914 , n50915 );
buf ( n50917 , n50916 );
buf ( n50918 , n50917 );
buf ( n50919 , n10613 );
buf ( n50920 , n10615 );
buf ( n50921 , n10613 );
not ( n50922 , n17451 );
and ( n50923 , n19079 , n17873 );
and ( n50924 , n39326 , n21330 );
and ( n50925 , n19079 , n21338 );
or ( n50926 , n50924 , n50925 );
and ( n50927 , n50926 , n21341 );
and ( n50928 , n39336 , n21330 );
and ( n50929 , n19079 , n21338 );
or ( n50930 , n50928 , n50929 );
and ( n50931 , n50930 , n23064 );
and ( n50932 , n39346 , n21330 );
and ( n50933 , n19079 , n21338 );
or ( n50934 , n50932 , n50933 );
and ( n50935 , n50934 , n23825 );
and ( n50936 , n22082 , n21330 );
and ( n50937 , n19079 , n21338 );
or ( n50938 , n50936 , n50937 );
and ( n50939 , n50938 , n23832 );
and ( n50940 , n19077 , n23834 );
and ( n50941 , n39356 , n21330 );
and ( n50942 , n19079 , n21338 );
or ( n50943 , n50941 , n50942 );
and ( n50944 , n50943 , n23917 );
or ( n50945 , n50923 , n50927 , n50931 , n50935 , n50939 , n50940 , n50944 );
and ( n50946 , n50922 , n50945 );
and ( n50947 , n19079 , n17451 );
or ( n50948 , n50946 , n50947 );
and ( n50949 , n50948 , n23924 );
and ( n50950 , n19079 , n23926 );
or ( n50951 , n50949 , n50950 );
buf ( n50952 , n50951 );
buf ( n50953 , n50952 );
buf ( n50954 , n10615 );
not ( n50955 , n34538 );
and ( n50956 , n50955 , n18915 );
and ( n50957 , n14759 , n34538 );
or ( n50958 , n50956 , n50957 );
and ( n50959 , n50958 , n23924 );
and ( n50960 , n14759 , n23926 );
or ( n50961 , n50959 , n50960 );
buf ( n50962 , n50961 );
buf ( n50963 , n50962 );
buf ( n50964 , n10613 );
buf ( n50965 , n10615 );
buf ( n50966 , n10615 );
and ( n50967 , n16720 , n23924 );
and ( n50968 , n21943 , n23926 );
or ( n50969 , n50967 , n50968 );
buf ( n50970 , n50969 );
buf ( n50971 , n50970 );
buf ( n50972 , n10613 );
buf ( n50973 , n10613 );
buf ( n50974 , n10615 );
not ( n50975 , n34821 );
and ( n50976 , n13263 , n14592 );
and ( n50977 , n45165 , n36350 );
and ( n50978 , n13263 , n43691 );
or ( n50979 , n50977 , n50978 );
and ( n50980 , n50979 , n14562 );
and ( n50981 , n45181 , n36350 );
and ( n50982 , n13263 , n43703 );
or ( n50983 , n50981 , n50982 );
and ( n50984 , n50983 , n14586 );
and ( n50985 , n45197 , n36345 );
and ( n50986 , n13263 , n43715 );
or ( n50987 , n50985 , n50986 );
and ( n50988 , n50987 , n14584 );
and ( n50989 , n45181 , n36345 );
and ( n50990 , n13263 , n43721 );
or ( n50991 , n50989 , n50990 );
and ( n50992 , n50991 , n37835 );
and ( n50993 , n45197 , n36345 );
and ( n50994 , n13263 , n43721 );
or ( n50995 , n50993 , n50994 );
and ( n50996 , n50995 , n37841 );
and ( n50997 , n15449 , n14564 );
and ( n50998 , n15449 , n36345 );
and ( n50999 , n13263 , n43721 );
or ( n51000 , n50998 , n50999 );
and ( n51001 , n51000 , n37847 );
or ( n51002 , n50976 , n50980 , n50984 , n50988 , n50992 , n50996 , n50997 , n51001 );
and ( n51003 , n50975 , n51002 );
and ( n51004 , n13263 , n34821 );
or ( n51005 , n51003 , n51004 );
and ( n51006 , n51005 , n16574 );
and ( n51007 , n12276 , n16576 );
or ( n51008 , n51006 , n51007 );
buf ( n51009 , n51008 );
buf ( n51010 , n51009 );
buf ( n51011 , n10615 );
buf ( n51012 , n10613 );
buf ( n51013 , n10613 );
buf ( n51014 , n10615 );
not ( n51015 , n34538 );
and ( n51016 , n51015 , n18813 );
and ( n51017 , n14777 , n34538 );
or ( n51018 , n51016 , n51017 );
and ( n51019 , n51018 , n23924 );
and ( n51020 , n14777 , n23926 );
or ( n51021 , n51019 , n51020 );
buf ( n51022 , n51021 );
buf ( n51023 , n51022 );
buf ( n51024 , n10615 );
buf ( n51025 , n10613 );
buf ( n51026 , n10615 );
buf ( n51027 , n10613 );
buf ( n51028 , n10615 );
not ( n51029 , n34821 );
and ( n51030 , n13191 , n14592 );
and ( n51031 , n49200 , n36350 );
and ( n51032 , n13191 , n43691 );
or ( n51033 , n51031 , n51032 );
and ( n51034 , n51033 , n14562 );
and ( n51035 , n49210 , n36350 );
and ( n51036 , n13191 , n43703 );
or ( n51037 , n51035 , n51036 );
and ( n51038 , n51037 , n14586 );
and ( n51039 , n49220 , n36345 );
and ( n51040 , n13191 , n43715 );
or ( n51041 , n51039 , n51040 );
and ( n51042 , n51041 , n14584 );
and ( n51043 , n49210 , n36345 );
and ( n51044 , n13191 , n43721 );
or ( n51045 , n51043 , n51044 );
and ( n51046 , n51045 , n37835 );
and ( n51047 , n49220 , n36345 );
and ( n51048 , n13191 , n43721 );
or ( n51049 , n51047 , n51048 );
and ( n51050 , n51049 , n37841 );
and ( n51051 , n15037 , n14564 );
and ( n51052 , n15037 , n36345 );
and ( n51053 , n13191 , n43721 );
or ( n51054 , n51052 , n51053 );
and ( n51055 , n51054 , n37847 );
or ( n51056 , n51030 , n51034 , n51038 , n51042 , n51046 , n51050 , n51051 , n51055 );
and ( n51057 , n51029 , n51056 );
and ( n51058 , n13191 , n34821 );
or ( n51059 , n51057 , n51058 );
and ( n51060 , n51059 , n16574 );
and ( n51061 , n12258 , n16576 );
or ( n51062 , n51060 , n51061 );
buf ( n51063 , n51062 );
buf ( n51064 , n51063 );
not ( n51065 , n24800 );
and ( n51066 , n45549 , n28587 );
and ( n51067 , n25989 , n39807 );
or ( n51068 , n51066 , n51067 );
and ( n51069 , n51068 , n28594 );
and ( n51070 , n45559 , n28587 );
and ( n51071 , n25989 , n39807 );
or ( n51072 , n51070 , n51071 );
and ( n51073 , n51072 , n30269 );
and ( n51074 , n45569 , n28587 );
and ( n51075 , n25989 , n39807 );
or ( n51076 , n51074 , n51075 );
and ( n51077 , n51076 , n30982 );
and ( n51078 , n29595 , n28587 );
and ( n51079 , n25989 , n39807 );
or ( n51080 , n51078 , n51079 );
and ( n51081 , n51080 , n30989 );
and ( n51082 , n45580 , n28587 );
and ( n51083 , n25989 , n39807 );
or ( n51084 , n51082 , n51083 );
and ( n51085 , n51084 , n31002 );
and ( n51086 , n25989 , n34607 );
or ( n51087 , n51069 , n51073 , n51077 , n51081 , n51085 , n51086 );
and ( n51088 , n51065 , n51087 );
and ( n51089 , n25989 , n24800 );
or ( n51090 , n51088 , n51089 );
and ( n51091 , n51090 , n31008 );
and ( n51092 , n25989 , n10618 );
or ( n51093 , n51091 , n51092 );
buf ( n51094 , n51093 );
buf ( n51095 , n51094 );
and ( n51096 , n11577 , n16574 );
and ( n51097 , n15528 , n16576 );
or ( n51098 , n51096 , n51097 );
buf ( n51099 , n51098 );
buf ( n51100 , n51099 );
and ( n51101 , n24190 , n31008 );
and ( n51102 , n29506 , n10618 );
or ( n51103 , n51101 , n51102 );
buf ( n51104 , n51103 );
buf ( n51105 , n51104 );
buf ( n51106 , n10615 );
buf ( n51107 , n10613 );
buf ( n51108 , n10615 );
buf ( n51109 , n10613 );
buf ( n51110 , n10615 );
not ( n51111 , n34804 );
and ( n51112 , n51111 , n25876 );
and ( n51113 , n14647 , n34804 );
or ( n51114 , n51112 , n51113 );
and ( n51115 , n51114 , n31008 );
and ( n51116 , n14647 , n10618 );
or ( n51117 , n51115 , n51116 );
buf ( n51118 , n51117 );
buf ( n51119 , n51118 );
buf ( n51120 , n10615 );
buf ( n51121 , n10613 );
buf ( n51122 , n10613 );
buf ( n51123 , n10615 );
buf ( n51124 , n10613 );
buf ( n51125 , n10613 );
not ( n51126 , n34538 );
and ( n51127 , n51126 , n19323 );
and ( n51128 , n14687 , n34538 );
or ( n51129 , n51127 , n51128 );
and ( n51130 , n51129 , n23924 );
and ( n51131 , n14687 , n23926 );
or ( n51132 , n51130 , n51131 );
buf ( n51133 , n51132 );
buf ( n51134 , n51133 );
not ( n51135 , n34821 );
not ( n51136 , n13916 );
and ( n51137 , n51136 , n13683 );
xor ( n51138 , n13684 , n13871 );
and ( n51139 , n51138 , n13916 );
or ( n51140 , n51137 , n51139 );
buf ( n51141 , n51140 );
and ( n51142 , n51141 , n14137 );
and ( n51143 , n51141 , n14143 );
not ( n51144 , n14139 );
and ( n51145 , n51144 , n35987 );
not ( n51146 , n36245 );
and ( n51147 , n51146 , n35999 );
xor ( n51148 , n45153 , n45154 );
and ( n51149 , n51148 , n36245 );
or ( n51150 , n51147 , n51149 );
buf ( n51151 , n51150 );
and ( n51152 , n51151 , n14139 );
or ( n51153 , n51145 , n51152 );
and ( n51154 , n51153 , n14140 );
and ( n51155 , n35987 , n14141 );
or ( n51156 , n51142 , n51143 , n51154 , n51155 );
and ( n51157 , n51156 , n36345 );
and ( n51158 , n13293 , n36352 );
or ( n51159 , n51157 , n51158 );
and ( n51160 , n51159 , n14562 );
not ( n51161 , n37048 );
and ( n51162 , n51161 , n36840 );
xor ( n51163 , n45174 , n45175 );
and ( n51164 , n51163 , n37048 );
or ( n51165 , n51162 , n51164 );
buf ( n51166 , n51165 );
and ( n51167 , n51166 , n36345 );
and ( n51168 , n13293 , n37073 );
or ( n51169 , n51167 , n51168 );
and ( n51170 , n51169 , n14586 );
not ( n51171 , n37801 );
and ( n51172 , n51171 , n37593 );
xor ( n51173 , n45190 , n45191 );
and ( n51174 , n51173 , n37801 );
or ( n51175 , n51172 , n51174 );
buf ( n51176 , n51175 );
and ( n51177 , n51176 , n36350 );
and ( n51178 , n13293 , n37825 );
or ( n51179 , n51177 , n51178 );
and ( n51180 , n51179 , n14584 );
and ( n51181 , n51166 , n36350 );
and ( n51182 , n13293 , n37831 );
or ( n51183 , n51181 , n51182 );
and ( n51184 , n51183 , n37835 );
and ( n51185 , n51176 , n36350 );
and ( n51186 , n13293 , n37831 );
or ( n51187 , n51185 , n51186 );
and ( n51188 , n51187 , n37841 );
and ( n51189 , n15493 , n36350 );
and ( n51190 , n13293 , n37831 );
or ( n51191 , n51189 , n51190 );
and ( n51192 , n51191 , n37847 );
and ( n51193 , n13293 , n37849 );
or ( n51194 , n51160 , n51170 , n51180 , n51184 , n51188 , n51192 , n51193 );
and ( n51195 , n51135 , n51194 );
and ( n51196 , n13293 , n34821 );
or ( n51197 , n51195 , n51196 );
and ( n51198 , n51197 , n16574 );
and ( n51199 , n13293 , n16576 );
or ( n51200 , n51198 , n51199 );
buf ( n51201 , n51200 );
buf ( n51202 , n51201 );
buf ( n51203 , n10613 );
buf ( n51204 , n10615 );
buf ( n51205 , n10613 );
not ( n51206 , n17451 );
and ( n51207 , n50716 , n21333 );
and ( n51208 , n18573 , n34758 );
or ( n51209 , n51207 , n51208 );
and ( n51210 , n51209 , n21341 );
and ( n51211 , n50726 , n21333 );
and ( n51212 , n18573 , n34758 );
or ( n51213 , n51211 , n51212 );
and ( n51214 , n51213 , n23064 );
and ( n51215 , n50736 , n21333 );
and ( n51216 , n18573 , n34758 );
or ( n51217 , n51215 , n51216 );
and ( n51218 , n51217 , n23825 );
and ( n51219 , n22382 , n21333 );
and ( n51220 , n18573 , n34758 );
or ( n51221 , n51219 , n51220 );
and ( n51222 , n51221 , n23832 );
and ( n51223 , n50747 , n21333 );
and ( n51224 , n18573 , n34758 );
or ( n51225 , n51223 , n51224 );
and ( n51226 , n51225 , n23917 );
and ( n51227 , n18573 , n34526 );
or ( n51228 , n51210 , n51214 , n51218 , n51222 , n51226 , n51227 );
and ( n51229 , n51206 , n51228 );
and ( n51230 , n18573 , n17451 );
or ( n51231 , n51229 , n51230 );
and ( n51232 , n51231 , n23924 );
and ( n51233 , n18573 , n23926 );
or ( n51234 , n51232 , n51233 );
buf ( n51235 , n51234 );
buf ( n51236 , n51235 );
buf ( n51237 , n10613 );
buf ( n51238 , n10613 );
not ( n51239 , n24511 );
not ( n51240 , n24799 );
and ( n51241 , n10655 , n40154 );
not ( n51242 , n40632 );
and ( n51243 , n51242 , n40577 );
xor ( n51244 , n43754 , n43755 );
and ( n51245 , n51244 , n40632 );
or ( n51246 , n51243 , n51245 );
buf ( n51247 , n51246 );
and ( n51248 , n51247 , n27046 );
not ( n51249 , n41147 );
and ( n51250 , n51249 , n41092 );
xor ( n51251 , n43769 , n43770 );
and ( n51252 , n51251 , n41147 );
or ( n51253 , n51250 , n51252 );
buf ( n51254 , n51253 );
and ( n51255 , n51254 , n27049 );
and ( n51256 , n29353 , n28506 );
and ( n51257 , n10655 , n28508 );
or ( n51258 , n51248 , n51255 , n51256 , n51257 );
and ( n51259 , n51258 , n41199 );
or ( n51260 , n51241 , n51259 );
and ( n51261 , n51240 , n51260 );
xor ( n51262 , n43847 , n43855 );
xor ( n51263 , n51262 , n43860 );
buf ( n51264 , n51263 );
and ( n51265 , n51264 , n27046 );
xor ( n51266 , n43914 , n43915 );
xor ( n51267 , n51266 , n43920 );
buf ( n51268 , n51267 );
and ( n51269 , n51268 , n27049 );
and ( n51270 , n29353 , n42306 );
or ( n51271 , n51265 , n51269 , n51270 );
buf ( n51272 , n51271 );
and ( n51273 , C1 , n51272 );
or ( n51274 , n51273 , C0 );
buf ( n51275 , n51274 );
not ( n51276 , n51275 );
buf ( n51277 , n51276 );
buf ( n51278 , n51277 );
not ( n51279 , n51278 );
and ( n51280 , C1 , n51279 );
or ( n51281 , n51280 , C0 );
buf ( n51282 , n51281 );
and ( n51283 , n51282 , n24799 );
or ( n51284 , n51261 , n51283 );
and ( n51285 , n51239 , n51284 );
and ( n51286 , n51258 , n24511 );
or ( n51287 , n51285 , n51286 );
and ( n51288 , n51287 , n31008 );
not ( n51289 , n42601 );
and ( n51290 , n51289 , n42555 );
xor ( n51291 , n43957 , n43958 );
and ( n51292 , n51291 , n42601 );
or ( n51293 , n51290 , n51292 );
buf ( n51294 , n51293 );
and ( n51295 , n51294 , n10618 );
or ( n51296 , n51288 , n51295 );
buf ( n51297 , n51296 );
buf ( n51298 , n51297 );
buf ( n51299 , n10613 );
not ( n51300 , n17162 );
not ( n51301 , n17450 );
and ( n51302 , n10648 , n37947 );
not ( n51303 , n38425 );
and ( n51304 , n51303 , n38387 );
xor ( n51305 , n38387 , n38099 );
xor ( n51306 , n38370 , n38099 );
and ( n51307 , n46211 , n46216 );
and ( n51308 , n51306 , n51307 );
xor ( n51309 , n51305 , n51308 );
and ( n51310 , n51309 , n38425 );
or ( n51311 , n51304 , n51310 );
buf ( n51312 , n51311 );
and ( n51313 , n51312 , n19745 );
not ( n51314 , n38934 );
and ( n51315 , n51314 , n38896 );
xor ( n51316 , n38896 , n38608 );
xor ( n51317 , n38879 , n38608 );
and ( n51318 , n46224 , n46229 );
and ( n51319 , n51317 , n51318 );
xor ( n51320 , n51316 , n51319 );
and ( n51321 , n51320 , n38934 );
or ( n51322 , n51315 , n51321 );
buf ( n51323 , n51322 );
and ( n51324 , n51323 , n19748 );
and ( n51325 , n22080 , n21253 );
and ( n51326 , n10648 , n21255 );
or ( n51327 , n51313 , n51324 , n51325 , n51326 );
and ( n51328 , n51327 , n38980 );
or ( n51329 , n51302 , n51328 );
and ( n51330 , n51301 , n51329 );
or ( n51331 , n51330 , C0 );
and ( n51332 , n51300 , n51331 );
and ( n51333 , n51327 , n17162 );
or ( n51334 , n51332 , n51333 );
and ( n51335 , n51334 , n23924 );
not ( n51336 , n39264 );
and ( n51337 , n51336 , n39232 );
xor ( n51338 , n39232 , n38995 );
xor ( n51339 , n39218 , n38995 );
and ( n51340 , n46248 , n46253 );
and ( n51341 , n51339 , n51340 );
xor ( n51342 , n51338 , n51341 );
and ( n51343 , n51342 , n39264 );
or ( n51344 , n51337 , n51343 );
buf ( n51345 , n51344 );
and ( n51346 , n51345 , n23926 );
or ( n51347 , n51335 , n51346 );
buf ( n51348 , n51347 );
buf ( n51349 , n51348 );
buf ( n51350 , n10613 );
not ( n51351 , n17451 );
and ( n51352 , n46077 , n21333 );
and ( n51353 , n19183 , n34758 );
or ( n51354 , n51352 , n51353 );
and ( n51355 , n51354 , n21341 );
and ( n51356 , n46087 , n21333 );
and ( n51357 , n19183 , n34758 );
or ( n51358 , n51356 , n51357 );
and ( n51359 , n51358 , n23064 );
and ( n51360 , n46097 , n21333 );
and ( n51361 , n19183 , n34758 );
or ( n51362 , n51360 , n51361 );
and ( n51363 , n51362 , n23825 );
and ( n51364 , n21984 , n21333 );
and ( n51365 , n19183 , n34758 );
or ( n51366 , n51364 , n51365 );
and ( n51367 , n51366 , n23832 );
and ( n51368 , n46108 , n21333 );
and ( n51369 , n19183 , n34758 );
or ( n51370 , n51368 , n51369 );
and ( n51371 , n51370 , n23917 );
and ( n51372 , n19183 , n34526 );
or ( n51373 , n51355 , n51359 , n51363 , n51367 , n51371 , n51372 );
and ( n51374 , n51351 , n51373 );
and ( n51375 , n19183 , n17451 );
or ( n51376 , n51374 , n51375 );
and ( n51377 , n51376 , n23924 );
and ( n51378 , n19183 , n23926 );
or ( n51379 , n51377 , n51378 );
buf ( n51380 , n51379 );
buf ( n51381 , n51380 );
buf ( n51382 , n10615 );
buf ( n51383 , n10613 );
buf ( n51384 , n10615 );
buf ( n51385 , n10613 );
buf ( n51386 , n10615 );
not ( n51387 , n34821 );
and ( n51388 , n47743 , n36347 );
and ( n51389 , n14960 , n39408 );
or ( n51390 , n51388 , n51389 );
and ( n51391 , n51390 , n14562 );
and ( n51392 , n47759 , n36348 );
and ( n51393 , n14960 , n39427 );
or ( n51394 , n51392 , n51393 );
and ( n51395 , n51394 , n14586 );
and ( n51396 , n47775 , n36347 );
and ( n51397 , n14960 , n39446 );
or ( n51398 , n51396 , n51397 );
and ( n51399 , n51398 , n14584 );
and ( n51400 , n47759 , n36348 );
and ( n51401 , n14960 , n39453 );
or ( n51402 , n51400 , n51401 );
and ( n51403 , n51402 , n37835 );
and ( n51404 , n47775 , n36348 );
and ( n51405 , n14960 , n39453 );
or ( n51406 , n51404 , n51405 );
and ( n51407 , n51406 , n37841 );
and ( n51408 , n14977 , n36348 );
and ( n51409 , n14960 , n39453 );
or ( n51410 , n51408 , n51409 );
and ( n51411 , n51410 , n37847 );
and ( n51412 , n14960 , n37849 );
or ( n51413 , n51391 , n51395 , n51399 , n51403 , n51407 , n51411 , n51412 );
and ( n51414 , n51387 , n51413 );
and ( n51415 , n14960 , n34821 );
or ( n51416 , n51414 , n51415 );
and ( n51417 , n51416 , n16574 );
and ( n51418 , n14960 , n16576 );
or ( n51419 , n51417 , n51418 );
buf ( n51420 , n51419 );
buf ( n51421 , n51420 );
buf ( n51422 , n10613 );
buf ( n51423 , n10613 );
and ( n51424 , n24349 , n31008 );
and ( n51425 , n29144 , n10618 );
or ( n51426 , n51424 , n51425 );
buf ( n51427 , n51426 );
buf ( n51428 , n51427 );
buf ( n51429 , n10615 );
not ( n51430 , n24800 );
and ( n51431 , n45874 , n28586 );
and ( n51432 , n26565 , n34573 );
or ( n51433 , n51431 , n51432 );
and ( n51434 , n51433 , n28594 );
and ( n51435 , n45884 , n28586 );
and ( n51436 , n26565 , n34573 );
or ( n51437 , n51435 , n51436 );
and ( n51438 , n51437 , n30269 );
and ( n51439 , n45894 , n28586 );
and ( n51440 , n26565 , n34573 );
or ( n51441 , n51439 , n51440 );
and ( n51442 , n51441 , n30982 );
and ( n51443 , n29224 , n28586 );
and ( n51444 , n26565 , n34573 );
or ( n51445 , n51443 , n51444 );
and ( n51446 , n51445 , n30989 );
and ( n51447 , n45905 , n28586 );
and ( n51448 , n26565 , n34573 );
or ( n51449 , n51447 , n51448 );
and ( n51450 , n51449 , n31002 );
and ( n51451 , n26565 , n34607 );
or ( n51452 , n51434 , n51438 , n51442 , n51446 , n51450 , n51451 );
and ( n51453 , n51430 , n51452 );
and ( n51454 , n26565 , n24800 );
or ( n51455 , n51453 , n51454 );
and ( n51456 , n51455 , n31008 );
and ( n51457 , n26565 , n10618 );
or ( n51458 , n51456 , n51457 );
buf ( n51459 , n51458 );
buf ( n51460 , n51459 );
buf ( n51461 , n10613 );
and ( n51462 , n24118 , n31008 );
and ( n51463 , n29326 , n10618 );
or ( n51464 , n51462 , n51463 );
buf ( n51465 , n51464 );
buf ( n51466 , n51465 );
buf ( n51467 , n10613 );
and ( n51468 , n16881 , n23924 );
and ( n51469 , n22353 , n23926 );
or ( n51470 , n51468 , n51469 );
buf ( n51471 , n51470 );
buf ( n51472 , n51471 );
not ( n51473 , n17451 );
and ( n51474 , n19113 , n17873 );
and ( n51475 , n39499 , n21330 );
and ( n51476 , n19113 , n21338 );
or ( n51477 , n51475 , n51476 );
and ( n51478 , n51477 , n21341 );
and ( n51479 , n39509 , n21330 );
and ( n51480 , n19113 , n21338 );
or ( n51481 , n51479 , n51480 );
and ( n51482 , n51481 , n23064 );
and ( n51483 , n39519 , n21330 );
and ( n51484 , n19113 , n21338 );
or ( n51485 , n51483 , n51484 );
and ( n51486 , n51485 , n23825 );
and ( n51487 , n22062 , n21330 );
and ( n51488 , n19113 , n21338 );
or ( n51489 , n51487 , n51488 );
and ( n51490 , n51489 , n23832 );
and ( n51491 , n19111 , n23834 );
and ( n51492 , n39529 , n21330 );
and ( n51493 , n19113 , n21338 );
or ( n51494 , n51492 , n51493 );
and ( n51495 , n51494 , n23917 );
or ( n51496 , n51474 , n51478 , n51482 , n51486 , n51490 , n51491 , n51495 );
and ( n51497 , n51473 , n51496 );
and ( n51498 , n19113 , n17451 );
or ( n51499 , n51497 , n51498 );
and ( n51500 , n51499 , n23924 );
and ( n51501 , n19113 , n23926 );
or ( n51502 , n51500 , n51501 );
buf ( n51503 , n51502 );
buf ( n51504 , n51503 );
buf ( n51505 , n10615 );
buf ( n51506 , n10613 );
buf ( n51507 , n10615 );
buf ( n51508 , n10615 );
not ( n51509 , n17451 );
and ( n51510 , n19416 , n17873 );
and ( n51511 , n48266 , n21336 );
and ( n51512 , n19416 , n42682 );
or ( n51513 , n51511 , n51512 );
and ( n51514 , n51513 , n21341 );
and ( n51515 , n48276 , n21336 );
and ( n51516 , n19416 , n42682 );
or ( n51517 , n51515 , n51516 );
and ( n51518 , n51517 , n23064 );
and ( n51519 , n48286 , n21336 );
and ( n51520 , n19416 , n42682 );
or ( n51521 , n51519 , n51520 );
and ( n51522 , n51521 , n23825 );
and ( n51523 , n21893 , n21336 );
and ( n51524 , n19416 , n42682 );
or ( n51525 , n51523 , n51524 );
and ( n51526 , n51525 , n23832 );
and ( n51527 , n21893 , n23834 );
and ( n51528 , n48297 , n21336 );
and ( n51529 , n19416 , n42682 );
or ( n51530 , n51528 , n51529 );
and ( n51531 , n51530 , n23917 );
or ( n51532 , n51510 , n51514 , n51518 , n51522 , n51526 , n51527 , n51531 );
and ( n51533 , n51509 , n51532 );
and ( n51534 , n19416 , n17451 );
or ( n51535 , n51533 , n51534 );
and ( n51536 , n51535 , n23924 );
and ( n51537 , n18275 , n23926 );
or ( n51538 , n51536 , n51537 );
buf ( n51539 , n51538 );
buf ( n51540 , n51539 );
not ( n51541 , n24800 );
not ( n51542 , n26823 );
and ( n51543 , n51542 , n26343 );
xor ( n51544 , n39634 , n39635 );
and ( n51545 , n51544 , n26823 );
or ( n51546 , n51543 , n51545 );
buf ( n51547 , n51546 );
and ( n51548 , n51547 , n27046 );
and ( n51549 , n51547 , n27049 );
not ( n51550 , n27051 );
and ( n51551 , n51550 , n28192 );
not ( n51552 , n28494 );
and ( n51553 , n51552 , n28204 );
xor ( n51554 , n39650 , n39651 );
and ( n51555 , n51554 , n28494 );
or ( n51556 , n51553 , n51555 );
buf ( n51557 , n51556 );
and ( n51558 , n51557 , n27051 );
or ( n51559 , n51551 , n51558 );
and ( n51560 , n51559 , n28506 );
and ( n51561 , n28192 , n28508 );
or ( n51562 , n51548 , n51549 , n51560 , n51561 );
and ( n51563 , n51562 , n28587 );
and ( n51564 , n26363 , n39807 );
or ( n51565 , n51563 , n51564 );
and ( n51566 , n51565 , n28594 );
not ( n51567 , n30249 );
and ( n51568 , n51567 , n30007 );
xor ( n51569 , n39671 , n39672 );
and ( n51570 , n51569 , n30249 );
or ( n51571 , n51568 , n51570 );
buf ( n51572 , n51571 );
and ( n51573 , n51572 , n28587 );
and ( n51574 , n26363 , n39807 );
or ( n51575 , n51573 , n51574 );
and ( n51576 , n51575 , n30269 );
not ( n51577 , n30963 );
and ( n51578 , n51577 , n30721 );
xor ( n51579 , n39687 , n39688 );
and ( n51580 , n51579 , n30963 );
or ( n51581 , n51578 , n51580 );
buf ( n51582 , n51581 );
and ( n51583 , n51582 , n28587 );
and ( n51584 , n26363 , n39807 );
or ( n51585 , n51583 , n51584 );
and ( n51586 , n51585 , n30982 );
and ( n51587 , n29375 , n28587 );
and ( n51588 , n26363 , n39807 );
or ( n51589 , n51587 , n51588 );
and ( n51590 , n51589 , n30989 );
xor ( n51591 , n39708 , n39709 );
buf ( n51592 , n51591 );
and ( n51593 , n51592 , n28587 );
and ( n51594 , n26363 , n39807 );
or ( n51595 , n51593 , n51594 );
and ( n51596 , n51595 , n31002 );
and ( n51597 , n26363 , n34607 );
or ( n51598 , n51566 , n51576 , n51586 , n51590 , n51596 , n51597 );
and ( n51599 , n51541 , n51598 );
and ( n51600 , n26363 , n24800 );
or ( n51601 , n51599 , n51600 );
and ( n51602 , n51601 , n31008 );
and ( n51603 , n26363 , n10618 );
or ( n51604 , n51602 , n51603 );
buf ( n51605 , n51604 );
buf ( n51606 , n51605 );
buf ( n51607 , n10613 );
not ( n51608 , n24800 );
and ( n51609 , n51562 , n28586 );
and ( n51610 , n26361 , n34573 );
or ( n51611 , n51609 , n51610 );
and ( n51612 , n51611 , n28594 );
and ( n51613 , n51572 , n28586 );
and ( n51614 , n26361 , n34573 );
or ( n51615 , n51613 , n51614 );
and ( n51616 , n51615 , n30269 );
and ( n51617 , n51582 , n28586 );
and ( n51618 , n26361 , n34573 );
or ( n51619 , n51617 , n51618 );
and ( n51620 , n51619 , n30982 );
and ( n51621 , n29375 , n28586 );
and ( n51622 , n26361 , n34573 );
or ( n51623 , n51621 , n51622 );
and ( n51624 , n51623 , n30989 );
and ( n51625 , n51592 , n28586 );
and ( n51626 , n26361 , n34573 );
or ( n51627 , n51625 , n51626 );
and ( n51628 , n51627 , n31002 );
and ( n51629 , n26361 , n34607 );
or ( n51630 , n51612 , n51616 , n51620 , n51624 , n51628 , n51629 );
and ( n51631 , n51608 , n51630 );
and ( n51632 , n26361 , n24800 );
or ( n51633 , n51631 , n51632 );
and ( n51634 , n51633 , n31008 );
and ( n51635 , n26361 , n10618 );
or ( n51636 , n51634 , n51635 );
buf ( n51637 , n51636 );
buf ( n51638 , n51637 );
buf ( n51639 , n10615 );
not ( n51640 , n34821 );
and ( n51641 , n13421 , n14592 );
and ( n51642 , n44068 , n36348 );
and ( n51643 , n13421 , n43530 );
or ( n51644 , n51642 , n51643 );
and ( n51645 , n51644 , n14562 );
and ( n51646 , n44078 , n36347 );
and ( n51647 , n13421 , n43543 );
or ( n51648 , n51646 , n51647 );
and ( n51649 , n51648 , n14586 );
and ( n51650 , n44088 , n36348 );
and ( n51651 , n13421 , n43556 );
or ( n51652 , n51650 , n51651 );
and ( n51653 , n51652 , n14584 );
and ( n51654 , n44078 , n36347 );
and ( n51655 , n13421 , n43563 );
or ( n51656 , n51654 , n51655 );
and ( n51657 , n51656 , n37835 );
and ( n51658 , n44088 , n36347 );
and ( n51659 , n13421 , n43563 );
or ( n51660 , n51658 , n51659 );
and ( n51661 , n51660 , n37841 );
and ( n51662 , n13419 , n14564 );
and ( n51663 , n15735 , n36347 );
and ( n51664 , n13421 , n43563 );
or ( n51665 , n51663 , n51664 );
and ( n51666 , n51665 , n37847 );
or ( n51667 , n51641 , n51645 , n51649 , n51653 , n51657 , n51661 , n51662 , n51666 );
and ( n51668 , n51640 , n51667 );
and ( n51669 , n13421 , n34821 );
or ( n51670 , n51668 , n51669 );
and ( n51671 , n51670 , n16574 );
and ( n51672 , n13421 , n16576 );
or ( n51673 , n51671 , n51672 );
buf ( n51674 , n51673 );
buf ( n51675 , n51674 );
buf ( n51676 , n10615 );
and ( n51677 , n16841 , n23924 );
and ( n51678 , n22253 , n23926 );
or ( n51679 , n51677 , n51678 );
buf ( n51680 , n51679 );
buf ( n51681 , n51680 );
buf ( n51682 , n10613 );
buf ( n51683 , n10615 );
buf ( n51684 , n10613 );
buf ( n51685 , n10615 );
not ( n51686 , n34821 );
and ( n51687 , n13193 , n14592 );
and ( n51688 , n49200 , n36348 );
and ( n51689 , n13193 , n43530 );
or ( n51690 , n51688 , n51689 );
and ( n51691 , n51690 , n14562 );
and ( n51692 , n49210 , n36347 );
and ( n51693 , n13193 , n43543 );
or ( n51694 , n51692 , n51693 );
and ( n51695 , n51694 , n14586 );
and ( n51696 , n49220 , n36348 );
and ( n51697 , n13193 , n43556 );
or ( n51698 , n51696 , n51697 );
and ( n51699 , n51698 , n14584 );
and ( n51700 , n49210 , n36347 );
and ( n51701 , n13193 , n43563 );
or ( n51702 , n51700 , n51701 );
and ( n51703 , n51702 , n37835 );
and ( n51704 , n49220 , n36347 );
and ( n51705 , n13193 , n43563 );
or ( n51706 , n51704 , n51705 );
and ( n51707 , n51706 , n37841 );
and ( n51708 , n13191 , n14564 );
and ( n51709 , n15037 , n36347 );
and ( n51710 , n13193 , n43563 );
or ( n51711 , n51709 , n51710 );
and ( n51712 , n51711 , n37847 );
or ( n51713 , n51687 , n51691 , n51695 , n51699 , n51703 , n51707 , n51708 , n51712 );
and ( n51714 , n51686 , n51713 );
and ( n51715 , n13193 , n34821 );
or ( n51716 , n51714 , n51715 );
and ( n51717 , n51716 , n16574 );
and ( n51718 , n13193 , n16576 );
or ( n51719 , n51717 , n51718 );
buf ( n51720 , n51719 );
buf ( n51721 , n51720 );
buf ( n51722 , n10615 );
buf ( n51723 , n10613 );
buf ( n51724 , n10613 );
buf ( n51725 , n10613 );
buf ( n51726 , n10613 );
buf ( n51727 , n10615 );
buf ( n51728 , n10615 );
buf ( n51729 , n10615 );
buf ( n51730 , n10615 );
and ( n51731 , n11800 , n16574 );
and ( n51732 , n15020 , n16576 );
or ( n51733 , n51731 , n51732 );
buf ( n51734 , n51733 );
buf ( n51735 , n51734 );
buf ( n51736 , n10613 );
buf ( n51737 , n10613 );
not ( n51738 , n17162 );
not ( n51739 , n17450 );
and ( n51740 , n10683 , n37947 );
not ( n51741 , n38425 );
and ( n51742 , n51741 , n38268 );
xor ( n51743 , n38430 , n38450 );
and ( n51744 , n51743 , n38425 );
or ( n51745 , n51742 , n51744 );
buf ( n51746 , n51745 );
and ( n51747 , n51746 , n19745 );
not ( n51748 , n38934 );
and ( n51749 , n51748 , n38777 );
xor ( n51750 , n38939 , n38959 );
and ( n51751 , n51750 , n38934 );
or ( n51752 , n51749 , n51751 );
buf ( n51753 , n51752 );
and ( n51754 , n51753 , n19748 );
and ( n51755 , n22220 , n21253 );
and ( n51756 , n10683 , n21255 );
or ( n51757 , n51747 , n51754 , n51755 , n51756 );
and ( n51758 , n51757 , n38980 );
or ( n51759 , n51740 , n51758 );
and ( n51760 , n51739 , n51759 );
or ( n51761 , n51760 , C0 );
and ( n51762 , n51738 , n51761 );
and ( n51763 , n51757 , n17162 );
or ( n51764 , n51762 , n51763 );
and ( n51765 , n51764 , n23924 );
not ( n51766 , n39264 );
and ( n51767 , n51766 , n39134 );
xor ( n51768 , n39269 , n39289 );
and ( n51769 , n51768 , n39264 );
or ( n51770 , n51767 , n51769 );
buf ( n51771 , n51770 );
and ( n51772 , n51771 , n23926 );
or ( n51773 , n51765 , n51772 );
buf ( n51774 , n51773 );
buf ( n51775 , n51774 );
not ( n51776 , n34821 );
and ( n51777 , n48669 , n36347 );
and ( n51778 , n13327 , n39408 );
or ( n51779 , n51777 , n51778 );
and ( n51780 , n51779 , n14562 );
and ( n51781 , n48679 , n36348 );
and ( n51782 , n13327 , n39427 );
or ( n51783 , n51781 , n51782 );
and ( n51784 , n51783 , n14586 );
and ( n51785 , n48689 , n36347 );
and ( n51786 , n13327 , n39446 );
or ( n51787 , n51785 , n51786 );
and ( n51788 , n51787 , n14584 );
and ( n51789 , n48679 , n36348 );
and ( n51790 , n13327 , n39453 );
or ( n51791 , n51789 , n51790 );
and ( n51792 , n51791 , n37835 );
and ( n51793 , n48689 , n36348 );
and ( n51794 , n13327 , n39453 );
or ( n51795 , n51793 , n51794 );
and ( n51796 , n51795 , n37841 );
and ( n51797 , n15559 , n36348 );
and ( n51798 , n13327 , n39453 );
or ( n51799 , n51797 , n51798 );
and ( n51800 , n51799 , n37847 );
and ( n51801 , n13327 , n37849 );
or ( n51802 , n51780 , n51784 , n51788 , n51792 , n51796 , n51800 , n51801 );
and ( n51803 , n51776 , n51802 );
and ( n51804 , n13327 , n34821 );
or ( n51805 , n51803 , n51804 );
and ( n51806 , n51805 , n16574 );
and ( n51807 , n13327 , n16576 );
or ( n51808 , n51806 , n51807 );
buf ( n51809 , n51808 );
buf ( n51810 , n51809 );
buf ( n51811 , n10613 );
not ( n51812 , n34821 );
and ( n51813 , n44068 , n36345 );
and ( n51814 , n13425 , n36352 );
or ( n51815 , n51813 , n51814 );
and ( n51816 , n51815 , n14562 );
and ( n51817 , n44078 , n36345 );
and ( n51818 , n13425 , n37073 );
or ( n51819 , n51817 , n51818 );
and ( n51820 , n51819 , n14586 );
and ( n51821 , n44088 , n36350 );
and ( n51822 , n13425 , n37825 );
or ( n51823 , n51821 , n51822 );
and ( n51824 , n51823 , n14584 );
and ( n51825 , n44078 , n36350 );
and ( n51826 , n13425 , n37831 );
or ( n51827 , n51825 , n51826 );
and ( n51828 , n51827 , n37835 );
and ( n51829 , n44088 , n36350 );
and ( n51830 , n13425 , n37831 );
or ( n51831 , n51829 , n51830 );
and ( n51832 , n51831 , n37841 );
and ( n51833 , n15735 , n36350 );
and ( n51834 , n13425 , n37831 );
or ( n51835 , n51833 , n51834 );
and ( n51836 , n51835 , n37847 );
and ( n51837 , n13425 , n37849 );
or ( n51838 , n51816 , n51820 , n51824 , n51828 , n51832 , n51836 , n51837 );
and ( n51839 , n51812 , n51838 );
and ( n51840 , n13425 , n34821 );
or ( n51841 , n51839 , n51840 );
and ( n51842 , n51841 , n16574 );
and ( n51843 , n13425 , n16576 );
or ( n51844 , n51842 , n51843 );
buf ( n51845 , n51844 );
buf ( n51846 , n51845 );
not ( n51847 , n17451 );
and ( n51848 , n19315 , n17873 );
and ( n51849 , n39576 , n21336 );
and ( n51850 , n19315 , n42682 );
or ( n51851 , n51849 , n51850 );
and ( n51852 , n51851 , n21341 );
and ( n51853 , n39586 , n21336 );
and ( n51854 , n19315 , n42682 );
or ( n51855 , n51853 , n51854 );
and ( n51856 , n51855 , n23064 );
and ( n51857 , n39596 , n21336 );
and ( n51858 , n19315 , n42682 );
or ( n51859 , n51857 , n51858 );
and ( n51860 , n51859 , n23825 );
and ( n51861 , n21932 , n21336 );
and ( n51862 , n19315 , n42682 );
or ( n51863 , n51861 , n51862 );
and ( n51864 , n51863 , n23832 );
and ( n51865 , n21932 , n23834 );
and ( n51866 , n39606 , n21336 );
and ( n51867 , n19315 , n42682 );
or ( n51868 , n51866 , n51867 );
and ( n51869 , n51868 , n23917 );
or ( n51870 , n51848 , n51852 , n51856 , n51860 , n51864 , n51865 , n51869 );
and ( n51871 , n51847 , n51870 );
and ( n51872 , n19315 , n17451 );
or ( n51873 , n51871 , n51872 );
and ( n51874 , n51873 , n23924 );
and ( n51875 , n18230 , n23926 );
or ( n51876 , n51874 , n51875 );
buf ( n51877 , n51876 );
buf ( n51878 , n51877 );
buf ( n51879 , n10615 );
buf ( n51880 , n10615 );
not ( n51881 , n34821 );
and ( n51882 , n49057 , n36347 );
and ( n51883 , n13171 , n39408 );
or ( n51884 , n51882 , n51883 );
and ( n51885 , n51884 , n14562 );
and ( n51886 , n49067 , n36348 );
and ( n51887 , n13171 , n39427 );
or ( n51888 , n51886 , n51887 );
and ( n51889 , n51888 , n14586 );
and ( n51890 , n49077 , n36347 );
and ( n51891 , n13171 , n39446 );
or ( n51892 , n51890 , n51891 );
and ( n51893 , n51892 , n14584 );
and ( n51894 , n49067 , n36348 );
and ( n51895 , n13171 , n39453 );
or ( n51896 , n51894 , n51895 );
and ( n51897 , n51896 , n37835 );
and ( n51898 , n49077 , n36348 );
and ( n51899 , n13171 , n39453 );
or ( n51900 , n51898 , n51899 );
and ( n51901 , n51900 , n37841 );
and ( n51902 , n15007 , n36348 );
and ( n51903 , n13171 , n39453 );
or ( n51904 , n51902 , n51903 );
and ( n51905 , n51904 , n37847 );
and ( n51906 , n13171 , n37849 );
or ( n51907 , n51885 , n51889 , n51893 , n51897 , n51901 , n51905 , n51906 );
and ( n51908 , n51881 , n51907 );
and ( n51909 , n13171 , n34821 );
or ( n51910 , n51908 , n51909 );
and ( n51911 , n51910 , n16574 );
and ( n51912 , n13171 , n16576 );
or ( n51913 , n51911 , n51912 );
buf ( n51914 , n51913 );
buf ( n51915 , n51914 );
buf ( n51916 , n10613 );
buf ( n51917 , n10613 );
not ( n51918 , n24800 );
and ( n51919 , n25917 , n25222 );
and ( n51920 , n34569 , n28589 );
and ( n51921 , n25917 , n31075 );
or ( n51922 , n51920 , n51921 );
and ( n51923 , n51922 , n28594 );
and ( n51924 , n34582 , n28589 );
and ( n51925 , n25917 , n31075 );
or ( n51926 , n51924 , n51925 );
and ( n51927 , n51926 , n30269 );
and ( n51928 , n34592 , n28589 );
and ( n51929 , n25917 , n31075 );
or ( n51930 , n51928 , n51929 );
and ( n51931 , n51930 , n30982 );
and ( n51932 , n29635 , n28589 );
and ( n51933 , n25917 , n31075 );
or ( n51934 , n51932 , n51933 );
and ( n51935 , n51934 , n30989 );
and ( n51936 , n29635 , n30991 );
and ( n51937 , n34602 , n28589 );
and ( n51938 , n25917 , n31075 );
or ( n51939 , n51937 , n51938 );
and ( n51940 , n51939 , n31002 );
or ( n51941 , n51919 , n51923 , n51927 , n51931 , n51935 , n51936 , n51940 );
and ( n51942 , n51918 , n51941 );
and ( n51943 , n25917 , n24800 );
or ( n51944 , n51942 , n51943 );
and ( n51945 , n51944 , n31008 );
and ( n51946 , n25249 , n10618 );
or ( n51947 , n51945 , n51946 );
buf ( n51948 , n51947 );
buf ( n51949 , n51948 );
buf ( n51950 , n10615 );
not ( n51951 , n17451 );
and ( n51952 , n18739 , n17873 );
not ( n51953 , n19474 );
and ( n51954 , n51953 , n18723 );
xor ( n51955 , n19495 , n19507 );
and ( n51956 , n51955 , n19474 );
or ( n51957 , n51954 , n51956 );
buf ( n51958 , n51957 );
and ( n51959 , n51958 , n19745 );
and ( n51960 , n51958 , n19748 );
not ( n51961 , n19750 );
and ( n51962 , n51961 , n20723 );
not ( n51963 , n21193 );
and ( n51964 , n51963 , n20735 );
xor ( n51965 , n21214 , n21228 );
and ( n51966 , n51965 , n21193 );
or ( n51967 , n51964 , n51966 );
buf ( n51968 , n51967 );
and ( n51969 , n51968 , n19750 );
or ( n51970 , n51962 , n51969 );
and ( n51971 , n51970 , n21253 );
and ( n51972 , n20723 , n21255 );
or ( n51973 , n51959 , n51960 , n51971 , n51972 );
and ( n51974 , n51973 , n21330 );
and ( n51975 , n18739 , n21338 );
or ( n51976 , n51974 , n51975 );
and ( n51977 , n51976 , n21341 );
not ( n51978 , n22996 );
and ( n51979 , n51978 , n22618 );
xor ( n51980 , n23017 , n23031 );
and ( n51981 , n51980 , n22996 );
or ( n51982 , n51979 , n51981 );
buf ( n51983 , n51982 );
and ( n51984 , n51983 , n21330 );
and ( n51985 , n18739 , n21338 );
or ( n51986 , n51984 , n51985 );
and ( n51987 , n51986 , n23064 );
not ( n51988 , n23758 );
and ( n51989 , n51988 , n23380 );
xor ( n51990 , n23779 , n23793 );
and ( n51991 , n51990 , n23758 );
or ( n51992 , n51989 , n51991 );
buf ( n51993 , n51992 );
and ( n51994 , n51993 , n21330 );
and ( n51995 , n18739 , n21338 );
or ( n51996 , n51994 , n51995 );
and ( n51997 , n51996 , n23825 );
and ( n51998 , n22282 , n21330 );
and ( n51999 , n18739 , n21338 );
or ( n52000 , n51998 , n51999 );
and ( n52001 , n52000 , n23832 );
and ( n52002 , n18737 , n23834 );
xor ( n52003 , n23873 , n23893 );
buf ( n52004 , n52003 );
and ( n52005 , n52004 , n21330 );
and ( n52006 , n18739 , n21338 );
or ( n52007 , n52005 , n52006 );
and ( n52008 , n52007 , n23917 );
or ( n52009 , n51952 , n51977 , n51987 , n51997 , n52001 , n52002 , n52008 );
and ( n52010 , n51951 , n52009 );
and ( n52011 , n18739 , n17451 );
or ( n52012 , n52010 , n52011 );
and ( n52013 , n52012 , n23924 );
and ( n52014 , n18739 , n23926 );
or ( n52015 , n52013 , n52014 );
buf ( n52016 , n52015 );
buf ( n52017 , n52016 );
not ( n52018 , n34804 );
and ( n52019 , n52018 , n26637 );
and ( n52020 , n14695 , n34804 );
or ( n52021 , n52019 , n52020 );
and ( n52022 , n52021 , n31008 );
and ( n52023 , n14695 , n10618 );
or ( n52024 , n52022 , n52023 );
buf ( n52025 , n52024 );
buf ( n52026 , n52025 );
buf ( n52027 , n10615 );
buf ( n52028 , n10615 );
buf ( n52029 , n10613 );
not ( n52030 , n17451 );
and ( n52031 , n19045 , n17873 );
and ( n52032 , n45943 , n21330 );
and ( n52033 , n19045 , n21338 );
or ( n52034 , n52032 , n52033 );
and ( n52035 , n52034 , n21341 );
and ( n52036 , n45953 , n21330 );
and ( n52037 , n19045 , n21338 );
or ( n52038 , n52036 , n52037 );
and ( n52039 , n52038 , n23064 );
and ( n52040 , n45963 , n21330 );
and ( n52041 , n19045 , n21338 );
or ( n52042 , n52040 , n52041 );
and ( n52043 , n52042 , n23825 );
and ( n52044 , n22102 , n21330 );
and ( n52045 , n19045 , n21338 );
or ( n52046 , n52044 , n52045 );
and ( n52047 , n52046 , n23832 );
and ( n52048 , n19043 , n23834 );
and ( n52049 , n45974 , n21330 );
and ( n52050 , n19045 , n21338 );
or ( n52051 , n52049 , n52050 );
and ( n52052 , n52051 , n23917 );
or ( n52053 , n52031 , n52035 , n52039 , n52043 , n52047 , n52048 , n52052 );
and ( n52054 , n52030 , n52053 );
and ( n52055 , n19045 , n17451 );
or ( n52056 , n52054 , n52055 );
and ( n52057 , n52056 , n23924 );
and ( n52058 , n19045 , n23926 );
or ( n52059 , n52057 , n52058 );
buf ( n52060 , n52059 );
buf ( n52061 , n52060 );
buf ( n52062 , n10613 );
not ( n52063 , n34538 );
and ( n52064 , n52063 , n19085 );
and ( n52065 , n14729 , n34538 );
or ( n52066 , n52064 , n52065 );
and ( n52067 , n52066 , n23924 );
and ( n52068 , n14729 , n23926 );
or ( n52069 , n52067 , n52068 );
buf ( n52070 , n52069 );
buf ( n52071 , n52070 );
buf ( n52072 , n10613 );
buf ( n52073 , n10613 );
not ( n52074 , n34821 );
and ( n52075 , n13140 , n14592 );
and ( n52076 , n47213 , n36348 );
and ( n52077 , n13140 , n43530 );
or ( n52078 , n52076 , n52077 );
and ( n52079 , n52078 , n14562 );
and ( n52080 , n13140 , n43543 );
or ( n52081 , C0 , n52080 );
and ( n52082 , n52081 , n14586 );
and ( n52083 , n13140 , n43556 );
or ( n52084 , C0 , n52083 );
and ( n52085 , n52084 , n14584 );
and ( n52086 , n13140 , n43563 );
or ( n52087 , C0 , n52086 );
and ( n52088 , n52087 , n37835 );
and ( n52089 , n13140 , n43563 );
or ( n52090 , C0 , n52089 );
and ( n52091 , n52090 , n37841 );
and ( n52092 , n12950 , n14564 );
and ( n52093 , n14934 , n36347 );
and ( n52094 , n13140 , n43563 );
or ( n52095 , n52093 , n52094 );
and ( n52096 , n52095 , n37847 );
or ( n52097 , n52075 , n52079 , n52082 , n52085 , n52088 , n52091 , n52092 , n52096 );
and ( n52098 , n52074 , n52097 );
and ( n52099 , n13140 , n34821 );
or ( n52100 , n52098 , n52099 );
and ( n52101 , n52100 , n16574 );
and ( n52102 , n13140 , n16576 );
or ( n52103 , n52101 , n52102 );
buf ( n52104 , n52103 );
buf ( n52105 , n52104 );
buf ( n52106 , n10615 );
buf ( n52107 , n10615 );
buf ( n52108 , n10613 );
buf ( n52109 , n10613 );
buf ( n52110 , n10615 );
buf ( n52111 , n10615 );
buf ( n52112 , n10613 );
and ( n52113 , n24069 , n31008 );
and ( n52114 , n29196 , n10618 );
or ( n52115 , n52113 , n52114 );
buf ( n52116 , n52115 );
buf ( n52117 , n52116 );
buf ( n52118 , n10613 );
buf ( n52119 , n10615 );
buf ( n52120 , n10615 );
buf ( n52121 , n10615 );
buf ( n52122 , n10613 );
buf ( n52123 , n10615 );
buf ( n52124 , n10613 );
buf ( n52125 , n10615 );
buf ( n52126 , n10613 );
not ( n52127 , n34538 );
and ( n52128 , n52127 , n18881 );
and ( n52129 , n14765 , n34538 );
or ( n52130 , n52128 , n52129 );
and ( n52131 , n52130 , n23924 );
and ( n52132 , n14765 , n23926 );
or ( n52133 , n52131 , n52132 );
buf ( n52134 , n52133 );
buf ( n52135 , n52134 );
buf ( n52136 , n10615 );
buf ( n52137 , n10613 );
not ( n52138 , n24800 );
and ( n52139 , n26767 , n25222 );
not ( n52140 , n26823 );
and ( n52141 , n52140 , n26751 );
xor ( n52142 , n45229 , n45232 );
and ( n52143 , n52142 , n26823 );
or ( n52144 , n52141 , n52143 );
buf ( n52145 , n52144 );
and ( n52146 , n52145 , n27046 );
and ( n52147 , n52145 , n27049 );
not ( n52148 , n27051 );
and ( n52149 , n52148 , n28456 );
not ( n52150 , n28494 );
and ( n52151 , n52150 , n28468 );
xor ( n52152 , n45245 , n45248 );
and ( n52153 , n52152 , n28494 );
or ( n52154 , n52151 , n52153 );
buf ( n52155 , n52154 );
and ( n52156 , n52155 , n27051 );
or ( n52157 , n52149 , n52156 );
and ( n52158 , n52157 , n28506 );
and ( n52159 , n28456 , n28508 );
or ( n52160 , n52146 , n52147 , n52158 , n52159 );
and ( n52161 , n52160 , n28583 );
and ( n52162 , n26767 , n28591 );
or ( n52163 , n52161 , n52162 );
and ( n52164 , n52163 , n28594 );
not ( n52165 , n30249 );
and ( n52166 , n52165 , n30211 );
xor ( n52167 , n45266 , n45269 );
and ( n52168 , n52167 , n30249 );
or ( n52169 , n52166 , n52168 );
buf ( n52170 , n52169 );
and ( n52171 , n52170 , n28583 );
and ( n52172 , n26767 , n28591 );
or ( n52173 , n52171 , n52172 );
and ( n52174 , n52173 , n30269 );
not ( n52175 , n30963 );
and ( n52176 , n52175 , n30925 );
xor ( n52177 , n45282 , n45285 );
and ( n52178 , n52177 , n30963 );
or ( n52179 , n52176 , n52178 );
buf ( n52180 , n52179 );
and ( n52181 , n52180 , n28583 );
and ( n52182 , n26767 , n28591 );
or ( n52183 , n52181 , n52182 );
and ( n52184 , n52183 , n30982 );
and ( n52185 , n29146 , n28583 );
and ( n52186 , n26767 , n28591 );
or ( n52187 , n52185 , n52186 );
and ( n52188 , n52187 , n30989 );
and ( n52189 , n26765 , n30991 );
xor ( n52190 , n45303 , n45307 );
buf ( n52191 , n52190 );
and ( n52192 , n52191 , n28583 );
and ( n52193 , n26767 , n28591 );
or ( n52194 , n52192 , n52193 );
and ( n52195 , n52194 , n31002 );
or ( n52196 , n52139 , n52164 , n52174 , n52184 , n52188 , n52189 , n52195 );
and ( n52197 , n52138 , n52196 );
and ( n52198 , n26767 , n24800 );
or ( n52199 , n52197 , n52198 );
and ( n52200 , n52199 , n31008 );
and ( n52201 , n26767 , n10618 );
or ( n52202 , n52200 , n52201 );
buf ( n52203 , n52202 );
buf ( n52204 , n52203 );
not ( n52205 , n17451 );
and ( n52206 , n47363 , n21333 );
and ( n52207 , n18639 , n34758 );
or ( n52208 , n52206 , n52207 );
and ( n52209 , n52208 , n21341 );
and ( n52210 , n47373 , n21333 );
and ( n52211 , n18639 , n34758 );
or ( n52212 , n52210 , n52211 );
and ( n52213 , n52212 , n23064 );
and ( n52214 , n47383 , n21333 );
and ( n52215 , n18639 , n34758 );
or ( n52216 , n52214 , n52215 );
and ( n52217 , n52216 , n23825 );
and ( n52218 , n22342 , n21333 );
and ( n52219 , n18639 , n34758 );
or ( n52220 , n52218 , n52219 );
and ( n52221 , n52220 , n23832 );
and ( n52222 , n47394 , n21333 );
and ( n52223 , n18639 , n34758 );
or ( n52224 , n52222 , n52223 );
and ( n52225 , n52224 , n23917 );
and ( n52226 , n18639 , n34526 );
or ( n52227 , n52209 , n52213 , n52217 , n52221 , n52225 , n52226 );
and ( n52228 , n52205 , n52227 );
and ( n52229 , n18639 , n17451 );
or ( n52230 , n52228 , n52229 );
and ( n52231 , n52230 , n23924 );
and ( n52232 , n18639 , n23926 );
or ( n52233 , n52231 , n52232 );
buf ( n52234 , n52233 );
buf ( n52235 , n52234 );
buf ( n52236 , n10613 );
not ( n52237 , n24800 );
and ( n52238 , n39944 , n28586 );
and ( n52239 , n25857 , n34573 );
or ( n52240 , n52238 , n52239 );
and ( n52241 , n52240 , n28594 );
and ( n52242 , n39954 , n28586 );
and ( n52243 , n25857 , n34573 );
or ( n52244 , n52242 , n52243 );
and ( n52245 , n52244 , n30269 );
and ( n52246 , n39964 , n28586 );
and ( n52247 , n25857 , n34573 );
or ( n52248 , n52246 , n52247 );
and ( n52249 , n52248 , n30982 );
and ( n52250 , n28892 , n28586 );
and ( n52251 , n25857 , n34573 );
or ( n52252 , n52250 , n52251 );
and ( n52253 , n52252 , n30989 );
and ( n52254 , n39974 , n28586 );
and ( n52255 , n25857 , n34573 );
or ( n52256 , n52254 , n52255 );
and ( n52257 , n52256 , n31002 );
and ( n52258 , n25857 , n34607 );
or ( n52259 , n52241 , n52245 , n52249 , n52253 , n52257 , n52258 );
and ( n52260 , n52237 , n52259 );
and ( n52261 , n25857 , n24800 );
or ( n52262 , n52260 , n52261 );
and ( n52263 , n52262 , n31008 );
and ( n52264 , n25857 , n10618 );
or ( n52265 , n52263 , n52264 );
buf ( n52266 , n52265 );
buf ( n52267 , n52266 );
buf ( n52268 , n10613 );
not ( n52269 , n17162 );
not ( n52270 , n17450 );
and ( n52271 , n10638 , n37947 );
not ( n52272 , n38425 );
and ( n52273 , n52272 , n38421 );
xor ( n52274 , n38421 , n38099 );
xor ( n52275 , n38404 , n38099 );
and ( n52276 , n51305 , n51308 );
and ( n52277 , n52275 , n52276 );
xor ( n52278 , n52274 , n52277 );
and ( n52279 , n52278 , n38425 );
or ( n52280 , n52273 , n52279 );
buf ( n52281 , n52280 );
and ( n52282 , n52281 , n19745 );
not ( n52283 , n38934 );
and ( n52284 , n52283 , n38930 );
xor ( n52285 , n38930 , n38608 );
xor ( n52286 , n38913 , n38608 );
and ( n52287 , n51316 , n51319 );
and ( n52288 , n52286 , n52287 );
xor ( n52289 , n52285 , n52288 );
and ( n52290 , n52289 , n38934 );
or ( n52291 , n52284 , n52290 );
buf ( n52292 , n52291 );
and ( n52293 , n52292 , n19748 );
and ( n52294 , n22040 , n21253 );
and ( n52295 , n10638 , n21255 );
or ( n52296 , n52282 , n52293 , n52294 , n52295 );
and ( n52297 , n52296 , n38980 );
or ( n52298 , n52271 , n52297 );
and ( n52299 , n52270 , n52298 );
or ( n52300 , n52299 , C0 );
and ( n52301 , n52269 , n52300 );
and ( n52302 , n52296 , n17162 );
or ( n52303 , n52301 , n52302 );
and ( n52304 , n52303 , n23924 );
not ( n52305 , n39264 );
and ( n52306 , n52305 , n39260 );
xor ( n52307 , n39260 , n38995 );
xor ( n52308 , n39246 , n38995 );
and ( n52309 , n51338 , n51341 );
and ( n52310 , n52308 , n52309 );
xor ( n52311 , n52307 , n52310 );
and ( n52312 , n52311 , n39264 );
or ( n52313 , n52306 , n52312 );
buf ( n52314 , n52313 );
and ( n52315 , n52314 , n23926 );
or ( n52316 , n52304 , n52315 );
buf ( n52317 , n52316 );
buf ( n52318 , n52317 );
buf ( n52319 , n10613 );
buf ( n52320 , n10613 );
buf ( n52321 , n10613 );
buf ( n52322 , n10613 );
buf ( n52323 , n10613 );
buf ( n52324 , n10613 );
not ( n52325 , n34538 );
and ( n52326 , n52325 , n18745 );
and ( n52327 , n14789 , n34538 );
or ( n52328 , n52326 , n52327 );
and ( n52329 , n52328 , n23924 );
and ( n52330 , n14789 , n23926 );
or ( n52331 , n52329 , n52330 );
buf ( n52332 , n52331 );
buf ( n52333 , n52332 );
not ( n52334 , n17451 );
and ( n52335 , n19382 , n17873 );
and ( n52336 , n39876 , n21336 );
and ( n52337 , n19382 , n42682 );
or ( n52338 , n52336 , n52337 );
and ( n52339 , n52338 , n21341 );
and ( n52340 , n39888 , n21336 );
and ( n52341 , n19382 , n42682 );
or ( n52342 , n52340 , n52341 );
and ( n52343 , n52342 , n23064 );
and ( n52344 , n39900 , n21336 );
and ( n52345 , n19382 , n42682 );
or ( n52346 , n52344 , n52345 );
and ( n52347 , n52346 , n23825 );
and ( n52348 , n21906 , n21336 );
and ( n52349 , n19382 , n42682 );
or ( n52350 , n52348 , n52349 );
and ( n52351 , n52350 , n23832 );
and ( n52352 , n21906 , n23834 );
and ( n52353 , n39913 , n21336 );
and ( n52354 , n19382 , n42682 );
or ( n52355 , n52353 , n52354 );
and ( n52356 , n52355 , n23917 );
or ( n52357 , n52335 , n52339 , n52343 , n52347 , n52351 , n52352 , n52356 );
and ( n52358 , n52334 , n52357 );
and ( n52359 , n19382 , n17451 );
or ( n52360 , n52358 , n52359 );
and ( n52361 , n52360 , n23924 );
and ( n52362 , n18260 , n23926 );
or ( n52363 , n52361 , n52362 );
buf ( n52364 , n52363 );
buf ( n52365 , n52364 );
not ( n52366 , n24800 );
and ( n52367 , n26289 , n25222 );
and ( n52368 , n45088 , n28589 );
and ( n52369 , n26289 , n31075 );
or ( n52370 , n52368 , n52369 );
and ( n52371 , n52370 , n28594 );
and ( n52372 , n45098 , n28589 );
and ( n52373 , n26289 , n31075 );
or ( n52374 , n52372 , n52373 );
and ( n52375 , n52374 , n30269 );
and ( n52376 , n45108 , n28589 );
and ( n52377 , n26289 , n31075 );
or ( n52378 , n52376 , n52377 );
and ( n52379 , n52378 , n30982 );
and ( n52380 , n29415 , n28589 );
and ( n52381 , n26289 , n31075 );
or ( n52382 , n52380 , n52381 );
and ( n52383 , n52382 , n30989 );
and ( n52384 , n29415 , n30991 );
and ( n52385 , n45119 , n28589 );
and ( n52386 , n26289 , n31075 );
or ( n52387 , n52385 , n52386 );
and ( n52388 , n52387 , n31002 );
or ( n52389 , n52367 , n52371 , n52375 , n52379 , n52383 , n52384 , n52388 );
and ( n52390 , n52366 , n52389 );
and ( n52391 , n26289 , n24800 );
or ( n52392 , n52390 , n52391 );
and ( n52393 , n52392 , n31008 );
and ( n52394 , n25414 , n10618 );
or ( n52395 , n52393 , n52394 );
buf ( n52396 , n52395 );
buf ( n52397 , n52396 );
and ( n52398 , n16729 , n23924 );
and ( n52399 , n21956 , n23926 );
or ( n52400 , n52398 , n52399 );
buf ( n52401 , n52400 );
buf ( n52402 , n52401 );
buf ( n52403 , n10615 );
not ( n52404 , n24800 );
and ( n52405 , n48113 , n28587 );
and ( n52406 , n26397 , n39807 );
or ( n52407 , n52405 , n52406 );
and ( n52408 , n52407 , n28594 );
and ( n52409 , n48123 , n28587 );
and ( n52410 , n26397 , n39807 );
or ( n52411 , n52409 , n52410 );
and ( n52412 , n52411 , n30269 );
and ( n52413 , n48133 , n28587 );
and ( n52414 , n26397 , n39807 );
or ( n52415 , n52413 , n52414 );
and ( n52416 , n52415 , n30982 );
and ( n52417 , n29355 , n28587 );
and ( n52418 , n26397 , n39807 );
or ( n52419 , n52417 , n52418 );
and ( n52420 , n52419 , n30989 );
and ( n52421 , n48144 , n28587 );
and ( n52422 , n26397 , n39807 );
or ( n52423 , n52421 , n52422 );
and ( n52424 , n52423 , n31002 );
and ( n52425 , n26397 , n34607 );
or ( n52426 , n52408 , n52412 , n52416 , n52420 , n52424 , n52425 );
and ( n52427 , n52404 , n52426 );
and ( n52428 , n26397 , n24800 );
or ( n52429 , n52427 , n52428 );
and ( n52430 , n52429 , n31008 );
and ( n52431 , n26397 , n10618 );
or ( n52432 , n52430 , n52431 );
buf ( n52433 , n52432 );
buf ( n52434 , n52433 );
not ( n52435 , n24800 );
and ( n52436 , n44989 , n28587 );
and ( n52437 , n26261 , n39807 );
or ( n52438 , n52436 , n52437 );
and ( n52439 , n52438 , n28594 );
and ( n52440 , n44999 , n28587 );
and ( n52441 , n26261 , n39807 );
or ( n52442 , n52440 , n52441 );
and ( n52443 , n52442 , n30269 );
and ( n52444 , n45009 , n28587 );
and ( n52445 , n26261 , n39807 );
or ( n52446 , n52444 , n52445 );
and ( n52447 , n52446 , n30982 );
and ( n52448 , n29435 , n28587 );
and ( n52449 , n26261 , n39807 );
or ( n52450 , n52448 , n52449 );
and ( n52451 , n52450 , n30989 );
and ( n52452 , n45019 , n28587 );
and ( n52453 , n26261 , n39807 );
or ( n52454 , n52452 , n52453 );
and ( n52455 , n52454 , n31002 );
and ( n52456 , n26261 , n34607 );
or ( n52457 , n52439 , n52443 , n52447 , n52451 , n52455 , n52456 );
and ( n52458 , n52435 , n52457 );
and ( n52459 , n26261 , n24800 );
or ( n52460 , n52458 , n52459 );
and ( n52461 , n52460 , n31008 );
and ( n52462 , n26261 , n10618 );
or ( n52463 , n52461 , n52462 );
buf ( n52464 , n52463 );
buf ( n52465 , n52464 );
and ( n52466 , n16769 , n23924 );
and ( n52467 , n22073 , n23926 );
or ( n52468 , n52466 , n52467 );
buf ( n52469 , n52468 );
buf ( n52470 , n52469 );
not ( n52471 , n17451 );
and ( n52472 , n19349 , n17873 );
and ( n52473 , n21257 , n21336 );
and ( n52474 , n19349 , n42682 );
or ( n52475 , n52473 , n52474 );
and ( n52476 , n52475 , n21341 );
and ( n52477 , n23053 , n21336 );
and ( n52478 , n19349 , n42682 );
or ( n52479 , n52477 , n52478 );
and ( n52480 , n52479 , n23064 );
and ( n52481 , n23815 , n21336 );
and ( n52482 , n19349 , n42682 );
or ( n52483 , n52481 , n52482 );
and ( n52484 , n52483 , n23825 );
and ( n52485 , n21919 , n21336 );
and ( n52486 , n19349 , n42682 );
or ( n52487 , n52485 , n52486 );
and ( n52488 , n52487 , n23832 );
and ( n52489 , n21919 , n23834 );
and ( n52490 , n23913 , n21336 );
and ( n52491 , n19349 , n42682 );
or ( n52492 , n52490 , n52491 );
and ( n52493 , n52492 , n23917 );
or ( n52494 , n52472 , n52476 , n52480 , n52484 , n52488 , n52489 , n52493 );
and ( n52495 , n52471 , n52494 );
and ( n52496 , n19349 , n17451 );
or ( n52497 , n52495 , n52496 );
and ( n52498 , n52497 , n23924 );
and ( n52499 , n18245 , n23926 );
or ( n52500 , n52498 , n52499 );
buf ( n52501 , n52500 );
buf ( n52502 , n52501 );
not ( n52503 , n24511 );
not ( n52504 , n24799 );
and ( n52505 , n10695 , n40154 );
not ( n52506 , n40632 );
and ( n52507 , n52506 , n40441 );
xor ( n52508 , n40642 , n40658 );
and ( n52509 , n52508 , n40632 );
or ( n52510 , n52507 , n52509 );
buf ( n52511 , n52510 );
and ( n52512 , n52511 , n27046 );
not ( n52513 , n41147 );
and ( n52514 , n52513 , n40956 );
xor ( n52515 , n41157 , n41173 );
and ( n52516 , n52515 , n41147 );
or ( n52517 , n52514 , n52516 );
buf ( n52518 , n52517 );
and ( n52519 , n52518 , n27049 );
and ( n52520 , n29513 , n28506 );
and ( n52521 , n10695 , n28508 );
or ( n52522 , n52512 , n52519 , n52520 , n52521 );
and ( n52523 , n52522 , n41199 );
or ( n52524 , n52505 , n52523 );
and ( n52525 , n52504 , n52524 );
xor ( n52526 , n41628 , n41636 );
xor ( n52527 , n52526 , n41785 );
buf ( n52528 , n52527 );
and ( n52529 , n52528 , n27046 );
xor ( n52530 , n42186 , n42187 );
xor ( n52531 , n52530 , n42281 );
buf ( n52532 , n52531 );
and ( n52533 , n52532 , n27049 );
and ( n52534 , n29513 , n42306 );
or ( n52535 , n52529 , n52533 , n52534 );
buf ( n52536 , n52535 );
and ( n52537 , C1 , n52536 );
or ( n52538 , n52537 , C0 );
buf ( n52539 , n52538 );
not ( n52540 , n52539 );
buf ( n52541 , n52540 );
buf ( n52542 , n52541 );
not ( n52543 , n52542 );
and ( n52544 , C1 , n52543 );
or ( n52545 , n52544 , C0 );
buf ( n52546 , n52545 );
and ( n52547 , n52546 , n24799 );
or ( n52548 , n52525 , n52547 );
and ( n52549 , n52503 , n52548 );
and ( n52550 , n52522 , n24511 );
or ( n52551 , n52549 , n52550 );
and ( n52552 , n52551 , n31008 );
not ( n52553 , n42601 );
and ( n52554 , n52553 , n42443 );
xor ( n52555 , n42611 , n42627 );
and ( n52556 , n52555 , n42601 );
or ( n52557 , n52554 , n52556 );
buf ( n52558 , n52557 );
and ( n52559 , n52558 , n10618 );
or ( n52560 , n52552 , n52559 );
buf ( n52561 , n52560 );
buf ( n52562 , n52561 );
buf ( n52563 , n10615 );
buf ( n52564 , n10613 );
not ( n52565 , n24800 );
and ( n52566 , n52160 , n28587 );
and ( n52567 , n26771 , n39807 );
or ( n52568 , n52566 , n52567 );
and ( n52569 , n52568 , n28594 );
and ( n52570 , n52170 , n28587 );
and ( n52571 , n26771 , n39807 );
or ( n52572 , n52570 , n52571 );
and ( n52573 , n52572 , n30269 );
and ( n52574 , n52180 , n28587 );
and ( n52575 , n26771 , n39807 );
or ( n52576 , n52574 , n52575 );
and ( n52577 , n52576 , n30982 );
and ( n52578 , n29146 , n28587 );
and ( n52579 , n26771 , n39807 );
or ( n52580 , n52578 , n52579 );
and ( n52581 , n52580 , n30989 );
and ( n52582 , n52191 , n28587 );
and ( n52583 , n26771 , n39807 );
or ( n52584 , n52582 , n52583 );
and ( n52585 , n52584 , n31002 );
and ( n52586 , n26771 , n34607 );
or ( n52587 , n52569 , n52573 , n52577 , n52581 , n52585 , n52586 );
and ( n52588 , n52565 , n52587 );
and ( n52589 , n26771 , n24800 );
or ( n52590 , n52588 , n52589 );
and ( n52591 , n52590 , n31008 );
and ( n52592 , n26771 , n10618 );
or ( n52593 , n52591 , n52592 );
buf ( n52594 , n52593 );
buf ( n52595 , n52594 );
buf ( n52596 , n10613 );
not ( n52597 , n34538 );
and ( n52598 , n52597 , n19255 );
and ( n52599 , n14699 , n34538 );
or ( n52600 , n52598 , n52599 );
and ( n52601 , n52600 , n23924 );
and ( n52602 , n14699 , n23926 );
or ( n52603 , n52601 , n52602 );
buf ( n52604 , n52603 );
buf ( n52605 , n52604 );
not ( n52606 , n24800 );
and ( n52607 , n50001 , n28586 );
and ( n52608 , n26157 , n34573 );
or ( n52609 , n52607 , n52608 );
and ( n52610 , n52609 , n28594 );
and ( n52611 , n50011 , n28586 );
and ( n52612 , n26157 , n34573 );
or ( n52613 , n52611 , n52612 );
and ( n52614 , n52613 , n30269 );
and ( n52615 , n50021 , n28586 );
and ( n52616 , n26157 , n34573 );
or ( n52617 , n52615 , n52616 );
and ( n52618 , n52617 , n30982 );
and ( n52619 , n29495 , n28586 );
and ( n52620 , n26157 , n34573 );
or ( n52621 , n52619 , n52620 );
and ( n52622 , n52621 , n30989 );
and ( n52623 , n50032 , n28586 );
and ( n52624 , n26157 , n34573 );
or ( n52625 , n52623 , n52624 );
and ( n52626 , n52625 , n31002 );
and ( n52627 , n26157 , n34607 );
or ( n52628 , n52610 , n52614 , n52618 , n52622 , n52626 , n52627 );
and ( n52629 , n52606 , n52628 );
and ( n52630 , n26157 , n24800 );
or ( n52631 , n52629 , n52630 );
and ( n52632 , n52631 , n31008 );
and ( n52633 , n26157 , n10618 );
or ( n52634 , n52632 , n52633 );
buf ( n52635 , n52634 );
buf ( n52636 , n52635 );
buf ( n52637 , n10613 );
buf ( n52638 , n10615 );
buf ( n52639 , n10615 );
buf ( n52640 , n10615 );
buf ( n52641 , n10615 );
buf ( n52642 , n10613 );
not ( n52643 , n34538 );
and ( n52644 , n52643 , n18847 );
and ( n52645 , n14771 , n34538 );
or ( n52646 , n52644 , n52645 );
and ( n52647 , n52646 , n23924 );
and ( n52648 , n14771 , n23926 );
or ( n52649 , n52647 , n52648 );
buf ( n52650 , n52649 );
buf ( n52651 , n52650 );
not ( n52652 , n34804 );
and ( n52653 , n52652 , n26501 );
and ( n52654 , n14719 , n34804 );
or ( n52655 , n52653 , n52654 );
and ( n52656 , n52655 , n31008 );
and ( n52657 , n14719 , n10618 );
or ( n52658 , n52656 , n52657 );
buf ( n52659 , n52658 );
buf ( n52660 , n52659 );
buf ( n52661 , n10615 );
not ( n52662 , n11333 );
and ( n52663 , n52662 , n11091 );
xor ( n52664 , n11346 , n11356 );
and ( n52665 , n52664 , n11333 );
or ( n52666 , n52663 , n52665 );
buf ( n52667 , n52666 );
buf ( n52668 , n52667 );
not ( n52669 , n34821 );
and ( n52670 , n46158 , n36347 );
and ( n52671 , n13279 , n39408 );
or ( n52672 , n52670 , n52671 );
and ( n52673 , n52672 , n14562 );
and ( n52674 , n46168 , n36348 );
and ( n52675 , n13279 , n39427 );
or ( n52676 , n52674 , n52675 );
and ( n52677 , n52676 , n14586 );
and ( n52678 , n46178 , n36347 );
and ( n52679 , n13279 , n39446 );
or ( n52680 , n52678 , n52679 );
and ( n52681 , n52680 , n14584 );
and ( n52682 , n46168 , n36348 );
and ( n52683 , n13279 , n39453 );
or ( n52684 , n52682 , n52683 );
and ( n52685 , n52684 , n37835 );
and ( n52686 , n46178 , n36348 );
and ( n52687 , n13279 , n39453 );
or ( n52688 , n52686 , n52687 );
and ( n52689 , n52688 , n37841 );
and ( n52690 , n15471 , n36348 );
and ( n52691 , n13279 , n39453 );
or ( n52692 , n52690 , n52691 );
and ( n52693 , n52692 , n37847 );
and ( n52694 , n13279 , n37849 );
or ( n52695 , n52673 , n52677 , n52681 , n52685 , n52689 , n52693 , n52694 );
and ( n52696 , n52669 , n52695 );
and ( n52697 , n13279 , n34821 );
or ( n52698 , n52696 , n52697 );
and ( n52699 , n52698 , n16574 );
and ( n52700 , n13279 , n16576 );
or ( n52701 , n52699 , n52700 );
buf ( n52702 , n52701 );
buf ( n52703 , n52702 );
not ( n52704 , n34821 );
and ( n52705 , n13313 , n14592 );
and ( n52706 , n45425 , n36348 );
and ( n52707 , n13313 , n43530 );
or ( n52708 , n52706 , n52707 );
and ( n52709 , n52708 , n14562 );
and ( n52710 , n45435 , n36347 );
and ( n52711 , n13313 , n43543 );
or ( n52712 , n52710 , n52711 );
and ( n52713 , n52712 , n14586 );
and ( n52714 , n45445 , n36348 );
and ( n52715 , n13313 , n43556 );
or ( n52716 , n52714 , n52715 );
and ( n52717 , n52716 , n14584 );
and ( n52718 , n45435 , n36347 );
and ( n52719 , n13313 , n43563 );
or ( n52720 , n52718 , n52719 );
and ( n52721 , n52720 , n37835 );
and ( n52722 , n45445 , n36347 );
and ( n52723 , n13313 , n43563 );
or ( n52724 , n52722 , n52723 );
and ( n52725 , n52724 , n37841 );
and ( n52726 , n13311 , n14564 );
and ( n52727 , n15537 , n36347 );
and ( n52728 , n13313 , n43563 );
or ( n52729 , n52727 , n52728 );
and ( n52730 , n52729 , n37847 );
or ( n52731 , n52705 , n52709 , n52713 , n52717 , n52721 , n52725 , n52726 , n52730 );
and ( n52732 , n52704 , n52731 );
and ( n52733 , n13313 , n34821 );
or ( n52734 , n52732 , n52733 );
and ( n52735 , n52734 , n16574 );
and ( n52736 , n13313 , n16576 );
or ( n52737 , n52735 , n52736 );
buf ( n52738 , n52737 );
buf ( n52739 , n52738 );
and ( n52740 , n16801 , n23924 );
and ( n52741 , n22153 , n23926 );
or ( n52742 , n52740 , n52741 );
buf ( n52743 , n52742 );
buf ( n52744 , n52743 );
buf ( n52745 , n10613 );
buf ( n52746 , n10615 );
buf ( n52747 , n10613 );
not ( n52748 , n34538 );
and ( n52749 , n52748 , n19424 );
and ( n52750 , n14669 , n34538 );
or ( n52751 , n52749 , n52750 );
and ( n52752 , n52751 , n23924 );
and ( n52753 , n14669 , n23926 );
or ( n52754 , n52752 , n52753 );
buf ( n52755 , n52754 );
buf ( n52756 , n52755 );
buf ( n52757 , n10613 );
buf ( n52758 , n10613 );
buf ( n52759 , n10615 );
buf ( n52760 , n10615 );
buf ( n52761 , n10613 );
buf ( n52762 , n10615 );
buf ( n52763 , n10613 );
buf ( n52764 , n10613 );
buf ( n52765 , n10613 );
not ( n52766 , n24800 );
and ( n52767 , n34569 , n28587 );
and ( n52768 , n25923 , n39807 );
or ( n52769 , n52767 , n52768 );
and ( n52770 , n52769 , n28594 );
and ( n52771 , n34582 , n28587 );
and ( n52772 , n25923 , n39807 );
or ( n52773 , n52771 , n52772 );
and ( n52774 , n52773 , n30269 );
and ( n52775 , n34592 , n28587 );
and ( n52776 , n25923 , n39807 );
or ( n52777 , n52775 , n52776 );
and ( n52778 , n52777 , n30982 );
and ( n52779 , n29635 , n28587 );
and ( n52780 , n25923 , n39807 );
or ( n52781 , n52779 , n52780 );
and ( n52782 , n52781 , n30989 );
and ( n52783 , n34602 , n28587 );
and ( n52784 , n25923 , n39807 );
or ( n52785 , n52783 , n52784 );
and ( n52786 , n52785 , n31002 );
and ( n52787 , n25923 , n34607 );
or ( n52788 , n52770 , n52774 , n52778 , n52782 , n52786 , n52787 );
and ( n52789 , n52766 , n52788 );
and ( n52790 , n25923 , n24800 );
or ( n52791 , n52789 , n52790 );
and ( n52792 , n52791 , n31008 );
and ( n52793 , n25923 , n10618 );
or ( n52794 , n52792 , n52793 );
buf ( n52795 , n52794 );
buf ( n52796 , n52795 );
and ( n52797 , n24214 , n31008 );
and ( n52798 , n29566 , n10618 );
or ( n52799 , n52797 , n52798 );
buf ( n52800 , n52799 );
buf ( n52801 , n52800 );
buf ( n52802 , n10613 );
buf ( n52803 , n10613 );
buf ( n52804 , n10613 );
buf ( n52805 , n10613 );
not ( n52806 , n17451 );
and ( n52807 , n47038 , n21334 );
and ( n52808 , n19287 , n34492 );
or ( n52809 , n52807 , n52808 );
and ( n52810 , n52809 , n21341 );
and ( n52811 , n47048 , n21334 );
and ( n52812 , n19287 , n34492 );
or ( n52813 , n52811 , n52812 );
and ( n52814 , n52813 , n23064 );
and ( n52815 , n47058 , n21334 );
and ( n52816 , n19287 , n34492 );
or ( n52817 , n52815 , n52816 );
and ( n52818 , n52817 , n23825 );
and ( n52819 , n21945 , n21334 );
and ( n52820 , n19287 , n34492 );
or ( n52821 , n52819 , n52820 );
and ( n52822 , n52821 , n23832 );
and ( n52823 , n47068 , n21334 );
and ( n52824 , n19287 , n34492 );
or ( n52825 , n52823 , n52824 );
and ( n52826 , n52825 , n23917 );
and ( n52827 , n19287 , n34526 );
or ( n52828 , n52810 , n52814 , n52818 , n52822 , n52826 , n52827 );
and ( n52829 , n52806 , n52828 );
and ( n52830 , n19287 , n17451 );
or ( n52831 , n52829 , n52830 );
and ( n52832 , n52831 , n23924 );
and ( n52833 , n19287 , n23926 );
or ( n52834 , n52832 , n52833 );
buf ( n52835 , n52834 );
buf ( n52836 , n52835 );
buf ( n52837 , n10615 );
not ( n52838 , n17162 );
buf ( n52839 , n21353 );
buf ( n52840 , n52839 );
and ( n52841 , n52840 , n38980 );
buf ( n52842 , n52841 );
not ( n52843 , n17450 );
and ( n52844 , n52842 , n52843 );
and ( n52845 , n52838 , n52844 );
and ( n52846 , n52840 , n17162 );
or ( n52847 , n52845 , n52846 );
and ( n52848 , n52847 , n23924 );
buf ( n52849 , n23926 );
or ( n52850 , n52848 , n52849 );
buf ( n52851 , n52850 );
buf ( n52852 , n52851 );
buf ( n52853 , n10615 );
buf ( n52854 , n10615 );
buf ( n52855 , n10615 );
buf ( n52856 , n10613 );
not ( n52857 , n24800 );
not ( n52858 , n26823 );
and ( n52859 , n52858 , n26513 );
xor ( n52860 , n42828 , n42833 );
and ( n52861 , n52860 , n26823 );
or ( n52862 , n52859 , n52861 );
buf ( n52863 , n52862 );
and ( n52864 , n52863 , n27046 );
and ( n52865 , n52863 , n27049 );
not ( n52866 , n27051 );
and ( n52867 , n52866 , n28302 );
not ( n52868 , n28494 );
and ( n52869 , n52868 , n28314 );
xor ( n52870 , n42848 , n42853 );
and ( n52871 , n52870 , n28494 );
or ( n52872 , n52869 , n52871 );
buf ( n52873 , n52872 );
and ( n52874 , n52873 , n27051 );
or ( n52875 , n52867 , n52874 );
and ( n52876 , n52875 , n28506 );
and ( n52877 , n28302 , n28508 );
or ( n52878 , n52864 , n52865 , n52876 , n52877 );
and ( n52879 , n52878 , n28587 );
and ( n52880 , n26533 , n39807 );
or ( n52881 , n52879 , n52880 );
and ( n52882 , n52881 , n28594 );
not ( n52883 , n30249 );
and ( n52884 , n52883 , n30092 );
xor ( n52885 , n42873 , n42878 );
and ( n52886 , n52885 , n30249 );
or ( n52887 , n52884 , n52886 );
buf ( n52888 , n52887 );
and ( n52889 , n52888 , n28587 );
and ( n52890 , n26533 , n39807 );
or ( n52891 , n52889 , n52890 );
and ( n52892 , n52891 , n30269 );
not ( n52893 , n30963 );
and ( n52894 , n52893 , n30806 );
xor ( n52895 , n42893 , n42898 );
and ( n52896 , n52895 , n30963 );
or ( n52897 , n52894 , n52896 );
buf ( n52898 , n52897 );
and ( n52899 , n52898 , n28587 );
and ( n52900 , n26533 , n39807 );
or ( n52901 , n52899 , n52900 );
and ( n52902 , n52901 , n30982 );
and ( n52903 , n29237 , n28587 );
and ( n52904 , n26533 , n39807 );
or ( n52905 , n52903 , n52904 );
and ( n52906 , n52905 , n30989 );
xor ( n52907 , n42918 , n42925 );
buf ( n52908 , n52907 );
and ( n52909 , n52908 , n28587 );
and ( n52910 , n26533 , n39807 );
or ( n52911 , n52909 , n52910 );
and ( n52912 , n52911 , n31002 );
and ( n52913 , n26533 , n34607 );
or ( n52914 , n52882 , n52892 , n52902 , n52906 , n52912 , n52913 );
and ( n52915 , n52857 , n52914 );
and ( n52916 , n26533 , n24800 );
or ( n52917 , n52915 , n52916 );
and ( n52918 , n52917 , n31008 );
and ( n52919 , n26533 , n10618 );
or ( n52920 , n52918 , n52919 );
buf ( n52921 , n52920 );
buf ( n52922 , n52921 );
buf ( n52923 , n10615 );
buf ( n52924 , n10615 );
and ( n52925 , n16873 , n23924 );
and ( n52926 , n22333 , n23926 );
or ( n52927 , n52925 , n52926 );
buf ( n52928 , n52927 );
buf ( n52929 , n52928 );
buf ( n52930 , n10613 );
buf ( n52931 , n10615 );
buf ( n52932 , n10615 );
not ( n52933 , n17451 );
and ( n52934 , n18521 , n17873 );
not ( n52935 , n19750 );
and ( n52936 , n52935 , n20581 );
or ( n52937 , n52936 , C0 );
and ( n52938 , n52937 , n21253 );
and ( n52939 , n20581 , n21255 );
or ( n52940 , C0 , C0 , n52938 , n52939 );
and ( n52941 , n52940 , n21330 );
and ( n52942 , n18521 , n21338 );
or ( n52943 , n52941 , n52942 );
and ( n52944 , n52943 , n21341 );
and ( n52945 , n18521 , n21338 );
buf ( n52946 , n52945 );
and ( n52947 , n52946 , n23064 );
and ( n52948 , n18521 , n21338 );
buf ( n52949 , n52948 );
and ( n52950 , n52949 , n23825 );
and ( n52951 , n21841 , n21330 );
and ( n52952 , n18521 , n21338 );
or ( n52953 , n52951 , n52952 );
and ( n52954 , n52953 , n23832 );
buf ( n52955 , n21841 );
not ( n52956 , n52955 );
and ( n52957 , n40122 , n40132 );
xor ( n52958 , n52956 , n52957 );
buf ( n52959 , n52958 );
and ( n52960 , n52959 , n21330 );
and ( n52961 , n18521 , n21338 );
or ( n52962 , n52960 , n52961 );
and ( n52963 , n52962 , n23917 );
or ( n52964 , n52934 , n52944 , n52947 , n52950 , n52954 , C0 , n52963 );
and ( n52965 , n52933 , n52964 );
and ( n52966 , n18521 , n17451 );
or ( n52967 , n52965 , n52966 );
and ( n52968 , n52967 , n23924 );
and ( n52969 , n18521 , n23926 );
or ( n52970 , n52968 , n52969 );
buf ( n52971 , n52970 );
buf ( n52972 , n52971 );
not ( n52973 , n24800 );
and ( n52974 , n26495 , n25222 );
and ( n52975 , n47500 , n28583 );
and ( n52976 , n26495 , n28591 );
or ( n52977 , n52975 , n52976 );
and ( n52978 , n52977 , n28594 );
and ( n52979 , n47510 , n28583 );
and ( n52980 , n26495 , n28591 );
or ( n52981 , n52979 , n52980 );
and ( n52982 , n52981 , n30269 );
and ( n52983 , n47520 , n28583 );
and ( n52984 , n26495 , n28591 );
or ( n52985 , n52983 , n52984 );
and ( n52986 , n52985 , n30982 );
and ( n52987 , n29295 , n28583 );
and ( n52988 , n26495 , n28591 );
or ( n52989 , n52987 , n52988 );
and ( n52990 , n52989 , n30989 );
and ( n52991 , n26493 , n30991 );
and ( n52992 , n47531 , n28583 );
and ( n52993 , n26495 , n28591 );
or ( n52994 , n52992 , n52993 );
and ( n52995 , n52994 , n31002 );
or ( n52996 , n52974 , n52978 , n52982 , n52986 , n52990 , n52991 , n52995 );
and ( n52997 , n52973 , n52996 );
and ( n52998 , n26495 , n24800 );
or ( n52999 , n52997 , n52998 );
and ( n53000 , n52999 , n31008 );
and ( n53001 , n26495 , n10618 );
or ( n53002 , n53000 , n53001 );
buf ( n53003 , n53002 );
buf ( n53004 , n53003 );
buf ( n53005 , n10615 );
buf ( n53006 , n10613 );
and ( n53007 , n16849 , n23924 );
and ( n53008 , n22273 , n23926 );
or ( n53009 , n53007 , n53008 );
buf ( n53010 , n53009 );
buf ( n53011 , n53010 );
and ( n53012 , n11689 , n16574 );
and ( n53013 , n15836 , n16576 );
or ( n53014 , n53012 , n53013 );
buf ( n53015 , n53014 );
buf ( n53016 , n53015 );
buf ( n53017 , n10613 );
not ( n53018 , n17451 );
and ( n53019 , n18909 , n17873 );
and ( n53020 , n43338 , n21330 );
and ( n53021 , n18909 , n21338 );
or ( n53022 , n53020 , n53021 );
and ( n53023 , n53022 , n21341 );
and ( n53024 , n43348 , n21330 );
and ( n53025 , n18909 , n21338 );
or ( n53026 , n53024 , n53025 );
and ( n53027 , n53026 , n23064 );
and ( n53028 , n43358 , n21330 );
and ( n53029 , n18909 , n21338 );
or ( n53030 , n53028 , n53029 );
and ( n53031 , n53030 , n23825 );
and ( n53032 , n22182 , n21330 );
and ( n53033 , n18909 , n21338 );
or ( n53034 , n53032 , n53033 );
and ( n53035 , n53034 , n23832 );
and ( n53036 , n18907 , n23834 );
and ( n53037 , n43368 , n21330 );
and ( n53038 , n18909 , n21338 );
or ( n53039 , n53037 , n53038 );
and ( n53040 , n53039 , n23917 );
or ( n53041 , n53019 , n53023 , n53027 , n53031 , n53035 , n53036 , n53040 );
and ( n53042 , n53018 , n53041 );
and ( n53043 , n18909 , n17451 );
or ( n53044 , n53042 , n53043 );
and ( n53045 , n53044 , n23924 );
and ( n53046 , n18909 , n23926 );
or ( n53047 , n53045 , n53046 );
buf ( n53048 , n53047 );
buf ( n53049 , n53048 );
buf ( n53050 , n10613 );
not ( n53051 , n17451 );
and ( n53052 , n47430 , n21333 );
and ( n53053 , n19251 , n34758 );
or ( n53054 , n53052 , n53053 );
and ( n53055 , n53054 , n21341 );
and ( n53056 , n47440 , n21333 );
and ( n53057 , n19251 , n34758 );
or ( n53058 , n53056 , n53057 );
and ( n53059 , n53058 , n23064 );
and ( n53060 , n47450 , n21333 );
and ( n53061 , n19251 , n34758 );
or ( n53062 , n53060 , n53061 );
and ( n53063 , n53062 , n23825 );
and ( n53064 , n21958 , n21333 );
and ( n53065 , n19251 , n34758 );
or ( n53066 , n53064 , n53065 );
and ( n53067 , n53066 , n23832 );
and ( n53068 , n47461 , n21333 );
and ( n53069 , n19251 , n34758 );
or ( n53070 , n53068 , n53069 );
and ( n53071 , n53070 , n23917 );
and ( n53072 , n19251 , n34526 );
or ( n53073 , n53055 , n53059 , n53063 , n53067 , n53071 , n53072 );
and ( n53074 , n53051 , n53073 );
and ( n53075 , n19251 , n17451 );
or ( n53076 , n53074 , n53075 );
and ( n53077 , n53076 , n23924 );
and ( n53078 , n19251 , n23926 );
or ( n53079 , n53077 , n53078 );
buf ( n53080 , n53079 );
buf ( n53081 , n53080 );
buf ( n53082 , n10613 );
not ( n53083 , n34538 );
and ( n53084 , n53083 , n18527 );
and ( n53085 , n14645 , n34538 );
or ( n53086 , n53084 , n53085 );
and ( n53087 , n53086 , n23924 );
and ( n53088 , n14645 , n23926 );
or ( n53089 , n53087 , n53088 );
buf ( n53090 , n53089 );
buf ( n53091 , n53090 );
buf ( n53092 , n10613 );
buf ( n53093 , n10615 );
and ( n53094 , n16745 , n23924 );
and ( n53095 , n21982 , n23926 );
or ( n53096 , n53094 , n53095 );
buf ( n53097 , n53096 );
buf ( n53098 , n53097 );
buf ( n53099 , n10615 );
buf ( n53100 , n10613 );
buf ( n53101 , n10615 );
not ( n53102 , n11954 );
not ( n53103 , n12243 );
and ( n53104 , n10941 , n31187 );
not ( n53105 , n31697 );
and ( n53106 , n53105 , n31387 );
xor ( n53107 , n50365 , n50366 );
and ( n53108 , n53107 , n31697 );
or ( n53109 , n53106 , n53108 );
buf ( n53110 , n53109 );
and ( n53111 , n53110 , n14140 );
not ( n53112 , n32214 );
and ( n53113 , n53112 , n31904 );
xor ( n53114 , n50392 , n50393 );
and ( n53115 , n53114 , n32214 );
or ( n53116 , n53113 , n53115 );
buf ( n53117 , n53116 );
and ( n53118 , n53117 , n14137 );
and ( n53119 , n15843 , n14143 );
and ( n53120 , n10941 , n14141 );
or ( n53121 , n53111 , n53118 , n53119 , n53120 );
and ( n53122 , n53121 , n32236 );
or ( n53123 , n53104 , n53122 );
and ( n53124 , n53103 , n53123 );
not ( n53125 , n34038 );
and ( n53126 , n53125 , n33602 );
xor ( n53127 , n50425 , n50426 );
and ( n53128 , n53127 , n34038 );
or ( n53129 , n53126 , n53128 );
buf ( n53130 , n53129 );
and ( n53131 , n53130 , n12243 );
or ( n53132 , n53124 , n53131 );
and ( n53133 , n53102 , n53132 );
and ( n53134 , n53121 , n11954 );
or ( n53135 , n53133 , n53134 );
and ( n53136 , n53135 , n16574 );
not ( n53137 , n34327 );
and ( n53138 , n53137 , n34071 );
xor ( n53139 , n50457 , n50458 );
and ( n53140 , n53139 , n34327 );
or ( n53141 , n53138 , n53140 );
buf ( n53142 , n53141 );
and ( n53143 , n53142 , n16576 );
or ( n53144 , n53136 , n53143 );
buf ( n53145 , n53144 );
buf ( n53146 , n53145 );
and ( n53147 , n16737 , n23924 );
and ( n53148 , n21969 , n23926 );
or ( n53149 , n53147 , n53148 );
buf ( n53150 , n53149 );
buf ( n53151 , n53150 );
not ( n53152 , n24800 );
and ( n53153 , n28510 , n28586 );
and ( n53154 , n25890 , n34573 );
or ( n53155 , n53153 , n53154 );
and ( n53156 , n53155 , n28594 );
and ( n53157 , n30258 , n28586 );
and ( n53158 , n25890 , n34573 );
or ( n53159 , n53157 , n53158 );
and ( n53160 , n53159 , n30269 );
and ( n53161 , n30972 , n28586 );
and ( n53162 , n25890 , n34573 );
or ( n53163 , n53161 , n53162 );
and ( n53164 , n53163 , n30982 );
and ( n53165 , n29655 , n28586 );
and ( n53166 , n25890 , n34573 );
or ( n53167 , n53165 , n53166 );
and ( n53168 , n53167 , n30989 );
and ( n53169 , n30998 , n28586 );
and ( n53170 , n25890 , n34573 );
or ( n53171 , n53169 , n53170 );
and ( n53172 , n53171 , n31002 );
and ( n53173 , n25890 , n34607 );
or ( n53174 , n53156 , n53160 , n53164 , n53168 , n53172 , n53173 );
and ( n53175 , n53152 , n53174 );
and ( n53176 , n25890 , n24800 );
or ( n53177 , n53175 , n53176 );
and ( n53178 , n53177 , n31008 );
and ( n53179 , n25890 , n10618 );
or ( n53180 , n53178 , n53179 );
buf ( n53181 , n53180 );
buf ( n53182 , n53181 );
buf ( n53183 , n10613 );
not ( n53184 , n17451 );
and ( n53185 , n40081 , n21334 );
and ( n53186 , n20482 , n34492 );
or ( n53187 , n53185 , n53186 );
and ( n53188 , n53187 , n21341 );
and ( n53189 , n40096 , n21334 );
and ( n53190 , n20482 , n34492 );
or ( n53191 , n53189 , n53190 );
and ( n53192 , n53191 , n23064 );
and ( n53193 , n40111 , n21334 );
and ( n53194 , n20482 , n34492 );
or ( n53195 , n53193 , n53194 );
and ( n53196 , n53195 , n23825 );
and ( n53197 , n21854 , n21334 );
and ( n53198 , n20482 , n34492 );
or ( n53199 , n53197 , n53198 );
and ( n53200 , n53199 , n23832 );
and ( n53201 , n40134 , n21334 );
and ( n53202 , n20482 , n34492 );
or ( n53203 , n53201 , n53202 );
and ( n53204 , n53203 , n23917 );
and ( n53205 , n20482 , n34526 );
or ( n53206 , n53188 , n53192 , n53196 , n53200 , n53204 , n53205 );
and ( n53207 , n53184 , n53206 );
and ( n53208 , n20482 , n17451 );
or ( n53209 , n53207 , n53208 );
and ( n53210 , n53209 , n23924 );
and ( n53211 , n20482 , n23926 );
or ( n53212 , n53210 , n53211 );
buf ( n53213 , n53212 );
buf ( n53214 , n53213 );
and ( n53215 , n24365 , n31008 );
and ( n53216 , n29170 , n10618 );
or ( n53217 , n53215 , n53216 );
buf ( n53218 , n53217 );
buf ( n53219 , n53218 );
buf ( n53220 , n10615 );
not ( n53221 , n17451 );
and ( n53222 , n21257 , n21333 );
and ( n53223 , n19352 , n34758 );
or ( n53224 , n53222 , n53223 );
and ( n53225 , n53224 , n21341 );
and ( n53226 , n23053 , n21333 );
and ( n53227 , n19352 , n34758 );
or ( n53228 , n53226 , n53227 );
and ( n53229 , n53228 , n23064 );
and ( n53230 , n23815 , n21333 );
and ( n53231 , n19352 , n34758 );
or ( n53232 , n53230 , n53231 );
and ( n53233 , n53232 , n23825 );
and ( n53234 , n21919 , n21333 );
and ( n53235 , n19352 , n34758 );
or ( n53236 , n53234 , n53235 );
and ( n53237 , n53236 , n23832 );
and ( n53238 , n23913 , n21333 );
and ( n53239 , n19352 , n34758 );
or ( n53240 , n53238 , n53239 );
and ( n53241 , n53240 , n23917 );
and ( n53242 , n19352 , n34526 );
or ( n53243 , n53225 , n53229 , n53233 , n53237 , n53241 , n53242 );
and ( n53244 , n53221 , n53243 );
and ( n53245 , n19352 , n17451 );
or ( n53246 , n53244 , n53245 );
and ( n53247 , n53246 , n23924 );
and ( n53248 , n19352 , n23926 );
or ( n53249 , n53247 , n53248 );
buf ( n53250 , n53249 );
buf ( n53251 , n53250 );
not ( n53252 , n34804 );
and ( n53253 , n53252 , n26161 );
and ( n53254 , n14779 , n34804 );
or ( n53255 , n53253 , n53254 );
and ( n53256 , n53255 , n31008 );
and ( n53257 , n14779 , n10618 );
or ( n53258 , n53256 , n53257 );
buf ( n53259 , n53258 );
buf ( n53260 , n53259 );
buf ( n53261 , n10615 );
buf ( n53262 , n10615 );
not ( n53263 , n34821 );
and ( n53264 , n13275 , n14592 );
and ( n53265 , n46158 , n36350 );
and ( n53266 , n13275 , n43691 );
or ( n53267 , n53265 , n53266 );
and ( n53268 , n53267 , n14562 );
and ( n53269 , n46168 , n36350 );
and ( n53270 , n13275 , n43703 );
or ( n53271 , n53269 , n53270 );
and ( n53272 , n53271 , n14586 );
and ( n53273 , n46178 , n36345 );
and ( n53274 , n13275 , n43715 );
or ( n53275 , n53273 , n53274 );
and ( n53276 , n53275 , n14584 );
and ( n53277 , n46168 , n36345 );
and ( n53278 , n13275 , n43721 );
or ( n53279 , n53277 , n53278 );
and ( n53280 , n53279 , n37835 );
and ( n53281 , n46178 , n36345 );
and ( n53282 , n13275 , n43721 );
or ( n53283 , n53281 , n53282 );
and ( n53284 , n53283 , n37841 );
and ( n53285 , n15471 , n14564 );
and ( n53286 , n15471 , n36345 );
and ( n53287 , n13275 , n43721 );
or ( n53288 , n53286 , n53287 );
and ( n53289 , n53288 , n37847 );
or ( n53290 , n53264 , n53268 , n53272 , n53276 , n53280 , n53284 , n53285 , n53289 );
and ( n53291 , n53263 , n53290 );
and ( n53292 , n13275 , n34821 );
or ( n53293 , n53291 , n53292 );
and ( n53294 , n53293 , n16574 );
and ( n53295 , n12279 , n16576 );
or ( n53296 , n53294 , n53295 );
buf ( n53297 , n53296 );
buf ( n53298 , n53297 );
buf ( n53299 , n10615 );
not ( n53300 , n17451 );
and ( n53301 , n18569 , n17873 );
and ( n53302 , n50716 , n21336 );
and ( n53303 , n18569 , n42682 );
or ( n53304 , n53302 , n53303 );
and ( n53305 , n53304 , n21341 );
and ( n53306 , n50726 , n21336 );
and ( n53307 , n18569 , n42682 );
or ( n53308 , n53306 , n53307 );
and ( n53309 , n53308 , n23064 );
and ( n53310 , n50736 , n21336 );
and ( n53311 , n18569 , n42682 );
or ( n53312 , n53310 , n53311 );
and ( n53313 , n53312 , n23825 );
and ( n53314 , n22382 , n21336 );
and ( n53315 , n18569 , n42682 );
or ( n53316 , n53314 , n53315 );
and ( n53317 , n53316 , n23832 );
and ( n53318 , n22382 , n23834 );
and ( n53319 , n50747 , n21336 );
and ( n53320 , n18569 , n42682 );
or ( n53321 , n53319 , n53320 );
and ( n53322 , n53321 , n23917 );
or ( n53323 , n53301 , n53305 , n53309 , n53313 , n53317 , n53318 , n53322 );
and ( n53324 , n53300 , n53323 );
and ( n53325 , n18569 , n17451 );
or ( n53326 , n53324 , n53325 );
and ( n53327 , n53326 , n23924 );
and ( n53328 , n17900 , n23926 );
or ( n53329 , n53327 , n53328 );
buf ( n53330 , n53329 );
buf ( n53331 , n53330 );
buf ( n53332 , n10613 );
buf ( n53333 , n10615 );
not ( n53334 , n17451 );
and ( n53335 , n48266 , n21334 );
and ( n53336 , n19422 , n34492 );
or ( n53337 , n53335 , n53336 );
and ( n53338 , n53337 , n21341 );
and ( n53339 , n48276 , n21334 );
and ( n53340 , n19422 , n34492 );
or ( n53341 , n53339 , n53340 );
and ( n53342 , n53341 , n23064 );
and ( n53343 , n48286 , n21334 );
and ( n53344 , n19422 , n34492 );
or ( n53345 , n53343 , n53344 );
and ( n53346 , n53345 , n23825 );
and ( n53347 , n21893 , n21334 );
and ( n53348 , n19422 , n34492 );
or ( n53349 , n53347 , n53348 );
and ( n53350 , n53349 , n23832 );
and ( n53351 , n48297 , n21334 );
and ( n53352 , n19422 , n34492 );
or ( n53353 , n53351 , n53352 );
and ( n53354 , n53353 , n23917 );
and ( n53355 , n19422 , n34526 );
or ( n53356 , n53338 , n53342 , n53346 , n53350 , n53354 , n53355 );
and ( n53357 , n53334 , n53356 );
and ( n53358 , n19422 , n17451 );
or ( n53359 , n53357 , n53358 );
and ( n53360 , n53359 , n23924 );
and ( n53361 , n19422 , n23926 );
or ( n53362 , n53360 , n53361 );
buf ( n53363 , n53362 );
buf ( n53364 , n53363 );
buf ( n53365 , n10613 );
buf ( n53366 , n10615 );
buf ( n53367 , n10613 );
not ( n53368 , n34821 );
and ( n53369 , n44916 , n36347 );
and ( n53370 , n13387 , n39408 );
or ( n53371 , n53369 , n53370 );
and ( n53372 , n53371 , n14562 );
and ( n53373 , n44926 , n36348 );
and ( n53374 , n13387 , n39427 );
or ( n53375 , n53373 , n53374 );
and ( n53376 , n53375 , n14586 );
and ( n53377 , n44936 , n36347 );
and ( n53378 , n13387 , n39446 );
or ( n53379 , n53377 , n53378 );
and ( n53380 , n53379 , n14584 );
and ( n53381 , n44926 , n36348 );
and ( n53382 , n13387 , n39453 );
or ( n53383 , n53381 , n53382 );
and ( n53384 , n53383 , n37835 );
and ( n53385 , n44936 , n36348 );
and ( n53386 , n13387 , n39453 );
or ( n53387 , n53385 , n53386 );
and ( n53388 , n53387 , n37841 );
and ( n53389 , n15669 , n36348 );
and ( n53390 , n13387 , n39453 );
or ( n53391 , n53389 , n53390 );
and ( n53392 , n53391 , n37847 );
and ( n53393 , n13387 , n37849 );
or ( n53394 , n53372 , n53376 , n53380 , n53384 , n53388 , n53392 , n53393 );
and ( n53395 , n53368 , n53394 );
and ( n53396 , n13387 , n34821 );
or ( n53397 , n53395 , n53396 );
and ( n53398 , n53397 , n16574 );
and ( n53399 , n13387 , n16576 );
or ( n53400 , n53398 , n53399 );
buf ( n53401 , n53400 );
buf ( n53402 , n53401 );
not ( n53403 , n34538 );
and ( n53404 , n53403 , n18514 );
and ( n53405 , n14831 , n34538 );
or ( n53406 , n53404 , n53405 );
and ( n53407 , n53406 , n23924 );
and ( n53408 , n14831 , n23926 );
or ( n53409 , n53407 , n53408 );
buf ( n53410 , n53409 );
buf ( n53411 , n53410 );
buf ( n53412 , n10615 );
and ( n53413 , n11673 , n16574 );
and ( n53414 , n15792 , n16576 );
or ( n53415 , n53413 , n53414 );
buf ( n53416 , n53415 );
buf ( n53417 , n53416 );
not ( n53418 , n17162 );
not ( n53419 , n17450 );
and ( n53420 , n10663 , n37947 );
not ( n53421 , n38425 );
and ( n53422 , n53421 , n38336 );
xor ( n53423 , n46212 , n46215 );
and ( n53424 , n53423 , n38425 );
or ( n53425 , n53422 , n53424 );
buf ( n53426 , n53425 );
and ( n53427 , n53426 , n19745 );
not ( n53428 , n38934 );
and ( n53429 , n53428 , n38845 );
xor ( n53430 , n46225 , n46228 );
and ( n53431 , n53430 , n38934 );
or ( n53432 , n53429 , n53431 );
buf ( n53433 , n53432 );
and ( n53434 , n53433 , n19748 );
and ( n53435 , n22140 , n21253 );
and ( n53436 , n10663 , n21255 );
or ( n53437 , n53427 , n53434 , n53435 , n53436 );
and ( n53438 , n53437 , n38980 );
or ( n53439 , n53420 , n53438 );
and ( n53440 , n53419 , n53439 );
or ( n53441 , n53440 , C0 );
and ( n53442 , n53418 , n53441 );
and ( n53443 , n53437 , n17162 );
or ( n53444 , n53442 , n53443 );
and ( n53445 , n53444 , n23924 );
not ( n53446 , n39264 );
and ( n53447 , n53446 , n39190 );
xor ( n53448 , n46249 , n46252 );
and ( n53449 , n53448 , n39264 );
or ( n53450 , n53447 , n53449 );
buf ( n53451 , n53450 );
and ( n53452 , n53451 , n23926 );
or ( n53453 , n53445 , n53452 );
buf ( n53454 , n53453 );
buf ( n53455 , n53454 );
not ( n53456 , n24800 );
and ( n53457 , n49354 , n28587 );
and ( n53458 , n26057 , n39807 );
or ( n53459 , n53457 , n53458 );
and ( n53460 , n53459 , n28594 );
and ( n53461 , n49364 , n28587 );
and ( n53462 , n26057 , n39807 );
or ( n53463 , n53461 , n53462 );
and ( n53464 , n53463 , n30269 );
and ( n53465 , n49374 , n28587 );
and ( n53466 , n26057 , n39807 );
or ( n53467 , n53465 , n53466 );
and ( n53468 , n53467 , n30982 );
and ( n53469 , n29555 , n28587 );
and ( n53470 , n26057 , n39807 );
or ( n53471 , n53469 , n53470 );
and ( n53472 , n53471 , n30989 );
and ( n53473 , n49385 , n28587 );
and ( n53474 , n26057 , n39807 );
or ( n53475 , n53473 , n53474 );
and ( n53476 , n53475 , n31002 );
and ( n53477 , n26057 , n34607 );
or ( n53478 , n53460 , n53464 , n53468 , n53472 , n53476 , n53477 );
and ( n53479 , n53456 , n53478 );
and ( n53480 , n26057 , n24800 );
or ( n53481 , n53479 , n53480 );
and ( n53482 , n53481 , n31008 );
and ( n53483 , n26057 , n10618 );
or ( n53484 , n53482 , n53483 );
buf ( n53485 , n53484 );
buf ( n53486 , n53485 );
not ( n53487 , n17451 );
and ( n53488 , n46077 , n21334 );
and ( n53489 , n19185 , n34492 );
or ( n53490 , n53488 , n53489 );
and ( n53491 , n53490 , n21341 );
and ( n53492 , n46087 , n21334 );
and ( n53493 , n19185 , n34492 );
or ( n53494 , n53492 , n53493 );
and ( n53495 , n53494 , n23064 );
and ( n53496 , n46097 , n21334 );
and ( n53497 , n19185 , n34492 );
or ( n53498 , n53496 , n53497 );
and ( n53499 , n53498 , n23825 );
and ( n53500 , n21984 , n21334 );
and ( n53501 , n19185 , n34492 );
or ( n53502 , n53500 , n53501 );
and ( n53503 , n53502 , n23832 );
and ( n53504 , n46108 , n21334 );
and ( n53505 , n19185 , n34492 );
or ( n53506 , n53504 , n53505 );
and ( n53507 , n53506 , n23917 );
and ( n53508 , n19185 , n34526 );
or ( n53509 , n53491 , n53495 , n53499 , n53503 , n53507 , n53508 );
and ( n53510 , n53487 , n53509 );
and ( n53511 , n19185 , n17451 );
or ( n53512 , n53510 , n53511 );
and ( n53513 , n53512 , n23924 );
and ( n53514 , n19185 , n23926 );
or ( n53515 , n53513 , n53514 );
buf ( n53516 , n53515 );
buf ( n53517 , n53516 );
not ( n53518 , n17451 );
and ( n53519 , n50716 , n21334 );
and ( n53520 , n18575 , n34492 );
or ( n53521 , n53519 , n53520 );
and ( n53522 , n53521 , n21341 );
and ( n53523 , n50726 , n21334 );
and ( n53524 , n18575 , n34492 );
or ( n53525 , n53523 , n53524 );
and ( n53526 , n53525 , n23064 );
and ( n53527 , n50736 , n21334 );
and ( n53528 , n18575 , n34492 );
or ( n53529 , n53527 , n53528 );
and ( n53530 , n53529 , n23825 );
and ( n53531 , n22382 , n21334 );
and ( n53532 , n18575 , n34492 );
or ( n53533 , n53531 , n53532 );
and ( n53534 , n53533 , n23832 );
and ( n53535 , n50747 , n21334 );
and ( n53536 , n18575 , n34492 );
or ( n53537 , n53535 , n53536 );
and ( n53538 , n53537 , n23917 );
and ( n53539 , n18575 , n34526 );
or ( n53540 , n53522 , n53526 , n53530 , n53534 , n53538 , n53539 );
and ( n53541 , n53518 , n53540 );
and ( n53542 , n18575 , n17451 );
or ( n53543 , n53541 , n53542 );
and ( n53544 , n53543 , n23924 );
and ( n53545 , n18575 , n23926 );
or ( n53546 , n53544 , n53545 );
buf ( n53547 , n53546 );
buf ( n53548 , n53547 );
buf ( n53549 , n10613 );
not ( n53550 , n24800 );
and ( n53551 , n48334 , n28586 );
and ( n53552 , n25954 , n34573 );
or ( n53553 , n53551 , n53552 );
and ( n53554 , n53553 , n28594 );
and ( n53555 , n48344 , n28586 );
and ( n53556 , n25954 , n34573 );
or ( n53557 , n53555 , n53556 );
and ( n53558 , n53557 , n30269 );
and ( n53559 , n48354 , n28586 );
and ( n53560 , n25954 , n34573 );
or ( n53561 , n53559 , n53560 );
and ( n53562 , n53561 , n30982 );
and ( n53563 , n29615 , n28586 );
and ( n53564 , n25954 , n34573 );
or ( n53565 , n53563 , n53564 );
and ( n53566 , n53565 , n30989 );
and ( n53567 , n48364 , n28586 );
and ( n53568 , n25954 , n34573 );
or ( n53569 , n53567 , n53568 );
and ( n53570 , n53569 , n31002 );
and ( n53571 , n25954 , n34607 );
or ( n53572 , n53554 , n53558 , n53562 , n53566 , n53570 , n53571 );
and ( n53573 , n53550 , n53572 );
and ( n53574 , n25954 , n24800 );
or ( n53575 , n53573 , n53574 );
and ( n53576 , n53575 , n31008 );
and ( n53577 , n25954 , n10618 );
or ( n53578 , n53576 , n53577 );
buf ( n53579 , n53578 );
buf ( n53580 , n53579 );
and ( n53581 , n11521 , n16574 );
and ( n53582 , n15080 , n16576 );
or ( n53583 , n53581 , n53582 );
buf ( n53584 , n53583 );
buf ( n53585 , n53584 );
buf ( n53586 , n10615 );
and ( n53587 , n11692 , n16574 );
and ( n53588 , n15857 , n16576 );
or ( n53589 , n53587 , n53588 );
buf ( n53590 , n53589 );
buf ( n53591 , n53590 );
not ( n53592 , n24800 );
and ( n53593 , n26223 , n25222 );
not ( n53594 , n26823 );
and ( n53595 , n53594 , n26207 );
xor ( n53596 , n34625 , n34626 );
and ( n53597 , n53596 , n26823 );
or ( n53598 , n53595 , n53597 );
buf ( n53599 , n53598 );
and ( n53600 , n53599 , n27046 );
and ( n53601 , n53599 , n27049 );
not ( n53602 , n27051 );
and ( n53603 , n53602 , n28104 );
not ( n53604 , n28494 );
and ( n53605 , n53604 , n28116 );
xor ( n53606 , n34643 , n34644 );
and ( n53607 , n53606 , n28494 );
or ( n53608 , n53605 , n53607 );
buf ( n53609 , n53608 );
and ( n53610 , n53609 , n27051 );
or ( n53611 , n53603 , n53610 );
and ( n53612 , n53611 , n28506 );
and ( n53613 , n28104 , n28508 );
or ( n53614 , n53600 , n53601 , n53612 , n53613 );
and ( n53615 , n53614 , n28583 );
and ( n53616 , n26223 , n28591 );
or ( n53617 , n53615 , n53616 );
and ( n53618 , n53617 , n28594 );
not ( n53619 , n30249 );
and ( n53620 , n53619 , n29939 );
xor ( n53621 , n34666 , n34667 );
and ( n53622 , n53621 , n30249 );
or ( n53623 , n53620 , n53622 );
buf ( n53624 , n53623 );
and ( n53625 , n53624 , n28583 );
and ( n53626 , n26223 , n28591 );
or ( n53627 , n53625 , n53626 );
and ( n53628 , n53627 , n30269 );
not ( n53629 , n30963 );
and ( n53630 , n53629 , n30653 );
xor ( n53631 , n34684 , n34685 );
and ( n53632 , n53631 , n30963 );
or ( n53633 , n53630 , n53632 );
buf ( n53634 , n53633 );
and ( n53635 , n53634 , n28583 );
and ( n53636 , n26223 , n28591 );
or ( n53637 , n53635 , n53636 );
and ( n53638 , n53637 , n30982 );
and ( n53639 , n29455 , n28583 );
and ( n53640 , n26223 , n28591 );
or ( n53641 , n53639 , n53640 );
and ( n53642 , n53641 , n30989 );
and ( n53643 , n26221 , n30991 );
xor ( n53644 , n34708 , n34709 );
buf ( n53645 , n53644 );
and ( n53646 , n53645 , n28583 );
and ( n53647 , n26223 , n28591 );
or ( n53648 , n53646 , n53647 );
and ( n53649 , n53648 , n31002 );
or ( n53650 , n53593 , n53618 , n53628 , n53638 , n53642 , n53643 , n53649 );
and ( n53651 , n53592 , n53650 );
and ( n53652 , n26223 , n24800 );
or ( n53653 , n53651 , n53652 );
and ( n53654 , n53653 , n31008 );
and ( n53655 , n26223 , n10618 );
or ( n53656 , n53654 , n53655 );
buf ( n53657 , n53656 );
buf ( n53658 , n53657 );
not ( n53659 , n24800 );
and ( n53660 , n26529 , n25222 );
and ( n53661 , n52878 , n28583 );
and ( n53662 , n26529 , n28591 );
or ( n53663 , n53661 , n53662 );
and ( n53664 , n53663 , n28594 );
and ( n53665 , n52888 , n28583 );
and ( n53666 , n26529 , n28591 );
or ( n53667 , n53665 , n53666 );
and ( n53668 , n53667 , n30269 );
and ( n53669 , n52898 , n28583 );
and ( n53670 , n26529 , n28591 );
or ( n53671 , n53669 , n53670 );
and ( n53672 , n53671 , n30982 );
and ( n53673 , n29237 , n28583 );
and ( n53674 , n26529 , n28591 );
or ( n53675 , n53673 , n53674 );
and ( n53676 , n53675 , n30989 );
and ( n53677 , n26527 , n30991 );
and ( n53678 , n52908 , n28583 );
and ( n53679 , n26529 , n28591 );
or ( n53680 , n53678 , n53679 );
and ( n53681 , n53680 , n31002 );
or ( n53682 , n53660 , n53664 , n53668 , n53672 , n53676 , n53677 , n53681 );
and ( n53683 , n53659 , n53682 );
and ( n53684 , n26529 , n24800 );
or ( n53685 , n53683 , n53684 );
and ( n53686 , n53685 , n31008 );
and ( n53687 , n26529 , n10618 );
or ( n53688 , n53686 , n53687 );
buf ( n53689 , n53688 );
buf ( n53690 , n53689 );
not ( n53691 , n34821 );
not ( n53692 , n13916 );
and ( n53693 , n53692 , n13639 );
xor ( n53694 , n13640 , n13875 );
and ( n53695 , n53694 , n13916 );
or ( n53696 , n53693 , n53695 );
buf ( n53697 , n53696 );
and ( n53698 , n53697 , n14137 );
and ( n53699 , n53697 , n14143 );
not ( n53700 , n14139 );
and ( n53701 , n53700 , n36075 );
not ( n53702 , n36245 );
and ( n53703 , n53702 , n36087 );
xor ( n53704 , n45733 , n45736 );
and ( n53705 , n53704 , n36245 );
or ( n53706 , n53703 , n53705 );
buf ( n53707 , n53706 );
and ( n53708 , n53707 , n14139 );
or ( n53709 , n53701 , n53708 );
and ( n53710 , n53709 , n14140 );
and ( n53711 , n36075 , n14141 );
or ( n53712 , n53698 , n53699 , n53710 , n53711 );
and ( n53713 , n53712 , n36347 );
and ( n53714 , n13243 , n39408 );
or ( n53715 , n53713 , n53714 );
and ( n53716 , n53715 , n14562 );
not ( n53717 , n37048 );
and ( n53718 , n53717 , n36908 );
xor ( n53719 , n45754 , n45757 );
and ( n53720 , n53719 , n37048 );
or ( n53721 , n53718 , n53720 );
buf ( n53722 , n53721 );
and ( n53723 , n53722 , n36348 );
and ( n53724 , n13243 , n39427 );
or ( n53725 , n53723 , n53724 );
and ( n53726 , n53725 , n14586 );
not ( n53727 , n37801 );
and ( n53728 , n53727 , n37661 );
xor ( n53729 , n45770 , n45773 );
and ( n53730 , n53729 , n37801 );
or ( n53731 , n53728 , n53730 );
buf ( n53732 , n53731 );
and ( n53733 , n53732 , n36347 );
and ( n53734 , n13243 , n39446 );
or ( n53735 , n53733 , n53734 );
and ( n53736 , n53735 , n14584 );
and ( n53737 , n53722 , n36348 );
and ( n53738 , n13243 , n39453 );
or ( n53739 , n53737 , n53738 );
and ( n53740 , n53739 , n37835 );
and ( n53741 , n53732 , n36348 );
and ( n53742 , n13243 , n39453 );
or ( n53743 , n53741 , n53742 );
and ( n53744 , n53743 , n37841 );
and ( n53745 , n15097 , n36348 );
and ( n53746 , n13243 , n39453 );
or ( n53747 , n53745 , n53746 );
and ( n53748 , n53747 , n37847 );
and ( n53749 , n13243 , n37849 );
or ( n53750 , n53716 , n53726 , n53736 , n53740 , n53744 , n53748 , n53749 );
and ( n53751 , n53691 , n53750 );
and ( n53752 , n13243 , n34821 );
or ( n53753 , n53751 , n53752 );
and ( n53754 , n53753 , n16574 );
and ( n53755 , n13243 , n16576 );
or ( n53756 , n53754 , n53755 );
buf ( n53757 , n53756 );
buf ( n53758 , n53757 );
not ( n53759 , n34821 );
not ( n53760 , n14139 );
and ( n53761 , n53760 , n35190 );
not ( n53762 , n36245 );
and ( n53763 , n53762 , n35196 );
xor ( n53764 , n36255 , n35634 );
and ( n53765 , n53764 , n36245 );
or ( n53766 , n53763 , n53765 );
buf ( n53767 , n53766 );
and ( n53768 , n53767 , n14139 );
or ( n53769 , n53761 , n53768 );
and ( n53770 , n53769 , n14140 );
and ( n53771 , n35190 , n14141 );
or ( n53772 , C0 , C0 , n53770 , n53771 );
and ( n53773 , n53772 , n36345 );
and ( n53774 , n13512 , n36352 );
or ( n53775 , n53773 , n53774 );
and ( n53776 , n53775 , n14562 );
not ( n53777 , n37048 );
and ( n53778 , n53777 , n36365 );
xor ( n53779 , n37058 , n36552 );
and ( n53780 , n53779 , n37048 );
or ( n53781 , n53778 , n53780 );
buf ( n53782 , n53781 );
and ( n53783 , n53782 , n36345 );
and ( n53784 , n13512 , n37073 );
or ( n53785 , n53783 , n53784 );
and ( n53786 , n53785 , n14586 );
not ( n53787 , n37801 );
and ( n53788 , n53787 , n37086 );
xor ( n53789 , n37811 , n37305 );
and ( n53790 , n53789 , n37801 );
or ( n53791 , n53788 , n53790 );
buf ( n53792 , n53791 );
and ( n53793 , n53792 , n36350 );
and ( n53794 , n13512 , n37825 );
or ( n53795 , n53793 , n53794 );
and ( n53796 , n53795 , n14584 );
and ( n53797 , n53782 , n36350 );
and ( n53798 , n13512 , n37831 );
or ( n53799 , n53797 , n53798 );
and ( n53800 , n53799 , n37835 );
and ( n53801 , n53792 , n36350 );
and ( n53802 , n13512 , n37831 );
or ( n53803 , n53801 , n53802 );
and ( n53804 , n53803 , n37841 );
and ( n53805 , n15866 , n36350 );
and ( n53806 , n13512 , n37831 );
or ( n53807 , n53805 , n53806 );
and ( n53808 , n53807 , n37847 );
and ( n53809 , n13512 , n37849 );
or ( n53810 , n53776 , n53786 , n53796 , n53800 , n53804 , n53808 , n53809 );
and ( n53811 , n53759 , n53810 );
and ( n53812 , n13512 , n34821 );
or ( n53813 , n53811 , n53812 );
and ( n53814 , n53813 , n16574 );
and ( n53815 , n13512 , n16576 );
or ( n53816 , n53814 , n53815 );
buf ( n53817 , n53816 );
buf ( n53818 , n53817 );
buf ( n53819 , n10615 );
buf ( n53820 , n10613 );
buf ( n53821 , n10613 );
buf ( n53822 , n10615 );
buf ( n53823 , n10615 );
and ( n53824 , n11545 , n16574 );
and ( n53825 , n15125 , n16576 );
or ( n53826 , n53824 , n53825 );
buf ( n53827 , n53826 );
buf ( n53828 , n53827 );
buf ( n53829 , n10613 );
buf ( n53830 , n10613 );
not ( n53831 , n11333 );
and ( n53832 , n53831 , n11210 );
xor ( n53833 , n11339 , n11363 );
and ( n53834 , n53833 , n11333 );
or ( n53835 , n53832 , n53834 );
buf ( n53836 , n53835 );
buf ( n53837 , n53836 );
buf ( n53838 , n10615 );
buf ( n53839 , n10613 );
buf ( n53840 , n10613 );
buf ( n53841 , n10615 );
buf ( n53842 , n10613 );
buf ( n53843 , n10615 );
buf ( n53844 , n10615 );
not ( n53845 , n34804 );
and ( n53846 , n53845 , n25925 );
and ( n53847 , n14821 , n34804 );
or ( n53848 , n53846 , n53847 );
and ( n53849 , n53848 , n31008 );
and ( n53850 , n14821 , n10618 );
or ( n53851 , n53849 , n53850 );
buf ( n53852 , n53851 );
buf ( n53853 , n53852 );
buf ( n53854 , n10615 );
not ( n53855 , n11333 );
and ( n53856 , n53855 , n11312 );
xor ( n53857 , n11312 , n11007 );
and ( n53858 , n50483 , n50484 );
xor ( n53859 , n53857 , n53858 );
and ( n53860 , n53859 , n11333 );
or ( n53861 , n53856 , n53860 );
buf ( n53862 , n53861 );
buf ( n53863 , n53862 );
buf ( n53864 , n10615 );
not ( n53865 , n11954 );
buf ( n53866 , n14932 );
buf ( n53867 , n53866 );
and ( n53868 , n53867 , n32236 );
buf ( n53869 , n53868 );
not ( n53870 , n12243 );
and ( n53871 , n53869 , n53870 );
and ( n53872 , n53865 , n53871 );
and ( n53873 , n53867 , n11954 );
or ( n53874 , n53872 , n53873 );
and ( n53875 , n53874 , n16574 );
buf ( n53876 , n16576 );
or ( n53877 , n53875 , n53876 );
buf ( n53878 , n53877 );
buf ( n53879 , n53878 );
buf ( n53880 , n10615 );
not ( n53881 , n24800 );
and ( n53882 , n26391 , n25222 );
and ( n53883 , n48113 , n28589 );
and ( n53884 , n26391 , n31075 );
or ( n53885 , n53883 , n53884 );
and ( n53886 , n53885 , n28594 );
and ( n53887 , n48123 , n28589 );
and ( n53888 , n26391 , n31075 );
or ( n53889 , n53887 , n53888 );
and ( n53890 , n53889 , n30269 );
and ( n53891 , n48133 , n28589 );
and ( n53892 , n26391 , n31075 );
or ( n53893 , n53891 , n53892 );
and ( n53894 , n53893 , n30982 );
and ( n53895 , n29355 , n28589 );
and ( n53896 , n26391 , n31075 );
or ( n53897 , n53895 , n53896 );
and ( n53898 , n53897 , n30989 );
and ( n53899 , n29355 , n30991 );
and ( n53900 , n48144 , n28589 );
and ( n53901 , n26391 , n31075 );
or ( n53902 , n53900 , n53901 );
and ( n53903 , n53902 , n31002 );
or ( n53904 , n53882 , n53886 , n53890 , n53894 , n53898 , n53899 , n53903 );
and ( n53905 , n53881 , n53904 );
and ( n53906 , n26391 , n24800 );
or ( n53907 , n53905 , n53906 );
and ( n53908 , n53907 , n31008 );
and ( n53909 , n25459 , n10618 );
or ( n53910 , n53908 , n53909 );
buf ( n53911 , n53910 );
buf ( n53912 , n53911 );
not ( n53913 , n17451 );
and ( n53914 , n46607 , n21333 );
and ( n53915 , n18775 , n34758 );
or ( n53916 , n53914 , n53915 );
and ( n53917 , n53916 , n21341 );
and ( n53918 , n46617 , n21333 );
and ( n53919 , n18775 , n34758 );
or ( n53920 , n53918 , n53919 );
and ( n53921 , n53920 , n23064 );
and ( n53922 , n46627 , n21333 );
and ( n53923 , n18775 , n34758 );
or ( n53924 , n53922 , n53923 );
and ( n53925 , n53924 , n23825 );
and ( n53926 , n22262 , n21333 );
and ( n53927 , n18775 , n34758 );
or ( n53928 , n53926 , n53927 );
and ( n53929 , n53928 , n23832 );
and ( n53930 , n46638 , n21333 );
and ( n53931 , n18775 , n34758 );
or ( n53932 , n53930 , n53931 );
and ( n53933 , n53932 , n23917 );
and ( n53934 , n18775 , n34526 );
or ( n53935 , n53917 , n53921 , n53925 , n53929 , n53933 , n53934 );
and ( n53936 , n53913 , n53935 );
and ( n53937 , n18775 , n17451 );
or ( n53938 , n53936 , n53937 );
and ( n53939 , n53938 , n23924 );
and ( n53940 , n18775 , n23926 );
or ( n53941 , n53939 , n53940 );
buf ( n53942 , n53941 );
buf ( n53943 , n53942 );
and ( n53944 , n24174 , n31008 );
and ( n53945 , n29466 , n10618 );
or ( n53946 , n53944 , n53945 );
buf ( n53947 , n53946 );
buf ( n53948 , n53947 );
and ( n53949 , n16865 , n23924 );
and ( n53950 , n22313 , n23926 );
or ( n53951 , n53949 , n53950 );
buf ( n53952 , n53951 );
buf ( n53953 , n53952 );
buf ( n53954 , n10613 );
buf ( n53955 , n10613 );
and ( n53956 , n16857 , n23924 );
and ( n53957 , n22293 , n23926 );
or ( n53958 , n53956 , n53957 );
buf ( n53959 , n53958 );
buf ( n53960 , n53959 );
buf ( n53961 , n10613 );
not ( n53962 , n17451 );
and ( n53963 , n18669 , n17873 );
and ( n53964 , n48886 , n21336 );
and ( n53965 , n18669 , n42682 );
or ( n53966 , n53964 , n53965 );
and ( n53967 , n53966 , n21341 );
and ( n53968 , n48896 , n21336 );
and ( n53969 , n18669 , n42682 );
or ( n53970 , n53968 , n53969 );
and ( n53971 , n53970 , n23064 );
and ( n53972 , n48906 , n21336 );
and ( n53973 , n18669 , n42682 );
or ( n53974 , n53972 , n53973 );
and ( n53975 , n53974 , n23825 );
and ( n53976 , n22322 , n21336 );
and ( n53977 , n18669 , n42682 );
or ( n53978 , n53976 , n53977 );
and ( n53979 , n53978 , n23832 );
and ( n53980 , n22322 , n23834 );
and ( n53981 , n48916 , n21336 );
and ( n53982 , n18669 , n42682 );
or ( n53983 , n53981 , n53982 );
and ( n53984 , n53983 , n23917 );
or ( n53985 , n53963 , n53967 , n53971 , n53975 , n53979 , n53980 , n53984 );
and ( n53986 , n53962 , n53985 );
and ( n53987 , n18669 , n17451 );
or ( n53988 , n53986 , n53987 );
and ( n53989 , n53988 , n23924 );
and ( n53990 , n17945 , n23926 );
or ( n53991 , n53989 , n53990 );
buf ( n53992 , n53991 );
buf ( n53993 , n53992 );
and ( n53994 , n24094 , n31008 );
and ( n53995 , n29235 , n10618 );
or ( n53996 , n53994 , n53995 );
buf ( n53997 , n53996 );
buf ( n53998 , n53997 );
buf ( n53999 , n10615 );
buf ( n54000 , n10615 );
buf ( n54001 , n10615 );
not ( n54002 , n24800 );
and ( n54003 , n47500 , n28586 );
and ( n54004 , n26497 , n34573 );
or ( n54005 , n54003 , n54004 );
and ( n54006 , n54005 , n28594 );
and ( n54007 , n47510 , n28586 );
and ( n54008 , n26497 , n34573 );
or ( n54009 , n54007 , n54008 );
and ( n54010 , n54009 , n30269 );
and ( n54011 , n47520 , n28586 );
and ( n54012 , n26497 , n34573 );
or ( n54013 , n54011 , n54012 );
and ( n54014 , n54013 , n30982 );
and ( n54015 , n29295 , n28586 );
and ( n54016 , n26497 , n34573 );
or ( n54017 , n54015 , n54016 );
and ( n54018 , n54017 , n30989 );
and ( n54019 , n47531 , n28586 );
and ( n54020 , n26497 , n34573 );
or ( n54021 , n54019 , n54020 );
and ( n54022 , n54021 , n31002 );
and ( n54023 , n26497 , n34607 );
or ( n54024 , n54006 , n54010 , n54014 , n54018 , n54022 , n54023 );
and ( n54025 , n54002 , n54024 );
and ( n54026 , n26497 , n24800 );
or ( n54027 , n54025 , n54026 );
and ( n54028 , n54027 , n31008 );
and ( n54029 , n26497 , n10618 );
or ( n54030 , n54028 , n54029 );
buf ( n54031 , n54030 );
buf ( n54032 , n54031 );
buf ( n54033 , n10613 );
buf ( n54034 , n10615 );
and ( n54035 , n11561 , n16574 );
and ( n54036 , n15484 , n16576 );
or ( n54037 , n54035 , n54036 );
buf ( n54038 , n54037 );
buf ( n54039 , n54038 );
buf ( n54040 , n10615 );
buf ( n54041 , n10615 );
not ( n54042 , n34804 );
and ( n54043 , n54042 , n27181 );
and ( n54044 , n14653 , n34804 );
or ( n54045 , n54043 , n54044 );
and ( n54046 , n54045 , n31008 );
and ( n54047 , n14653 , n10618 );
or ( n54048 , n54046 , n54047 );
buf ( n54049 , n54048 );
buf ( n54050 , n54049 );
buf ( n54051 , n10613 );
buf ( n54052 , n10613 );
buf ( n54053 , n10615 );
buf ( n54054 , n10615 );
buf ( n54055 , n10615 );
buf ( n54056 , RI210cdf40_249);
buf ( n54057 , RI2107db58_464);
not ( n54058 , n54057 );
xor ( n54059 , n54056 , n54058 );
buf ( n54060 , RI21069950_647);
or ( n54061 , n54059 , n54060 );
buf ( n54062 , n54061 );
buf ( n54063 , n54062 );
not ( n54064 , n34821 );
and ( n54065 , n13239 , n14592 );
and ( n54066 , n53712 , n36350 );
and ( n54067 , n13239 , n43691 );
or ( n54068 , n54066 , n54067 );
and ( n54069 , n54068 , n14562 );
and ( n54070 , n53722 , n36350 );
and ( n54071 , n13239 , n43703 );
or ( n54072 , n54070 , n54071 );
and ( n54073 , n54072 , n14586 );
and ( n54074 , n53732 , n36345 );
and ( n54075 , n13239 , n43715 );
or ( n54076 , n54074 , n54075 );
and ( n54077 , n54076 , n14584 );
and ( n54078 , n53722 , n36345 );
and ( n54079 , n13239 , n43721 );
or ( n54080 , n54078 , n54079 );
and ( n54081 , n54080 , n37835 );
and ( n54082 , n53732 , n36345 );
and ( n54083 , n13239 , n43721 );
or ( n54084 , n54082 , n54083 );
and ( n54085 , n54084 , n37841 );
and ( n54086 , n15097 , n14564 );
and ( n54087 , n15097 , n36345 );
and ( n54088 , n13239 , n43721 );
or ( n54089 , n54087 , n54088 );
and ( n54090 , n54089 , n37847 );
or ( n54091 , n54065 , n54069 , n54073 , n54077 , n54081 , n54085 , n54086 , n54090 );
and ( n54092 , n54064 , n54091 );
and ( n54093 , n13239 , n34821 );
or ( n54094 , n54092 , n54093 );
and ( n54095 , n54094 , n16574 );
and ( n54096 , n12270 , n16576 );
or ( n54097 , n54095 , n54096 );
buf ( n54098 , n54097 );
buf ( n54099 , n54098 );
buf ( n54100 , n10613 );
buf ( n54101 , n10613 );
not ( n54102 , n24800 );
and ( n54103 , n26697 , n25222 );
and ( n54104 , n43420 , n28589 );
and ( n54105 , n26697 , n31075 );
or ( n54106 , n54104 , n54105 );
and ( n54107 , n54106 , n28594 );
and ( n54108 , n43436 , n28589 );
and ( n54109 , n26697 , n31075 );
or ( n54110 , n54108 , n54109 );
and ( n54111 , n54110 , n30269 );
and ( n54112 , n43452 , n28589 );
and ( n54113 , n26697 , n31075 );
or ( n54114 , n54112 , n54113 );
and ( n54115 , n54114 , n30982 );
and ( n54116 , n29172 , n28589 );
and ( n54117 , n26697 , n31075 );
or ( n54118 , n54116 , n54117 );
and ( n54119 , n54118 , n30989 );
and ( n54120 , n29172 , n30991 );
and ( n54121 , n43471 , n28589 );
and ( n54122 , n26697 , n31075 );
or ( n54123 , n54121 , n54122 );
and ( n54124 , n54123 , n31002 );
or ( n54125 , n54103 , n54107 , n54111 , n54115 , n54119 , n54120 , n54124 );
and ( n54126 , n54102 , n54125 );
and ( n54127 , n26697 , n24800 );
or ( n54128 , n54126 , n54127 );
and ( n54129 , n54128 , n31008 );
and ( n54130 , n25594 , n10618 );
or ( n54131 , n54129 , n54130 );
buf ( n54132 , n54131 );
buf ( n54133 , n54132 );
not ( n54134 , n24800 );
and ( n54135 , n25950 , n25222 );
and ( n54136 , n48334 , n28589 );
and ( n54137 , n25950 , n31075 );
or ( n54138 , n54136 , n54137 );
and ( n54139 , n54138 , n28594 );
and ( n54140 , n48344 , n28589 );
and ( n54141 , n25950 , n31075 );
or ( n54142 , n54140 , n54141 );
and ( n54143 , n54142 , n30269 );
and ( n54144 , n48354 , n28589 );
and ( n54145 , n25950 , n31075 );
or ( n54146 , n54144 , n54145 );
and ( n54147 , n54146 , n30982 );
and ( n54148 , n29615 , n28589 );
and ( n54149 , n25950 , n31075 );
or ( n54150 , n54148 , n54149 );
and ( n54151 , n54150 , n30989 );
and ( n54152 , n29615 , n30991 );
and ( n54153 , n48364 , n28589 );
and ( n54154 , n25950 , n31075 );
or ( n54155 , n54153 , n54154 );
and ( n54156 , n54155 , n31002 );
or ( n54157 , n54135 , n54139 , n54143 , n54147 , n54151 , n54152 , n54156 );
and ( n54158 , n54134 , n54157 );
and ( n54159 , n25950 , n24800 );
or ( n54160 , n54158 , n54159 );
and ( n54161 , n54160 , n31008 );
and ( n54162 , n25264 , n10618 );
or ( n54163 , n54161 , n54162 );
buf ( n54164 , n54163 );
buf ( n54165 , n54164 );
buf ( n54166 , n10615 );
buf ( n54167 , n10615 );
buf ( n54168 , n10615 );
buf ( n54169 , n10615 );
buf ( n54170 , n10613 );
not ( n54171 , n34821 );
and ( n54172 , n13445 , n14592 );
and ( n54173 , n43142 , n36348 );
and ( n54174 , n13445 , n43530 );
or ( n54175 , n54173 , n54174 );
and ( n54176 , n54175 , n14562 );
and ( n54177 , n43152 , n36347 );
and ( n54178 , n13445 , n43543 );
or ( n54179 , n54177 , n54178 );
and ( n54180 , n54179 , n14586 );
and ( n54181 , n43162 , n36348 );
and ( n54182 , n13445 , n43556 );
or ( n54183 , n54181 , n54182 );
and ( n54184 , n54183 , n14584 );
and ( n54185 , n43152 , n36347 );
and ( n54186 , n13445 , n43563 );
or ( n54187 , n54185 , n54186 );
and ( n54188 , n54187 , n37835 );
and ( n54189 , n43162 , n36347 );
and ( n54190 , n13445 , n43563 );
or ( n54191 , n54189 , n54190 );
and ( n54192 , n54191 , n37841 );
and ( n54193 , n13443 , n14564 );
and ( n54194 , n15779 , n36347 );
and ( n54195 , n13445 , n43563 );
or ( n54196 , n54194 , n54195 );
and ( n54197 , n54196 , n37847 );
or ( n54198 , n54172 , n54176 , n54180 , n54184 , n54188 , n54192 , n54193 , n54197 );
and ( n54199 , n54171 , n54198 );
and ( n54200 , n13445 , n34821 );
or ( n54201 , n54199 , n54200 );
and ( n54202 , n54201 , n16574 );
and ( n54203 , n13445 , n16576 );
or ( n54204 , n54202 , n54203 );
buf ( n54205 , n54204 );
buf ( n54206 , n54205 );
buf ( n54207 , n10613 );
buf ( n54208 , n10613 );
buf ( n54209 , n10613 );
buf ( n54210 , n10613 );
buf ( n54211 , n10613 );
and ( n54212 , n24126 , n31008 );
and ( n54213 , n29346 , n10618 );
or ( n54214 , n54212 , n54213 );
buf ( n54215 , n54214 );
buf ( n54216 , n54215 );
buf ( n54217 , n10613 );
buf ( n54218 , n10615 );
not ( n54219 , n34821 );
and ( n54220 , n53712 , n36345 );
and ( n54221 , n13245 , n36352 );
or ( n54222 , n54220 , n54221 );
and ( n54223 , n54222 , n14562 );
and ( n54224 , n53722 , n36345 );
and ( n54225 , n13245 , n37073 );
or ( n54226 , n54224 , n54225 );
and ( n54227 , n54226 , n14586 );
and ( n54228 , n53732 , n36350 );
and ( n54229 , n13245 , n37825 );
or ( n54230 , n54228 , n54229 );
and ( n54231 , n54230 , n14584 );
and ( n54232 , n53722 , n36350 );
and ( n54233 , n13245 , n37831 );
or ( n54234 , n54232 , n54233 );
and ( n54235 , n54234 , n37835 );
and ( n54236 , n53732 , n36350 );
and ( n54237 , n13245 , n37831 );
or ( n54238 , n54236 , n54237 );
and ( n54239 , n54238 , n37841 );
and ( n54240 , n15097 , n36350 );
and ( n54241 , n13245 , n37831 );
or ( n54242 , n54240 , n54241 );
and ( n54243 , n54242 , n37847 );
and ( n54244 , n13245 , n37849 );
or ( n54245 , n54223 , n54227 , n54231 , n54235 , n54239 , n54243 , n54244 );
and ( n54246 , n54219 , n54245 );
and ( n54247 , n13245 , n34821 );
or ( n54248 , n54246 , n54247 );
and ( n54249 , n54248 , n16574 );
and ( n54250 , n13245 , n16576 );
or ( n54251 , n54249 , n54250 );
buf ( n54252 , n54251 );
buf ( n54253 , n54252 );
and ( n54254 , n11792 , n16574 );
and ( n54255 , n15005 , n16576 );
or ( n54256 , n54254 , n54255 );
buf ( n54257 , n54256 );
buf ( n54258 , n54257 );
buf ( n54259 , n10615 );
buf ( n54260 , n10613 );
not ( n54261 , n17451 );
and ( n54262 , n19077 , n17873 );
and ( n54263 , n39326 , n21336 );
and ( n54264 , n19077 , n42682 );
or ( n54265 , n54263 , n54264 );
and ( n54266 , n54265 , n21341 );
and ( n54267 , n39336 , n21336 );
and ( n54268 , n19077 , n42682 );
or ( n54269 , n54267 , n54268 );
and ( n54270 , n54269 , n23064 );
and ( n54271 , n39346 , n21336 );
and ( n54272 , n19077 , n42682 );
or ( n54273 , n54271 , n54272 );
and ( n54274 , n54273 , n23825 );
and ( n54275 , n22082 , n21336 );
and ( n54276 , n19077 , n42682 );
or ( n54277 , n54275 , n54276 );
and ( n54278 , n54277 , n23832 );
and ( n54279 , n22082 , n23834 );
and ( n54280 , n39356 , n21336 );
and ( n54281 , n19077 , n42682 );
or ( n54282 , n54280 , n54281 );
and ( n54283 , n54282 , n23917 );
or ( n54284 , n54262 , n54266 , n54270 , n54274 , n54278 , n54279 , n54283 );
and ( n54285 , n54261 , n54284 );
and ( n54286 , n19077 , n17451 );
or ( n54287 , n54285 , n54286 );
and ( n54288 , n54287 , n23924 );
and ( n54289 , n18125 , n23926 );
or ( n54290 , n54288 , n54289 );
buf ( n54291 , n54290 );
buf ( n54292 , n54291 );
buf ( n54293 , n10615 );
not ( n54294 , n24511 );
not ( n54295 , n24799 );
and ( n54296 , n10710 , n40154 );
not ( n54297 , n40632 );
and ( n54298 , n54297 , n40390 );
xor ( n54299 , n40645 , n40655 );
and ( n54300 , n54299 , n40632 );
or ( n54301 , n54298 , n54300 );
buf ( n54302 , n54301 );
and ( n54303 , n54302 , n27046 );
not ( n54304 , n41147 );
and ( n54305 , n54304 , n40905 );
xor ( n54306 , n41160 , n41170 );
and ( n54307 , n54306 , n41147 );
or ( n54308 , n54305 , n54307 );
buf ( n54309 , n54308 );
and ( n54310 , n54309 , n27049 );
and ( n54311 , n29573 , n28506 );
and ( n54312 , n10710 , n28508 );
or ( n54313 , n54303 , n54310 , n54311 , n54312 );
and ( n54314 , n54313 , n41199 );
or ( n54315 , n54296 , n54314 );
and ( n54316 , n54295 , n54315 );
xor ( n54317 , n41676 , n41684 );
xor ( n54318 , n54317 , n41776 );
buf ( n54319 , n54318 );
and ( n54320 , n54319 , n27046 );
xor ( n54321 , n42213 , n42214 );
xor ( n54322 , n54321 , n42272 );
buf ( n54323 , n54322 );
and ( n54324 , n54323 , n27049 );
and ( n54325 , n29573 , n42306 );
or ( n54326 , n54320 , n54324 , n54325 );
buf ( n54327 , n54326 );
and ( n54328 , C1 , n54327 );
or ( n54329 , n54328 , C0 );
buf ( n54330 , n54329 );
not ( n54331 , n54330 );
buf ( n54332 , n54331 );
buf ( n54333 , n54332 );
not ( n54334 , n54333 );
and ( n54335 , C1 , n54334 );
or ( n54336 , n54335 , C0 );
buf ( n54337 , n54336 );
and ( n54338 , n54337 , n24799 );
or ( n54339 , n54316 , n54338 );
and ( n54340 , n54294 , n54339 );
and ( n54341 , n54313 , n24511 );
or ( n54342 , n54340 , n54341 );
and ( n54343 , n54342 , n31008 );
not ( n54344 , n42601 );
and ( n54345 , n54344 , n42401 );
xor ( n54346 , n42614 , n42624 );
and ( n54347 , n54346 , n42601 );
or ( n54348 , n54345 , n54347 );
buf ( n54349 , n54348 );
and ( n54350 , n54349 , n10618 );
or ( n54351 , n54343 , n54350 );
buf ( n54352 , n54351 );
buf ( n54353 , n54352 );
buf ( n54354 , n10613 );
not ( n54355 , n34821 );
and ( n54356 , n43049 , n36345 );
and ( n54357 , n13305 , n36352 );
or ( n54358 , n54356 , n54357 );
and ( n54359 , n54358 , n14562 );
and ( n54360 , n43071 , n36345 );
and ( n54361 , n13305 , n37073 );
or ( n54362 , n54360 , n54361 );
and ( n54363 , n54362 , n14586 );
and ( n54364 , n43093 , n36350 );
and ( n54365 , n13305 , n37825 );
or ( n54366 , n54364 , n54365 );
and ( n54367 , n54366 , n14584 );
and ( n54368 , n43071 , n36350 );
and ( n54369 , n13305 , n37831 );
or ( n54370 , n54368 , n54369 );
and ( n54371 , n54370 , n37835 );
and ( n54372 , n43093 , n36350 );
and ( n54373 , n13305 , n37831 );
or ( n54374 , n54372 , n54373 );
and ( n54375 , n54374 , n37841 );
and ( n54376 , n15515 , n36350 );
and ( n54377 , n13305 , n37831 );
or ( n54378 , n54376 , n54377 );
and ( n54379 , n54378 , n37847 );
and ( n54380 , n13305 , n37849 );
or ( n54381 , n54359 , n54363 , n54367 , n54371 , n54375 , n54379 , n54380 );
and ( n54382 , n54355 , n54381 );
and ( n54383 , n13305 , n34821 );
or ( n54384 , n54382 , n54383 );
and ( n54385 , n54384 , n16574 );
and ( n54386 , n13305 , n16576 );
or ( n54387 , n54385 , n54386 );
buf ( n54388 , n54387 );
buf ( n54389 , n54388 );
not ( n54390 , n11954 );
not ( n54391 , n12243 );
and ( n54392 , n10861 , n31187 );
not ( n54393 , n31697 );
and ( n54394 , n54393 , n31557 );
xor ( n54395 , n31557 , n31371 );
and ( n54396 , n50356 , n50375 );
xor ( n54397 , n54395 , n54396 );
and ( n54398 , n54397 , n31697 );
or ( n54399 , n54394 , n54398 );
buf ( n54400 , n54399 );
and ( n54401 , n54400 , n14140 );
not ( n54402 , n32214 );
and ( n54403 , n54402 , n32074 );
xor ( n54404 , n32074 , n31888 );
and ( n54405 , n50383 , n50402 );
xor ( n54406 , n54404 , n54405 );
and ( n54407 , n54406 , n32214 );
or ( n54408 , n54403 , n54407 );
buf ( n54409 , n54408 );
and ( n54410 , n54409 , n14137 );
and ( n54411 , n15623 , n14143 );
and ( n54412 , n10861 , n14141 );
or ( n54413 , n54401 , n54410 , n54411 , n54412 );
and ( n54414 , n54413 , n32236 );
or ( n54415 , n54392 , n54414 );
and ( n54416 , n54391 , n54415 );
not ( n54417 , n34038 );
and ( n54418 , n54417 , n33842 );
xor ( n54419 , n33842 , n33579 );
and ( n54420 , n50416 , n50435 );
xor ( n54421 , n54419 , n54420 );
and ( n54422 , n54421 , n34038 );
or ( n54423 , n54418 , n54422 );
buf ( n54424 , n54423 );
and ( n54425 , n54424 , n12243 );
or ( n54426 , n54416 , n54425 );
and ( n54427 , n54390 , n54426 );
and ( n54428 , n54413 , n11954 );
or ( n54429 , n54427 , n54428 );
and ( n54430 , n54429 , n16574 );
not ( n54431 , n34327 );
and ( n54432 , n54431 , n34211 );
xor ( n54433 , n34211 , n34058 );
and ( n54434 , n50448 , n50467 );
xor ( n54435 , n54433 , n54434 );
and ( n54436 , n54435 , n34327 );
or ( n54437 , n54432 , n54436 );
buf ( n54438 , n54437 );
and ( n54439 , n54438 , n16576 );
or ( n54440 , n54430 , n54439 );
buf ( n54441 , n54440 );
buf ( n54442 , n54441 );
buf ( n54443 , n10615 );
not ( n54444 , n34821 );
and ( n54445 , n13407 , n14592 );
and ( n54446 , n36271 , n36350 );
and ( n54447 , n13407 , n43691 );
or ( n54448 , n54446 , n54447 );
and ( n54449 , n54448 , n14562 );
and ( n54450 , n37069 , n36350 );
and ( n54451 , n13407 , n43703 );
or ( n54452 , n54450 , n54451 );
and ( n54453 , n54452 , n14586 );
and ( n54454 , n37822 , n36345 );
and ( n54455 , n13407 , n43715 );
or ( n54456 , n54454 , n54455 );
and ( n54457 , n54456 , n14584 );
and ( n54458 , n37069 , n36345 );
and ( n54459 , n13407 , n43721 );
or ( n54460 , n54458 , n54459 );
and ( n54461 , n54460 , n37835 );
and ( n54462 , n37822 , n36345 );
and ( n54463 , n13407 , n43721 );
or ( n54464 , n54462 , n54463 );
and ( n54465 , n54464 , n37841 );
and ( n54466 , n15713 , n14564 );
and ( n54467 , n15713 , n36345 );
and ( n54468 , n13407 , n43721 );
or ( n54469 , n54467 , n54468 );
and ( n54470 , n54469 , n37847 );
or ( n54471 , n54445 , n54449 , n54453 , n54457 , n54461 , n54465 , n54466 , n54470 );
and ( n54472 , n54444 , n54471 );
and ( n54473 , n13407 , n34821 );
or ( n54474 , n54472 , n54473 );
and ( n54475 , n54474 , n16574 );
and ( n54476 , n12312 , n16576 );
or ( n54477 , n54475 , n54476 );
buf ( n54478 , n54477 );
buf ( n54479 , n54478 );
buf ( n54480 , n10613 );
buf ( n54481 , n10613 );
buf ( n54482 , n10615 );
and ( n54483 , n11681 , n16574 );
and ( n54484 , n15814 , n16576 );
or ( n54485 , n54483 , n54484 );
buf ( n54486 , n54485 );
buf ( n54487 , n54486 );
buf ( n54488 , n10615 );
not ( n54489 , n17162 );
not ( n54490 , n17450 );
and ( n54491 , n10621 , n37947 );
not ( n54492 , n38425 );
and ( n54493 , n54492 , n37958 );
xor ( n54494 , n38440 , n38099 );
and ( n54495 , n54494 , n38425 );
or ( n54496 , n54493 , n54495 );
buf ( n54497 , n54496 );
and ( n54498 , n54497 , n19745 );
not ( n54499 , n38934 );
and ( n54500 , n54499 , n38467 );
xor ( n54501 , n38949 , n38608 );
and ( n54502 , n54501 , n38934 );
or ( n54503 , n54500 , n54502 );
buf ( n54504 , n54503 );
and ( n54505 , n54504 , n19748 );
and ( n54506 , n21637 , n21253 );
and ( n54507 , n10621 , n21255 );
or ( n54508 , n54498 , n54505 , n54506 , n54507 );
and ( n54509 , n54508 , n38980 );
or ( n54510 , n54491 , n54509 );
and ( n54511 , n54490 , n54510 );
or ( n54512 , n54511 , C0 );
and ( n54513 , n54489 , n54512 );
and ( n54514 , n54508 , n17162 );
or ( n54515 , n54513 , n54514 );
and ( n54516 , n54515 , n23924 );
not ( n54517 , n39264 );
and ( n54518 , n54517 , n38994 );
xor ( n54519 , n39279 , n38995 );
and ( n54520 , n54519 , n39264 );
or ( n54521 , n54518 , n54520 );
buf ( n54522 , n54521 );
and ( n54523 , n54522 , n23926 );
or ( n54524 , n54516 , n54523 );
buf ( n54525 , n54524 );
buf ( n54526 , n54525 );
buf ( n54527 , n10615 );
buf ( n54528 , n10613 );
buf ( n54529 , n10613 );
buf ( n54530 , n10613 );
buf ( n54531 , n10615 );
buf ( n54532 , n10613 );
buf ( n54533 , n10615 );
buf ( n54534 , n10615 );
buf ( n54535 , n10615 );
not ( n54536 , n34804 );
and ( n54537 , n54536 , n26671 );
and ( n54538 , n14689 , n34804 );
or ( n54539 , n54537 , n54538 );
and ( n54540 , n54539 , n31008 );
and ( n54541 , n14689 , n10618 );
or ( n54542 , n54540 , n54541 );
buf ( n54543 , n54542 );
buf ( n54544 , n54543 );
buf ( n54545 , n10613 );
not ( n54546 , n24511 );
buf ( n54547 , n28606 );
buf ( n54548 , n54547 );
and ( n54549 , n54548 , n41199 );
buf ( n54550 , n54549 );
not ( n54551 , n24799 );
and ( n54552 , n54550 , n54551 );
and ( n54553 , n54546 , n54552 );
and ( n54554 , n54548 , n24511 );
or ( n54555 , n54553 , n54554 );
and ( n54556 , n54555 , n31008 );
buf ( n54557 , n10618 );
or ( n54558 , n54556 , n54557 );
buf ( n54559 , n54558 );
buf ( n54560 , n54559 );
buf ( n54561 , n10613 );
buf ( n54562 , n10613 );
buf ( n54563 , n10613 );
buf ( n54564 , n10615 );
buf ( n54565 , n10613 );
not ( n54566 , n17451 );
and ( n54567 , n48952 , n21333 );
and ( n54568 , n18606 , n34758 );
or ( n54569 , n54567 , n54568 );
and ( n54570 , n54569 , n21341 );
and ( n54571 , n48962 , n21333 );
and ( n54572 , n18606 , n34758 );
or ( n54573 , n54571 , n54572 );
and ( n54574 , n54573 , n23064 );
and ( n54575 , n48972 , n21333 );
and ( n54576 , n18606 , n34758 );
or ( n54577 , n54575 , n54576 );
and ( n54578 , n54577 , n23825 );
and ( n54579 , n22362 , n21333 );
and ( n54580 , n18606 , n34758 );
or ( n54581 , n54579 , n54580 );
and ( n54582 , n54581 , n23832 );
and ( n54583 , n48982 , n21333 );
and ( n54584 , n18606 , n34758 );
or ( n54585 , n54583 , n54584 );
and ( n54586 , n54585 , n23917 );
and ( n54587 , n18606 , n34526 );
or ( n54588 , n54570 , n54574 , n54578 , n54582 , n54586 , n54587 );
and ( n54589 , n54566 , n54588 );
and ( n54590 , n18606 , n17451 );
or ( n54591 , n54589 , n54590 );
and ( n54592 , n54591 , n23924 );
and ( n54593 , n18606 , n23926 );
or ( n54594 , n54592 , n54593 );
buf ( n54595 , n54594 );
buf ( n54596 , n54595 );
not ( n54597 , n34821 );
and ( n54598 , n13383 , n14592 );
and ( n54599 , n44916 , n36350 );
and ( n54600 , n13383 , n43691 );
or ( n54601 , n54599 , n54600 );
and ( n54602 , n54601 , n14562 );
and ( n54603 , n44926 , n36350 );
and ( n54604 , n13383 , n43703 );
or ( n54605 , n54603 , n54604 );
and ( n54606 , n54605 , n14586 );
and ( n54607 , n44936 , n36345 );
and ( n54608 , n13383 , n43715 );
or ( n54609 , n54607 , n54608 );
and ( n54610 , n54609 , n14584 );
and ( n54611 , n44926 , n36345 );
and ( n54612 , n13383 , n43721 );
or ( n54613 , n54611 , n54612 );
and ( n54614 , n54613 , n37835 );
and ( n54615 , n44936 , n36345 );
and ( n54616 , n13383 , n43721 );
or ( n54617 , n54615 , n54616 );
and ( n54618 , n54617 , n37841 );
and ( n54619 , n15669 , n14564 );
and ( n54620 , n15669 , n36345 );
and ( n54621 , n13383 , n43721 );
or ( n54622 , n54620 , n54621 );
and ( n54623 , n54622 , n37847 );
or ( n54624 , n54598 , n54602 , n54606 , n54610 , n54614 , n54618 , n54619 , n54623 );
and ( n54625 , n54597 , n54624 );
and ( n54626 , n13383 , n34821 );
or ( n54627 , n54625 , n54626 );
and ( n54628 , n54627 , n16574 );
and ( n54629 , n12306 , n16576 );
or ( n54630 , n54628 , n54629 );
buf ( n54631 , n54630 );
buf ( n54632 , n54631 );
not ( n54633 , n24800 );
and ( n54634 , n26595 , n25222 );
and ( n54635 , n42864 , n28589 );
and ( n54636 , n26595 , n31075 );
or ( n54637 , n54635 , n54636 );
and ( n54638 , n54637 , n28594 );
and ( n54639 , n42884 , n28589 );
and ( n54640 , n26595 , n31075 );
or ( n54641 , n54639 , n54640 );
and ( n54642 , n54641 , n30269 );
and ( n54643 , n42904 , n28589 );
and ( n54644 , n26595 , n31075 );
or ( n54645 , n54643 , n54644 );
and ( n54646 , n54645 , n30982 );
and ( n54647 , n29211 , n28589 );
and ( n54648 , n26595 , n31075 );
or ( n54649 , n54647 , n54648 );
and ( n54650 , n54649 , n30989 );
and ( n54651 , n29211 , n30991 );
and ( n54652 , n42929 , n28589 );
and ( n54653 , n26595 , n31075 );
or ( n54654 , n54652 , n54653 );
and ( n54655 , n54654 , n31002 );
or ( n54656 , n54634 , n54638 , n54642 , n54646 , n54650 , n54651 , n54655 );
and ( n54657 , n54633 , n54656 );
and ( n54658 , n26595 , n24800 );
or ( n54659 , n54657 , n54658 );
and ( n54660 , n54659 , n31008 );
and ( n54661 , n25549 , n10618 );
or ( n54662 , n54660 , n54661 );
buf ( n54663 , n54662 );
buf ( n54664 , n54663 );
buf ( n54665 , n10613 );
buf ( n54666 , n10615 );
buf ( n54667 , n10613 );
buf ( n54668 , n10615 );
not ( n54669 , n34821 );
and ( n54670 , n13506 , n14592 );
and ( n54671 , n53772 , n36350 );
and ( n54672 , n13506 , n43691 );
or ( n54673 , n54671 , n54672 );
and ( n54674 , n54673 , n14562 );
and ( n54675 , n53782 , n36350 );
and ( n54676 , n13506 , n43703 );
or ( n54677 , n54675 , n54676 );
and ( n54678 , n54677 , n14586 );
and ( n54679 , n53792 , n36345 );
and ( n54680 , n13506 , n43715 );
or ( n54681 , n54679 , n54680 );
and ( n54682 , n54681 , n14584 );
and ( n54683 , n53782 , n36345 );
and ( n54684 , n13506 , n43721 );
or ( n54685 , n54683 , n54684 );
and ( n54686 , n54685 , n37835 );
and ( n54687 , n53792 , n36345 );
and ( n54688 , n13506 , n43721 );
or ( n54689 , n54687 , n54688 );
and ( n54690 , n54689 , n37841 );
and ( n54691 , n15866 , n14564 );
and ( n54692 , n15866 , n36345 );
and ( n54693 , n13506 , n43721 );
or ( n54694 , n54692 , n54693 );
and ( n54695 , n54694 , n37847 );
or ( n54696 , n54670 , n54674 , n54678 , n54682 , n54686 , n54690 , n54691 , n54695 );
and ( n54697 , n54669 , n54696 );
and ( n54698 , n13506 , n34821 );
or ( n54699 , n54697 , n54698 );
and ( n54700 , n54699 , n16574 );
and ( n54701 , n12333 , n16576 );
or ( n54702 , n54700 , n54701 );
buf ( n54703 , n54702 );
buf ( n54704 , n54703 );
buf ( n54705 , n10613 );
buf ( n54706 , n10613 );
buf ( n54707 , n10613 );
not ( n54708 , n17162 );
not ( n54709 , n17450 );
and ( n54710 , n10698 , n37947 );
not ( n54711 , n38425 );
and ( n54712 , n54711 , n38217 );
xor ( n54713 , n38433 , n38447 );
and ( n54714 , n54713 , n38425 );
or ( n54715 , n54712 , n54714 );
buf ( n54716 , n54715 );
and ( n54717 , n54716 , n19745 );
not ( n54718 , n38934 );
and ( n54719 , n54718 , n38726 );
xor ( n54720 , n38942 , n38956 );
and ( n54721 , n54720 , n38934 );
or ( n54722 , n54719 , n54721 );
buf ( n54723 , n54722 );
and ( n54724 , n54723 , n19748 );
and ( n54725 , n22280 , n21253 );
and ( n54726 , n10698 , n21255 );
or ( n54727 , n54717 , n54724 , n54725 , n54726 );
and ( n54728 , n54727 , n38980 );
or ( n54729 , n54710 , n54728 );
and ( n54730 , n54709 , n54729 );
or ( n54731 , n54730 , C0 );
and ( n54732 , n54708 , n54731 );
and ( n54733 , n54727 , n17162 );
or ( n54734 , n54732 , n54733 );
and ( n54735 , n54734 , n23924 );
not ( n54736 , n39264 );
and ( n54737 , n54736 , n39092 );
xor ( n54738 , n39272 , n39286 );
and ( n54739 , n54738 , n39264 );
or ( n54740 , n54737 , n54739 );
buf ( n54741 , n54740 );
and ( n54742 , n54741 , n23926 );
or ( n54743 , n54735 , n54742 );
buf ( n54744 , n54743 );
buf ( n54745 , n54744 );
not ( n54746 , n24800 );
and ( n54747 , n26461 , n25222 );
and ( n54748 , n47642 , n28583 );
and ( n54749 , n26461 , n28591 );
or ( n54750 , n54748 , n54749 );
and ( n54751 , n54750 , n28594 );
and ( n54752 , n47652 , n28583 );
and ( n54753 , n26461 , n28591 );
or ( n54754 , n54752 , n54753 );
and ( n54755 , n54754 , n30269 );
and ( n54756 , n47662 , n28583 );
and ( n54757 , n26461 , n28591 );
or ( n54758 , n54756 , n54757 );
and ( n54759 , n54758 , n30982 );
and ( n54760 , n29315 , n28583 );
and ( n54761 , n26461 , n28591 );
or ( n54762 , n54760 , n54761 );
and ( n54763 , n54762 , n30989 );
and ( n54764 , n26459 , n30991 );
and ( n54765 , n47672 , n28583 );
and ( n54766 , n26461 , n28591 );
or ( n54767 , n54765 , n54766 );
and ( n54768 , n54767 , n31002 );
or ( n54769 , n54747 , n54751 , n54755 , n54759 , n54763 , n54764 , n54768 );
and ( n54770 , n54746 , n54769 );
and ( n54771 , n26461 , n24800 );
or ( n54772 , n54770 , n54771 );
and ( n54773 , n54772 , n31008 );
and ( n54774 , n26461 , n10618 );
or ( n54775 , n54773 , n54774 );
buf ( n54776 , n54775 );
buf ( n54777 , n54776 );
buf ( n54778 , n10615 );
not ( n54779 , n17451 );
and ( n54780 , n21257 , n21334 );
and ( n54781 , n19354 , n34492 );
or ( n54782 , n54780 , n54781 );
and ( n54783 , n54782 , n21341 );
and ( n54784 , n23053 , n21334 );
and ( n54785 , n19354 , n34492 );
or ( n54786 , n54784 , n54785 );
and ( n54787 , n54786 , n23064 );
and ( n54788 , n23815 , n21334 );
and ( n54789 , n19354 , n34492 );
or ( n54790 , n54788 , n54789 );
and ( n54791 , n54790 , n23825 );
and ( n54792 , n21919 , n21334 );
and ( n54793 , n19354 , n34492 );
or ( n54794 , n54792 , n54793 );
and ( n54795 , n54794 , n23832 );
and ( n54796 , n23913 , n21334 );
and ( n54797 , n19354 , n34492 );
or ( n54798 , n54796 , n54797 );
and ( n54799 , n54798 , n23917 );
and ( n54800 , n19354 , n34526 );
or ( n54801 , n54783 , n54787 , n54791 , n54795 , n54799 , n54800 );
and ( n54802 , n54779 , n54801 );
and ( n54803 , n19354 , n17451 );
or ( n54804 , n54802 , n54803 );
and ( n54805 , n54804 , n23924 );
and ( n54806 , n19354 , n23926 );
or ( n54807 , n54805 , n54806 );
buf ( n54808 , n54807 );
buf ( n54809 , n54808 );
buf ( n54810 , n10615 );
buf ( n54811 , n10613 );
not ( n54812 , n24800 );
not ( n54813 , n26823 );
and ( n54814 , n54813 , n26615 );
xor ( n54815 , n43392 , n43393 );
and ( n54816 , n54815 , n26823 );
or ( n54817 , n54814 , n54816 );
buf ( n54818 , n54817 );
and ( n54819 , n54818 , n27046 );
and ( n54820 , n54818 , n27049 );
not ( n54821 , n27051 );
and ( n54822 , n54821 , n28368 );
not ( n54823 , n28494 );
and ( n54824 , n54823 , n28380 );
xor ( n54825 , n43408 , n43409 );
and ( n54826 , n54825 , n28494 );
or ( n54827 , n54824 , n54826 );
buf ( n54828 , n54827 );
and ( n54829 , n54828 , n27051 );
or ( n54830 , n54822 , n54829 );
and ( n54831 , n54830 , n28506 );
and ( n54832 , n28368 , n28508 );
or ( n54833 , n54819 , n54820 , n54831 , n54832 );
and ( n54834 , n54833 , n28587 );
and ( n54835 , n26635 , n39807 );
or ( n54836 , n54834 , n54835 );
and ( n54837 , n54836 , n28594 );
not ( n54838 , n30249 );
and ( n54839 , n54838 , n30143 );
xor ( n54840 , n43429 , n43430 );
and ( n54841 , n54840 , n30249 );
or ( n54842 , n54839 , n54841 );
buf ( n54843 , n54842 );
and ( n54844 , n54843 , n28587 );
and ( n54845 , n26635 , n39807 );
or ( n54846 , n54844 , n54845 );
and ( n54847 , n54846 , n30269 );
not ( n54848 , n30963 );
and ( n54849 , n54848 , n30857 );
xor ( n54850 , n43445 , n43446 );
and ( n54851 , n54850 , n30963 );
or ( n54852 , n54849 , n54851 );
buf ( n54853 , n54852 );
and ( n54854 , n54853 , n28587 );
and ( n54855 , n26635 , n39807 );
or ( n54856 , n54854 , n54855 );
and ( n54857 , n54856 , n30982 );
and ( n54858 , n29198 , n28587 );
and ( n54859 , n26635 , n39807 );
or ( n54860 , n54858 , n54859 );
and ( n54861 , n54860 , n30989 );
xor ( n54862 , n43466 , n43467 );
buf ( n54863 , n54862 );
and ( n54864 , n54863 , n28587 );
and ( n54865 , n26635 , n39807 );
or ( n54866 , n54864 , n54865 );
and ( n54867 , n54866 , n31002 );
and ( n54868 , n26635 , n34607 );
or ( n54869 , n54837 , n54847 , n54857 , n54861 , n54867 , n54868 );
and ( n54870 , n54812 , n54869 );
and ( n54871 , n26635 , n24800 );
or ( n54872 , n54870 , n54871 );
and ( n54873 , n54872 , n31008 );
and ( n54874 , n26635 , n10618 );
or ( n54875 , n54873 , n54874 );
buf ( n54876 , n54875 );
buf ( n54877 , n54876 );
buf ( n54878 , n10615 );
buf ( n54879 , n10613 );
buf ( n54880 , n10615 );
buf ( n54881 , n10613 );
not ( n54882 , n24800 );
and ( n54883 , n45258 , n28587 );
and ( n54884 , n26805 , n39807 );
or ( n54885 , n54883 , n54884 );
and ( n54886 , n54885 , n28594 );
and ( n54887 , n45274 , n28587 );
and ( n54888 , n26805 , n39807 );
or ( n54889 , n54887 , n54888 );
and ( n54890 , n54889 , n30269 );
and ( n54891 , n45290 , n28587 );
and ( n54892 , n26805 , n39807 );
or ( n54893 , n54891 , n54892 );
and ( n54894 , n54893 , n30982 );
and ( n54895 , n29133 , n28587 );
and ( n54896 , n26805 , n39807 );
or ( n54897 , n54895 , n54896 );
and ( n54898 , n54897 , n30989 );
and ( n54899 , n45310 , n28587 );
and ( n54900 , n26805 , n39807 );
or ( n54901 , n54899 , n54900 );
and ( n54902 , n54901 , n31002 );
and ( n54903 , n26805 , n34607 );
or ( n54904 , n54886 , n54890 , n54894 , n54898 , n54902 , n54903 );
and ( n54905 , n54882 , n54904 );
and ( n54906 , n26805 , n24800 );
or ( n54907 , n54905 , n54906 );
and ( n54908 , n54907 , n31008 );
and ( n54909 , n26805 , n10618 );
or ( n54910 , n54908 , n54909 );
buf ( n54911 , n54910 );
buf ( n54912 , n54911 );
buf ( n54913 , n10613 );
buf ( n54914 , n10615 );
not ( n54915 , n34804 );
and ( n54916 , n54915 , n26229 );
and ( n54917 , n14767 , n34804 );
or ( n54918 , n54916 , n54917 );
and ( n54919 , n54918 , n31008 );
and ( n54920 , n14767 , n10618 );
or ( n54921 , n54919 , n54920 );
buf ( n54922 , n54921 );
buf ( n54923 , n54922 );
not ( n54924 , n34821 );
and ( n54925 , n13287 , n14592 );
and ( n54926 , n51156 , n36350 );
and ( n54927 , n13287 , n43691 );
or ( n54928 , n54926 , n54927 );
and ( n54929 , n54928 , n14562 );
and ( n54930 , n51166 , n36350 );
and ( n54931 , n13287 , n43703 );
or ( n54932 , n54930 , n54931 );
and ( n54933 , n54932 , n14586 );
and ( n54934 , n51176 , n36345 );
and ( n54935 , n13287 , n43715 );
or ( n54936 , n54934 , n54935 );
and ( n54937 , n54936 , n14584 );
and ( n54938 , n51166 , n36345 );
and ( n54939 , n13287 , n43721 );
or ( n54940 , n54938 , n54939 );
and ( n54941 , n54940 , n37835 );
and ( n54942 , n51176 , n36345 );
and ( n54943 , n13287 , n43721 );
or ( n54944 , n54942 , n54943 );
and ( n54945 , n54944 , n37841 );
and ( n54946 , n15493 , n14564 );
and ( n54947 , n15493 , n36345 );
and ( n54948 , n13287 , n43721 );
or ( n54949 , n54947 , n54948 );
and ( n54950 , n54949 , n37847 );
or ( n54951 , n54925 , n54929 , n54933 , n54937 , n54941 , n54945 , n54946 , n54950 );
and ( n54952 , n54924 , n54951 );
and ( n54953 , n13287 , n34821 );
or ( n54954 , n54952 , n54953 );
and ( n54955 , n54954 , n16574 );
and ( n54956 , n12282 , n16576 );
or ( n54957 , n54955 , n54956 );
buf ( n54958 , n54957 );
buf ( n54959 , n54958 );
not ( n54960 , n34821 );
and ( n54961 , n13361 , n14592 );
and ( n54962 , n45647 , n36348 );
and ( n54963 , n13361 , n43530 );
or ( n54964 , n54962 , n54963 );
and ( n54965 , n54964 , n14562 );
and ( n54966 , n45657 , n36347 );
and ( n54967 , n13361 , n43543 );
or ( n54968 , n54966 , n54967 );
and ( n54969 , n54968 , n14586 );
and ( n54970 , n45667 , n36348 );
and ( n54971 , n13361 , n43556 );
or ( n54972 , n54970 , n54971 );
and ( n54973 , n54972 , n14584 );
and ( n54974 , n45657 , n36347 );
and ( n54975 , n13361 , n43563 );
or ( n54976 , n54974 , n54975 );
and ( n54977 , n54976 , n37835 );
and ( n54978 , n45667 , n36347 );
and ( n54979 , n13361 , n43563 );
or ( n54980 , n54978 , n54979 );
and ( n54981 , n54980 , n37841 );
and ( n54982 , n13359 , n14564 );
and ( n54983 , n15625 , n36347 );
and ( n54984 , n13361 , n43563 );
or ( n54985 , n54983 , n54984 );
and ( n54986 , n54985 , n37847 );
or ( n54987 , n54961 , n54965 , n54969 , n54973 , n54977 , n54981 , n54982 , n54986 );
and ( n54988 , n54960 , n54987 );
and ( n54989 , n13361 , n34821 );
or ( n54990 , n54988 , n54989 );
and ( n54991 , n54990 , n16574 );
and ( n54992 , n13361 , n16576 );
or ( n54993 , n54991 , n54992 );
buf ( n54994 , n54993 );
buf ( n54995 , n54994 );
not ( n54996 , n34821 );
and ( n54997 , n43617 , n36347 );
and ( n54998 , n13339 , n39408 );
or ( n54999 , n54997 , n54998 );
and ( n55000 , n54999 , n14562 );
and ( n55001 , n43627 , n36348 );
and ( n55002 , n13339 , n39427 );
or ( n55003 , n55001 , n55002 );
and ( n55004 , n55003 , n14586 );
and ( n55005 , n43637 , n36347 );
and ( n55006 , n13339 , n39446 );
or ( n55007 , n55005 , n55006 );
and ( n55008 , n55007 , n14584 );
and ( n55009 , n43627 , n36348 );
and ( n55010 , n13339 , n39453 );
or ( n55011 , n55009 , n55010 );
and ( n55012 , n55011 , n37835 );
and ( n55013 , n43637 , n36348 );
and ( n55014 , n13339 , n39453 );
or ( n55015 , n55013 , n55014 );
and ( n55016 , n55015 , n37841 );
and ( n55017 , n15581 , n36348 );
and ( n55018 , n13339 , n39453 );
or ( n55019 , n55017 , n55018 );
and ( n55020 , n55019 , n37847 );
and ( n55021 , n13339 , n37849 );
or ( n55022 , n55000 , n55004 , n55008 , n55012 , n55016 , n55020 , n55021 );
and ( n55023 , n54996 , n55022 );
and ( n55024 , n13339 , n34821 );
or ( n55025 , n55023 , n55024 );
and ( n55026 , n55025 , n16574 );
and ( n55027 , n13339 , n16576 );
or ( n55028 , n55026 , n55027 );
buf ( n55029 , n55028 );
buf ( n55030 , n55029 );
not ( n55031 , n17451 );
and ( n55032 , n40081 , n21333 );
and ( n55033 , n20480 , n34758 );
or ( n55034 , n55032 , n55033 );
and ( n55035 , n55034 , n21341 );
and ( n55036 , n40096 , n21333 );
and ( n55037 , n20480 , n34758 );
or ( n55038 , n55036 , n55037 );
and ( n55039 , n55038 , n23064 );
and ( n55040 , n40111 , n21333 );
and ( n55041 , n20480 , n34758 );
or ( n55042 , n55040 , n55041 );
and ( n55043 , n55042 , n23825 );
and ( n55044 , n21854 , n21333 );
and ( n55045 , n20480 , n34758 );
or ( n55046 , n55044 , n55045 );
and ( n55047 , n55046 , n23832 );
and ( n55048 , n40134 , n21333 );
and ( n55049 , n20480 , n34758 );
or ( n55050 , n55048 , n55049 );
and ( n55051 , n55050 , n23917 );
and ( n55052 , n20480 , n34526 );
or ( n55053 , n55035 , n55039 , n55043 , n55047 , n55051 , n55052 );
and ( n55054 , n55031 , n55053 );
and ( n55055 , n20480 , n17451 );
or ( n55056 , n55054 , n55055 );
and ( n55057 , n55056 , n23924 );
and ( n55058 , n20480 , n23926 );
or ( n55059 , n55057 , n55058 );
buf ( n55060 , n55059 );
buf ( n55061 , n55060 );
buf ( n55062 , n10613 );
buf ( n55063 , n10615 );
buf ( n55064 , n10613 );
not ( n55065 , n34821 );
and ( n55066 , n13301 , n14592 );
and ( n55067 , n43049 , n36348 );
and ( n55068 , n13301 , n43530 );
or ( n55069 , n55067 , n55068 );
and ( n55070 , n55069 , n14562 );
and ( n55071 , n43071 , n36347 );
and ( n55072 , n13301 , n43543 );
or ( n55073 , n55071 , n55072 );
and ( n55074 , n55073 , n14586 );
and ( n55075 , n43093 , n36348 );
and ( n55076 , n13301 , n43556 );
or ( n55077 , n55075 , n55076 );
and ( n55078 , n55077 , n14584 );
and ( n55079 , n43071 , n36347 );
and ( n55080 , n13301 , n43563 );
or ( n55081 , n55079 , n55080 );
and ( n55082 , n55081 , n37835 );
and ( n55083 , n43093 , n36347 );
and ( n55084 , n13301 , n43563 );
or ( n55085 , n55083 , n55084 );
and ( n55086 , n55085 , n37841 );
and ( n55087 , n13299 , n14564 );
and ( n55088 , n15515 , n36347 );
and ( n55089 , n13301 , n43563 );
or ( n55090 , n55088 , n55089 );
and ( n55091 , n55090 , n37847 );
or ( n55092 , n55066 , n55070 , n55074 , n55078 , n55082 , n55086 , n55087 , n55091 );
and ( n55093 , n55065 , n55092 );
and ( n55094 , n13301 , n34821 );
or ( n55095 , n55093 , n55094 );
and ( n55096 , n55095 , n16574 );
and ( n55097 , n13301 , n16576 );
or ( n55098 , n55096 , n55097 );
buf ( n55099 , n55098 );
buf ( n55100 , n55099 );
buf ( n55101 , n10613 );
not ( n55102 , n24800 );
and ( n55103 , n26359 , n25222 );
and ( n55104 , n51562 , n28583 );
and ( n55105 , n26359 , n28591 );
or ( n55106 , n55104 , n55105 );
and ( n55107 , n55106 , n28594 );
and ( n55108 , n51572 , n28583 );
and ( n55109 , n26359 , n28591 );
or ( n55110 , n55108 , n55109 );
and ( n55111 , n55110 , n30269 );
and ( n55112 , n51582 , n28583 );
and ( n55113 , n26359 , n28591 );
or ( n55114 , n55112 , n55113 );
and ( n55115 , n55114 , n30982 );
and ( n55116 , n29375 , n28583 );
and ( n55117 , n26359 , n28591 );
or ( n55118 , n55116 , n55117 );
and ( n55119 , n55118 , n30989 );
and ( n55120 , n26357 , n30991 );
and ( n55121 , n51592 , n28583 );
and ( n55122 , n26359 , n28591 );
or ( n55123 , n55121 , n55122 );
and ( n55124 , n55123 , n31002 );
or ( n55125 , n55103 , n55107 , n55111 , n55115 , n55119 , n55120 , n55124 );
and ( n55126 , n55102 , n55125 );
and ( n55127 , n26359 , n24800 );
or ( n55128 , n55126 , n55127 );
and ( n55129 , n55128 , n31008 );
and ( n55130 , n26359 , n10618 );
or ( n55131 , n55129 , n55130 );
buf ( n55132 , n55131 );
buf ( n55133 , n55132 );
buf ( n55134 , n10613 );
buf ( n55135 , n10615 );
not ( n55136 , n34821 );
and ( n55137 , n13474 , n14592 );
and ( n55138 , n44175 , n36348 );
and ( n55139 , n13474 , n43530 );
or ( n55140 , n55138 , n55139 );
and ( n55141 , n55140 , n14562 );
and ( n55142 , n44185 , n36347 );
and ( n55143 , n13474 , n43543 );
or ( n55144 , n55142 , n55143 );
and ( n55145 , n55144 , n14586 );
and ( n55146 , n44195 , n36348 );
and ( n55147 , n13474 , n43556 );
or ( n55148 , n55146 , n55147 );
and ( n55149 , n55148 , n14584 );
and ( n55150 , n44185 , n36347 );
and ( n55151 , n13474 , n43563 );
or ( n55152 , n55150 , n55151 );
and ( n55153 , n55152 , n37835 );
and ( n55154 , n44195 , n36347 );
and ( n55155 , n13474 , n43563 );
or ( n55156 , n55154 , n55155 );
and ( n55157 , n55156 , n37841 );
and ( n55158 , n13472 , n14564 );
and ( n55159 , n15823 , n36347 );
and ( n55160 , n13474 , n43563 );
or ( n55161 , n55159 , n55160 );
and ( n55162 , n55161 , n37847 );
or ( n55163 , n55137 , n55141 , n55145 , n55149 , n55153 , n55157 , n55158 , n55162 );
and ( n55164 , n55136 , n55163 );
and ( n55165 , n13474 , n34821 );
or ( n55166 , n55164 , n55165 );
and ( n55167 , n55166 , n16574 );
and ( n55168 , n13474 , n16576 );
or ( n55169 , n55167 , n55168 );
buf ( n55170 , n55169 );
buf ( n55171 , n55170 );
buf ( n55172 , n10615 );
buf ( n55173 , n10613 );
and ( n55174 , n11609 , n16574 );
and ( n55175 , n15616 , n16576 );
or ( n55176 , n55174 , n55175 );
buf ( n55177 , n55176 );
buf ( n55178 , n55177 );
not ( n55179 , n34821 );
and ( n55180 , n49057 , n36345 );
and ( n55181 , n13173 , n36352 );
or ( n55182 , n55180 , n55181 );
and ( n55183 , n55182 , n14562 );
and ( n55184 , n49067 , n36345 );
and ( n55185 , n13173 , n37073 );
or ( n55186 , n55184 , n55185 );
and ( n55187 , n55186 , n14586 );
and ( n55188 , n49077 , n36350 );
and ( n55189 , n13173 , n37825 );
or ( n55190 , n55188 , n55189 );
and ( n55191 , n55190 , n14584 );
and ( n55192 , n49067 , n36350 );
and ( n55193 , n13173 , n37831 );
or ( n55194 , n55192 , n55193 );
and ( n55195 , n55194 , n37835 );
and ( n55196 , n49077 , n36350 );
and ( n55197 , n13173 , n37831 );
or ( n55198 , n55196 , n55197 );
and ( n55199 , n55198 , n37841 );
and ( n55200 , n15007 , n36350 );
and ( n55201 , n13173 , n37831 );
or ( n55202 , n55200 , n55201 );
and ( n55203 , n55202 , n37847 );
and ( n55204 , n13173 , n37849 );
or ( n55205 , n55183 , n55187 , n55191 , n55195 , n55199 , n55203 , n55204 );
and ( n55206 , n55179 , n55205 );
and ( n55207 , n13173 , n34821 );
or ( n55208 , n55206 , n55207 );
and ( n55209 , n55208 , n16574 );
and ( n55210 , n13173 , n16576 );
or ( n55211 , n55209 , n55210 );
buf ( n55212 , n55211 );
buf ( n55213 , n55212 );
not ( n55214 , n17451 );
and ( n55215 , n19283 , n17873 );
and ( n55216 , n47038 , n21330 );
and ( n55217 , n19283 , n21338 );
or ( n55218 , n55216 , n55217 );
and ( n55219 , n55218 , n21341 );
and ( n55220 , n47048 , n21330 );
and ( n55221 , n19283 , n21338 );
or ( n55222 , n55220 , n55221 );
and ( n55223 , n55222 , n23064 );
and ( n55224 , n47058 , n21330 );
and ( n55225 , n19283 , n21338 );
or ( n55226 , n55224 , n55225 );
and ( n55227 , n55226 , n23825 );
and ( n55228 , n21945 , n21330 );
and ( n55229 , n19283 , n21338 );
or ( n55230 , n55228 , n55229 );
and ( n55231 , n55230 , n23832 );
and ( n55232 , n19281 , n23834 );
and ( n55233 , n47068 , n21330 );
and ( n55234 , n19283 , n21338 );
or ( n55235 , n55233 , n55234 );
and ( n55236 , n55235 , n23917 );
or ( n55237 , n55215 , n55219 , n55223 , n55227 , n55231 , n55232 , n55236 );
and ( n55238 , n55214 , n55237 );
and ( n55239 , n19283 , n17451 );
or ( n55240 , n55238 , n55239 );
and ( n55241 , n55240 , n23924 );
and ( n55242 , n19283 , n23926 );
or ( n55243 , n55241 , n55242 );
buf ( n55244 , n55243 );
buf ( n55245 , n55244 );
buf ( n55246 , n10613 );
buf ( n55247 , n10615 );
buf ( n55248 , n10615 );
buf ( n55249 , n10615 );
buf ( n55250 , n10613 );
buf ( n55251 , n10615 );
buf ( n55252 , n10613 );
buf ( n55253 , n10615 );
buf ( n55254 , n10613 );
not ( n55255 , n24800 );
and ( n55256 , n49846 , n28587 );
and ( n55257 , n26125 , n39807 );
or ( n55258 , n55256 , n55257 );
and ( n55259 , n55258 , n28594 );
and ( n55260 , n49856 , n28587 );
and ( n55261 , n26125 , n39807 );
or ( n55262 , n55260 , n55261 );
and ( n55263 , n55262 , n30269 );
and ( n55264 , n49866 , n28587 );
and ( n55265 , n26125 , n39807 );
or ( n55266 , n55264 , n55265 );
and ( n55267 , n55266 , n30982 );
and ( n55268 , n29515 , n28587 );
and ( n55269 , n26125 , n39807 );
or ( n55270 , n55268 , n55269 );
and ( n55271 , n55270 , n30989 );
and ( n55272 , n49876 , n28587 );
and ( n55273 , n26125 , n39807 );
or ( n55274 , n55272 , n55273 );
and ( n55275 , n55274 , n31002 );
and ( n55276 , n26125 , n34607 );
or ( n55277 , n55259 , n55263 , n55267 , n55271 , n55275 , n55276 );
and ( n55278 , n55255 , n55277 );
and ( n55279 , n26125 , n24800 );
or ( n55280 , n55278 , n55279 );
and ( n55281 , n55280 , n31008 );
and ( n55282 , n26125 , n10618 );
or ( n55283 , n55281 , n55282 );
buf ( n55284 , n55283 );
buf ( n55285 , n55284 );
not ( n55286 , n17451 );
and ( n55287 , n34353 , n21333 );
and ( n55288 , n18508 , n34758 );
or ( n55289 , n55287 , n55288 );
and ( n55290 , n55289 , n21341 );
and ( n55291 , n34363 , n21333 );
and ( n55292 , n18508 , n34758 );
or ( n55293 , n55291 , n55292 );
and ( n55294 , n55293 , n23064 );
and ( n55295 , n34373 , n21333 );
and ( n55296 , n18508 , n34758 );
or ( n55297 , n55295 , n55296 );
and ( n55298 , n55297 , n23825 );
and ( n55299 , n21639 , n21333 );
and ( n55300 , n18508 , n34758 );
or ( n55301 , n55299 , n55300 );
and ( n55302 , n55301 , n23832 );
and ( n55303 , n34383 , n21333 );
and ( n55304 , n18508 , n34758 );
or ( n55305 , n55303 , n55304 );
and ( n55306 , n55305 , n23917 );
and ( n55307 , n18508 , n34526 );
or ( n55308 , n55290 , n55294 , n55298 , n55302 , n55306 , n55307 );
and ( n55309 , n55286 , n55308 );
and ( n55310 , n18508 , n17451 );
or ( n55311 , n55309 , n55310 );
and ( n55312 , n55311 , n23924 );
and ( n55313 , n18508 , n23926 );
or ( n55314 , n55312 , n55313 );
buf ( n55315 , n55314 );
buf ( n55316 , n55315 );
buf ( n55317 , n10615 );
buf ( n55318 , n10613 );
not ( n55319 , n24800 );
and ( n55320 , n45088 , n28586 );
and ( n55321 , n26293 , n34573 );
or ( n55322 , n55320 , n55321 );
and ( n55323 , n55322 , n28594 );
and ( n55324 , n45098 , n28586 );
and ( n55325 , n26293 , n34573 );
or ( n55326 , n55324 , n55325 );
and ( n55327 , n55326 , n30269 );
and ( n55328 , n45108 , n28586 );
and ( n55329 , n26293 , n34573 );
or ( n55330 , n55328 , n55329 );
and ( n55331 , n55330 , n30982 );
and ( n55332 , n29415 , n28586 );
and ( n55333 , n26293 , n34573 );
or ( n55334 , n55332 , n55333 );
and ( n55335 , n55334 , n30989 );
and ( n55336 , n45119 , n28586 );
and ( n55337 , n26293 , n34573 );
or ( n55338 , n55336 , n55337 );
and ( n55339 , n55338 , n31002 );
and ( n55340 , n26293 , n34607 );
or ( n55341 , n55323 , n55327 , n55331 , n55335 , n55339 , n55340 );
and ( n55342 , n55319 , n55341 );
and ( n55343 , n26293 , n24800 );
or ( n55344 , n55342 , n55343 );
and ( n55345 , n55344 , n31008 );
and ( n55346 , n26293 , n10618 );
or ( n55347 , n55345 , n55346 );
buf ( n55348 , n55347 );
buf ( n55349 , n55348 );
not ( n55350 , n34821 );
and ( n55351 , n13205 , n14592 );
and ( n55352 , n47932 , n36348 );
and ( n55353 , n13205 , n43530 );
or ( n55354 , n55352 , n55353 );
and ( n55355 , n55354 , n14562 );
and ( n55356 , n47942 , n36347 );
and ( n55357 , n13205 , n43543 );
or ( n55358 , n55356 , n55357 );
and ( n55359 , n55358 , n14586 );
and ( n55360 , n47952 , n36348 );
and ( n55361 , n13205 , n43556 );
or ( n55362 , n55360 , n55361 );
and ( n55363 , n55362 , n14584 );
and ( n55364 , n47942 , n36347 );
and ( n55365 , n13205 , n43563 );
or ( n55366 , n55364 , n55365 );
and ( n55367 , n55366 , n37835 );
and ( n55368 , n47952 , n36347 );
and ( n55369 , n13205 , n43563 );
or ( n55370 , n55368 , n55369 );
and ( n55371 , n55370 , n37841 );
and ( n55372 , n13203 , n14564 );
and ( n55373 , n15052 , n36347 );
and ( n55374 , n13205 , n43563 );
or ( n55375 , n55373 , n55374 );
and ( n55376 , n55375 , n37847 );
or ( n55377 , n55351 , n55355 , n55359 , n55363 , n55367 , n55371 , n55372 , n55376 );
and ( n55378 , n55350 , n55377 );
and ( n55379 , n13205 , n34821 );
or ( n55380 , n55378 , n55379 );
and ( n55381 , n55380 , n16574 );
and ( n55382 , n13205 , n16576 );
or ( n55383 , n55381 , n55382 );
buf ( n55384 , n55383 );
buf ( n55385 , n55384 );
not ( n55386 , n34821 );
and ( n55387 , n13508 , n14592 );
and ( n55388 , n53772 , n36348 );
and ( n55389 , n13508 , n43530 );
or ( n55390 , n55388 , n55389 );
and ( n55391 , n55390 , n14562 );
and ( n55392 , n53782 , n36347 );
and ( n55393 , n13508 , n43543 );
or ( n55394 , n55392 , n55393 );
and ( n55395 , n55394 , n14586 );
and ( n55396 , n53792 , n36348 );
and ( n55397 , n13508 , n43556 );
or ( n55398 , n55396 , n55397 );
and ( n55399 , n55398 , n14584 );
and ( n55400 , n53782 , n36347 );
and ( n55401 , n13508 , n43563 );
or ( n55402 , n55400 , n55401 );
and ( n55403 , n55402 , n37835 );
and ( n55404 , n53792 , n36347 );
and ( n55405 , n13508 , n43563 );
or ( n55406 , n55404 , n55405 );
and ( n55407 , n55406 , n37841 );
and ( n55408 , n13506 , n14564 );
and ( n55409 , n15866 , n36347 );
and ( n55410 , n13508 , n43563 );
or ( n55411 , n55409 , n55410 );
and ( n55412 , n55411 , n37847 );
or ( n55413 , n55387 , n55391 , n55395 , n55399 , n55403 , n55407 , n55408 , n55412 );
and ( n55414 , n55386 , n55413 );
and ( n55415 , n13508 , n34821 );
or ( n55416 , n55414 , n55415 );
and ( n55417 , n55416 , n16574 );
and ( n55418 , n13508 , n16576 );
or ( n55419 , n55417 , n55418 );
buf ( n55420 , n55419 );
buf ( n55421 , n55420 );
not ( n55422 , n34821 );
and ( n55423 , n48401 , n36345 );
and ( n55424 , n13401 , n36352 );
or ( n55425 , n55423 , n55424 );
and ( n55426 , n55425 , n14562 );
and ( n55427 , n48411 , n36345 );
and ( n55428 , n13401 , n37073 );
or ( n55429 , n55427 , n55428 );
and ( n55430 , n55429 , n14586 );
and ( n55431 , n48421 , n36350 );
and ( n55432 , n13401 , n37825 );
or ( n55433 , n55431 , n55432 );
and ( n55434 , n55433 , n14584 );
and ( n55435 , n48411 , n36350 );
and ( n55436 , n13401 , n37831 );
or ( n55437 , n55435 , n55436 );
and ( n55438 , n55437 , n37835 );
and ( n55439 , n48421 , n36350 );
and ( n55440 , n13401 , n37831 );
or ( n55441 , n55439 , n55440 );
and ( n55442 , n55441 , n37841 );
and ( n55443 , n15691 , n36350 );
and ( n55444 , n13401 , n37831 );
or ( n55445 , n55443 , n55444 );
and ( n55446 , n55445 , n37847 );
and ( n55447 , n13401 , n37849 );
or ( n55448 , n55426 , n55430 , n55434 , n55438 , n55442 , n55446 , n55447 );
and ( n55449 , n55422 , n55448 );
and ( n55450 , n13401 , n34821 );
or ( n55451 , n55449 , n55450 );
and ( n55452 , n55451 , n16574 );
and ( n55453 , n13401 , n16576 );
or ( n55454 , n55452 , n55453 );
buf ( n55455 , n55454 );
buf ( n55456 , n55455 );
buf ( n55457 , n10613 );
buf ( n55458 , n10613 );
buf ( n55459 , n10613 );
and ( n55460 , n16761 , n23924 );
and ( n55461 , n22053 , n23926 );
or ( n55462 , n55460 , n55461 );
buf ( n55463 , n55462 );
buf ( n55464 , n55463 );
not ( n55465 , n24800 );
and ( n55466 , n37895 , n28587 );
and ( n55467 , n26091 , n39807 );
or ( n55468 , n55466 , n55467 );
and ( n55469 , n55468 , n28594 );
and ( n55470 , n37905 , n28587 );
and ( n55471 , n26091 , n39807 );
or ( n55472 , n55470 , n55471 );
and ( n55473 , n55472 , n30269 );
and ( n55474 , n37915 , n28587 );
and ( n55475 , n26091 , n39807 );
or ( n55476 , n55474 , n55475 );
and ( n55477 , n55476 , n30982 );
and ( n55478 , n29535 , n28587 );
and ( n55479 , n26091 , n39807 );
or ( n55480 , n55478 , n55479 );
and ( n55481 , n55480 , n30989 );
and ( n55482 , n37925 , n28587 );
and ( n55483 , n26091 , n39807 );
or ( n55484 , n55482 , n55483 );
and ( n55485 , n55484 , n31002 );
and ( n55486 , n26091 , n34607 );
or ( n55487 , n55469 , n55473 , n55477 , n55481 , n55485 , n55486 );
and ( n55488 , n55465 , n55487 );
and ( n55489 , n26091 , n24800 );
or ( n55490 , n55488 , n55489 );
and ( n55491 , n55490 , n31008 );
and ( n55492 , n26091 , n10618 );
or ( n55493 , n55491 , n55492 );
buf ( n55494 , n55493 );
buf ( n55495 , n55494 );
not ( n55496 , n17451 );
and ( n55497 , n48746 , n21333 );
and ( n55498 , n20492 , n34758 );
or ( n55499 , n55497 , n55498 );
and ( n55500 , n55499 , n21341 );
and ( n55501 , n48756 , n21333 );
and ( n55502 , n20492 , n34758 );
or ( n55503 , n55501 , n55502 );
and ( n55504 , n55503 , n23064 );
and ( n55505 , n48766 , n21333 );
and ( n55506 , n20492 , n34758 );
or ( n55507 , n55505 , n55506 );
and ( n55508 , n55507 , n23825 );
and ( n55509 , n21867 , n21333 );
and ( n55510 , n20492 , n34758 );
or ( n55511 , n55509 , n55510 );
and ( n55512 , n55511 , n23832 );
and ( n55513 , n48776 , n21333 );
and ( n55514 , n20492 , n34758 );
or ( n55515 , n55513 , n55514 );
and ( n55516 , n55515 , n23917 );
and ( n55517 , n20492 , n34526 );
or ( n55518 , n55500 , n55504 , n55508 , n55512 , n55516 , n55517 );
and ( n55519 , n55496 , n55518 );
and ( n55520 , n20492 , n17451 );
or ( n55521 , n55519 , n55520 );
and ( n55522 , n55521 , n23924 );
and ( n55523 , n20492 , n23926 );
or ( n55524 , n55522 , n55523 );
buf ( n55525 , n55524 );
buf ( n55526 , n55525 );
not ( n55527 , n34821 );
and ( n55528 , n13156 , n14592 );
not ( n55529 , n13916 );
and ( n55530 , n55529 , n13562 );
xor ( n55531 , n13563 , n13882 );
and ( n55532 , n55531 , n13916 );
or ( n55533 , n55530 , n55532 );
buf ( n55534 , n55533 );
and ( n55535 , n55534 , n14137 );
and ( n55536 , n55534 , n14143 );
not ( n55537 , n14139 );
and ( n55538 , n55537 , n36229 );
not ( n55539 , n36245 );
and ( n55540 , n55539 , n36241 );
xor ( n55541 , n47730 , n47733 );
and ( n55542 , n55541 , n36245 );
or ( n55543 , n55540 , n55542 );
buf ( n55544 , n55543 );
and ( n55545 , n55544 , n14139 );
or ( n55546 , n55538 , n55545 );
and ( n55547 , n55546 , n14140 );
and ( n55548 , n36229 , n14141 );
or ( n55549 , n55535 , n55536 , n55547 , n55548 );
and ( n55550 , n55549 , n36348 );
and ( n55551 , n13156 , n43530 );
or ( n55552 , n55550 , n55551 );
and ( n55553 , n55552 , n14562 );
not ( n55554 , n37048 );
and ( n55555 , n55554 , n37027 );
xor ( n55556 , n47751 , n47754 );
and ( n55557 , n55556 , n37048 );
or ( n55558 , n55555 , n55557 );
buf ( n55559 , n55558 );
and ( n55560 , n55559 , n36347 );
and ( n55561 , n13156 , n43543 );
or ( n55562 , n55560 , n55561 );
and ( n55563 , n55562 , n14586 );
not ( n55564 , n37801 );
and ( n55565 , n55564 , n37780 );
xor ( n55566 , n47767 , n47770 );
and ( n55567 , n55566 , n37801 );
or ( n55568 , n55565 , n55567 );
buf ( n55569 , n55568 );
and ( n55570 , n55569 , n36348 );
and ( n55571 , n13156 , n43556 );
or ( n55572 , n55570 , n55571 );
and ( n55573 , n55572 , n14584 );
and ( n55574 , n55559 , n36347 );
and ( n55575 , n13156 , n43563 );
or ( n55576 , n55574 , n55575 );
and ( n55577 , n55576 , n37835 );
and ( n55578 , n55569 , n36347 );
and ( n55579 , n13156 , n43563 );
or ( n55580 , n55578 , n55579 );
and ( n55581 , n55580 , n37841 );
and ( n55582 , n13154 , n14564 );
and ( n55583 , n14992 , n36347 );
and ( n55584 , n13156 , n43563 );
or ( n55585 , n55583 , n55584 );
and ( n55586 , n55585 , n37847 );
or ( n55587 , n55528 , n55553 , n55563 , n55573 , n55577 , n55581 , n55582 , n55586 );
and ( n55588 , n55527 , n55587 );
and ( n55589 , n13156 , n34821 );
or ( n55590 , n55588 , n55589 );
and ( n55591 , n55590 , n16574 );
and ( n55592 , n13156 , n16576 );
or ( n55593 , n55591 , n55592 );
buf ( n55594 , n55593 );
buf ( n55595 , n55594 );
buf ( n55596 , n10615 );
and ( n55597 , n11625 , n16574 );
and ( n55598 , n15660 , n16576 );
or ( n55599 , n55597 , n55598 );
buf ( n55600 , n55599 );
buf ( n55601 , n55600 );
buf ( n55602 , n10615 );
not ( n55603 , n34821 );
and ( n55604 , n13919 , n14137 );
and ( n55605 , n13919 , n14143 );
not ( n55606 , n14139 );
xor ( n55607 , n35275 , n35627 );
buf ( n55608 , n55607 );
and ( n55609 , n55608 , n34833 );
or ( n55610 , C0 , n55609 );
buf ( n55611 , n55610 );
and ( n55612 , n55606 , n55611 );
or ( n55613 , n55612 , C0 );
and ( n55614 , n55613 , n14140 );
and ( n55615 , n55611 , n14141 );
or ( n55616 , n55604 , n55605 , n55614 , n55615 );
and ( n55617 , n55616 , n36345 );
and ( n55618 , n14609 , n36352 );
or ( n55619 , n55617 , n55618 );
and ( n55620 , n55619 , n14562 );
and ( n55621 , n47750 , n47755 );
xor ( n55622 , C0 , n55621 );
and ( n55623 , n55622 , n37048 );
or ( n55624 , C0 , n55623 );
buf ( n55625 , n55624 );
and ( n55626 , n55625 , n36345 );
and ( n55627 , n14609 , n37073 );
or ( n55628 , n55626 , n55627 );
and ( n55629 , n55628 , n14586 );
and ( n55630 , n47766 , n47771 );
xor ( n55631 , C0 , n55630 );
and ( n55632 , n55631 , n37801 );
or ( n55633 , C0 , n55632 );
buf ( n55634 , n55633 );
and ( n55635 , n55634 , n36350 );
and ( n55636 , n14609 , n37825 );
or ( n55637 , n55635 , n55636 );
and ( n55638 , n55637 , n14584 );
and ( n55639 , n55625 , n36350 );
and ( n55640 , n14609 , n37831 );
or ( n55641 , n55639 , n55640 );
and ( n55642 , n55641 , n37835 );
and ( n55643 , n55634 , n36350 );
and ( n55644 , n14609 , n37831 );
or ( n55645 , n55643 , n55644 );
and ( n55646 , n55645 , n37841 );
and ( n55647 , n14952 , n36350 );
and ( n55648 , n14609 , n37831 );
or ( n55649 , n55647 , n55648 );
and ( n55650 , n55649 , n37847 );
and ( n55651 , n14609 , n37849 );
or ( n55652 , n55620 , n55629 , n55638 , n55642 , n55646 , n55650 , n55651 );
and ( n55653 , n55603 , n55652 );
and ( n55654 , n14609 , n34821 );
or ( n55655 , n55653 , n55654 );
and ( n55656 , n55655 , n16574 );
and ( n55657 , n14609 , n16576 );
or ( n55658 , n55656 , n55657 );
buf ( n55659 , n55658 );
buf ( n55660 , n55659 );
buf ( n55661 , n10615 );
not ( n55662 , n11333 );
and ( n55663 , n55662 , n11108 );
xor ( n55664 , n11345 , n11357 );
and ( n55665 , n55664 , n11333 );
or ( n55666 , n55663 , n55665 );
buf ( n55667 , n55666 );
buf ( n55668 , n55667 );
not ( n55669 , n24800 );
and ( n55670 , n26733 , n25222 );
and ( n55671 , n49562 , n28583 );
and ( n55672 , n26733 , n28591 );
or ( n55673 , n55671 , n55672 );
and ( n55674 , n55673 , n28594 );
and ( n55675 , n49572 , n28583 );
and ( n55676 , n26733 , n28591 );
or ( n55677 , n55675 , n55676 );
and ( n55678 , n55677 , n30269 );
and ( n55679 , n49582 , n28583 );
and ( n55680 , n26733 , n28591 );
or ( n55681 , n55679 , n55680 );
and ( n55682 , n55681 , n30982 );
and ( n55683 , n29159 , n28583 );
and ( n55684 , n26733 , n28591 );
or ( n55685 , n55683 , n55684 );
and ( n55686 , n55685 , n30989 );
and ( n55687 , n26731 , n30991 );
and ( n55688 , n49592 , n28583 );
and ( n55689 , n26733 , n28591 );
or ( n55690 , n55688 , n55689 );
and ( n55691 , n55690 , n31002 );
or ( n55692 , n55670 , n55674 , n55678 , n55682 , n55686 , n55687 , n55691 );
and ( n55693 , n55669 , n55692 );
and ( n55694 , n26733 , n24800 );
or ( n55695 , n55693 , n55694 );
and ( n55696 , n55695 , n31008 );
and ( n55697 , n26733 , n10618 );
or ( n55698 , n55696 , n55697 );
buf ( n55699 , n55698 );
buf ( n55700 , n55699 );
buf ( n55701 , n10613 );
buf ( n55702 , n10615 );
buf ( n55703 , n10613 );
buf ( n55704 , n10613 );
buf ( n55705 , n10615 );
buf ( n55706 , n10613 );
buf ( n55707 , n10615 );
buf ( n55708 , n10613 );
buf ( n55709 , n10615 );
buf ( n55710 , n10613 );
buf ( n55711 , n10613 );
buf ( n55712 , n10613 );
not ( n55713 , n17451 );
and ( n55714 , n18705 , n17873 );
and ( n55715 , n40011 , n21330 );
and ( n55716 , n18705 , n21338 );
or ( n55717 , n55715 , n55716 );
and ( n55718 , n55717 , n21341 );
and ( n55719 , n40021 , n21330 );
and ( n55720 , n18705 , n21338 );
or ( n55721 , n55719 , n55720 );
and ( n55722 , n55721 , n23064 );
and ( n55723 , n40031 , n21330 );
and ( n55724 , n18705 , n21338 );
or ( n55725 , n55723 , n55724 );
and ( n55726 , n55725 , n23825 );
and ( n55727 , n22302 , n21330 );
and ( n55728 , n18705 , n21338 );
or ( n55729 , n55727 , n55728 );
and ( n55730 , n55729 , n23832 );
and ( n55731 , n18703 , n23834 );
and ( n55732 , n40041 , n21330 );
and ( n55733 , n18705 , n21338 );
or ( n55734 , n55732 , n55733 );
and ( n55735 , n55734 , n23917 );
or ( n55736 , n55714 , n55718 , n55722 , n55726 , n55730 , n55731 , n55735 );
and ( n55737 , n55713 , n55736 );
and ( n55738 , n18705 , n17451 );
or ( n55739 , n55737 , n55738 );
and ( n55740 , n55739 , n23924 );
and ( n55741 , n18705 , n23926 );
or ( n55742 , n55740 , n55741 );
buf ( n55743 , n55742 );
buf ( n55744 , n55743 );
buf ( n55745 , n10613 );
buf ( n55746 , n10615 );
buf ( n55747 , n10613 );
not ( n55748 , n34804 );
and ( n55749 , n55748 , n25863 );
and ( n55750 , n14833 , n34804 );
or ( n55751 , n55749 , n55750 );
and ( n55752 , n55751 , n31008 );
and ( n55753 , n14833 , n10618 );
or ( n55754 , n55752 , n55753 );
buf ( n55755 , n55754 );
buf ( n55756 , n55755 );
buf ( n55757 , n10613 );
buf ( n55758 , n10613 );
buf ( n55759 , n10615 );
buf ( n55760 , n10613 );
not ( n55761 , n34804 );
and ( n55762 , n55761 , n26025 );
and ( n55763 , n14803 , n34804 );
or ( n55764 , n55762 , n55763 );
and ( n55765 , n55764 , n31008 );
and ( n55766 , n14803 , n10618 );
or ( n55767 , n55765 , n55766 );
buf ( n55768 , n55767 );
buf ( n55769 , n55768 );
not ( n55770 , n24800 );
not ( n55771 , n26823 );
and ( n55772 , n55771 , n26819 );
xor ( n55773 , n26819 , n25877 );
and ( n55774 , n45228 , n45233 );
xor ( n55775 , n55773 , n55774 );
and ( n55776 , n55775 , n26823 );
or ( n55777 , n55772 , n55776 );
buf ( n55778 , n55777 );
and ( n55779 , n55778 , n27046 );
and ( n55780 , n55778 , n27049 );
not ( n55781 , n27051 );
not ( n55782 , n27054 );
buf ( n55783 , n27298 );
and ( n55784 , n55782 , n55783 );
xor ( n55785 , n27300 , n27875 );
buf ( n55786 , n55785 );
and ( n55787 , n55786 , n27054 );
or ( n55788 , n55784 , n55787 );
buf ( n55789 , n55788 );
and ( n55790 , n55781 , n55789 );
and ( n55791 , n45244 , n45249 );
buf ( n55792 , n55791 );
and ( n55793 , n55792 , n28494 );
or ( n55794 , C0 , n55793 );
buf ( n55795 , n55794 );
and ( n55796 , n55795 , n27051 );
or ( n55797 , n55790 , n55796 );
and ( n55798 , n55797 , n28506 );
and ( n55799 , n55789 , n28508 );
or ( n55800 , n55779 , n55780 , n55798 , n55799 );
and ( n55801 , n55800 , n28586 );
and ( n55802 , n27189 , n34573 );
or ( n55803 , n55801 , n55802 );
and ( n55804 , n55803 , n28594 );
not ( n55805 , n30249 );
and ( n55806 , n55805 , n30245 );
xor ( n55807 , n30245 , n29753 );
and ( n55808 , n45265 , n45270 );
xor ( n55809 , n55807 , n55808 );
and ( n55810 , n55809 , n30249 );
or ( n55811 , n55806 , n55810 );
buf ( n55812 , n55811 );
and ( n55813 , n55812 , n28586 );
and ( n55814 , n27189 , n34573 );
or ( n55815 , n55813 , n55814 );
and ( n55816 , n55815 , n30269 );
not ( n55817 , n30963 );
and ( n55818 , n55817 , n30959 );
xor ( n55819 , n30959 , n30467 );
and ( n55820 , n45281 , n45286 );
xor ( n55821 , n55819 , n55820 );
and ( n55822 , n55821 , n30963 );
or ( n55823 , n55818 , n55822 );
buf ( n55824 , n55823 );
and ( n55825 , n55824 , n28586 );
and ( n55826 , n27189 , n34573 );
or ( n55827 , n55825 , n55826 );
and ( n55828 , n55827 , n30982 );
and ( n55829 , n29120 , n28586 );
and ( n55830 , n27189 , n34573 );
or ( n55831 , n55829 , n55830 );
and ( n55832 , n55831 , n30989 );
xor ( n55833 , n48520 , n48521 );
buf ( n55834 , n55833 );
and ( n55835 , n55834 , n28586 );
and ( n55836 , n27189 , n34573 );
or ( n55837 , n55835 , n55836 );
and ( n55838 , n55837 , n31002 );
and ( n55839 , n27189 , n34607 );
or ( n55840 , n55804 , n55816 , n55828 , n55832 , n55838 , n55839 );
and ( n55841 , n55770 , n55840 );
and ( n55842 , n27189 , n24800 );
or ( n55843 , n55841 , n55842 );
and ( n55844 , n55843 , n31008 );
and ( n55845 , n27189 , n10618 );
or ( n55846 , n55844 , n55845 );
buf ( n55847 , n55846 );
buf ( n55848 , n55847 );
buf ( n55849 , n10613 );
buf ( n55850 , n10613 );
buf ( n55851 , n10613 );
buf ( n55852 , n10613 );
buf ( n55853 , n10615 );
buf ( n55854 , n10615 );
buf ( n55855 , n10615 );
and ( n55856 , n11784 , n16574 );
and ( n55857 , n14990 , n16576 );
or ( n55858 , n55856 , n55857 );
buf ( n55859 , n55858 );
buf ( n55860 , n55859 );
buf ( n55861 , n10615 );
not ( n55862 , n24800 );
and ( n55863 , n53614 , n28586 );
and ( n55864 , n26225 , n34573 );
or ( n55865 , n55863 , n55864 );
and ( n55866 , n55865 , n28594 );
and ( n55867 , n53624 , n28586 );
and ( n55868 , n26225 , n34573 );
or ( n55869 , n55867 , n55868 );
and ( n55870 , n55869 , n30269 );
and ( n55871 , n53634 , n28586 );
and ( n55872 , n26225 , n34573 );
or ( n55873 , n55871 , n55872 );
and ( n55874 , n55873 , n30982 );
and ( n55875 , n29455 , n28586 );
and ( n55876 , n26225 , n34573 );
or ( n55877 , n55875 , n55876 );
and ( n55878 , n55877 , n30989 );
and ( n55879 , n53645 , n28586 );
and ( n55880 , n26225 , n34573 );
or ( n55881 , n55879 , n55880 );
and ( n55882 , n55881 , n31002 );
and ( n55883 , n26225 , n34607 );
or ( n55884 , n55866 , n55870 , n55874 , n55878 , n55882 , n55883 );
and ( n55885 , n55862 , n55884 );
and ( n55886 , n26225 , n24800 );
or ( n55887 , n55885 , n55886 );
and ( n55888 , n55887 , n31008 );
and ( n55889 , n26225 , n10618 );
or ( n55890 , n55888 , n55889 );
buf ( n55891 , n55890 );
buf ( n55892 , n55891 );
buf ( n55893 , n10615 );
buf ( n55894 , n10615 );
not ( n55895 , n17162 );
not ( n55896 , n17450 );
and ( n55897 , n10713 , n37947 );
not ( n55898 , n38425 );
and ( n55899 , n55898 , n38166 );
xor ( n55900 , n38436 , n38444 );
and ( n55901 , n55900 , n38425 );
or ( n55902 , n55899 , n55901 );
buf ( n55903 , n55902 );
and ( n55904 , n55903 , n19745 );
not ( n55905 , n38934 );
and ( n55906 , n55905 , n38675 );
xor ( n55907 , n38945 , n38953 );
and ( n55908 , n55907 , n38934 );
or ( n55909 , n55906 , n55908 );
buf ( n55910 , n55909 );
and ( n55911 , n55910 , n19748 );
and ( n55912 , n22340 , n21253 );
and ( n55913 , n10713 , n21255 );
or ( n55914 , n55904 , n55911 , n55912 , n55913 );
and ( n55915 , n55914 , n38980 );
or ( n55916 , n55897 , n55915 );
and ( n55917 , n55896 , n55916 );
xor ( n55918 , C0 , n44840 );
buf ( n55919 , n55918 );
and ( n55920 , n55919 , n17450 );
or ( n55921 , n55917 , n55920 );
and ( n55922 , n55895 , n55921 );
and ( n55923 , n55914 , n17162 );
or ( n55924 , n55922 , n55923 );
and ( n55925 , n55924 , n23924 );
not ( n55926 , n39264 );
and ( n55927 , n55926 , n39050 );
xor ( n55928 , n39275 , n39283 );
and ( n55929 , n55928 , n39264 );
or ( n55930 , n55927 , n55929 );
buf ( n55931 , n55930 );
and ( n55932 , n55931 , n23926 );
or ( n55933 , n55925 , n55932 );
buf ( n55934 , n55933 );
buf ( n55935 , n55934 );
buf ( n55936 , n10615 );
not ( n55937 , n24800 );
and ( n55938 , n25887 , n25222 );
and ( n55939 , n28510 , n28589 );
and ( n55940 , n25887 , n31075 );
or ( n55941 , n55939 , n55940 );
and ( n55942 , n55941 , n28594 );
and ( n55943 , n30258 , n28589 );
and ( n55944 , n25887 , n31075 );
or ( n55945 , n55943 , n55944 );
and ( n55946 , n55945 , n30269 );
and ( n55947 , n30972 , n28589 );
and ( n55948 , n25887 , n31075 );
or ( n55949 , n55947 , n55948 );
and ( n55950 , n55949 , n30982 );
and ( n55951 , n29655 , n28589 );
and ( n55952 , n25887 , n31075 );
or ( n55953 , n55951 , n55952 );
and ( n55954 , n55953 , n30989 );
and ( n55955 , n29655 , n30991 );
and ( n55956 , n30998 , n28589 );
and ( n55957 , n25887 , n31075 );
or ( n55958 , n55956 , n55957 );
and ( n55959 , n55958 , n31002 );
or ( n55960 , n55938 , n55942 , n55946 , n55950 , n55954 , n55955 , n55959 );
and ( n55961 , n55937 , n55960 );
and ( n55962 , n25887 , n24800 );
or ( n55963 , n55961 , n55962 );
and ( n55964 , n55963 , n31008 );
and ( n55965 , n25234 , n10618 );
or ( n55966 , n55964 , n55965 );
buf ( n55967 , n55966 );
buf ( n55968 , n55967 );
buf ( n55969 , n10615 );
not ( n55970 , n17451 );
and ( n55971 , n48266 , n21333 );
and ( n55972 , n19420 , n34758 );
or ( n55973 , n55971 , n55972 );
and ( n55974 , n55973 , n21341 );
and ( n55975 , n48276 , n21333 );
and ( n55976 , n19420 , n34758 );
or ( n55977 , n55975 , n55976 );
and ( n55978 , n55977 , n23064 );
and ( n55979 , n48286 , n21333 );
and ( n55980 , n19420 , n34758 );
or ( n55981 , n55979 , n55980 );
and ( n55982 , n55981 , n23825 );
and ( n55983 , n21893 , n21333 );
and ( n55984 , n19420 , n34758 );
or ( n55985 , n55983 , n55984 );
and ( n55986 , n55985 , n23832 );
and ( n55987 , n48297 , n21333 );
and ( n55988 , n19420 , n34758 );
or ( n55989 , n55987 , n55988 );
and ( n55990 , n55989 , n23917 );
and ( n55991 , n19420 , n34526 );
or ( n55992 , n55974 , n55978 , n55982 , n55986 , n55990 , n55991 );
and ( n55993 , n55970 , n55992 );
and ( n55994 , n19420 , n17451 );
or ( n55995 , n55993 , n55994 );
and ( n55996 , n55995 , n23924 );
and ( n55997 , n19420 , n23926 );
or ( n55998 , n55996 , n55997 );
buf ( n55999 , n55998 );
buf ( n56000 , n55999 );
buf ( n56001 , n10615 );
and ( n56002 , n24166 , n31008 );
and ( n56003 , n29446 , n10618 );
or ( n56004 , n56002 , n56003 );
buf ( n56005 , n56004 );
buf ( n56006 , n56005 );
buf ( n56007 , n10615 );
not ( n56008 , n24800 );
and ( n56009 , n25870 , n25222 );
and ( n56010 , n48500 , n28583 );
and ( n56011 , n25870 , n28591 );
or ( n56012 , n56010 , n56011 );
and ( n56013 , n56012 , n28594 );
and ( n56014 , n25870 , n28591 );
buf ( n56015 , n56014 );
and ( n56016 , n56015 , n30269 );
and ( n56017 , n25870 , n28591 );
buf ( n56018 , n56017 );
and ( n56019 , n56018 , n30982 );
and ( n56020 , n29094 , n28583 );
and ( n56021 , n25870 , n28591 );
or ( n56022 , n56020 , n56021 );
and ( n56023 , n56022 , n30989 );
and ( n56024 , n48525 , n28583 );
and ( n56025 , n25870 , n28591 );
or ( n56026 , n56024 , n56025 );
and ( n56027 , n56026 , n31002 );
or ( n56028 , n56009 , n56013 , n56016 , n56019 , n56023 , C0 , n56027 );
and ( n56029 , n56008 , n56028 );
and ( n56030 , n25870 , n24800 );
or ( n56031 , n56029 , n56030 );
and ( n56032 , n56031 , n31008 );
and ( n56033 , n25870 , n10618 );
or ( n56034 , n56032 , n56033 );
buf ( n56035 , n56034 );
buf ( n56036 , n56035 );
not ( n56037 , n17451 );
and ( n56038 , n18873 , n17873 );
and ( n56039 , n42969 , n21336 );
and ( n56040 , n18873 , n42682 );
or ( n56041 , n56039 , n56040 );
and ( n56042 , n56041 , n21341 );
and ( n56043 , n42979 , n21336 );
and ( n56044 , n18873 , n42682 );
or ( n56045 , n56043 , n56044 );
and ( n56046 , n56045 , n23064 );
and ( n56047 , n42989 , n21336 );
and ( n56048 , n18873 , n42682 );
or ( n56049 , n56047 , n56048 );
and ( n56050 , n56049 , n23825 );
and ( n56051 , n22202 , n21336 );
and ( n56052 , n18873 , n42682 );
or ( n56053 , n56051 , n56052 );
and ( n56054 , n56053 , n23832 );
and ( n56055 , n22202 , n23834 );
and ( n56056 , n42999 , n21336 );
and ( n56057 , n18873 , n42682 );
or ( n56058 , n56056 , n56057 );
and ( n56059 , n56058 , n23917 );
or ( n56060 , n56038 , n56042 , n56046 , n56050 , n56054 , n56055 , n56059 );
and ( n56061 , n56037 , n56060 );
and ( n56062 , n18873 , n17451 );
or ( n56063 , n56061 , n56062 );
and ( n56064 , n56063 , n23924 );
and ( n56065 , n18035 , n23926 );
or ( n56066 , n56064 , n56065 );
buf ( n56067 , n56066 );
buf ( n56068 , n56067 );
buf ( n56069 , n10613 );
buf ( n56070 , n10613 );
buf ( n56071 , n10615 );
buf ( n56072 , n10613 );
buf ( n56073 , n10613 );
buf ( n56074 , n10613 );
not ( n56075 , n24800 );
and ( n56076 , n26051 , n25222 );
and ( n56077 , n49354 , n28589 );
and ( n56078 , n26051 , n31075 );
or ( n56079 , n56077 , n56078 );
and ( n56080 , n56079 , n28594 );
and ( n56081 , n49364 , n28589 );
and ( n56082 , n26051 , n31075 );
or ( n56083 , n56081 , n56082 );
and ( n56084 , n56083 , n30269 );
and ( n56085 , n49374 , n28589 );
and ( n56086 , n26051 , n31075 );
or ( n56087 , n56085 , n56086 );
and ( n56088 , n56087 , n30982 );
and ( n56089 , n29555 , n28589 );
and ( n56090 , n26051 , n31075 );
or ( n56091 , n56089 , n56090 );
and ( n56092 , n56091 , n30989 );
and ( n56093 , n29555 , n30991 );
and ( n56094 , n49385 , n28589 );
and ( n56095 , n26051 , n31075 );
or ( n56096 , n56094 , n56095 );
and ( n56097 , n56096 , n31002 );
or ( n56098 , n56076 , n56080 , n56084 , n56088 , n56092 , n56093 , n56097 );
and ( n56099 , n56075 , n56098 );
and ( n56100 , n26051 , n24800 );
or ( n56101 , n56099 , n56100 );
and ( n56102 , n56101 , n31008 );
and ( n56103 , n25309 , n10618 );
or ( n56104 , n56102 , n56103 );
buf ( n56105 , n56104 );
buf ( n56106 , n56105 );
buf ( n56107 , n10613 );
not ( n56108 , n34804 );
and ( n56109 , n56108 , n27193 );
and ( n56110 , n14659 , n34804 );
or ( n56111 , n56109 , n56110 );
and ( n56112 , n56111 , n31008 );
and ( n56113 , n14659 , n10618 );
or ( n56114 , n56112 , n56113 );
buf ( n56115 , n56114 );
buf ( n56116 , n56115 );
buf ( n56117 , n10615 );
not ( n56118 , n24800 );
and ( n56119 , n48500 , n28587 );
and ( n56120 , n25874 , n39807 );
or ( n56121 , n56119 , n56120 );
and ( n56122 , n56121 , n28594 );
and ( n56123 , n25874 , n39807 );
buf ( n56124 , n56123 );
and ( n56125 , n56124 , n30269 );
and ( n56126 , n25874 , n39807 );
buf ( n56127 , n56126 );
and ( n56128 , n56127 , n30982 );
and ( n56129 , n29094 , n28587 );
and ( n56130 , n25874 , n39807 );
or ( n56131 , n56129 , n56130 );
and ( n56132 , n56131 , n30989 );
and ( n56133 , n48525 , n28587 );
and ( n56134 , n25874 , n39807 );
or ( n56135 , n56133 , n56134 );
and ( n56136 , n56135 , n31002 );
and ( n56137 , n25874 , n34607 );
or ( n56138 , n56122 , n56125 , n56128 , n56132 , n56136 , n56137 );
and ( n56139 , n56118 , n56138 );
and ( n56140 , n25874 , n24800 );
or ( n56141 , n56139 , n56140 );
and ( n56142 , n56141 , n31008 );
and ( n56143 , n25874 , n10618 );
or ( n56144 , n56142 , n56143 );
buf ( n56145 , n56144 );
buf ( n56146 , n56145 );
buf ( n56147 , n10613 );
and ( n56148 , n24134 , n31008 );
and ( n56149 , n29366 , n10618 );
or ( n56150 , n56148 , n56149 );
buf ( n56151 , n56150 );
buf ( n56152 , n56151 );
buf ( n56153 , n10615 );
buf ( n56154 , n10615 );
buf ( n56155 , n10615 );
and ( n56156 , n17000 , n23924 );
and ( n56157 , n21891 , n23926 );
or ( n56158 , n56156 , n56157 );
buf ( n56159 , n56158 );
buf ( n56160 , n56159 );
buf ( n56161 , n10613 );
buf ( n56162 , n10615 );
buf ( n56163 , n10613 );
buf ( n56164 , n10613 );
not ( n56165 , n17451 );
and ( n56166 , n18943 , n17873 );
and ( n56167 , n42746 , n21330 );
and ( n56168 , n18943 , n21338 );
or ( n56169 , n56167 , n56168 );
and ( n56170 , n56169 , n21341 );
and ( n56171 , n42756 , n21330 );
and ( n56172 , n18943 , n21338 );
or ( n56173 , n56171 , n56172 );
and ( n56174 , n56173 , n23064 );
and ( n56175 , n42766 , n21330 );
and ( n56176 , n18943 , n21338 );
or ( n56177 , n56175 , n56176 );
and ( n56178 , n56177 , n23825 );
and ( n56179 , n22162 , n21330 );
and ( n56180 , n18943 , n21338 );
or ( n56181 , n56179 , n56180 );
and ( n56182 , n56181 , n23832 );
and ( n56183 , n18941 , n23834 );
and ( n56184 , n42776 , n21330 );
and ( n56185 , n18943 , n21338 );
or ( n56186 , n56184 , n56185 );
and ( n56187 , n56186 , n23917 );
or ( n56188 , n56166 , n56170 , n56174 , n56178 , n56182 , n56183 , n56187 );
and ( n56189 , n56165 , n56188 );
and ( n56190 , n18943 , n17451 );
or ( n56191 , n56189 , n56190 );
and ( n56192 , n56191 , n23924 );
and ( n56193 , n18943 , n23926 );
or ( n56194 , n56192 , n56193 );
buf ( n56195 , n56194 );
buf ( n56196 , n56195 );
buf ( n56197 , n10615 );
buf ( n56198 , n10615 );
buf ( n56199 , n10615 );
buf ( n56200 , n10613 );
buf ( n56201 , n10615 );
not ( n56202 , n34821 );
and ( n56203 , n47932 , n36347 );
and ( n56204 , n13207 , n39408 );
or ( n56205 , n56203 , n56204 );
and ( n56206 , n56205 , n14562 );
and ( n56207 , n47942 , n36348 );
and ( n56208 , n13207 , n39427 );
or ( n56209 , n56207 , n56208 );
and ( n56210 , n56209 , n14586 );
and ( n56211 , n47952 , n36347 );
and ( n56212 , n13207 , n39446 );
or ( n56213 , n56211 , n56212 );
and ( n56214 , n56213 , n14584 );
and ( n56215 , n47942 , n36348 );
and ( n56216 , n13207 , n39453 );
or ( n56217 , n56215 , n56216 );
and ( n56218 , n56217 , n37835 );
and ( n56219 , n47952 , n36348 );
and ( n56220 , n13207 , n39453 );
or ( n56221 , n56219 , n56220 );
and ( n56222 , n56221 , n37841 );
and ( n56223 , n15052 , n36348 );
and ( n56224 , n13207 , n39453 );
or ( n56225 , n56223 , n56224 );
and ( n56226 , n56225 , n37847 );
and ( n56227 , n13207 , n37849 );
or ( n56228 , n56206 , n56210 , n56214 , n56218 , n56222 , n56226 , n56227 );
and ( n56229 , n56202 , n56228 );
and ( n56230 , n13207 , n34821 );
or ( n56231 , n56229 , n56230 );
and ( n56232 , n56231 , n16574 );
and ( n56233 , n13207 , n16576 );
or ( n56234 , n56232 , n56233 );
buf ( n56235 , n56234 );
buf ( n56236 , n56235 );
buf ( n56237 , n10615 );
buf ( n56238 , n10615 );
buf ( n56239 , n10615 );
buf ( n56240 , n10615 );
buf ( n56241 , n10613 );
not ( n56242 , n24800 );
and ( n56243 , n55800 , n28587 );
and ( n56244 , n27191 , n39807 );
or ( n56245 , n56243 , n56244 );
and ( n56246 , n56245 , n28594 );
and ( n56247 , n55812 , n28587 );
and ( n56248 , n27191 , n39807 );
or ( n56249 , n56247 , n56248 );
and ( n56250 , n56249 , n30269 );
and ( n56251 , n55824 , n28587 );
and ( n56252 , n27191 , n39807 );
or ( n56253 , n56251 , n56252 );
and ( n56254 , n56253 , n30982 );
and ( n56255 , n29120 , n28587 );
and ( n56256 , n27191 , n39807 );
or ( n56257 , n56255 , n56256 );
and ( n56258 , n56257 , n30989 );
and ( n56259 , n55834 , n28587 );
and ( n56260 , n27191 , n39807 );
or ( n56261 , n56259 , n56260 );
and ( n56262 , n56261 , n31002 );
and ( n56263 , n27191 , n34607 );
or ( n56264 , n56246 , n56250 , n56254 , n56258 , n56262 , n56263 );
and ( n56265 , n56242 , n56264 );
and ( n56266 , n27191 , n24800 );
or ( n56267 , n56265 , n56266 );
and ( n56268 , n56267 , n31008 );
and ( n56269 , n27191 , n10618 );
or ( n56270 , n56268 , n56269 );
buf ( n56271 , n56270 );
buf ( n56272 , n56271 );
buf ( n56273 , n10615 );
buf ( n56274 , n10613 );
not ( n56275 , n17451 );
and ( n56276 , n19384 , n17873 );
and ( n56277 , n39876 , n21330 );
and ( n56278 , n19384 , n21338 );
or ( n56279 , n56277 , n56278 );
and ( n56280 , n56279 , n21341 );
and ( n56281 , n39888 , n21330 );
and ( n56282 , n19384 , n21338 );
or ( n56283 , n56281 , n56282 );
and ( n56284 , n56283 , n23064 );
and ( n56285 , n39900 , n21330 );
and ( n56286 , n19384 , n21338 );
or ( n56287 , n56285 , n56286 );
and ( n56288 , n56287 , n23825 );
and ( n56289 , n21906 , n21330 );
and ( n56290 , n19384 , n21338 );
or ( n56291 , n56289 , n56290 );
and ( n56292 , n56291 , n23832 );
and ( n56293 , n19382 , n23834 );
and ( n56294 , n39913 , n21330 );
and ( n56295 , n19384 , n21338 );
or ( n56296 , n56294 , n56295 );
and ( n56297 , n56296 , n23917 );
or ( n56298 , n56276 , n56280 , n56284 , n56288 , n56292 , n56293 , n56297 );
and ( n56299 , n56275 , n56298 );
and ( n56300 , n19384 , n17451 );
or ( n56301 , n56299 , n56300 );
and ( n56302 , n56301 , n23924 );
and ( n56303 , n19384 , n23926 );
or ( n56304 , n56302 , n56303 );
buf ( n56305 , n56304 );
buf ( n56306 , n56305 );
buf ( n56307 , n10613 );
buf ( n56308 , n10615 );
buf ( n56309 , n10615 );
buf ( n56310 , n10613 );
buf ( n56311 , n10613 );
buf ( n56312 , n10613 );
not ( n56313 , n34804 );
and ( n56314 , n56313 , n26705 );
and ( n56315 , n14683 , n34804 );
or ( n56316 , n56314 , n56315 );
and ( n56317 , n56316 , n31008 );
and ( n56318 , n14683 , n10618 );
or ( n56319 , n56317 , n56318 );
buf ( n56320 , n56319 );
buf ( n56321 , n56320 );
buf ( n56322 , n10615 );
buf ( n56323 , n10615 );
xor ( n56324 , n14628 , n14639 );
buf ( n56325 , RI210699c8_646);
or ( n56326 , n56324 , n56325 );
buf ( n56327 , n56326 );
buf ( n56328 , n56327 );
not ( n56329 , n34821 );
and ( n56330 , n13154 , n14592 );
and ( n56331 , n55549 , n36350 );
and ( n56332 , n13154 , n43691 );
or ( n56333 , n56331 , n56332 );
and ( n56334 , n56333 , n14562 );
and ( n56335 , n55559 , n36350 );
and ( n56336 , n13154 , n43703 );
or ( n56337 , n56335 , n56336 );
and ( n56338 , n56337 , n14586 );
and ( n56339 , n55569 , n36345 );
and ( n56340 , n13154 , n43715 );
or ( n56341 , n56339 , n56340 );
and ( n56342 , n56341 , n14584 );
and ( n56343 , n55559 , n36345 );
and ( n56344 , n13154 , n43721 );
or ( n56345 , n56343 , n56344 );
and ( n56346 , n56345 , n37835 );
and ( n56347 , n55569 , n36345 );
and ( n56348 , n13154 , n43721 );
or ( n56349 , n56347 , n56348 );
and ( n56350 , n56349 , n37841 );
and ( n56351 , n14992 , n14564 );
and ( n56352 , n14992 , n36345 );
and ( n56353 , n13154 , n43721 );
or ( n56354 , n56352 , n56353 );
and ( n56355 , n56354 , n37847 );
or ( n56356 , n56330 , n56334 , n56338 , n56342 , n56346 , n56350 , n56351 , n56355 );
and ( n56357 , n56329 , n56356 );
and ( n56358 , n13154 , n34821 );
or ( n56359 , n56357 , n56358 );
and ( n56360 , n56359 , n16574 );
and ( n56361 , n12248 , n16576 );
or ( n56362 , n56360 , n56361 );
buf ( n56363 , n56362 );
buf ( n56364 , n56363 );
buf ( n56365 , n10613 );
buf ( n56366 , n10615 );
buf ( n56367 , n10615 );
buf ( n56368 , n10613 );
buf ( n56369 , n10613 );
buf ( n56370 , n10613 );
buf ( n56371 , n10615 );
buf ( n56372 , n10613 );
buf ( n56373 , n10613 );
buf ( n56374 , n10615 );
not ( n56375 , n24800 );
and ( n56376 , n55773 , n55774 );
buf ( n56377 , n56376 );
and ( n56378 , n56377 , n26823 );
or ( n56379 , C0 , n56378 );
buf ( n56380 , n56379 );
and ( n56381 , n56380 , n27046 );
and ( n56382 , n56380 , n27049 );
not ( n56383 , n27051 );
xor ( n56384 , n27287 , n27876 );
buf ( n56385 , n56384 );
and ( n56386 , n56385 , n27054 );
or ( n56387 , C0 , n56386 );
buf ( n56388 , n56387 );
and ( n56389 , n56383 , n56388 );
or ( n56390 , n56389 , C0 );
and ( n56391 , n56390 , n28506 );
and ( n56392 , n56388 , n28508 );
or ( n56393 , n56381 , n56382 , n56391 , n56392 );
and ( n56394 , n56393 , n28587 );
and ( n56395 , n27179 , n39807 );
or ( n56396 , n56394 , n56395 );
and ( n56397 , n56396 , n28594 );
and ( n56398 , n55807 , n55808 );
buf ( n56399 , n56398 );
and ( n56400 , n56399 , n30249 );
or ( n56401 , C0 , n56400 );
buf ( n56402 , n56401 );
and ( n56403 , n56402 , n28587 );
and ( n56404 , n27179 , n39807 );
or ( n56405 , n56403 , n56404 );
and ( n56406 , n56405 , n30269 );
and ( n56407 , n55819 , n55820 );
buf ( n56408 , n56407 );
and ( n56409 , n56408 , n30963 );
or ( n56410 , C0 , n56409 );
buf ( n56411 , n56410 );
and ( n56412 , n56411 , n28587 );
and ( n56413 , n27179 , n39807 );
or ( n56414 , n56412 , n56413 );
and ( n56415 , n56414 , n30982 );
and ( n56416 , n29107 , n28587 );
and ( n56417 , n27179 , n39807 );
or ( n56418 , n56416 , n56417 );
and ( n56419 , n56418 , n30989 );
xor ( n56420 , n48518 , n48522 );
buf ( n56421 , n56420 );
and ( n56422 , n56421 , n28587 );
and ( n56423 , n27179 , n39807 );
or ( n56424 , n56422 , n56423 );
and ( n56425 , n56424 , n31002 );
and ( n56426 , n27179 , n34607 );
or ( n56427 , n56397 , n56406 , n56415 , n56419 , n56425 , n56426 );
and ( n56428 , n56375 , n56427 );
and ( n56429 , n27179 , n24800 );
or ( n56430 , n56428 , n56429 );
and ( n56431 , n56430 , n31008 );
and ( n56432 , n27179 , n10618 );
or ( n56433 , n56431 , n56432 );
buf ( n56434 , n56433 );
buf ( n56435 , n56434 );
not ( n56436 , n17162 );
not ( n56437 , n17450 );
and ( n56438 , n10688 , n37947 );
not ( n56439 , n38425 );
and ( n56440 , n56439 , n38251 );
xor ( n56441 , n38431 , n38449 );
and ( n56442 , n56441 , n38425 );
or ( n56443 , n56440 , n56442 );
buf ( n56444 , n56443 );
and ( n56445 , n56444 , n19745 );
not ( n56446 , n38934 );
and ( n56447 , n56446 , n38760 );
xor ( n56448 , n38940 , n38958 );
and ( n56449 , n56448 , n38934 );
or ( n56450 , n56447 , n56449 );
buf ( n56451 , n56450 );
and ( n56452 , n56451 , n19748 );
and ( n56453 , n22240 , n21253 );
and ( n56454 , n10688 , n21255 );
or ( n56455 , n56445 , n56452 , n56453 , n56454 );
and ( n56456 , n56455 , n38980 );
or ( n56457 , n56438 , n56456 );
and ( n56458 , n56437 , n56457 );
or ( n56459 , n56458 , C0 );
and ( n56460 , n56436 , n56459 );
and ( n56461 , n56455 , n17162 );
or ( n56462 , n56460 , n56461 );
and ( n56463 , n56462 , n23924 );
not ( n56464 , n39264 );
and ( n56465 , n56464 , n39120 );
xor ( n56466 , n39270 , n39288 );
and ( n56467 , n56466 , n39264 );
or ( n56468 , n56465 , n56467 );
buf ( n56469 , n56468 );
and ( n56470 , n56469 , n23926 );
or ( n56471 , n56463 , n56470 );
buf ( n56472 , n56471 );
buf ( n56473 , n56472 );
buf ( n56474 , n10613 );
buf ( n56475 , n10613 );
and ( n56476 , n11776 , n16574 );
and ( n56477 , n14975 , n16576 );
or ( n56478 , n56476 , n56477 );
buf ( n56479 , n56478 );
buf ( n56480 , n56479 );
not ( n56481 , n24800 );
and ( n56482 , n25985 , n25222 );
and ( n56483 , n45549 , n28583 );
and ( n56484 , n25985 , n28591 );
or ( n56485 , n56483 , n56484 );
and ( n56486 , n56485 , n28594 );
and ( n56487 , n45559 , n28583 );
and ( n56488 , n25985 , n28591 );
or ( n56489 , n56487 , n56488 );
and ( n56490 , n56489 , n30269 );
and ( n56491 , n45569 , n28583 );
and ( n56492 , n25985 , n28591 );
or ( n56493 , n56491 , n56492 );
and ( n56494 , n56493 , n30982 );
and ( n56495 , n29595 , n28583 );
and ( n56496 , n25985 , n28591 );
or ( n56497 , n56495 , n56496 );
and ( n56498 , n56497 , n30989 );
and ( n56499 , n25983 , n30991 );
and ( n56500 , n45580 , n28583 );
and ( n56501 , n25985 , n28591 );
or ( n56502 , n56500 , n56501 );
and ( n56503 , n56502 , n31002 );
or ( n56504 , n56482 , n56486 , n56490 , n56494 , n56498 , n56499 , n56503 );
and ( n56505 , n56481 , n56504 );
and ( n56506 , n25985 , n24800 );
or ( n56507 , n56505 , n56506 );
and ( n56508 , n56507 , n31008 );
and ( n56509 , n25985 , n10618 );
or ( n56510 , n56508 , n56509 );
buf ( n56511 , n56510 );
buf ( n56512 , n56511 );
not ( n56513 , n24511 );
not ( n56514 , n24799 );
and ( n56515 , n10650 , n40154 );
not ( n56516 , n40632 );
and ( n56517 , n56516 , n40594 );
xor ( n56518 , n43753 , n43756 );
and ( n56519 , n56518 , n40632 );
or ( n56520 , n56517 , n56519 );
buf ( n56521 , n56520 );
and ( n56522 , n56521 , n27046 );
not ( n56523 , n41147 );
and ( n56524 , n56523 , n41109 );
xor ( n56525 , n43768 , n43771 );
and ( n56526 , n56525 , n41147 );
or ( n56527 , n56524 , n56526 );
buf ( n56528 , n56527 );
and ( n56529 , n56528 , n27049 );
and ( n56530 , n29333 , n28506 );
and ( n56531 , n10650 , n28508 );
or ( n56532 , n56522 , n56529 , n56530 , n56531 );
and ( n56533 , n56532 , n41199 );
or ( n56534 , n56515 , n56533 );
and ( n56535 , n56514 , n56534 );
xor ( n56536 , n43831 , n43839 );
xor ( n56537 , n56536 , n43863 );
buf ( n56538 , n56537 );
and ( n56539 , n56538 , n27046 );
xor ( n56540 , n43905 , n43906 );
xor ( n56541 , n56540 , n43923 );
buf ( n56542 , n56541 );
and ( n56543 , n56542 , n27049 );
and ( n56544 , n29333 , n42306 );
or ( n56545 , n56539 , n56543 , n56544 );
buf ( n56546 , n56545 );
and ( n56547 , C1 , n56546 );
or ( n56548 , n56547 , C0 );
buf ( n56549 , n56548 );
not ( n56550 , n56549 );
buf ( n56551 , n56550 );
buf ( n56552 , n56551 );
not ( n56553 , n56552 );
and ( n56554 , C1 , n56553 );
or ( n56555 , n56554 , C0 );
buf ( n56556 , n56555 );
and ( n56557 , n56556 , n24799 );
or ( n56558 , n56535 , n56557 );
and ( n56559 , n56513 , n56558 );
and ( n56560 , n56532 , n24511 );
or ( n56561 , n56559 , n56560 );
and ( n56562 , n56561 , n31008 );
not ( n56563 , n42601 );
and ( n56564 , n56563 , n42569 );
xor ( n56565 , n43956 , n43959 );
and ( n56566 , n56565 , n42601 );
or ( n56567 , n56564 , n56566 );
buf ( n56568 , n56567 );
and ( n56569 , n56568 , n10618 );
or ( n56570 , n56562 , n56569 );
buf ( n56571 , n56570 );
buf ( n56572 , n56571 );
not ( n56573 , n34821 );
and ( n56574 , n45425 , n36345 );
and ( n56575 , n13317 , n36352 );
or ( n56576 , n56574 , n56575 );
and ( n56577 , n56576 , n14562 );
and ( n56578 , n45435 , n36345 );
and ( n56579 , n13317 , n37073 );
or ( n56580 , n56578 , n56579 );
and ( n56581 , n56580 , n14586 );
and ( n56582 , n45445 , n36350 );
and ( n56583 , n13317 , n37825 );
or ( n56584 , n56582 , n56583 );
and ( n56585 , n56584 , n14584 );
and ( n56586 , n45435 , n36350 );
and ( n56587 , n13317 , n37831 );
or ( n56588 , n56586 , n56587 );
and ( n56589 , n56588 , n37835 );
and ( n56590 , n45445 , n36350 );
and ( n56591 , n13317 , n37831 );
or ( n56592 , n56590 , n56591 );
and ( n56593 , n56592 , n37841 );
and ( n56594 , n15537 , n36350 );
and ( n56595 , n13317 , n37831 );
or ( n56596 , n56594 , n56595 );
and ( n56597 , n56596 , n37847 );
and ( n56598 , n13317 , n37849 );
or ( n56599 , n56577 , n56581 , n56585 , n56589 , n56593 , n56597 , n56598 );
and ( n56600 , n56573 , n56599 );
and ( n56601 , n13317 , n34821 );
or ( n56602 , n56600 , n56601 );
and ( n56603 , n56602 , n16574 );
and ( n56604 , n13317 , n16576 );
or ( n56605 , n56603 , n56604 );
buf ( n56606 , n56605 );
buf ( n56607 , n56606 );
not ( n56608 , n11954 );
not ( n56609 , n12243 );
and ( n56610 , n10933 , n31187 );
not ( n56611 , n31697 );
and ( n56612 , n56611 , n31404 );
xor ( n56613 , n50364 , n50367 );
and ( n56614 , n56613 , n31697 );
or ( n56615 , n56612 , n56614 );
buf ( n56616 , n56615 );
and ( n56617 , n56616 , n14140 );
not ( n56618 , n32214 );
and ( n56619 , n56618 , n31921 );
xor ( n56620 , n50391 , n50394 );
and ( n56621 , n56620 , n32214 );
or ( n56622 , n56619 , n56621 );
buf ( n56623 , n56622 );
and ( n56624 , n56623 , n14137 );
and ( n56625 , n15821 , n14143 );
and ( n56626 , n10933 , n14141 );
or ( n56627 , n56617 , n56624 , n56625 , n56626 );
and ( n56628 , n56627 , n32236 );
or ( n56629 , n56610 , n56628 );
and ( n56630 , n56609 , n56629 );
not ( n56631 , n34038 );
and ( n56632 , n56631 , n33626 );
xor ( n56633 , n50424 , n50427 );
and ( n56634 , n56633 , n34038 );
or ( n56635 , n56632 , n56634 );
buf ( n56636 , n56635 );
and ( n56637 , n56636 , n12243 );
or ( n56638 , n56630 , n56637 );
and ( n56639 , n56608 , n56638 );
and ( n56640 , n56627 , n11954 );
or ( n56641 , n56639 , n56640 );
and ( n56642 , n56641 , n16574 );
not ( n56643 , n34327 );
and ( n56644 , n56643 , n34085 );
xor ( n56645 , n50456 , n50459 );
and ( n56646 , n56645 , n34327 );
or ( n56647 , n56644 , n56646 );
buf ( n56648 , n56647 );
and ( n56649 , n56648 , n16576 );
or ( n56650 , n56642 , n56649 );
buf ( n56651 , n56650 );
buf ( n56652 , n56651 );
buf ( n56653 , n10613 );
buf ( n56654 , n10613 );
buf ( n56655 , n10615 );
not ( n56656 , n24511 );
not ( n56657 , n24799 );
and ( n56658 , n10690 , n40154 );
not ( n56659 , n40632 );
and ( n56660 , n56659 , n40458 );
xor ( n56661 , n40641 , n40659 );
and ( n56662 , n56661 , n40632 );
or ( n56663 , n56660 , n56662 );
buf ( n56664 , n56663 );
and ( n56665 , n56664 , n27046 );
not ( n56666 , n41147 );
and ( n56667 , n56666 , n40973 );
xor ( n56668 , n41156 , n41174 );
and ( n56669 , n56668 , n41147 );
or ( n56670 , n56667 , n56669 );
buf ( n56671 , n56670 );
and ( n56672 , n56671 , n27049 );
and ( n56673 , n29493 , n28506 );
and ( n56674 , n10690 , n28508 );
or ( n56675 , n56665 , n56672 , n56673 , n56674 );
and ( n56676 , n56675 , n41199 );
or ( n56677 , n56658 , n56676 );
and ( n56678 , n56657 , n56677 );
xor ( n56679 , n41612 , n41620 );
xor ( n56680 , n56679 , n41788 );
buf ( n56681 , n56680 );
and ( n56682 , n56681 , n27046 );
xor ( n56683 , n42177 , n42178 );
xor ( n56684 , n56683 , n42284 );
buf ( n56685 , n56684 );
and ( n56686 , n56685 , n27049 );
and ( n56687 , n29493 , n42306 );
or ( n56688 , n56682 , n56686 , n56687 );
buf ( n56689 , n56688 );
and ( n56690 , C1 , n56689 );
or ( n56691 , n56690 , C0 );
buf ( n56692 , n56691 );
not ( n56693 , n56692 );
buf ( n56694 , n56693 );
buf ( n56695 , n56694 );
not ( n56696 , n56695 );
and ( n56697 , C1 , n56696 );
or ( n56698 , n56697 , C0 );
buf ( n56699 , n56698 );
and ( n56700 , n56699 , n24799 );
or ( n56701 , n56678 , n56700 );
and ( n56702 , n56656 , n56701 );
and ( n56703 , n56675 , n24511 );
or ( n56704 , n56702 , n56703 );
and ( n56705 , n56704 , n31008 );
not ( n56706 , n42601 );
and ( n56707 , n56706 , n42457 );
xor ( n56708 , n42610 , n42628 );
and ( n56709 , n56708 , n42601 );
or ( n56710 , n56707 , n56709 );
buf ( n56711 , n56710 );
and ( n56712 , n56711 , n10618 );
or ( n56713 , n56705 , n56712 );
buf ( n56714 , n56713 );
buf ( n56715 , n56714 );
buf ( n56716 , n10613 );
buf ( n56717 , n10615 );
buf ( n56718 , n10615 );
buf ( n56719 , n10613 );
not ( n56720 , n24800 );
and ( n56721 , n26255 , n25222 );
and ( n56722 , n44989 , n28589 );
and ( n56723 , n26255 , n31075 );
or ( n56724 , n56722 , n56723 );
and ( n56725 , n56724 , n28594 );
and ( n56726 , n44999 , n28589 );
and ( n56727 , n26255 , n31075 );
or ( n56728 , n56726 , n56727 );
and ( n56729 , n56728 , n30269 );
and ( n56730 , n45009 , n28589 );
and ( n56731 , n26255 , n31075 );
or ( n56732 , n56730 , n56731 );
and ( n56733 , n56732 , n30982 );
and ( n56734 , n29435 , n28589 );
and ( n56735 , n26255 , n31075 );
or ( n56736 , n56734 , n56735 );
and ( n56737 , n56736 , n30989 );
and ( n56738 , n29435 , n30991 );
and ( n56739 , n45019 , n28589 );
and ( n56740 , n26255 , n31075 );
or ( n56741 , n56739 , n56740 );
and ( n56742 , n56741 , n31002 );
or ( n56743 , n56721 , n56725 , n56729 , n56733 , n56737 , n56738 , n56742 );
and ( n56744 , n56720 , n56743 );
and ( n56745 , n26255 , n24800 );
or ( n56746 , n56744 , n56745 );
and ( n56747 , n56746 , n31008 );
and ( n56748 , n25399 , n10618 );
or ( n56749 , n56747 , n56748 );
buf ( n56750 , n56749 );
buf ( n56751 , n56750 );
buf ( n56752 , n10613 );
not ( n56753 , n34821 );
and ( n56754 , n39404 , n36345 );
and ( n56755 , n13377 , n36352 );
or ( n56756 , n56754 , n56755 );
and ( n56757 , n56756 , n14562 );
and ( n56758 , n39423 , n36345 );
and ( n56759 , n13377 , n37073 );
or ( n56760 , n56758 , n56759 );
and ( n56761 , n56760 , n14586 );
and ( n56762 , n39442 , n36350 );
and ( n56763 , n13377 , n37825 );
or ( n56764 , n56762 , n56763 );
and ( n56765 , n56764 , n14584 );
and ( n56766 , n39423 , n36350 );
and ( n56767 , n13377 , n37831 );
or ( n56768 , n56766 , n56767 );
and ( n56769 , n56768 , n37835 );
and ( n56770 , n39442 , n36350 );
and ( n56771 , n13377 , n37831 );
or ( n56772 , n56770 , n56771 );
and ( n56773 , n56772 , n37841 );
and ( n56774 , n15647 , n36350 );
and ( n56775 , n13377 , n37831 );
or ( n56776 , n56774 , n56775 );
and ( n56777 , n56776 , n37847 );
and ( n56778 , n13377 , n37849 );
or ( n56779 , n56757 , n56761 , n56765 , n56769 , n56773 , n56777 , n56778 );
and ( n56780 , n56753 , n56779 );
and ( n56781 , n13377 , n34821 );
or ( n56782 , n56780 , n56781 );
and ( n56783 , n56782 , n16574 );
and ( n56784 , n13377 , n16576 );
or ( n56785 , n56783 , n56784 );
buf ( n56786 , n56785 );
buf ( n56787 , n56786 );
not ( n56788 , n11333 );
and ( n56789 , n56788 , n11227 );
xor ( n56790 , n11338 , n11364 );
and ( n56791 , n56790 , n11333 );
or ( n56792 , n56789 , n56791 );
buf ( n56793 , n56792 );
buf ( n56794 , n56793 );
buf ( n56795 , n10613 );
buf ( n56796 , n10615 );
buf ( n56797 , n10615 );
not ( n56798 , n17451 );
and ( n56799 , n34488 , n21333 );
and ( n56800 , n18843 , n34758 );
or ( n56801 , n56799 , n56800 );
and ( n56802 , n56801 , n21341 );
and ( n56803 , n34501 , n21333 );
and ( n56804 , n18843 , n34758 );
or ( n56805 , n56803 , n56804 );
and ( n56806 , n56805 , n23064 );
and ( n56807 , n34511 , n21333 );
and ( n56808 , n18843 , n34758 );
or ( n56809 , n56807 , n56808 );
and ( n56810 , n56809 , n23825 );
and ( n56811 , n22222 , n21333 );
and ( n56812 , n18843 , n34758 );
or ( n56813 , n56811 , n56812 );
and ( n56814 , n56813 , n23832 );
and ( n56815 , n34521 , n21333 );
and ( n56816 , n18843 , n34758 );
or ( n56817 , n56815 , n56816 );
and ( n56818 , n56817 , n23917 );
and ( n56819 , n18843 , n34526 );
or ( n56820 , n56802 , n56806 , n56810 , n56814 , n56818 , n56819 );
and ( n56821 , n56798 , n56820 );
and ( n56822 , n18843 , n17451 );
or ( n56823 , n56821 , n56822 );
and ( n56824 , n56823 , n23924 );
and ( n56825 , n18843 , n23926 );
or ( n56826 , n56824 , n56825 );
buf ( n56827 , n56826 );
buf ( n56828 , n56827 );
buf ( n56829 , n10613 );
buf ( n56830 , n10613 );
buf ( n56831 , n10613 );
not ( n56832 , n24800 );
and ( n56833 , n52878 , n28586 );
and ( n56834 , n26531 , n34573 );
or ( n56835 , n56833 , n56834 );
and ( n56836 , n56835 , n28594 );
and ( n56837 , n52888 , n28586 );
and ( n56838 , n26531 , n34573 );
or ( n56839 , n56837 , n56838 );
and ( n56840 , n56839 , n30269 );
and ( n56841 , n52898 , n28586 );
and ( n56842 , n26531 , n34573 );
or ( n56843 , n56841 , n56842 );
and ( n56844 , n56843 , n30982 );
and ( n56845 , n29237 , n28586 );
and ( n56846 , n26531 , n34573 );
or ( n56847 , n56845 , n56846 );
and ( n56848 , n56847 , n30989 );
and ( n56849 , n52908 , n28586 );
and ( n56850 , n26531 , n34573 );
or ( n56851 , n56849 , n56850 );
and ( n56852 , n56851 , n31002 );
and ( n56853 , n26531 , n34607 );
or ( n56854 , n56836 , n56840 , n56844 , n56848 , n56852 , n56853 );
and ( n56855 , n56832 , n56854 );
and ( n56856 , n26531 , n24800 );
or ( n56857 , n56855 , n56856 );
and ( n56858 , n56857 , n31008 );
and ( n56859 , n26531 , n10618 );
or ( n56860 , n56858 , n56859 );
buf ( n56861 , n56860 );
buf ( n56862 , n56861 );
buf ( n56863 , n10613 );
buf ( n56864 , n10615 );
buf ( n56865 , n10615 );
buf ( n56866 , n10615 );
buf ( n56867 , n10615 );
buf ( n56868 , n10615 );
buf ( n56869 , n10613 );
buf ( n56870 , n10615 );
buf ( n56871 , n10613 );
not ( n56872 , n11954 );
not ( n56873 , n12243 );
and ( n56874 , n10797 , n31187 );
not ( n56875 , n31697 );
and ( n56876 , n56875 , n31693 );
xor ( n56877 , n31693 , n31371 );
xor ( n56878 , n31676 , n31371 );
xor ( n56879 , n31659 , n31371 );
xor ( n56880 , n31642 , n31371 );
xor ( n56881 , n31625 , n31371 );
xor ( n56882 , n31608 , n31371 );
xor ( n56883 , n31591 , n31371 );
xor ( n56884 , n31574 , n31371 );
and ( n56885 , n54395 , n54396 );
and ( n56886 , n56884 , n56885 );
and ( n56887 , n56883 , n56886 );
and ( n56888 , n56882 , n56887 );
and ( n56889 , n56881 , n56888 );
and ( n56890 , n56880 , n56889 );
and ( n56891 , n56879 , n56890 );
and ( n56892 , n56878 , n56891 );
xor ( n56893 , n56877 , n56892 );
and ( n56894 , n56893 , n31697 );
or ( n56895 , n56876 , n56894 );
buf ( n56896 , n56895 );
and ( n56897 , n56896 , n14140 );
not ( n56898 , n32214 );
and ( n56899 , n56898 , n32210 );
xor ( n56900 , n32210 , n31888 );
xor ( n56901 , n32193 , n31888 );
xor ( n56902 , n32176 , n31888 );
xor ( n56903 , n32159 , n31888 );
xor ( n56904 , n32142 , n31888 );
xor ( n56905 , n32125 , n31888 );
xor ( n56906 , n32108 , n31888 );
xor ( n56907 , n32091 , n31888 );
and ( n56908 , n54404 , n54405 );
and ( n56909 , n56907 , n56908 );
and ( n56910 , n56906 , n56909 );
and ( n56911 , n56905 , n56910 );
and ( n56912 , n56904 , n56911 );
and ( n56913 , n56903 , n56912 );
and ( n56914 , n56902 , n56913 );
and ( n56915 , n56901 , n56914 );
xor ( n56916 , n56900 , n56915 );
and ( n56917 , n56916 , n32214 );
or ( n56918 , n56899 , n56917 );
buf ( n56919 , n56918 );
and ( n56920 , n56919 , n14137 );
and ( n56921 , n15447 , n14143 );
and ( n56922 , n10797 , n14141 );
or ( n56923 , n56897 , n56920 , n56921 , n56922 );
and ( n56924 , n56923 , n32236 );
or ( n56925 , n56874 , n56924 );
and ( n56926 , n56873 , n56925 );
not ( n56927 , n34038 );
and ( n56928 , n56927 , n34034 );
xor ( n56929 , n34034 , n33579 );
xor ( n56930 , n34010 , n33579 );
xor ( n56931 , n33986 , n33579 );
xor ( n56932 , n33962 , n33579 );
xor ( n56933 , n33938 , n33579 );
xor ( n56934 , n33914 , n33579 );
xor ( n56935 , n33890 , n33579 );
xor ( n56936 , n33866 , n33579 );
and ( n56937 , n54419 , n54420 );
and ( n56938 , n56936 , n56937 );
and ( n56939 , n56935 , n56938 );
and ( n56940 , n56934 , n56939 );
and ( n56941 , n56933 , n56940 );
nand ( n56942 , n56932 , n56941 );
nand ( n56943 , n56931 , n56942 );
and ( n56944 , n56930 , n56943 );
xor ( n56945 , n56929 , n56944 );
and ( n56946 , n56945 , n34038 );
or ( n56947 , n56928 , n56946 );
buf ( n56948 , n56947 );
and ( n56949 , n56948 , n12243 );
or ( n56950 , n56926 , n56949 );
and ( n56951 , n56872 , n56950 );
and ( n56952 , n56923 , n11954 );
or ( n56953 , n56951 , n56952 );
and ( n56954 , n56953 , n16574 );
not ( n56955 , n34327 );
and ( n56956 , n56955 , n34323 );
xor ( n56957 , n34323 , n34058 );
xor ( n56958 , n34309 , n34058 );
xor ( n56959 , n34295 , n34058 );
xor ( n56960 , n34281 , n34058 );
xor ( n56961 , n34267 , n34058 );
xor ( n56962 , n34253 , n34058 );
xor ( n56963 , n34239 , n34058 );
xor ( n56964 , n34225 , n34058 );
and ( n56965 , n54433 , n54434 );
and ( n56966 , n56964 , n56965 );
and ( n56967 , n56963 , n56966 );
and ( n56968 , n56962 , n56967 );
and ( n56969 , n56961 , n56968 );
and ( n56970 , n56960 , n56969 );
and ( n56971 , n56959 , n56970 );
and ( n56972 , n56958 , n56971 );
xor ( n56973 , n56957 , n56972 );
and ( n56974 , n56973 , n34327 );
or ( n56975 , n56956 , n56974 );
buf ( n56976 , n56975 );
and ( n56977 , n56976 , n16576 );
or ( n56978 , n56954 , n56977 );
buf ( n56979 , n56978 );
buf ( n56980 , n56979 );
buf ( n56981 , n10613 );
and ( n56982 , n24158 , n31008 );
and ( n56983 , n29426 , n10618 );
or ( n56984 , n56982 , n56983 );
buf ( n56985 , n56984 );
buf ( n56986 , n56985 );
buf ( n56987 , n10615 );
not ( n56988 , n34538 );
and ( n56989 , n56988 , n19051 );
and ( n56990 , n14735 , n34538 );
or ( n56991 , n56989 , n56990 );
and ( n56992 , n56991 , n23924 );
and ( n56993 , n14735 , n23926 );
or ( n56994 , n56992 , n56993 );
buf ( n56995 , n56994 );
buf ( n56996 , n56995 );
buf ( n56997 , n10613 );
buf ( n56998 , n10615 );
buf ( n56999 , n10615 );
buf ( n57000 , n10613 );
buf ( n57001 , n10615 );
buf ( n57002 , n10615 );
buf ( n57003 , n10613 );
not ( n57004 , n24800 );
and ( n57005 , n54833 , n28586 );
and ( n57006 , n26633 , n34573 );
or ( n57007 , n57005 , n57006 );
and ( n57008 , n57007 , n28594 );
and ( n57009 , n54843 , n28586 );
and ( n57010 , n26633 , n34573 );
or ( n57011 , n57009 , n57010 );
and ( n57012 , n57011 , n30269 );
and ( n57013 , n54853 , n28586 );
and ( n57014 , n26633 , n34573 );
or ( n57015 , n57013 , n57014 );
and ( n57016 , n57015 , n30982 );
and ( n57017 , n29198 , n28586 );
and ( n57018 , n26633 , n34573 );
or ( n57019 , n57017 , n57018 );
and ( n57020 , n57019 , n30989 );
and ( n57021 , n54863 , n28586 );
and ( n57022 , n26633 , n34573 );
or ( n57023 , n57021 , n57022 );
and ( n57024 , n57023 , n31002 );
and ( n57025 , n26633 , n34607 );
or ( n57026 , n57008 , n57012 , n57016 , n57020 , n57024 , n57025 );
and ( n57027 , n57004 , n57026 );
and ( n57028 , n26633 , n24800 );
or ( n57029 , n57027 , n57028 );
and ( n57030 , n57029 , n31008 );
and ( n57031 , n26633 , n10618 );
or ( n57032 , n57030 , n57031 );
buf ( n57033 , n57032 );
buf ( n57034 , n57033 );
and ( n57035 , n24142 , n31008 );
and ( n57036 , n29386 , n10618 );
or ( n57037 , n57035 , n57036 );
buf ( n57038 , n57037 );
buf ( n57039 , n57038 );
not ( n57040 , n11333 );
and ( n57041 , n57040 , n11329 );
xor ( n57042 , n11329 , n11007 );
and ( n57043 , n53857 , n53858 );
xor ( n57044 , n57042 , n57043 );
and ( n57045 , n57044 , n11333 );
or ( n57046 , n57041 , n57045 );
buf ( n57047 , n57046 );
buf ( n57048 , n57047 );
buf ( n57049 , n10615 );
not ( n57050 , n24800 );
and ( n57051 , n26459 , n25222 );
and ( n57052 , n47642 , n28589 );
and ( n57053 , n26459 , n31075 );
or ( n57054 , n57052 , n57053 );
and ( n57055 , n57054 , n28594 );
and ( n57056 , n47652 , n28589 );
and ( n57057 , n26459 , n31075 );
or ( n57058 , n57056 , n57057 );
and ( n57059 , n57058 , n30269 );
and ( n57060 , n47662 , n28589 );
and ( n57061 , n26459 , n31075 );
or ( n57062 , n57060 , n57061 );
and ( n57063 , n57062 , n30982 );
and ( n57064 , n29315 , n28589 );
and ( n57065 , n26459 , n31075 );
or ( n57066 , n57064 , n57065 );
and ( n57067 , n57066 , n30989 );
and ( n57068 , n29315 , n30991 );
and ( n57069 , n47672 , n28589 );
and ( n57070 , n26459 , n31075 );
or ( n57071 , n57069 , n57070 );
and ( n57072 , n57071 , n31002 );
or ( n57073 , n57051 , n57055 , n57059 , n57063 , n57067 , n57068 , n57072 );
and ( n57074 , n57050 , n57073 );
and ( n57075 , n26459 , n24800 );
or ( n57076 , n57074 , n57075 );
and ( n57077 , n57076 , n31008 );
and ( n57078 , n25489 , n10618 );
or ( n57079 , n57077 , n57078 );
buf ( n57080 , n57079 );
buf ( n57081 , n57080 );
buf ( n57082 , n10613 );
not ( n57083 , n24511 );
not ( n57084 , n24799 );
and ( n57085 , n10665 , n40154 );
not ( n57086 , n40632 );
and ( n57087 , n57086 , n40543 );
xor ( n57088 , n40636 , n40664 );
and ( n57089 , n57088 , n40632 );
or ( n57090 , n57087 , n57089 );
buf ( n57091 , n57090 );
and ( n57092 , n57091 , n27046 );
not ( n57093 , n41147 );
and ( n57094 , n57093 , n41058 );
xor ( n57095 , n41151 , n41179 );
and ( n57096 , n57095 , n41147 );
or ( n57097 , n57094 , n57096 );
buf ( n57098 , n57097 );
and ( n57099 , n57098 , n27049 );
and ( n57100 , n29393 , n28506 );
and ( n57101 , n10665 , n28508 );
or ( n57102 , n57092 , n57099 , n57100 , n57101 );
and ( n57103 , n57102 , n41199 );
or ( n57104 , n57085 , n57103 );
and ( n57105 , n57084 , n57104 );
xor ( n57106 , n41532 , n41540 );
xor ( n57107 , n57106 , n41803 );
buf ( n57108 , n57107 );
and ( n57109 , n57108 , n27046 );
xor ( n57110 , n42132 , n42133 );
xor ( n57111 , n57110 , n42299 );
buf ( n57112 , n57111 );
and ( n57113 , n57112 , n27049 );
and ( n57114 , n29393 , n42306 );
or ( n57115 , n57109 , n57113 , n57114 );
buf ( n57116 , n57115 );
and ( n57117 , C1 , n57116 );
or ( n57118 , n57117 , C0 );
buf ( n57119 , n57118 );
not ( n57120 , n57119 );
buf ( n57121 , n57120 );
buf ( n57122 , n57121 );
not ( n57123 , n57122 );
and ( n57124 , C1 , n57123 );
or ( n57125 , n57124 , C0 );
buf ( n57126 , n57125 );
and ( n57127 , n57126 , n24799 );
or ( n57128 , n57105 , n57127 );
and ( n57129 , n57083 , n57128 );
and ( n57130 , n57102 , n24511 );
or ( n57131 , n57129 , n57130 );
and ( n57132 , n57131 , n31008 );
not ( n57133 , n42601 );
and ( n57134 , n57133 , n42527 );
xor ( n57135 , n42605 , n42633 );
and ( n57136 , n57135 , n42601 );
or ( n57137 , n57134 , n57136 );
buf ( n57138 , n57137 );
and ( n57139 , n57138 , n10618 );
or ( n57140 , n57132 , n57139 );
buf ( n57141 , n57140 );
buf ( n57142 , n57141 );
buf ( n57143 , n10615 );
buf ( n57144 , n10613 );
and ( n57145 , n16753 , n23924 );
and ( n57146 , n21995 , n23926 );
or ( n57147 , n57145 , n57146 );
buf ( n57148 , n57147 );
buf ( n57149 , n57148 );
buf ( n57150 , n10613 );
not ( n57151 , n34804 );
and ( n57152 , n57151 , n26807 );
and ( n57153 , n14665 , n34804 );
or ( n57154 , n57152 , n57153 );
and ( n57155 , n57154 , n31008 );
and ( n57156 , n14665 , n10618 );
or ( n57157 , n57155 , n57156 );
buf ( n57158 , n57157 );
buf ( n57159 , n57158 );
buf ( n57160 , n10613 );
buf ( n57161 , n10613 );
buf ( n57162 , n10615 );
buf ( n57163 , n10613 );
buf ( n57164 , n10615 );
buf ( n57165 , n10615 );
buf ( n57166 , n10615 );
buf ( n57167 , n10615 );
buf ( n57168 , n10615 );
buf ( n57169 , n10615 );
not ( n57170 , n11954 );
not ( n57171 , n12243 );
and ( n57172 , n10853 , n31187 );
not ( n57173 , n31697 );
and ( n57174 , n57173 , n31574 );
xor ( n57175 , n56884 , n56885 );
and ( n57176 , n57175 , n31697 );
or ( n57177 , n57174 , n57176 );
buf ( n57178 , n57177 );
and ( n57179 , n57178 , n14140 );
not ( n57180 , n32214 );
and ( n57181 , n57180 , n32091 );
xor ( n57182 , n56907 , n56908 );
and ( n57183 , n57182 , n32214 );
or ( n57184 , n57181 , n57183 );
buf ( n57185 , n57184 );
and ( n57186 , n57185 , n14137 );
and ( n57187 , n15601 , n14143 );
and ( n57188 , n10853 , n14141 );
or ( n57189 , n57179 , n57186 , n57187 , n57188 );
and ( n57190 , n57189 , n32236 );
or ( n57191 , n57172 , n57190 );
and ( n57192 , n57171 , n57191 );
not ( n57193 , n34038 );
and ( n57194 , n57193 , n33866 );
xor ( n57195 , n56936 , n56937 );
and ( n57196 , n57195 , n34038 );
or ( n57197 , n57194 , n57196 );
buf ( n57198 , n57197 );
and ( n57199 , n57198 , n12243 );
or ( n57200 , n57192 , n57199 );
and ( n57201 , n57170 , n57200 );
and ( n57202 , n57189 , n11954 );
or ( n57203 , n57201 , n57202 );
and ( n57204 , n57203 , n16574 );
not ( n57205 , n34327 );
and ( n57206 , n57205 , n34225 );
xor ( n57207 , n56964 , n56965 );
and ( n57208 , n57207 , n34327 );
or ( n57209 , n57206 , n57208 );
buf ( n57210 , n57209 );
and ( n57211 , n57210 , n16576 );
or ( n57212 , n57204 , n57211 );
buf ( n57213 , n57212 );
buf ( n57214 , n57213 );
buf ( n57215 , n10613 );
not ( n57216 , n34821 );
and ( n57217 , n13419 , n14592 );
and ( n57218 , n44068 , n36350 );
and ( n57219 , n13419 , n43691 );
or ( n57220 , n57218 , n57219 );
and ( n57221 , n57220 , n14562 );
and ( n57222 , n44078 , n36350 );
and ( n57223 , n13419 , n43703 );
or ( n57224 , n57222 , n57223 );
and ( n57225 , n57224 , n14586 );
and ( n57226 , n44088 , n36345 );
and ( n57227 , n13419 , n43715 );
or ( n57228 , n57226 , n57227 );
and ( n57229 , n57228 , n14584 );
and ( n57230 , n44078 , n36345 );
and ( n57231 , n13419 , n43721 );
or ( n57232 , n57230 , n57231 );
and ( n57233 , n57232 , n37835 );
and ( n57234 , n44088 , n36345 );
and ( n57235 , n13419 , n43721 );
or ( n57236 , n57234 , n57235 );
and ( n57237 , n57236 , n37841 );
and ( n57238 , n15735 , n14564 );
and ( n57239 , n15735 , n36345 );
and ( n57240 , n13419 , n43721 );
or ( n57241 , n57239 , n57240 );
and ( n57242 , n57241 , n37847 );
or ( n57243 , n57217 , n57221 , n57225 , n57229 , n57233 , n57237 , n57238 , n57242 );
and ( n57244 , n57216 , n57243 );
and ( n57245 , n13419 , n34821 );
or ( n57246 , n57244 , n57245 );
and ( n57247 , n57246 , n16574 );
and ( n57248 , n12315 , n16576 );
or ( n57249 , n57247 , n57248 );
buf ( n57250 , n57249 );
buf ( n57251 , n57250 );
buf ( n57252 , n10615 );
buf ( n57253 , n10615 );
buf ( n57254 , n10615 );
buf ( n57255 , n10615 );
buf ( n57256 , n10613 );
not ( n57257 , n24800 );
and ( n57258 , n26527 , n25222 );
and ( n57259 , n52878 , n28589 );
and ( n57260 , n26527 , n31075 );
or ( n57261 , n57259 , n57260 );
and ( n57262 , n57261 , n28594 );
and ( n57263 , n52888 , n28589 );
and ( n57264 , n26527 , n31075 );
or ( n57265 , n57263 , n57264 );
and ( n57266 , n57265 , n30269 );
and ( n57267 , n52898 , n28589 );
and ( n57268 , n26527 , n31075 );
or ( n57269 , n57267 , n57268 );
and ( n57270 , n57269 , n30982 );
and ( n57271 , n29237 , n28589 );
and ( n57272 , n26527 , n31075 );
or ( n57273 , n57271 , n57272 );
and ( n57274 , n57273 , n30989 );
and ( n57275 , n29237 , n30991 );
and ( n57276 , n52908 , n28589 );
and ( n57277 , n26527 , n31075 );
or ( n57278 , n57276 , n57277 );
and ( n57279 , n57278 , n31002 );
or ( n57280 , n57258 , n57262 , n57266 , n57270 , n57274 , n57275 , n57279 );
and ( n57281 , n57257 , n57280 );
and ( n57282 , n26527 , n24800 );
or ( n57283 , n57281 , n57282 );
and ( n57284 , n57283 , n31008 );
and ( n57285 , n25519 , n10618 );
or ( n57286 , n57284 , n57285 );
buf ( n57287 , n57286 );
buf ( n57288 , n57287 );
buf ( n57289 , n10613 );
not ( n57290 , n34804 );
and ( n57291 , n57290 , n26739 );
and ( n57292 , n14677 , n34804 );
or ( n57293 , n57291 , n57292 );
and ( n57294 , n57293 , n31008 );
and ( n57295 , n14677 , n10618 );
or ( n57296 , n57294 , n57295 );
buf ( n57297 , n57296 );
buf ( n57298 , n57297 );
buf ( n57299 , n10615 );
not ( n57300 , n24800 );
and ( n57301 , n49354 , n28586 );
and ( n57302 , n26055 , n34573 );
or ( n57303 , n57301 , n57302 );
and ( n57304 , n57303 , n28594 );
and ( n57305 , n49364 , n28586 );
and ( n57306 , n26055 , n34573 );
or ( n57307 , n57305 , n57306 );
and ( n57308 , n57307 , n30269 );
and ( n57309 , n49374 , n28586 );
and ( n57310 , n26055 , n34573 );
or ( n57311 , n57309 , n57310 );
and ( n57312 , n57311 , n30982 );
and ( n57313 , n29555 , n28586 );
and ( n57314 , n26055 , n34573 );
or ( n57315 , n57313 , n57314 );
and ( n57316 , n57315 , n30989 );
and ( n57317 , n49385 , n28586 );
and ( n57318 , n26055 , n34573 );
or ( n57319 , n57317 , n57318 );
and ( n57320 , n57319 , n31002 );
and ( n57321 , n26055 , n34607 );
or ( n57322 , n57304 , n57308 , n57312 , n57316 , n57320 , n57321 );
and ( n57323 , n57300 , n57322 );
and ( n57324 , n26055 , n24800 );
or ( n57325 , n57323 , n57324 );
and ( n57326 , n57325 , n31008 );
and ( n57327 , n26055 , n10618 );
or ( n57328 , n57326 , n57327 );
buf ( n57329 , n57328 );
buf ( n57330 , n57329 );
and ( n57331 , n24150 , n31008 );
and ( n57332 , n29406 , n10618 );
or ( n57333 , n57331 , n57332 );
buf ( n57334 , n57333 );
buf ( n57335 , n57334 );
not ( n57336 , n34821 );
not ( n57337 , n13916 );
and ( n57338 , n57337 , n13650 );
xor ( n57339 , n13651 , n13874 );
and ( n57340 , n57339 , n13916 );
or ( n57341 , n57338 , n57340 );
buf ( n57342 , n57341 );
and ( n57343 , n57342 , n14137 );
and ( n57344 , n57342 , n14143 );
not ( n57345 , n14139 );
and ( n57346 , n57345 , n36053 );
not ( n57347 , n36245 );
and ( n57348 , n57347 , n36065 );
xor ( n57349 , n45734 , n45735 );
and ( n57350 , n57349 , n36245 );
or ( n57351 , n57348 , n57350 );
buf ( n57352 , n57351 );
and ( n57353 , n57352 , n14139 );
or ( n57354 , n57346 , n57353 );
and ( n57355 , n57354 , n14140 );
and ( n57356 , n36053 , n14141 );
or ( n57357 , n57343 , n57344 , n57355 , n57356 );
and ( n57358 , n57357 , n36347 );
and ( n57359 , n13255 , n39408 );
or ( n57360 , n57358 , n57359 );
and ( n57361 , n57360 , n14562 );
not ( n57362 , n37048 );
and ( n57363 , n57362 , n36891 );
xor ( n57364 , n45755 , n45756 );
and ( n57365 , n57364 , n37048 );
or ( n57366 , n57363 , n57365 );
buf ( n57367 , n57366 );
and ( n57368 , n57367 , n36348 );
and ( n57369 , n13255 , n39427 );
or ( n57370 , n57368 , n57369 );
and ( n57371 , n57370 , n14586 );
not ( n57372 , n37801 );
and ( n57373 , n57372 , n37644 );
xor ( n57374 , n45771 , n45772 );
and ( n57375 , n57374 , n37801 );
or ( n57376 , n57373 , n57375 );
buf ( n57377 , n57376 );
and ( n57378 , n57377 , n36347 );
and ( n57379 , n13255 , n39446 );
or ( n57380 , n57378 , n57379 );
and ( n57381 , n57380 , n14584 );
and ( n57382 , n57367 , n36348 );
and ( n57383 , n13255 , n39453 );
or ( n57384 , n57382 , n57383 );
and ( n57385 , n57384 , n37835 );
and ( n57386 , n57377 , n36348 );
and ( n57387 , n13255 , n39453 );
or ( n57388 , n57386 , n57387 );
and ( n57389 , n57388 , n37841 );
and ( n57390 , n15112 , n36348 );
and ( n57391 , n13255 , n39453 );
or ( n57392 , n57390 , n57391 );
and ( n57393 , n57392 , n37847 );
and ( n57394 , n13255 , n37849 );
or ( n57395 , n57361 , n57371 , n57381 , n57385 , n57389 , n57393 , n57394 );
and ( n57396 , n57336 , n57395 );
and ( n57397 , n13255 , n34821 );
or ( n57398 , n57396 , n57397 );
and ( n57399 , n57398 , n16574 );
and ( n57400 , n13255 , n16576 );
or ( n57401 , n57399 , n57400 );
buf ( n57402 , n57401 );
buf ( n57403 , n57402 );
buf ( n57404 , n10615 );
buf ( n57405 , n10615 );
not ( n57406 , n24800 );
and ( n57407 , n25952 , n25222 );
and ( n57408 , n48334 , n28583 );
and ( n57409 , n25952 , n28591 );
or ( n57410 , n57408 , n57409 );
and ( n57411 , n57410 , n28594 );
and ( n57412 , n48344 , n28583 );
and ( n57413 , n25952 , n28591 );
or ( n57414 , n57412 , n57413 );
and ( n57415 , n57414 , n30269 );
and ( n57416 , n48354 , n28583 );
and ( n57417 , n25952 , n28591 );
or ( n57418 , n57416 , n57417 );
and ( n57419 , n57418 , n30982 );
and ( n57420 , n29615 , n28583 );
and ( n57421 , n25952 , n28591 );
or ( n57422 , n57420 , n57421 );
and ( n57423 , n57422 , n30989 );
and ( n57424 , n25950 , n30991 );
and ( n57425 , n48364 , n28583 );
and ( n57426 , n25952 , n28591 );
or ( n57427 , n57425 , n57426 );
and ( n57428 , n57427 , n31002 );
or ( n57429 , n57407 , n57411 , n57415 , n57419 , n57423 , n57424 , n57428 );
and ( n57430 , n57406 , n57429 );
and ( n57431 , n25952 , n24800 );
or ( n57432 , n57430 , n57431 );
and ( n57433 , n57432 , n31008 );
and ( n57434 , n25952 , n10618 );
or ( n57435 , n57433 , n57434 );
buf ( n57436 , n57435 );
buf ( n57437 , n57436 );
not ( n57438 , n24511 );
not ( n57439 , n24799 );
and ( n57440 , n10623 , n40154 );
not ( n57441 , n40632 );
and ( n57442 , n57441 , n40165 );
xor ( n57443 , n40650 , n40306 );
and ( n57444 , n57443 , n40632 );
or ( n57445 , n57442 , n57444 );
buf ( n57446 , n57445 );
and ( n57447 , n57446 , n27046 );
not ( n57448 , n41147 );
and ( n57449 , n57448 , n40680 );
xor ( n57450 , n41165 , n40821 );
and ( n57451 , n57450 , n41147 );
or ( n57452 , n57449 , n57451 );
buf ( n57453 , n57452 );
and ( n57454 , n57453 , n27049 );
and ( n57455 , n28890 , n28506 );
and ( n57456 , n10623 , n28508 );
or ( n57457 , n57447 , n57454 , n57455 , n57456 );
and ( n57458 , n57457 , n41199 );
or ( n57459 , n57440 , n57458 );
and ( n57460 , n57439 , n57459 );
xor ( n57461 , n41756 , n41763 );
buf ( n57462 , n57461 );
and ( n57463 , n57462 , n27046 );
xor ( n57464 , n42258 , n42259 );
buf ( n57465 , n57464 );
and ( n57466 , n57465 , n27049 );
and ( n57467 , n28890 , n42306 );
or ( n57468 , n57463 , n57466 , n57467 );
buf ( n57469 , n57468 );
buf ( n57470 , n57469 );
not ( n57471 , n57470 );
buf ( n57472 , n57471 );
buf ( n57473 , n57472 );
not ( n57474 , n57473 );
and ( n57475 , C1 , n57474 );
or ( n57476 , n57475 , C0 );
buf ( n57477 , n57476 );
and ( n57478 , n57477 , n24799 );
or ( n57479 , n57460 , n57478 );
and ( n57480 , n57438 , n57479 );
and ( n57481 , n57457 , n24511 );
or ( n57482 , n57480 , n57481 );
and ( n57483 , n57482 , n31008 );
not ( n57484 , n42601 );
and ( n57485 , n57484 , n42331 );
xor ( n57486 , n42619 , n42332 );
and ( n57487 , n57486 , n42601 );
or ( n57488 , n57485 , n57487 );
buf ( n57489 , n57488 );
and ( n57490 , n57489 , n10618 );
or ( n57491 , n57483 , n57490 );
buf ( n57492 , n57491 );
buf ( n57493 , n57492 );
buf ( n57494 , n10615 );
buf ( n57495 , n10615 );
buf ( n57496 , n10615 );
buf ( n57497 , n10613 );
not ( n57498 , n24800 );
and ( n57499 , n53614 , n28587 );
and ( n57500 , n26227 , n39807 );
or ( n57501 , n57499 , n57500 );
and ( n57502 , n57501 , n28594 );
and ( n57503 , n53624 , n28587 );
and ( n57504 , n26227 , n39807 );
or ( n57505 , n57503 , n57504 );
and ( n57506 , n57505 , n30269 );
and ( n57507 , n53634 , n28587 );
and ( n57508 , n26227 , n39807 );
or ( n57509 , n57507 , n57508 );
and ( n57510 , n57509 , n30982 );
and ( n57511 , n29455 , n28587 );
and ( n57512 , n26227 , n39807 );
or ( n57513 , n57511 , n57512 );
and ( n57514 , n57513 , n30989 );
and ( n57515 , n53645 , n28587 );
and ( n57516 , n26227 , n39807 );
or ( n57517 , n57515 , n57516 );
and ( n57518 , n57517 , n31002 );
and ( n57519 , n26227 , n34607 );
or ( n57520 , n57502 , n57506 , n57510 , n57514 , n57518 , n57519 );
and ( n57521 , n57498 , n57520 );
and ( n57522 , n26227 , n24800 );
or ( n57523 , n57521 , n57522 );
and ( n57524 , n57523 , n31008 );
and ( n57525 , n26227 , n10618 );
or ( n57526 , n57524 , n57525 );
buf ( n57527 , n57526 );
buf ( n57528 , n57527 );
not ( n57529 , n34821 );
not ( n57530 , n13916 );
and ( n57531 , n57530 , n13617 );
xor ( n57532 , n13618 , n13877 );
and ( n57533 , n57532 , n13916 );
or ( n57534 , n57531 , n57533 );
buf ( n57535 , n57534 );
and ( n57536 , n57535 , n14137 );
and ( n57537 , n57535 , n14143 );
not ( n57538 , n14139 );
and ( n57539 , n57538 , n36119 );
not ( n57540 , n36245 );
and ( n57541 , n57540 , n36131 );
xor ( n57542 , n46405 , n46406 );
and ( n57543 , n57542 , n36245 );
or ( n57544 , n57541 , n57543 );
buf ( n57545 , n57544 );
and ( n57546 , n57545 , n14139 );
or ( n57547 , n57539 , n57546 );
and ( n57548 , n57547 , n14140 );
and ( n57549 , n36119 , n14141 );
or ( n57550 , n57536 , n57537 , n57548 , n57549 );
and ( n57551 , n57550 , n36345 );
and ( n57552 , n13221 , n36352 );
or ( n57553 , n57551 , n57552 );
and ( n57554 , n57553 , n14562 );
not ( n57555 , n37048 );
and ( n57556 , n57555 , n36942 );
xor ( n57557 , n46428 , n46429 );
and ( n57558 , n57557 , n37048 );
or ( n57559 , n57556 , n57558 );
buf ( n57560 , n57559 );
and ( n57561 , n57560 , n36345 );
and ( n57562 , n13221 , n37073 );
or ( n57563 , n57561 , n57562 );
and ( n57564 , n57563 , n14586 );
not ( n57565 , n37801 );
and ( n57566 , n57565 , n37695 );
xor ( n57567 , n46446 , n46447 );
and ( n57568 , n57567 , n37801 );
or ( n57569 , n57566 , n57568 );
buf ( n57570 , n57569 );
and ( n57571 , n57570 , n36350 );
and ( n57572 , n13221 , n37825 );
or ( n57573 , n57571 , n57572 );
and ( n57574 , n57573 , n14584 );
and ( n57575 , n57560 , n36350 );
and ( n57576 , n13221 , n37831 );
or ( n57577 , n57575 , n57576 );
and ( n57578 , n57577 , n37835 );
and ( n57579 , n57570 , n36350 );
and ( n57580 , n13221 , n37831 );
or ( n57581 , n57579 , n57580 );
and ( n57582 , n57581 , n37841 );
and ( n57583 , n15067 , n36350 );
and ( n57584 , n13221 , n37831 );
or ( n57585 , n57583 , n57584 );
and ( n57586 , n57585 , n37847 );
and ( n57587 , n13221 , n37849 );
or ( n57588 , n57554 , n57564 , n57574 , n57578 , n57582 , n57586 , n57587 );
and ( n57589 , n57529 , n57588 );
and ( n57590 , n13221 , n34821 );
or ( n57591 , n57589 , n57590 );
and ( n57592 , n57591 , n16574 );
and ( n57593 , n13221 , n16576 );
or ( n57594 , n57592 , n57593 );
buf ( n57595 , n57594 );
buf ( n57596 , n57595 );
buf ( n57597 , n10613 );
buf ( n57598 , n10613 );
buf ( n57599 , n10615 );
buf ( n57600 , n10613 );
buf ( n57601 , n10615 );
not ( n57602 , n34821 );
and ( n57603 , n13409 , n14592 );
and ( n57604 , n36271 , n36348 );
and ( n57605 , n13409 , n43530 );
or ( n57606 , n57604 , n57605 );
and ( n57607 , n57606 , n14562 );
and ( n57608 , n37069 , n36347 );
and ( n57609 , n13409 , n43543 );
or ( n57610 , n57608 , n57609 );
and ( n57611 , n57610 , n14586 );
and ( n57612 , n37822 , n36348 );
and ( n57613 , n13409 , n43556 );
or ( n57614 , n57612 , n57613 );
and ( n57615 , n57614 , n14584 );
and ( n57616 , n37069 , n36347 );
and ( n57617 , n13409 , n43563 );
or ( n57618 , n57616 , n57617 );
and ( n57619 , n57618 , n37835 );
and ( n57620 , n37822 , n36347 );
and ( n57621 , n13409 , n43563 );
or ( n57622 , n57620 , n57621 );
and ( n57623 , n57622 , n37841 );
and ( n57624 , n13407 , n14564 );
and ( n57625 , n15713 , n36347 );
and ( n57626 , n13409 , n43563 );
or ( n57627 , n57625 , n57626 );
and ( n57628 , n57627 , n37847 );
or ( n57629 , n57603 , n57607 , n57611 , n57615 , n57619 , n57623 , n57624 , n57628 );
and ( n57630 , n57602 , n57629 );
and ( n57631 , n13409 , n34821 );
or ( n57632 , n57630 , n57631 );
and ( n57633 , n57632 , n16574 );
and ( n57634 , n13409 , n16576 );
or ( n57635 , n57633 , n57634 );
buf ( n57636 , n57635 );
buf ( n57637 , n57636 );
not ( n57638 , n34821 );
and ( n57639 , n13457 , n14592 );
and ( n57640 , n46341 , n36348 );
and ( n57641 , n13457 , n43530 );
or ( n57642 , n57640 , n57641 );
and ( n57643 , n57642 , n14562 );
and ( n57644 , n46351 , n36347 );
and ( n57645 , n13457 , n43543 );
or ( n57646 , n57644 , n57645 );
and ( n57647 , n57646 , n14586 );
and ( n57648 , n46361 , n36348 );
and ( n57649 , n13457 , n43556 );
or ( n57650 , n57648 , n57649 );
and ( n57651 , n57650 , n14584 );
and ( n57652 , n46351 , n36347 );
and ( n57653 , n13457 , n43563 );
or ( n57654 , n57652 , n57653 );
and ( n57655 , n57654 , n37835 );
and ( n57656 , n46361 , n36347 );
and ( n57657 , n13457 , n43563 );
or ( n57658 , n57656 , n57657 );
and ( n57659 , n57658 , n37841 );
and ( n57660 , n13455 , n14564 );
and ( n57661 , n15801 , n36347 );
and ( n57662 , n13457 , n43563 );
or ( n57663 , n57661 , n57662 );
and ( n57664 , n57663 , n37847 );
or ( n57665 , n57639 , n57643 , n57647 , n57651 , n57655 , n57659 , n57660 , n57664 );
and ( n57666 , n57638 , n57665 );
and ( n57667 , n13457 , n34821 );
or ( n57668 , n57666 , n57667 );
and ( n57669 , n57668 , n16574 );
and ( n57670 , n13457 , n16576 );
or ( n57671 , n57669 , n57670 );
buf ( n57672 , n57671 );
buf ( n57673 , n57672 );
buf ( n57674 , n10613 );
buf ( n57675 , n10613 );
buf ( n57676 , n10613 );
buf ( n57677 , n10613 );
not ( n57678 , n24800 );
and ( n57679 , n57678 , n28550 );
and ( n57680 , n28525 , n24800 );
or ( n57681 , n57679 , n57680 );
and ( n57682 , n57681 , n31008 );
and ( n57683 , n28525 , n10618 );
or ( n57684 , n57682 , n57683 );
buf ( n57685 , n57684 );
buf ( n57686 , n57685 );
not ( n57687 , n34804 );
and ( n57688 , n57687 , n26773 );
and ( n57689 , n14671 , n34804 );
or ( n57690 , n57688 , n57689 );
and ( n57691 , n57690 , n31008 );
and ( n57692 , n14671 , n10618 );
or ( n57693 , n57691 , n57692 );
buf ( n57694 , n57693 );
buf ( n57695 , n57694 );
buf ( n57696 , n10613 );
buf ( n57697 , n10615 );
buf ( n57698 , n10613 );
buf ( n57699 , n10615 );
and ( n57700 , n16817 , n23924 );
and ( n57701 , n22193 , n23926 );
or ( n57702 , n57700 , n57701 );
buf ( n57703 , n57702 );
buf ( n57704 , n57703 );
buf ( n57705 , n10615 );
not ( n57706 , n17162 );
not ( n57707 , n17450 );
buf ( n57708 , n40068 );
and ( n57709 , n57708 , n19745 );
or ( n57710 , n21253 , n21255 );
or ( n57711 , n57710 , n19748 );
and ( n57712 , n19750 , n57711 );
or ( n57713 , n57709 , n57712 );
and ( n57714 , n57713 , n21341 );
or ( n57715 , n23834 , n23917 );
or ( n57716 , n57715 , n23830 );
or ( n57717 , n57716 , n23831 );
or ( n57718 , n57717 , n23819 );
or ( n57719 , n57718 , n23820 );
or ( n57720 , n57719 , n23058 );
or ( n57721 , n57720 , n23059 );
or ( n57722 , n57721 , n23822 );
or ( n57723 , n57722 , n23061 );
or ( n57724 , n57723 , n23824 );
or ( n57725 , n57724 , n23063 );
or ( n57726 , n57725 , n17873 );
and ( n57727 , n19750 , n57726 );
or ( n57728 , n57714 , n57727 );
and ( n57729 , n57707 , n57728 );
and ( n57730 , n19750 , n17450 );
or ( n57731 , n57729 , n57730 );
and ( n57732 , n57706 , n57731 );
buf ( n57733 , n18527 );
not ( n57734 , n57733 );
buf ( n57735 , n20484 );
and ( n57736 , n57734 , n57735 );
buf ( n57737 , n57736 );
not ( n57738 , n57737 );
and ( n57739 , n57738 , n18527 );
or ( n57740 , n57739 , C0 );
buf ( n57741 , n57740 );
buf ( n57742 , n21841 );
xor ( n57743 , n57741 , n57742 );
not ( n57744 , n57743 );
not ( n57745 , n57737 );
and ( n57746 , n57745 , n20484 );
or ( n57747 , n57746 , C0 );
buf ( n57748 , n57747 );
not ( n57749 , n57748 );
buf ( n57750 , n21854 );
and ( n57751 , n57749 , n57750 );
buf ( n57752 , n20496 );
buf ( n57753 , n57752 );
not ( n57754 , n57753 );
buf ( n57755 , n21867 );
and ( n57756 , n57754 , n57755 );
buf ( n57757 , n19458 );
buf ( n57758 , n57757 );
not ( n57759 , n57758 );
buf ( n57760 , n21880 );
and ( n57761 , n57759 , n57760 );
buf ( n57762 , n19424 );
buf ( n57763 , n57762 );
not ( n57764 , n57763 );
buf ( n57765 , n21893 );
and ( n57766 , n57764 , n57765 );
buf ( n57767 , n19390 );
buf ( n57768 , n57767 );
not ( n57769 , n57768 );
buf ( n57770 , n21906 );
and ( n57771 , n57769 , n57770 );
buf ( n57772 , n19356 );
buf ( n57773 , n57772 );
not ( n57774 , n57773 );
buf ( n57775 , n21919 );
and ( n57776 , n57774 , n57775 );
buf ( n57777 , n19323 );
buf ( n57778 , n57777 );
not ( n57779 , n57778 );
buf ( n57780 , n21932 );
and ( n57781 , n57779 , n57780 );
buf ( n57782 , n19289 );
buf ( n57783 , n57782 );
not ( n57784 , n57783 );
buf ( n57785 , n21945 );
and ( n57786 , n57784 , n57785 );
buf ( n57787 , n19255 );
buf ( n57788 , n57787 );
not ( n57789 , n57788 );
buf ( n57790 , n21958 );
and ( n57791 , n57789 , n57790 );
buf ( n57792 , n19221 );
buf ( n57793 , n57792 );
not ( n57794 , n57793 );
buf ( n57795 , n21971 );
and ( n57796 , n57794 , n57795 );
buf ( n57797 , n19187 );
buf ( n57798 , n57797 );
not ( n57799 , n57798 );
buf ( n57800 , n21984 );
and ( n57801 , n57799 , n57800 );
buf ( n57802 , n19153 );
buf ( n57803 , n57802 );
not ( n57804 , n57803 );
buf ( n57805 , n22042 );
and ( n57806 , n57804 , n57805 );
buf ( n57807 , n19119 );
buf ( n57808 , n57807 );
not ( n57809 , n57808 );
buf ( n57810 , n22062 );
and ( n57811 , n57809 , n57810 );
buf ( n57812 , n19085 );
buf ( n57813 , n57812 );
not ( n57814 , n57813 );
buf ( n57815 , n22082 );
and ( n57816 , n57814 , n57815 );
buf ( n57817 , n19051 );
buf ( n57818 , n57817 );
not ( n57819 , n57818 );
buf ( n57820 , n22102 );
and ( n57821 , n57819 , n57820 );
buf ( n57822 , n19017 );
buf ( n57823 , n57822 );
not ( n57824 , n57823 );
buf ( n57825 , n22122 );
and ( n57826 , n57824 , n57825 );
buf ( n57827 , n18983 );
buf ( n57828 , n57827 );
not ( n57829 , n57828 );
buf ( n57830 , n22142 );
and ( n57831 , n57829 , n57830 );
buf ( n57832 , n18949 );
buf ( n57833 , n57832 );
not ( n57834 , n57833 );
buf ( n57835 , n22162 );
and ( n57836 , n57834 , n57835 );
buf ( n57837 , n18915 );
buf ( n57838 , n57837 );
not ( n57839 , n57838 );
buf ( n57840 , n22182 );
and ( n57841 , n57839 , n57840 );
buf ( n57842 , n18881 );
buf ( n57843 , n57842 );
not ( n57844 , n57843 );
buf ( n57845 , n22202 );
and ( n57846 , n57844 , n57845 );
buf ( n57847 , n18847 );
buf ( n57848 , n57847 );
not ( n57849 , n57848 );
buf ( n57850 , n22222 );
and ( n57851 , n57849 , n57850 );
buf ( n57852 , n18813 );
buf ( n57853 , n57852 );
not ( n57854 , n57853 );
buf ( n57855 , n22242 );
and ( n57856 , n57854 , n57855 );
buf ( n57857 , n18779 );
buf ( n57858 , n57857 );
not ( n57859 , n57858 );
buf ( n57860 , n22262 );
and ( n57861 , n57859 , n57860 );
buf ( n57862 , n18745 );
buf ( n57863 , n57862 );
not ( n57864 , n57863 );
buf ( n57865 , n22282 );
and ( n57866 , n57864 , n57865 );
buf ( n57867 , n18711 );
buf ( n57868 , n57867 );
not ( n57869 , n57868 );
buf ( n57870 , n22302 );
and ( n57871 , n57869 , n57870 );
buf ( n57872 , n18677 );
buf ( n57873 , n57872 );
not ( n57874 , n57873 );
buf ( n57875 , n22322 );
and ( n57876 , n57874 , n57875 );
buf ( n57877 , n18643 );
buf ( n57878 , n57877 );
not ( n57879 , n57878 );
buf ( n57880 , n22342 );
and ( n57881 , n57879 , n57880 );
buf ( n57882 , n18610 );
buf ( n57883 , n57882 );
not ( n57884 , n57883 );
buf ( n57885 , n22362 );
and ( n57886 , n57884 , n57885 );
buf ( n57887 , n18577 );
buf ( n57888 , n57887 );
not ( n57889 , n57888 );
buf ( n57890 , n22382 );
and ( n57891 , n57889 , n57890 );
buf ( n57892 , n18546 );
buf ( n57893 , n57892 );
not ( n57894 , n57893 );
buf ( n57895 , n22402 );
and ( n57896 , n57894 , n57895 );
buf ( n57897 , n18514 );
buf ( n57898 , n57897 );
not ( n57899 , n57898 );
buf ( n57900 , n21639 );
and ( n57901 , n57899 , n57900 );
xnor ( n57902 , n57893 , n57895 );
and ( n57903 , n57901 , n57902 );
or ( n57904 , n57896 , n57903 );
xnor ( n57905 , n57888 , n57890 );
and ( n57906 , n57904 , n57905 );
or ( n57907 , n57891 , n57906 );
xnor ( n57908 , n57883 , n57885 );
and ( n57909 , n57907 , n57908 );
or ( n57910 , n57886 , n57909 );
xnor ( n57911 , n57878 , n57880 );
and ( n57912 , n57910 , n57911 );
or ( n57913 , n57881 , n57912 );
nor ( n57914 , n57873 , n57875 );
and ( n57915 , n57913 , n57914 );
or ( n57916 , n57876 , n57915 );
xnor ( n57917 , n57868 , n57870 );
and ( n57918 , n57916 , n57917 );
or ( n57919 , n57871 , n57918 );
xnor ( n57920 , n57863 , n57865 );
and ( n57921 , n57919 , n57920 );
or ( n57922 , n57866 , n57921 );
xnor ( n57923 , n57858 , n57860 );
and ( n57924 , n57922 , n57923 );
or ( n57925 , n57861 , n57924 );
xnor ( n57926 , n57853 , n57855 );
and ( n57927 , n57925 , n57926 );
or ( n57928 , n57856 , n57927 );
xnor ( n57929 , n57848 , n57850 );
and ( n57930 , n57928 , n57929 );
or ( n57931 , n57851 , n57930 );
xnor ( n57932 , n57843 , n57845 );
and ( n57933 , n57931 , n57932 );
or ( n57934 , n57846 , n57933 );
xnor ( n57935 , n57838 , n57840 );
and ( n57936 , n57934 , n57935 );
or ( n57937 , n57841 , n57936 );
xnor ( n57938 , n57833 , n57835 );
and ( n57939 , n57937 , n57938 );
or ( n57940 , n57836 , n57939 );
xnor ( n57941 , n57828 , n57830 );
and ( n57942 , n57940 , n57941 );
or ( n57943 , n57831 , n57942 );
xnor ( n57944 , n57823 , n57825 );
and ( n57945 , n57943 , n57944 );
or ( n57946 , n57826 , n57945 );
xnor ( n57947 , n57818 , n57820 );
and ( n57948 , n57946 , n57947 );
or ( n57949 , n57821 , n57948 );
xnor ( n57950 , n57813 , n57815 );
and ( n57951 , n57949 , n57950 );
or ( n57952 , n57816 , n57951 );
xnor ( n57953 , n57808 , n57810 );
and ( n57954 , n57952 , n57953 );
or ( n57955 , n57811 , n57954 );
xnor ( n57956 , n57803 , n57805 );
and ( n57957 , n57955 , n57956 );
or ( n57958 , n57806 , n57957 );
xnor ( n57959 , n57798 , n57800 );
and ( n57960 , n57958 , n57959 );
or ( n57961 , n57801 , n57960 );
xnor ( n57962 , n57793 , n57795 );
and ( n57963 , n57961 , n57962 );
or ( n57964 , n57796 , n57963 );
xnor ( n57965 , n57788 , n57790 );
and ( n57966 , n57964 , n57965 );
or ( n57967 , n57791 , n57966 );
xnor ( n57968 , n57783 , n57785 );
and ( n57969 , n57967 , n57968 );
or ( n57970 , n57786 , n57969 );
xnor ( n57971 , n57778 , n57780 );
and ( n57972 , n57970 , n57971 );
or ( n57973 , n57781 , n57972 );
xnor ( n57974 , n57773 , n57775 );
and ( n57975 , n57973 , n57974 );
or ( n57976 , n57776 , n57975 );
xnor ( n57977 , n57768 , n57770 );
and ( n57978 , n57976 , n57977 );
or ( n57979 , n57771 , n57978 );
xnor ( n57980 , n57763 , n57765 );
and ( n57981 , n57979 , n57980 );
or ( n57982 , n57766 , n57981 );
xnor ( n57983 , n57758 , n57760 );
and ( n57984 , n57982 , n57983 );
or ( n57985 , n57761 , n57984 );
xnor ( n57986 , n57753 , n57755 );
and ( n57987 , n57985 , n57986 );
or ( n57988 , n57756 , n57987 );
xnor ( n57989 , n57748 , n57750 );
and ( n57990 , n57988 , n57989 );
or ( n57991 , n57751 , n57990 );
and ( n57992 , n57744 , n57991 );
not ( n57993 , n57742 );
and ( n57994 , n57993 , n57741 );
and ( n57995 , n57994 , n57743 );
or ( n57996 , n57992 , n57995 );
buf ( n57997 , n57996 );
not ( n57998 , n57997 );
or ( n57999 , n57998 , n19750 );
and ( n58000 , n57999 , n17872 );
or ( n58001 , n57997 , n19750 );
and ( n58002 , n58001 , n17870 );
buf ( n58003 , n18527 );
buf ( n58004 , n21841 );
xor ( n58005 , n58003 , n58004 );
not ( n58006 , n58005 );
buf ( n58007 , n21854 );
not ( n58008 , n58007 );
buf ( n58009 , n20484 );
and ( n58010 , n58008 , n58009 );
buf ( n58011 , n21867 );
not ( n58012 , n58011 );
buf ( n58013 , n20496 );
and ( n58014 , n58012 , n58013 );
buf ( n58015 , n21880 );
not ( n58016 , n58015 );
buf ( n58017 , n19458 );
and ( n58018 , n58016 , n58017 );
buf ( n58019 , n21893 );
not ( n58020 , n58019 );
buf ( n58021 , n19424 );
and ( n58022 , n58020 , n58021 );
buf ( n58023 , n21906 );
not ( n58024 , n58023 );
buf ( n58025 , n19390 );
and ( n58026 , n58024 , n58025 );
buf ( n58027 , n21919 );
not ( n58028 , n58027 );
buf ( n58029 , n19356 );
and ( n58030 , n58028 , n58029 );
buf ( n58031 , n21932 );
not ( n58032 , n58031 );
buf ( n58033 , n19323 );
and ( n58034 , n58032 , n58033 );
buf ( n58035 , n21945 );
not ( n58036 , n58035 );
buf ( n58037 , n19289 );
and ( n58038 , n58036 , n58037 );
buf ( n58039 , n21958 );
not ( n58040 , n58039 );
buf ( n58041 , n19255 );
and ( n58042 , n58040 , n58041 );
buf ( n58043 , n21971 );
not ( n58044 , n58043 );
buf ( n58045 , n19221 );
and ( n58046 , n58044 , n58045 );
buf ( n58047 , n21984 );
not ( n58048 , n58047 );
buf ( n58049 , n19187 );
and ( n58050 , n58048 , n58049 );
buf ( n58051 , n22042 );
not ( n58052 , n58051 );
buf ( n58053 , n19153 );
and ( n58054 , n58052 , n58053 );
buf ( n58055 , n22062 );
not ( n58056 , n58055 );
buf ( n58057 , n19119 );
and ( n58058 , n58056 , n58057 );
buf ( n58059 , n22082 );
not ( n58060 , n58059 );
buf ( n58061 , n19085 );
and ( n58062 , n58060 , n58061 );
buf ( n58063 , n22102 );
not ( n58064 , n58063 );
buf ( n58065 , n19051 );
and ( n58066 , n58064 , n58065 );
buf ( n58067 , n22122 );
not ( n58068 , n58067 );
buf ( n58069 , n19017 );
and ( n58070 , n58068 , n58069 );
buf ( n58071 , n22142 );
not ( n58072 , n58071 );
buf ( n58073 , n18983 );
and ( n58074 , n58072 , n58073 );
buf ( n58075 , n22162 );
not ( n58076 , n58075 );
buf ( n58077 , n18949 );
and ( n58078 , n58076 , n58077 );
buf ( n58079 , n22182 );
not ( n58080 , n58079 );
buf ( n58081 , n18915 );
and ( n58082 , n58080 , n58081 );
buf ( n58083 , n22202 );
not ( n58084 , n58083 );
buf ( n58085 , n18881 );
and ( n58086 , n58084 , n58085 );
buf ( n58087 , n22222 );
not ( n58088 , n58087 );
buf ( n58089 , n18847 );
and ( n58090 , n58088 , n58089 );
buf ( n58091 , n22242 );
not ( n58092 , n58091 );
buf ( n58093 , n18813 );
and ( n58094 , n58092 , n58093 );
buf ( n58095 , n22262 );
not ( n58096 , n58095 );
buf ( n58097 , n18779 );
and ( n58098 , n58096 , n58097 );
buf ( n58099 , n22282 );
not ( n58100 , n58099 );
buf ( n58101 , n18745 );
and ( n58102 , n58100 , n58101 );
buf ( n58103 , n22302 );
not ( n58104 , n58103 );
buf ( n58105 , n18711 );
and ( n58106 , n58104 , n58105 );
buf ( n58107 , n22322 );
not ( n58108 , n58107 );
buf ( n58109 , n18677 );
and ( n58110 , n58108 , n58109 );
buf ( n58111 , n22342 );
not ( n58112 , n58111 );
buf ( n58113 , n18643 );
and ( n58114 , n58112 , n58113 );
buf ( n58115 , n22362 );
not ( n58116 , n58115 );
buf ( n58117 , n18610 );
and ( n58118 , n58116 , n58117 );
buf ( n58119 , n22382 );
not ( n58120 , n58119 );
buf ( n58121 , n18577 );
and ( n58122 , n58120 , n58121 );
buf ( n58123 , n22402 );
not ( n58124 , n58123 );
buf ( n58125 , n18546 );
and ( n58126 , n58124 , n58125 );
buf ( n58127 , n21639 );
not ( n58128 , n58127 );
buf ( n58129 , n18514 );
and ( n58130 , n58128 , n58129 );
xnor ( n58131 , n58125 , n58123 );
and ( n58132 , n58130 , n58131 );
or ( n58133 , n58126 , n58132 );
xnor ( n58134 , n58121 , n58119 );
and ( n58135 , n58133 , n58134 );
or ( n58136 , n58122 , n58135 );
xnor ( n58137 , n58117 , n58115 );
and ( n58138 , n58136 , n58137 );
or ( n58139 , n58118 , n58138 );
xnor ( n58140 , n58113 , n58111 );
and ( n58141 , n58139 , n58140 );
or ( n58142 , n58114 , n58141 );
xnor ( n58143 , n58109 , n58107 );
and ( n58144 , n58142 , n58143 );
or ( n58145 , n58110 , n58144 );
xnor ( n58146 , n58105 , n58103 );
and ( n58147 , n58145 , n58146 );
or ( n58148 , n58106 , n58147 );
xnor ( n58149 , n58101 , n58099 );
and ( n58150 , n58148 , n58149 );
or ( n58151 , n58102 , n58150 );
xnor ( n58152 , n58097 , n58095 );
and ( n58153 , n58151 , n58152 );
or ( n58154 , n58098 , n58153 );
xnor ( n58155 , n58093 , n58091 );
and ( n58156 , n58154 , n58155 );
or ( n58157 , n58094 , n58156 );
xnor ( n58158 , n58089 , n58087 );
and ( n58159 , n58157 , n58158 );
or ( n58160 , n58090 , n58159 );
xnor ( n58161 , n58085 , n58083 );
and ( n58162 , n58160 , n58161 );
or ( n58163 , n58086 , n58162 );
xnor ( n58164 , n58081 , n58079 );
and ( n58165 , n58163 , n58164 );
or ( n58166 , n58082 , n58165 );
xnor ( n58167 , n58077 , n58075 );
and ( n58168 , n58166 , n58167 );
or ( n58169 , n58078 , n58168 );
xnor ( n58170 , n58073 , n58071 );
and ( n58171 , n58169 , n58170 );
or ( n58172 , n58074 , n58171 );
xnor ( n58173 , n58069 , n58067 );
and ( n58174 , n58172 , n58173 );
or ( n58175 , n58070 , n58174 );
xnor ( n58176 , n58065 , n58063 );
and ( n58177 , n58175 , n58176 );
or ( n58178 , n58066 , n58177 );
xnor ( n58179 , n58061 , n58059 );
and ( n58180 , n58178 , n58179 );
or ( n58181 , n58062 , n58180 );
xnor ( n58182 , n58057 , n58055 );
and ( n58183 , n58181 , n58182 );
or ( n58184 , n58058 , n58183 );
xnor ( n58185 , n58053 , n58051 );
and ( n58186 , n58184 , n58185 );
or ( n58187 , n58054 , n58186 );
xnor ( n58188 , n58049 , n58047 );
and ( n58189 , n58187 , n58188 );
or ( n58190 , n58050 , n58189 );
xnor ( n58191 , n58045 , n58043 );
and ( n58192 , n58190 , n58191 );
or ( n58193 , n58046 , n58192 );
xnor ( n58194 , n58041 , n58039 );
and ( n58195 , n58193 , n58194 );
or ( n58196 , n58042 , n58195 );
xnor ( n58197 , n58037 , n58035 );
and ( n58198 , n58196 , n58197 );
or ( n58199 , n58038 , n58198 );
xnor ( n58200 , n58033 , n58031 );
and ( n58201 , n58199 , n58200 );
or ( n58202 , n58034 , n58201 );
xnor ( n58203 , n58029 , n58027 );
and ( n58204 , n58202 , n58203 );
or ( n58205 , n58030 , n58204 );
xnor ( n58206 , n58025 , n58023 );
and ( n58207 , n58205 , n58206 );
or ( n58208 , n58026 , n58207 );
xnor ( n58209 , n58021 , n58019 );
and ( n58210 , n58208 , n58209 );
or ( n58211 , n58022 , n58210 );
xnor ( n58212 , n58017 , n58015 );
and ( n58213 , n58211 , n58212 );
or ( n58214 , n58018 , n58213 );
xnor ( n58215 , n58013 , n58011 );
and ( n58216 , n58214 , n58215 );
or ( n58217 , n58014 , n58216 );
xnor ( n58218 , n58009 , n58007 );
and ( n58219 , n58217 , n58218 );
or ( n58220 , n58010 , n58219 );
and ( n58221 , n58006 , n58220 );
not ( n58222 , n58003 );
and ( n58223 , n58222 , n58004 );
and ( n58224 , n58223 , n58005 );
or ( n58225 , n58221 , n58224 );
buf ( n58226 , n58225 );
or ( n58227 , n58226 , n19750 );
and ( n58228 , n58227 , n17868 );
not ( n58229 , n58226 );
or ( n58230 , n58229 , n19750 );
and ( n58231 , n58230 , n21341 );
buf ( n58232 , n18527 );
buf ( n58233 , n21841 );
xor ( n58234 , n58232 , n58233 );
buf ( n58235 , n20484 );
buf ( n58236 , n21854 );
xor ( n58237 , n58235 , n58236 );
or ( n58238 , n58234 , n58237 );
buf ( n58239 , n20496 );
buf ( n58240 , n21867 );
xor ( n58241 , n58239 , n58240 );
or ( n58242 , n58238 , n58241 );
buf ( n58243 , n19458 );
buf ( n58244 , n21880 );
xor ( n58245 , n58243 , n58244 );
or ( n58246 , n58242 , n58245 );
buf ( n58247 , n19424 );
buf ( n58248 , n21893 );
xor ( n58249 , n58247 , n58248 );
or ( n58250 , n58246 , n58249 );
buf ( n58251 , n19390 );
buf ( n58252 , n21906 );
xor ( n58253 , n58251 , n58252 );
or ( n58254 , n58250 , n58253 );
buf ( n58255 , n19356 );
buf ( n58256 , n21919 );
xor ( n58257 , n58255 , n58256 );
or ( n58258 , n58254 , n58257 );
buf ( n58259 , n19323 );
buf ( n58260 , n21932 );
xor ( n58261 , n58259 , n58260 );
or ( n58262 , n58258 , n58261 );
buf ( n58263 , n19289 );
buf ( n58264 , n21945 );
xor ( n58265 , n58263 , n58264 );
or ( n58266 , n58262 , n58265 );
buf ( n58267 , n19255 );
buf ( n58268 , n21958 );
xor ( n58269 , n58267 , n58268 );
or ( n58270 , n58266 , n58269 );
buf ( n58271 , n19221 );
buf ( n58272 , n21971 );
xor ( n58273 , n58271 , n58272 );
or ( n58274 , n58270 , n58273 );
buf ( n58275 , n19187 );
buf ( n58276 , n21984 );
xor ( n58277 , n58275 , n58276 );
or ( n58278 , n58274 , n58277 );
buf ( n58279 , n19153 );
buf ( n58280 , n22042 );
xor ( n58281 , n58279 , n58280 );
or ( n58282 , n58278 , n58281 );
buf ( n58283 , n19119 );
buf ( n58284 , n22062 );
xor ( n58285 , n58283 , n58284 );
or ( n58286 , n58282 , n58285 );
buf ( n58287 , n19085 );
buf ( n58288 , n22082 );
xor ( n58289 , n58287 , n58288 );
or ( n58290 , n58286 , n58289 );
buf ( n58291 , n19051 );
buf ( n58292 , n22102 );
xor ( n58293 , n58291 , n58292 );
or ( n58294 , n58290 , n58293 );
buf ( n58295 , n19017 );
buf ( n58296 , n22122 );
xor ( n58297 , n58295 , n58296 );
or ( n58298 , n58294 , n58297 );
buf ( n58299 , n18983 );
buf ( n58300 , n22142 );
xor ( n58301 , n58299 , n58300 );
or ( n58302 , n58298 , n58301 );
buf ( n58303 , n18949 );
buf ( n58304 , n22162 );
xor ( n58305 , n58303 , n58304 );
or ( n58306 , n58302 , n58305 );
buf ( n58307 , n18915 );
buf ( n58308 , n22182 );
xor ( n58309 , n58307 , n58308 );
or ( n58310 , n58306 , n58309 );
buf ( n58311 , n18881 );
buf ( n58312 , n22202 );
xor ( n58313 , n58311 , n58312 );
or ( n58314 , n58310 , n58313 );
buf ( n58315 , n18847 );
buf ( n58316 , n22222 );
xor ( n58317 , n58315 , n58316 );
or ( n58318 , n58314 , n58317 );
buf ( n58319 , n18813 );
buf ( n58320 , n22242 );
xor ( n58321 , n58319 , n58320 );
or ( n58322 , n58318 , n58321 );
buf ( n58323 , n18779 );
buf ( n58324 , n22262 );
xor ( n58325 , n58323 , n58324 );
or ( n58326 , n58322 , n58325 );
buf ( n58327 , n18745 );
buf ( n58328 , n22282 );
xor ( n58329 , n58327 , n58328 );
or ( n58330 , n58326 , n58329 );
buf ( n58331 , n18711 );
buf ( n58332 , n22302 );
xor ( n58333 , n58331 , n58332 );
or ( n58334 , n58330 , n58333 );
buf ( n58335 , n18677 );
buf ( n58336 , n22322 );
xor ( n58337 , n58335 , n58336 );
or ( n58338 , n58334 , n58337 );
buf ( n58339 , n18643 );
buf ( n58340 , n22342 );
xor ( n58341 , n58339 , n58340 );
or ( n58342 , n58338 , n58341 );
buf ( n58343 , n18610 );
buf ( n58344 , n22362 );
xor ( n58345 , n58343 , n58344 );
or ( n58346 , n58342 , n58345 );
buf ( n58347 , n18577 );
buf ( n58348 , n22382 );
xor ( n58349 , n58347 , n58348 );
or ( n58350 , n58346 , n58349 );
buf ( n58351 , n18546 );
buf ( n58352 , n22402 );
xor ( n58353 , n58351 , n58352 );
or ( n58354 , n58350 , n58353 );
buf ( n58355 , n18514 );
buf ( n58356 , n21639 );
xor ( n58357 , n58355 , n58356 );
or ( n58358 , n58354 , n58357 );
not ( n58359 , n58358 );
buf ( n58360 , n58359 );
not ( n58361 , n58360 );
or ( n58362 , n58361 , n19750 );
and ( n58363 , n58362 , n23063 );
or ( n58364 , n58360 , n19750 );
and ( n58365 , n58364 , n23824 );
buf ( n58366 , n18527 );
buf ( n58367 , n21841 );
xor ( n58368 , n58366 , n58367 );
not ( n58369 , n58368 );
buf ( n58370 , n20484 );
not ( n58371 , n58370 );
buf ( n58372 , n21854 );
and ( n58373 , n58371 , n58372 );
buf ( n58374 , n20496 );
not ( n58375 , n58374 );
buf ( n58376 , n21867 );
and ( n58377 , n58375 , n58376 );
buf ( n58378 , n19458 );
not ( n58379 , n58378 );
buf ( n58380 , n21880 );
and ( n58381 , n58379 , n58380 );
buf ( n58382 , n19424 );
not ( n58383 , n58382 );
buf ( n58384 , n21893 );
and ( n58385 , n58383 , n58384 );
buf ( n58386 , n19390 );
not ( n58387 , n58386 );
buf ( n58388 , n21906 );
and ( n58389 , n58387 , n58388 );
buf ( n58390 , n19356 );
not ( n58391 , n58390 );
buf ( n58392 , n21919 );
and ( n58393 , n58391 , n58392 );
buf ( n58394 , n19323 );
not ( n58395 , n58394 );
buf ( n58396 , n21932 );
and ( n58397 , n58395 , n58396 );
buf ( n58398 , n19289 );
not ( n58399 , n58398 );
buf ( n58400 , n21945 );
and ( n58401 , n58399 , n58400 );
buf ( n58402 , n19255 );
not ( n58403 , n58402 );
buf ( n58404 , n21958 );
and ( n58405 , n58403 , n58404 );
buf ( n58406 , n19221 );
not ( n58407 , n58406 );
buf ( n58408 , n21971 );
and ( n58409 , n58407 , n58408 );
buf ( n58410 , n19187 );
not ( n58411 , n58410 );
buf ( n58412 , n21984 );
and ( n58413 , n58411 , n58412 );
buf ( n58414 , n19153 );
not ( n58415 , n58414 );
buf ( n58416 , n22042 );
and ( n58417 , n58415 , n58416 );
buf ( n58418 , n19119 );
not ( n58419 , n58418 );
buf ( n58420 , n22062 );
and ( n58421 , n58419 , n58420 );
buf ( n58422 , n19085 );
not ( n58423 , n58422 );
buf ( n58424 , n22082 );
and ( n58425 , n58423 , n58424 );
buf ( n58426 , n19051 );
not ( n58427 , n58426 );
buf ( n58428 , n22102 );
and ( n58429 , n58427 , n58428 );
buf ( n58430 , n19017 );
not ( n58431 , n58430 );
buf ( n58432 , n22122 );
and ( n58433 , n58431 , n58432 );
buf ( n58434 , n18983 );
not ( n58435 , n58434 );
buf ( n58436 , n22142 );
and ( n58437 , n58435 , n58436 );
buf ( n58438 , n18949 );
not ( n58439 , n58438 );
buf ( n58440 , n22162 );
and ( n58441 , n58439 , n58440 );
buf ( n58442 , n18915 );
not ( n58443 , n58442 );
buf ( n58444 , n22182 );
and ( n58445 , n58443 , n58444 );
buf ( n58446 , n18881 );
not ( n58447 , n58446 );
buf ( n58448 , n22202 );
and ( n58449 , n58447 , n58448 );
buf ( n58450 , n18847 );
not ( n58451 , n58450 );
buf ( n58452 , n22222 );
and ( n58453 , n58451 , n58452 );
buf ( n58454 , n18813 );
not ( n58455 , n58454 );
buf ( n58456 , n22242 );
and ( n58457 , n58455 , n58456 );
buf ( n58458 , n18779 );
not ( n58459 , n58458 );
buf ( n58460 , n22262 );
and ( n58461 , n58459 , n58460 );
buf ( n58462 , n18745 );
not ( n58463 , n58462 );
buf ( n58464 , n22282 );
and ( n58465 , n58463 , n58464 );
buf ( n58466 , n18711 );
not ( n58467 , n58466 );
buf ( n58468 , n22302 );
and ( n58469 , n58467 , n58468 );
buf ( n58470 , n18677 );
not ( n58471 , n58470 );
buf ( n58472 , n22322 );
and ( n58473 , n58471 , n58472 );
buf ( n58474 , n18643 );
not ( n58475 , n58474 );
buf ( n58476 , n22342 );
nand ( n58477 , n58475 , n58476 );
buf ( n58478 , n18610 );
not ( n58479 , n58478 );
buf ( n58480 , n22362 );
and ( n58481 , n58479 , n58480 );
buf ( n58482 , n18577 );
not ( n58483 , n58482 );
buf ( n58484 , n22382 );
and ( n58485 , n58483 , n58484 );
buf ( n58486 , n18546 );
not ( n58487 , n58486 );
buf ( n58488 , n22402 );
and ( n58489 , n58487 , n58488 );
buf ( n58490 , n18514 );
not ( n58491 , n58490 );
buf ( n58492 , n21639 );
and ( n58493 , n58491 , n58492 );
xnor ( n58494 , n58486 , n58488 );
and ( n58495 , n58493 , n58494 );
or ( n58496 , n58489 , n58495 );
xnor ( n58497 , n58482 , n58484 );
and ( n58498 , n58496 , n58497 );
or ( n58499 , n58485 , n58498 );
xnor ( n58500 , n58478 , n58480 );
and ( n58501 , n58499 , n58500 );
or ( n58502 , n58481 , n58501 );
xnor ( n58503 , n58474 , n58476 );
and ( n58504 , n58502 , n58503 );
or ( n58505 , n58477 , n58504 );
xnor ( n58506 , n58470 , n58472 );
and ( n58507 , n58505 , n58506 );
or ( n58508 , n58473 , n58507 );
xnor ( n58509 , n58466 , n58468 );
and ( n58510 , n58508 , n58509 );
or ( n58511 , n58469 , n58510 );
xnor ( n58512 , n58462 , n58464 );
and ( n58513 , n58511 , n58512 );
or ( n58514 , n58465 , n58513 );
xnor ( n58515 , n58458 , n58460 );
and ( n58516 , n58514 , n58515 );
or ( n58517 , n58461 , n58516 );
xnor ( n58518 , n58454 , n58456 );
and ( n58519 , n58517 , n58518 );
or ( n58520 , n58457 , n58519 );
xnor ( n58521 , n58450 , n58452 );
and ( n58522 , n58520 , n58521 );
or ( n58523 , n58453 , n58522 );
xnor ( n58524 , n58446 , n58448 );
and ( n58525 , n58523 , n58524 );
or ( n58526 , n58449 , n58525 );
xnor ( n58527 , n58442 , n58444 );
and ( n58528 , n58526 , n58527 );
or ( n58529 , n58445 , n58528 );
xnor ( n58530 , n58438 , n58440 );
and ( n58531 , n58529 , n58530 );
or ( n58532 , n58441 , n58531 );
xnor ( n58533 , n58434 , n58436 );
and ( n58534 , n58532 , n58533 );
or ( n58535 , n58437 , n58534 );
xnor ( n58536 , n58430 , n58432 );
and ( n58537 , n58535 , n58536 );
or ( n58538 , n58433 , n58537 );
xnor ( n58539 , n58426 , n58428 );
and ( n58540 , n58538 , n58539 );
or ( n58541 , n58429 , n58540 );
xnor ( n58542 , n58422 , n58424 );
and ( n58543 , n58541 , n58542 );
or ( n58544 , n58425 , n58543 );
xnor ( n58545 , n58418 , n58420 );
and ( n58546 , n58544 , n58545 );
or ( n58547 , n58421 , n58546 );
xnor ( n58548 , n58414 , n58416 );
and ( n58549 , n58547 , n58548 );
or ( n58550 , n58417 , n58549 );
xnor ( n58551 , n58410 , n58412 );
and ( n58552 , n58550 , n58551 );
or ( n58553 , n58413 , n58552 );
xnor ( n58554 , n58406 , n58408 );
and ( n58555 , n58553 , n58554 );
or ( n58556 , n58409 , n58555 );
xnor ( n58557 , n58402 , n58404 );
and ( n58558 , n58556 , n58557 );
or ( n58559 , n58405 , n58558 );
xnor ( n58560 , n58398 , n58400 );
and ( n58561 , n58559 , n58560 );
or ( n58562 , n58401 , n58561 );
xnor ( n58563 , n58394 , n58396 );
and ( n58564 , n58562 , n58563 );
or ( n58565 , n58397 , n58564 );
xnor ( n58566 , n58390 , n58392 );
and ( n58567 , n58565 , n58566 );
or ( n58568 , n58393 , n58567 );
xnor ( n58569 , n58386 , n58388 );
and ( n58570 , n58568 , n58569 );
or ( n58571 , n58389 , n58570 );
xnor ( n58572 , n58382 , n58384 );
and ( n58573 , n58571 , n58572 );
or ( n58574 , n58385 , n58573 );
xnor ( n58575 , n58378 , n58380 );
and ( n58576 , n58574 , n58575 );
or ( n58577 , n58381 , n58576 );
xnor ( n58578 , n58374 , n58376 );
and ( n58579 , n58577 , n58578 );
or ( n58580 , n58377 , n58579 );
xnor ( n58581 , n58370 , n58372 );
and ( n58582 , n58580 , n58581 );
or ( n58583 , n58373 , n58582 );
and ( n58584 , n58369 , n58583 );
not ( n58585 , n58367 );
and ( n58586 , n58585 , n58366 );
and ( n58587 , n58586 , n58368 );
or ( n58588 , n58584 , n58587 );
buf ( n58589 , n58588 );
not ( n58590 , n58589 );
or ( n58591 , n58590 , n19750 );
and ( n58592 , n58591 , n23061 );
or ( n58593 , n58589 , n19750 );
and ( n58594 , n58593 , n23822 );
and ( n58595 , n57998 , n23059 );
and ( n58596 , n57997 , n23058 );
and ( n58597 , n58226 , n23820 );
and ( n58598 , n58229 , n23819 );
and ( n58599 , n58361 , n23831 );
and ( n58600 , n58360 , n23830 );
and ( n58601 , n58590 , n23834 );
and ( n58602 , n58589 , n23917 );
or ( n58603 , n58000 , n58002 , n58228 , n58231 , n58363 , n58365 , n58592 , n58594 , n58595 , n58596 , n58597 , n58598 , n58599 , n58600 , n58601 , n58602 );
and ( n58604 , n58603 , n17162 );
or ( n58605 , n57732 , n58604 );
and ( n58606 , n58605 , n23924 );
and ( n58607 , n19750 , n23926 );
or ( n58608 , n58606 , n58607 );
buf ( n58609 , n58608 );
buf ( n58610 , n58609 );
buf ( n58611 , n10615 );
buf ( n58612 , n10613 );
buf ( n58613 , n10615 );
not ( n58614 , n24800 );
and ( n58615 , n26699 , n25222 );
and ( n58616 , n43420 , n28583 );
and ( n58617 , n26699 , n28591 );
or ( n58618 , n58616 , n58617 );
and ( n58619 , n58618 , n28594 );
and ( n58620 , n43436 , n28583 );
and ( n58621 , n26699 , n28591 );
or ( n58622 , n58620 , n58621 );
and ( n58623 , n58622 , n30269 );
and ( n58624 , n43452 , n28583 );
and ( n58625 , n26699 , n28591 );
or ( n58626 , n58624 , n58625 );
and ( n58627 , n58626 , n30982 );
and ( n58628 , n29172 , n28583 );
and ( n58629 , n26699 , n28591 );
or ( n58630 , n58628 , n58629 );
and ( n58631 , n58630 , n30989 );
and ( n58632 , n26697 , n30991 );
and ( n58633 , n43471 , n28583 );
and ( n58634 , n26699 , n28591 );
or ( n58635 , n58633 , n58634 );
and ( n58636 , n58635 , n31002 );
or ( n58637 , n58615 , n58619 , n58623 , n58627 , n58631 , n58632 , n58636 );
and ( n58638 , n58614 , n58637 );
and ( n58639 , n26699 , n24800 );
or ( n58640 , n58638 , n58639 );
and ( n58641 , n58640 , n31008 );
and ( n58642 , n26699 , n10618 );
or ( n58643 , n58641 , n58642 );
buf ( n58644 , n58643 );
buf ( n58645 , n58644 );
buf ( n58646 , n10615 );
buf ( n58647 , n10613 );
not ( n58648 , n24800 );
and ( n58649 , n26153 , n25222 );
and ( n58650 , n50001 , n28589 );
and ( n58651 , n26153 , n31075 );
or ( n58652 , n58650 , n58651 );
and ( n58653 , n58652 , n28594 );
and ( n58654 , n50011 , n28589 );
and ( n58655 , n26153 , n31075 );
or ( n58656 , n58654 , n58655 );
and ( n58657 , n58656 , n30269 );
and ( n58658 , n50021 , n28589 );
and ( n58659 , n26153 , n31075 );
or ( n58660 , n58658 , n58659 );
and ( n58661 , n58660 , n30982 );
and ( n58662 , n29495 , n28589 );
and ( n58663 , n26153 , n31075 );
or ( n58664 , n58662 , n58663 );
and ( n58665 , n58664 , n30989 );
and ( n58666 , n29495 , n30991 );
and ( n58667 , n50032 , n28589 );
and ( n58668 , n26153 , n31075 );
or ( n58669 , n58667 , n58668 );
and ( n58670 , n58669 , n31002 );
or ( n58671 , n58649 , n58653 , n58657 , n58661 , n58665 , n58666 , n58670 );
and ( n58672 , n58648 , n58671 );
and ( n58673 , n26153 , n24800 );
or ( n58674 , n58672 , n58673 );
and ( n58675 , n58674 , n31008 );
and ( n58676 , n25354 , n10618 );
or ( n58677 , n58675 , n58676 );
buf ( n58678 , n58677 );
buf ( n58679 , n58678 );
buf ( n58680 , n10615 );
buf ( n58681 , n10615 );
not ( n58682 , n24511 );
not ( n58683 , n24799 );
and ( n58684 , n10720 , n40154 );
not ( n58685 , n40632 );
and ( n58686 , n58685 , n40356 );
xor ( n58687 , n40647 , n40653 );
and ( n58688 , n58687 , n40632 );
or ( n58689 , n58686 , n58688 );
buf ( n58690 , n58689 );
and ( n58691 , n58690 , n27046 );
not ( n58692 , n41147 );
and ( n58693 , n58692 , n40871 );
xor ( n58694 , n41162 , n41168 );
and ( n58695 , n58694 , n41147 );
or ( n58696 , n58693 , n58695 );
buf ( n58697 , n58696 );
and ( n58698 , n58697 , n27049 );
and ( n58699 , n29613 , n28506 );
and ( n58700 , n10720 , n28508 );
or ( n58701 , n58691 , n58698 , n58699 , n58700 );
and ( n58702 , n58701 , n41199 );
or ( n58703 , n58684 , n58702 );
and ( n58704 , n58683 , n58703 );
xor ( n58705 , n41708 , n41716 );
xor ( n58706 , n58705 , n41770 );
buf ( n58707 , n58706 );
and ( n58708 , n58707 , n27046 );
xor ( n58709 , n42231 , n42232 );
xor ( n58710 , n58709 , n42266 );
buf ( n58711 , n58710 );
and ( n58712 , n58711 , n27049 );
and ( n58713 , n29613 , n42306 );
or ( n58714 , n58708 , n58712 , n58713 );
buf ( n58715 , n58714 );
and ( n58716 , C1 , n58715 );
or ( n58717 , n58716 , C0 );
buf ( n58718 , n58717 );
not ( n58719 , n58718 );
buf ( n58720 , n58719 );
buf ( n58721 , n58720 );
not ( n58722 , n58721 );
and ( n58723 , C1 , n58722 );
or ( n58724 , n58723 , C0 );
buf ( n58725 , n58724 );
and ( n58726 , n58725 , n24799 );
or ( n58727 , n58704 , n58726 );
and ( n58728 , n58682 , n58727 );
and ( n58729 , n58701 , n24511 );
or ( n58730 , n58728 , n58729 );
and ( n58731 , n58730 , n31008 );
not ( n58732 , n42601 );
and ( n58733 , n58732 , n42373 );
xor ( n58734 , n42616 , n42622 );
and ( n58735 , n58734 , n42601 );
or ( n58736 , n58733 , n58735 );
buf ( n58737 , n58736 );
and ( n58738 , n58737 , n10618 );
or ( n58739 , n58731 , n58738 );
buf ( n58740 , n58739 );
buf ( n58741 , n58740 );
not ( n58742 , n17451 );
and ( n58743 , n34421 , n21333 );
and ( n58744 , n19217 , n34758 );
or ( n58745 , n58743 , n58744 );
and ( n58746 , n58745 , n21341 );
and ( n58747 , n34431 , n21333 );
and ( n58748 , n19217 , n34758 );
or ( n58749 , n58747 , n58748 );
and ( n58750 , n58749 , n23064 );
and ( n58751 , n34441 , n21333 );
and ( n58752 , n19217 , n34758 );
or ( n58753 , n58751 , n58752 );
and ( n58754 , n58753 , n23825 );
and ( n58755 , n21971 , n21333 );
and ( n58756 , n19217 , n34758 );
or ( n58757 , n58755 , n58756 );
and ( n58758 , n58757 , n23832 );
and ( n58759 , n34452 , n21333 );
and ( n58760 , n19217 , n34758 );
or ( n58761 , n58759 , n58760 );
and ( n58762 , n58761 , n23917 );
and ( n58763 , n19217 , n34526 );
or ( n58764 , n58746 , n58750 , n58754 , n58758 , n58762 , n58763 );
and ( n58765 , n58742 , n58764 );
and ( n58766 , n19217 , n17451 );
or ( n58767 , n58765 , n58766 );
and ( n58768 , n58767 , n23924 );
and ( n58769 , n19217 , n23926 );
or ( n58770 , n58768 , n58769 );
buf ( n58771 , n58770 );
buf ( n58772 , n58771 );
not ( n58773 , n34804 );
and ( n58774 , n58773 , n26433 );
and ( n58775 , n14731 , n34804 );
or ( n58776 , n58774 , n58775 );
and ( n58777 , n58776 , n31008 );
and ( n58778 , n14731 , n10618 );
or ( n58779 , n58777 , n58778 );
buf ( n58780 , n58779 );
buf ( n58781 , n58780 );
and ( n58782 , n11649 , n16574 );
and ( n58783 , n15726 , n16576 );
or ( n58784 , n58782 , n58783 );
buf ( n58785 , n58784 );
buf ( n58786 , n58785 );
not ( n58787 , n17451 );
and ( n58788 , n51973 , n21334 );
and ( n58789 , n18743 , n34492 );
or ( n58790 , n58788 , n58789 );
and ( n58791 , n58790 , n21341 );
and ( n58792 , n51983 , n21334 );
and ( n58793 , n18743 , n34492 );
or ( n58794 , n58792 , n58793 );
and ( n58795 , n58794 , n23064 );
and ( n58796 , n51993 , n21334 );
and ( n58797 , n18743 , n34492 );
or ( n58798 , n58796 , n58797 );
and ( n58799 , n58798 , n23825 );
and ( n58800 , n22282 , n21334 );
and ( n58801 , n18743 , n34492 );
or ( n58802 , n58800 , n58801 );
and ( n58803 , n58802 , n23832 );
and ( n58804 , n52004 , n21334 );
and ( n58805 , n18743 , n34492 );
or ( n58806 , n58804 , n58805 );
and ( n58807 , n58806 , n23917 );
and ( n58808 , n18743 , n34526 );
or ( n58809 , n58791 , n58795 , n58799 , n58803 , n58807 , n58808 );
and ( n58810 , n58787 , n58809 );
and ( n58811 , n18743 , n17451 );
or ( n58812 , n58810 , n58811 );
and ( n58813 , n58812 , n23924 );
and ( n58814 , n18743 , n23926 );
or ( n58815 , n58813 , n58814 );
buf ( n58816 , n58815 );
buf ( n58817 , n58816 );
buf ( n58818 , n10613 );
not ( n58819 , n17451 );
and ( n58820 , n19009 , n17873 );
not ( n58821 , n19474 );
and ( n58822 , n58821 , n18995 );
xor ( n58823 , n19487 , n19515 );
and ( n58824 , n58823 , n19474 );
or ( n58825 , n58822 , n58824 );
buf ( n58826 , n58825 );
and ( n58827 , n58826 , n19745 );
and ( n58828 , n58826 , n19748 );
not ( n58829 , n19750 );
and ( n58830 , n58829 , n20899 );
not ( n58831 , n21193 );
and ( n58832 , n58831 , n20911 );
xor ( n58833 , n21206 , n21236 );
and ( n58834 , n58833 , n21193 );
or ( n58835 , n58832 , n58834 );
buf ( n58836 , n58835 );
and ( n58837 , n58836 , n19750 );
or ( n58838 , n58830 , n58837 );
and ( n58839 , n58838 , n21253 );
and ( n58840 , n20899 , n21255 );
or ( n58841 , n58827 , n58828 , n58839 , n58840 );
and ( n58842 , n58841 , n21336 );
and ( n58843 , n19009 , n42682 );
or ( n58844 , n58842 , n58843 );
and ( n58845 , n58844 , n21341 );
not ( n58846 , n22996 );
and ( n58847 , n58846 , n22754 );
xor ( n58848 , n23009 , n23039 );
and ( n58849 , n58848 , n22996 );
or ( n58850 , n58847 , n58849 );
buf ( n58851 , n58850 );
and ( n58852 , n58851 , n21336 );
and ( n58853 , n19009 , n42682 );
or ( n58854 , n58852 , n58853 );
and ( n58855 , n58854 , n23064 );
not ( n58856 , n23758 );
and ( n58857 , n58856 , n23516 );
xor ( n58858 , n23771 , n23801 );
and ( n58859 , n58858 , n23758 );
or ( n58860 , n58857 , n58859 );
buf ( n58861 , n58860 );
and ( n58862 , n58861 , n21336 );
and ( n58863 , n19009 , n42682 );
or ( n58864 , n58862 , n58863 );
and ( n58865 , n58864 , n23825 );
and ( n58866 , n22122 , n21336 );
and ( n58867 , n19009 , n42682 );
or ( n58868 , n58866 , n58867 );
and ( n58869 , n58868 , n23832 );
and ( n58870 , n22122 , n23834 );
xor ( n58871 , n23857 , n23901 );
buf ( n58872 , n58871 );
and ( n58873 , n58872 , n21336 );
and ( n58874 , n19009 , n42682 );
or ( n58875 , n58873 , n58874 );
and ( n58876 , n58875 , n23917 );
or ( n58877 , n58820 , n58845 , n58855 , n58865 , n58869 , n58870 , n58876 );
and ( n58878 , n58819 , n58877 );
and ( n58879 , n19009 , n17451 );
or ( n58880 , n58878 , n58879 );
and ( n58881 , n58880 , n23924 );
and ( n58882 , n18095 , n23926 );
or ( n58883 , n58881 , n58882 );
buf ( n58884 , n58883 );
buf ( n58885 , n58884 );
not ( n58886 , n34821 );
and ( n58887 , n49200 , n36345 );
and ( n58888 , n13197 , n36352 );
or ( n58889 , n58887 , n58888 );
and ( n58890 , n58889 , n14562 );
and ( n58891 , n49210 , n36345 );
and ( n58892 , n13197 , n37073 );
or ( n58893 , n58891 , n58892 );
and ( n58894 , n58893 , n14586 );
and ( n58895 , n49220 , n36350 );
and ( n58896 , n13197 , n37825 );
or ( n58897 , n58895 , n58896 );
and ( n58898 , n58897 , n14584 );
and ( n58899 , n49210 , n36350 );
and ( n58900 , n13197 , n37831 );
or ( n58901 , n58899 , n58900 );
and ( n58902 , n58901 , n37835 );
and ( n58903 , n49220 , n36350 );
and ( n58904 , n13197 , n37831 );
or ( n58905 , n58903 , n58904 );
and ( n58906 , n58905 , n37841 );
and ( n58907 , n15037 , n36350 );
and ( n58908 , n13197 , n37831 );
or ( n58909 , n58907 , n58908 );
and ( n58910 , n58909 , n37847 );
and ( n58911 , n13197 , n37849 );
or ( n58912 , n58890 , n58894 , n58898 , n58902 , n58906 , n58910 , n58911 );
and ( n58913 , n58886 , n58912 );
and ( n58914 , n13197 , n34821 );
or ( n58915 , n58913 , n58914 );
and ( n58916 , n58915 , n16574 );
and ( n58917 , n13197 , n16576 );
or ( n58918 , n58916 , n58917 );
buf ( n58919 , n58918 );
buf ( n58920 , n58919 );
buf ( n58921 , n10615 );
buf ( n58922 , n10615 );
and ( n58923 , n11585 , n16574 );
and ( n58924 , n15550 , n16576 );
or ( n58925 , n58923 , n58924 );
buf ( n58926 , n58925 );
buf ( n58927 , n58926 );
not ( n58928 , n34821 );
and ( n58929 , n13217 , n14592 );
and ( n58930 , n57550 , n36348 );
and ( n58931 , n13217 , n43530 );
or ( n58932 , n58930 , n58931 );
and ( n58933 , n58932 , n14562 );
and ( n58934 , n57560 , n36347 );
and ( n58935 , n13217 , n43543 );
or ( n58936 , n58934 , n58935 );
and ( n58937 , n58936 , n14586 );
and ( n58938 , n57570 , n36348 );
and ( n58939 , n13217 , n43556 );
or ( n58940 , n58938 , n58939 );
and ( n58941 , n58940 , n14584 );
and ( n58942 , n57560 , n36347 );
and ( n58943 , n13217 , n43563 );
or ( n58944 , n58942 , n58943 );
and ( n58945 , n58944 , n37835 );
and ( n58946 , n57570 , n36347 );
and ( n58947 , n13217 , n43563 );
or ( n58948 , n58946 , n58947 );
and ( n58949 , n58948 , n37841 );
and ( n58950 , n13215 , n14564 );
and ( n58951 , n15067 , n36347 );
and ( n58952 , n13217 , n43563 );
or ( n58953 , n58951 , n58952 );
and ( n58954 , n58953 , n37847 );
or ( n58955 , n58929 , n58933 , n58937 , n58941 , n58945 , n58949 , n58950 , n58954 );
and ( n58956 , n58928 , n58955 );
and ( n58957 , n13217 , n34821 );
or ( n58958 , n58956 , n58957 );
and ( n58959 , n58958 , n16574 );
and ( n58960 , n13217 , n16576 );
or ( n58961 , n58959 , n58960 );
buf ( n58962 , n58961 );
buf ( n58963 , n58962 );
buf ( n58964 , n10613 );
buf ( n58965 , n10615 );
buf ( n58966 , n10615 );
buf ( n58967 , n10615 );
not ( n58968 , n24800 );
and ( n58969 , n48113 , n28586 );
and ( n58970 , n26395 , n34573 );
or ( n58971 , n58969 , n58970 );
and ( n58972 , n58971 , n28594 );
and ( n58973 , n48123 , n28586 );
and ( n58974 , n26395 , n34573 );
or ( n58975 , n58973 , n58974 );
and ( n58976 , n58975 , n30269 );
and ( n58977 , n48133 , n28586 );
and ( n58978 , n26395 , n34573 );
or ( n58979 , n58977 , n58978 );
and ( n58980 , n58979 , n30982 );
and ( n58981 , n29355 , n28586 );
and ( n58982 , n26395 , n34573 );
or ( n58983 , n58981 , n58982 );
and ( n58984 , n58983 , n30989 );
and ( n58985 , n48144 , n28586 );
and ( n58986 , n26395 , n34573 );
or ( n58987 , n58985 , n58986 );
and ( n58988 , n58987 , n31002 );
and ( n58989 , n26395 , n34607 );
or ( n58990 , n58972 , n58976 , n58980 , n58984 , n58988 , n58989 );
and ( n58991 , n58968 , n58990 );
and ( n58992 , n26395 , n24800 );
or ( n58993 , n58991 , n58992 );
and ( n58994 , n58993 , n31008 );
and ( n58995 , n26395 , n10618 );
or ( n58996 , n58994 , n58995 );
buf ( n58997 , n58996 );
buf ( n58998 , n58997 );
buf ( n58999 , n10615 );
buf ( n59000 , n10613 );
and ( n59001 , n16897 , n23924 );
and ( n59002 , n22393 , n23926 );
or ( n59003 , n59001 , n59002 );
buf ( n59004 , n59003 );
buf ( n59005 , n59004 );
buf ( n59006 , n10613 );
buf ( n59007 , n10615 );
not ( n59008 , n17451 );
and ( n59009 , n45943 , n21334 );
and ( n59010 , n19049 , n34492 );
or ( n59011 , n59009 , n59010 );
and ( n59012 , n59011 , n21341 );
and ( n59013 , n45953 , n21334 );
and ( n59014 , n19049 , n34492 );
or ( n59015 , n59013 , n59014 );
and ( n59016 , n59015 , n23064 );
and ( n59017 , n45963 , n21334 );
and ( n59018 , n19049 , n34492 );
or ( n59019 , n59017 , n59018 );
and ( n59020 , n59019 , n23825 );
and ( n59021 , n22102 , n21334 );
and ( n59022 , n19049 , n34492 );
or ( n59023 , n59021 , n59022 );
and ( n59024 , n59023 , n23832 );
and ( n59025 , n45974 , n21334 );
and ( n59026 , n19049 , n34492 );
or ( n59027 , n59025 , n59026 );
and ( n59028 , n59027 , n23917 );
and ( n59029 , n19049 , n34526 );
or ( n59030 , n59012 , n59016 , n59020 , n59024 , n59028 , n59029 );
and ( n59031 , n59008 , n59030 );
and ( n59032 , n19049 , n17451 );
or ( n59033 , n59031 , n59032 );
and ( n59034 , n59033 , n23924 );
and ( n59035 , n19049 , n23926 );
or ( n59036 , n59034 , n59035 );
buf ( n59037 , n59036 );
buf ( n59038 , n59037 );
buf ( n59039 , n10615 );
buf ( n59040 , n10615 );
not ( n59041 , n34538 );
and ( n59042 , n59041 , n19458 );
and ( n59043 , n14663 , n34538 );
or ( n59044 , n59042 , n59043 );
and ( n59045 , n59044 , n23924 );
and ( n59046 , n14663 , n23926 );
or ( n59047 , n59045 , n59046 );
buf ( n59048 , n59047 );
buf ( n59049 , n59048 );
not ( n59050 , n34821 );
and ( n59051 , n48401 , n36347 );
and ( n59052 , n13399 , n39408 );
or ( n59053 , n59051 , n59052 );
and ( n59054 , n59053 , n14562 );
and ( n59055 , n48411 , n36348 );
and ( n59056 , n13399 , n39427 );
or ( n59057 , n59055 , n59056 );
and ( n59058 , n59057 , n14586 );
and ( n59059 , n48421 , n36347 );
and ( n59060 , n13399 , n39446 );
or ( n59061 , n59059 , n59060 );
and ( n59062 , n59061 , n14584 );
and ( n59063 , n48411 , n36348 );
and ( n59064 , n13399 , n39453 );
or ( n59065 , n59063 , n59064 );
and ( n59066 , n59065 , n37835 );
and ( n59067 , n48421 , n36348 );
and ( n59068 , n13399 , n39453 );
or ( n59069 , n59067 , n59068 );
and ( n59070 , n59069 , n37841 );
and ( n59071 , n15691 , n36348 );
and ( n59072 , n13399 , n39453 );
or ( n59073 , n59071 , n59072 );
and ( n59074 , n59073 , n37847 );
and ( n59075 , n13399 , n37849 );
or ( n59076 , n59054 , n59058 , n59062 , n59066 , n59070 , n59074 , n59075 );
and ( n59077 , n59050 , n59076 );
and ( n59078 , n13399 , n34821 );
or ( n59079 , n59077 , n59078 );
and ( n59080 , n59079 , n16574 );
and ( n59081 , n13399 , n16576 );
or ( n59082 , n59080 , n59081 );
buf ( n59083 , n59082 );
buf ( n59084 , n59083 );
buf ( n59085 , n10615 );
buf ( n59086 , n10615 );
buf ( n59087 , n10613 );
buf ( n59088 , n10615 );
buf ( n59089 , n10613 );
not ( n59090 , n34538 );
and ( n59091 , n59090 , n18643 );
and ( n59092 , n14807 , n34538 );
or ( n59093 , n59091 , n59092 );
and ( n59094 , n59093 , n23924 );
and ( n59095 , n14807 , n23926 );
or ( n59096 , n59094 , n59095 );
buf ( n59097 , n59096 );
buf ( n59098 , n59097 );
buf ( n59099 , n10615 );
buf ( n59100 , n10615 );
not ( n59101 , n11333 );
and ( n59102 , n59101 , n11125 );
xor ( n59103 , n11344 , n11358 );
and ( n59104 , n59103 , n11333 );
or ( n59105 , n59102 , n59104 );
buf ( n59106 , n59105 );
buf ( n59107 , n59106 );
buf ( n59108 , n10615 );
buf ( n59109 , n10615 );
buf ( n59110 , n10615 );
buf ( n59111 , n10613 );
not ( n59112 , n34821 );
and ( n59113 , n51156 , n36347 );
and ( n59114 , n13291 , n39408 );
or ( n59115 , n59113 , n59114 );
and ( n59116 , n59115 , n14562 );
and ( n59117 , n51166 , n36348 );
and ( n59118 , n13291 , n39427 );
or ( n59119 , n59117 , n59118 );
and ( n59120 , n59119 , n14586 );
and ( n59121 , n51176 , n36347 );
and ( n59122 , n13291 , n39446 );
or ( n59123 , n59121 , n59122 );
and ( n59124 , n59123 , n14584 );
and ( n59125 , n51166 , n36348 );
and ( n59126 , n13291 , n39453 );
or ( n59127 , n59125 , n59126 );
and ( n59128 , n59127 , n37835 );
and ( n59129 , n51176 , n36348 );
and ( n59130 , n13291 , n39453 );
or ( n59131 , n59129 , n59130 );
and ( n59132 , n59131 , n37841 );
and ( n59133 , n15493 , n36348 );
and ( n59134 , n13291 , n39453 );
or ( n59135 , n59133 , n59134 );
and ( n59136 , n59135 , n37847 );
and ( n59137 , n13291 , n37849 );
or ( n59138 , n59116 , n59120 , n59124 , n59128 , n59132 , n59136 , n59137 );
and ( n59139 , n59112 , n59138 );
and ( n59140 , n13291 , n34821 );
or ( n59141 , n59139 , n59140 );
and ( n59142 , n59141 , n16574 );
and ( n59143 , n13291 , n16576 );
or ( n59144 , n59142 , n59143 );
buf ( n59145 , n59144 );
buf ( n59146 , n59145 );
buf ( n59147 , n10615 );
buf ( n59148 , n10615 );
buf ( n59149 , n10613 );
buf ( n59150 , n10613 );
not ( n59151 , n17451 );
and ( n59152 , n52940 , n21334 );
and ( n59153 , n18525 , n34492 );
or ( n59154 , n59152 , n59153 );
and ( n59155 , n59154 , n21341 );
and ( n59156 , n18525 , n34492 );
buf ( n59157 , n59156 );
and ( n59158 , n59157 , n23064 );
and ( n59159 , n18525 , n34492 );
buf ( n59160 , n59159 );
and ( n59161 , n59160 , n23825 );
and ( n59162 , n21841 , n21334 );
and ( n59163 , n18525 , n34492 );
or ( n59164 , n59162 , n59163 );
and ( n59165 , n59164 , n23832 );
and ( n59166 , n52959 , n21334 );
and ( n59167 , n18525 , n34492 );
or ( n59168 , n59166 , n59167 );
and ( n59169 , n59168 , n23917 );
and ( n59170 , n18525 , n34526 );
or ( n59171 , n59155 , n59158 , n59161 , n59165 , n59169 , n59170 );
and ( n59172 , n59151 , n59171 );
and ( n59173 , n18525 , n17451 );
or ( n59174 , n59172 , n59173 );
and ( n59175 , n59174 , n23924 );
and ( n59176 , n18525 , n23926 );
or ( n59177 , n59175 , n59176 );
buf ( n59178 , n59177 );
buf ( n59179 , n59178 );
buf ( n59180 , n10615 );
buf ( n59181 , n10613 );
not ( n59182 , n34821 );
and ( n59183 , n48669 , n36345 );
and ( n59184 , n13329 , n36352 );
or ( n59185 , n59183 , n59184 );
and ( n59186 , n59185 , n14562 );
and ( n59187 , n48679 , n36345 );
and ( n59188 , n13329 , n37073 );
or ( n59189 , n59187 , n59188 );
and ( n59190 , n59189 , n14586 );
and ( n59191 , n48689 , n36350 );
and ( n59192 , n13329 , n37825 );
or ( n59193 , n59191 , n59192 );
and ( n59194 , n59193 , n14584 );
and ( n59195 , n48679 , n36350 );
and ( n59196 , n13329 , n37831 );
or ( n59197 , n59195 , n59196 );
and ( n59198 , n59197 , n37835 );
and ( n59199 , n48689 , n36350 );
and ( n59200 , n13329 , n37831 );
or ( n59201 , n59199 , n59200 );
and ( n59202 , n59201 , n37841 );
and ( n59203 , n15559 , n36350 );
and ( n59204 , n13329 , n37831 );
or ( n59205 , n59203 , n59204 );
and ( n59206 , n59205 , n37847 );
and ( n59207 , n13329 , n37849 );
or ( n59208 , n59186 , n59190 , n59194 , n59198 , n59202 , n59206 , n59207 );
and ( n59209 , n59182 , n59208 );
and ( n59210 , n13329 , n34821 );
or ( n59211 , n59209 , n59210 );
and ( n59212 , n59211 , n16574 );
and ( n59213 , n13329 , n16576 );
or ( n59214 , n59212 , n59213 );
buf ( n59215 , n59214 );
buf ( n59216 , n59215 );
buf ( n59217 , n10615 );
buf ( n59218 , n10615 );
buf ( n59219 , n10613 );
and ( n59220 , n16712 , n23924 );
and ( n59221 , n21839 , n23926 );
or ( n59222 , n59220 , n59221 );
buf ( n59223 , n59222 );
buf ( n59224 , n59223 );
not ( n59225 , n34804 );
and ( n59226 , n24799 , n59225 );
and ( n59227 , n59226 , n31008 );
buf ( n59228 , n59227 );
buf ( n59229 , n59228 );
buf ( n59230 , n10613 );
not ( n59231 , n34821 );
and ( n59232 , n45647 , n36345 );
and ( n59233 , n13365 , n36352 );
or ( n59234 , n59232 , n59233 );
and ( n59235 , n59234 , n14562 );
and ( n59236 , n45657 , n36345 );
and ( n59237 , n13365 , n37073 );
or ( n59238 , n59236 , n59237 );
and ( n59239 , n59238 , n14586 );
and ( n59240 , n45667 , n36350 );
and ( n59241 , n13365 , n37825 );
or ( n59242 , n59240 , n59241 );
and ( n59243 , n59242 , n14584 );
and ( n59244 , n45657 , n36350 );
and ( n59245 , n13365 , n37831 );
or ( n59246 , n59244 , n59245 );
and ( n59247 , n59246 , n37835 );
and ( n59248 , n45667 , n36350 );
and ( n59249 , n13365 , n37831 );
or ( n59250 , n59248 , n59249 );
and ( n59251 , n59250 , n37841 );
and ( n59252 , n15625 , n36350 );
and ( n59253 , n13365 , n37831 );
or ( n59254 , n59252 , n59253 );
and ( n59255 , n59254 , n37847 );
and ( n59256 , n13365 , n37849 );
or ( n59257 , n59235 , n59239 , n59243 , n59247 , n59251 , n59255 , n59256 );
and ( n59258 , n59231 , n59257 );
and ( n59259 , n13365 , n34821 );
or ( n59260 , n59258 , n59259 );
and ( n59261 , n59260 , n16574 );
and ( n59262 , n13365 , n16576 );
or ( n59263 , n59261 , n59262 );
buf ( n59264 , n59263 );
buf ( n59265 , n59264 );
and ( n59266 , n24222 , n31008 );
and ( n59267 , n29586 , n10618 );
or ( n59268 , n59266 , n59267 );
buf ( n59269 , n59268 );
buf ( n59270 , n59269 );
not ( n59271 , n34538 );
and ( n59272 , n59271 , n19153 );
and ( n59273 , n14717 , n34538 );
or ( n59274 , n59272 , n59273 );
and ( n59275 , n59274 , n23924 );
and ( n59276 , n14717 , n23926 );
or ( n59277 , n59275 , n59276 );
buf ( n59278 , n59277 );
buf ( n59279 , n59278 );
not ( n59280 , n34821 );
and ( n59281 , n13251 , n14592 );
and ( n59282 , n57357 , n36350 );
and ( n59283 , n13251 , n43691 );
or ( n59284 , n59282 , n59283 );
and ( n59285 , n59284 , n14562 );
and ( n59286 , n57367 , n36350 );
and ( n59287 , n13251 , n43703 );
or ( n59288 , n59286 , n59287 );
and ( n59289 , n59288 , n14586 );
and ( n59290 , n57377 , n36345 );
and ( n59291 , n13251 , n43715 );
or ( n59292 , n59290 , n59291 );
and ( n59293 , n59292 , n14584 );
and ( n59294 , n57367 , n36345 );
and ( n59295 , n13251 , n43721 );
or ( n59296 , n59294 , n59295 );
and ( n59297 , n59296 , n37835 );
and ( n59298 , n57377 , n36345 );
and ( n59299 , n13251 , n43721 );
or ( n59300 , n59298 , n59299 );
and ( n59301 , n59300 , n37841 );
and ( n59302 , n15112 , n14564 );
and ( n59303 , n15112 , n36345 );
and ( n59304 , n13251 , n43721 );
or ( n59305 , n59303 , n59304 );
and ( n59306 , n59305 , n37847 );
or ( n59307 , n59281 , n59285 , n59289 , n59293 , n59297 , n59301 , n59302 , n59306 );
and ( n59308 , n59280 , n59307 );
and ( n59309 , n13251 , n34821 );
or ( n59310 , n59308 , n59309 );
and ( n59311 , n59310 , n16574 );
and ( n59312 , n12273 , n16576 );
or ( n59313 , n59311 , n59312 );
buf ( n59314 , n59313 );
buf ( n59315 , n59314 );
not ( n59316 , n17451 );
and ( n59317 , n18977 , n17873 );
and ( n59318 , n49126 , n21330 );
and ( n59319 , n18977 , n21338 );
or ( n59320 , n59318 , n59319 );
and ( n59321 , n59320 , n21341 );
and ( n59322 , n49136 , n21330 );
and ( n59323 , n18977 , n21338 );
or ( n59324 , n59322 , n59323 );
and ( n59325 , n59324 , n23064 );
and ( n59326 , n49146 , n21330 );
and ( n59327 , n18977 , n21338 );
or ( n59328 , n59326 , n59327 );
and ( n59329 , n59328 , n23825 );
and ( n59330 , n22142 , n21330 );
and ( n59331 , n18977 , n21338 );
or ( n59332 , n59330 , n59331 );
and ( n59333 , n59332 , n23832 );
and ( n59334 , n18975 , n23834 );
and ( n59335 , n49157 , n21330 );
and ( n59336 , n18977 , n21338 );
or ( n59337 , n59335 , n59336 );
and ( n59338 , n59337 , n23917 );
or ( n59339 , n59317 , n59321 , n59325 , n59329 , n59333 , n59334 , n59338 );
and ( n59340 , n59316 , n59339 );
and ( n59341 , n18977 , n17451 );
or ( n59342 , n59340 , n59341 );
and ( n59343 , n59342 , n23924 );
and ( n59344 , n18977 , n23926 );
or ( n59345 , n59343 , n59344 );
buf ( n59346 , n59345 );
buf ( n59347 , n59346 );
not ( n59348 , n17451 );
and ( n59349 , n18671 , n17873 );
and ( n59350 , n48886 , n21330 );
and ( n59351 , n18671 , n21338 );
or ( n59352 , n59350 , n59351 );
and ( n59353 , n59352 , n21341 );
and ( n59354 , n48896 , n21330 );
and ( n59355 , n18671 , n21338 );
or ( n59356 , n59354 , n59355 );
and ( n59357 , n59356 , n23064 );
and ( n59358 , n48906 , n21330 );
and ( n59359 , n18671 , n21338 );
or ( n59360 , n59358 , n59359 );
and ( n59361 , n59360 , n23825 );
and ( n59362 , n22322 , n21330 );
and ( n59363 , n18671 , n21338 );
or ( n59364 , n59362 , n59363 );
and ( n59365 , n59364 , n23832 );
and ( n59366 , n18669 , n23834 );
and ( n59367 , n48916 , n21330 );
and ( n59368 , n18671 , n21338 );
or ( n59369 , n59367 , n59368 );
and ( n59370 , n59369 , n23917 );
or ( n59371 , n59349 , n59353 , n59357 , n59361 , n59365 , n59366 , n59370 );
and ( n59372 , n59348 , n59371 );
and ( n59373 , n18671 , n17451 );
or ( n59374 , n59372 , n59373 );
and ( n59375 , n59374 , n23924 );
and ( n59376 , n18671 , n23926 );
or ( n59377 , n59375 , n59376 );
buf ( n59378 , n59377 );
buf ( n59379 , n59378 );
buf ( n59380 , n10615 );
buf ( n59381 , n10615 );
not ( n59382 , n24511 );
not ( n59383 , n24799 );
and ( n59384 , n10730 , n40154 );
not ( n59385 , n40632 );
and ( n59386 , n59385 , n40322 );
xor ( n59387 , n40649 , n40651 );
and ( n59388 , n59387 , n40632 );
or ( n59389 , n59386 , n59388 );
buf ( n59390 , n59389 );
and ( n59391 , n59390 , n27046 );
not ( n59392 , n41147 );
and ( n59393 , n59392 , n40837 );
xor ( n59394 , n41164 , n41166 );
and ( n59395 , n59394 , n41147 );
or ( n59396 , n59393 , n59395 );
buf ( n59397 , n59396 );
and ( n59398 , n59397 , n27049 );
and ( n59399 , n29653 , n28506 );
and ( n59400 , n10730 , n28508 );
or ( n59401 , n59391 , n59398 , n59399 , n59400 );
and ( n59402 , n59401 , n41199 );
or ( n59403 , n59384 , n59402 );
and ( n59404 , n59383 , n59403 );
xor ( n59405 , n41740 , n41748 );
xor ( n59406 , n59405 , n41764 );
buf ( n59407 , n59406 );
and ( n59408 , n59407 , n27046 );
xor ( n59409 , n42249 , n42250 );
xor ( n59410 , n59409 , n42260 );
buf ( n59411 , n59410 );
and ( n59412 , n59411 , n27049 );
and ( n59413 , n29653 , n42306 );
or ( n59414 , n59408 , n59412 , n59413 );
buf ( n59415 , n59414 );
and ( n59416 , C1 , n59415 );
or ( n59417 , n59416 , C0 );
buf ( n59418 , n59417 );
not ( n59419 , n59418 );
buf ( n59420 , n59419 );
buf ( n59421 , n59420 );
not ( n59422 , n59421 );
and ( n59423 , C1 , n59422 );
or ( n59424 , n59423 , C0 );
buf ( n59425 , n59424 );
and ( n59426 , n59425 , n24799 );
or ( n59427 , n59404 , n59426 );
and ( n59428 , n59382 , n59427 );
and ( n59429 , n59401 , n24511 );
or ( n59430 , n59428 , n59429 );
and ( n59431 , n59430 , n31008 );
not ( n59432 , n42601 );
and ( n59433 , n59432 , n42345 );
xor ( n59434 , n42618 , n42620 );
and ( n59435 , n59434 , n42601 );
or ( n59436 , n59433 , n59435 );
buf ( n59437 , n59436 );
and ( n59438 , n59437 , n10618 );
or ( n59439 , n59431 , n59438 );
buf ( n59440 , n59439 );
buf ( n59441 , n59440 );
buf ( n59442 , n10615 );
buf ( n59443 , n10613 );
not ( n59444 , n34804 );
and ( n59445 , n59444 , n26535 );
and ( n59446 , n14713 , n34804 );
or ( n59447 , n59445 , n59446 );
and ( n59448 , n59447 , n31008 );
and ( n59449 , n14713 , n10618 );
or ( n59450 , n59448 , n59449 );
buf ( n59451 , n59450 );
buf ( n59452 , n59451 );
buf ( n59453 , n10615 );
buf ( n59454 , n10613 );
buf ( n59455 , n10613 );
buf ( n59456 , n10615 );
buf ( n59457 , n10615 );
buf ( n59458 , n10613 );
buf ( n59459 , n10613 );
buf ( n59460 , n10615 );
buf ( n59461 , n10615 );
not ( n59462 , n34821 );
not ( n59463 , n13916 );
and ( n59464 , n59463 , n13815 );
xor ( n59465 , n13816 , n13859 );
and ( n59466 , n59465 , n13916 );
or ( n59467 , n59464 , n59466 );
buf ( n59468 , n59467 );
and ( n59469 , n59468 , n14137 );
and ( n59470 , n59468 , n14143 );
not ( n59471 , n14139 );
and ( n59472 , n59471 , n35731 );
not ( n59473 , n36245 );
and ( n59474 , n59473 , n35743 );
xor ( n59475 , n36250 , n36260 );
and ( n59476 , n59475 , n36245 );
or ( n59477 , n59474 , n59476 );
buf ( n59478 , n59477 );
and ( n59479 , n59478 , n14139 );
or ( n59480 , n59472 , n59479 );
and ( n59481 , n59480 , n14140 );
and ( n59482 , n35731 , n14141 );
or ( n59483 , n59469 , n59470 , n59481 , n59482 );
and ( n59484 , n59483 , n36345 );
and ( n59485 , n13437 , n36352 );
or ( n59486 , n59484 , n59485 );
and ( n59487 , n59486 , n14562 );
not ( n59488 , n37048 );
and ( n59489 , n59488 , n36636 );
xor ( n59490 , n37053 , n37063 );
and ( n59491 , n59490 , n37048 );
or ( n59492 , n59489 , n59491 );
buf ( n59493 , n59492 );
and ( n59494 , n59493 , n36345 );
and ( n59495 , n13437 , n37073 );
or ( n59496 , n59494 , n59495 );
and ( n59497 , n59496 , n14586 );
not ( n59498 , n37801 );
and ( n59499 , n59498 , n37389 );
xor ( n59500 , n37806 , n37816 );
and ( n59501 , n59500 , n37801 );
or ( n59502 , n59499 , n59501 );
buf ( n59503 , n59502 );
and ( n59504 , n59503 , n36350 );
and ( n59505 , n13437 , n37825 );
or ( n59506 , n59504 , n59505 );
and ( n59507 , n59506 , n14584 );
and ( n59508 , n59493 , n36350 );
and ( n59509 , n13437 , n37831 );
or ( n59510 , n59508 , n59509 );
and ( n59511 , n59510 , n37835 );
and ( n59512 , n59503 , n36350 );
and ( n59513 , n13437 , n37831 );
or ( n59514 , n59512 , n59513 );
and ( n59515 , n59514 , n37841 );
and ( n59516 , n15757 , n36350 );
and ( n59517 , n13437 , n37831 );
or ( n59518 , n59516 , n59517 );
and ( n59519 , n59518 , n37847 );
and ( n59520 , n13437 , n37849 );
or ( n59521 , n59487 , n59497 , n59507 , n59511 , n59515 , n59519 , n59520 );
and ( n59522 , n59462 , n59521 );
and ( n59523 , n13437 , n34821 );
or ( n59524 , n59522 , n59523 );
and ( n59525 , n59524 , n16574 );
and ( n59526 , n13437 , n16576 );
or ( n59527 , n59525 , n59526 );
buf ( n59528 , n59527 );
buf ( n59529 , n59528 );
not ( n59530 , n17451 );
and ( n59531 , n18941 , n17873 );
and ( n59532 , n42746 , n21336 );
and ( n59533 , n18941 , n42682 );
or ( n59534 , n59532 , n59533 );
and ( n59535 , n59534 , n21341 );
and ( n59536 , n42756 , n21336 );
and ( n59537 , n18941 , n42682 );
or ( n59538 , n59536 , n59537 );
and ( n59539 , n59538 , n23064 );
and ( n59540 , n42766 , n21336 );
and ( n59541 , n18941 , n42682 );
or ( n59542 , n59540 , n59541 );
and ( n59543 , n59542 , n23825 );
and ( n59544 , n22162 , n21336 );
and ( n59545 , n18941 , n42682 );
or ( n59546 , n59544 , n59545 );
and ( n59547 , n59546 , n23832 );
and ( n59548 , n22162 , n23834 );
and ( n59549 , n42776 , n21336 );
and ( n59550 , n18941 , n42682 );
or ( n59551 , n59549 , n59550 );
and ( n59552 , n59551 , n23917 );
or ( n59553 , n59531 , n59535 , n59539 , n59543 , n59547 , n59548 , n59552 );
and ( n59554 , n59530 , n59553 );
and ( n59555 , n18941 , n17451 );
or ( n59556 , n59554 , n59555 );
and ( n59557 , n59556 , n23924 );
and ( n59558 , n18065 , n23926 );
or ( n59559 , n59557 , n59558 );
buf ( n59560 , n59559 );
buf ( n59561 , n59560 );
buf ( n59562 , n10615 );
buf ( n59563 , n10613 );
buf ( n59564 , n10615 );
buf ( n59565 , n10613 );
buf ( n59566 , n10613 );
buf ( n59567 , n10613 );
not ( n59568 , n17451 );
and ( n59569 , n45943 , n21333 );
and ( n59570 , n19047 , n34758 );
or ( n59571 , n59569 , n59570 );
and ( n59572 , n59571 , n21341 );
and ( n59573 , n45953 , n21333 );
and ( n59574 , n19047 , n34758 );
or ( n59575 , n59573 , n59574 );
and ( n59576 , n59575 , n23064 );
and ( n59577 , n45963 , n21333 );
and ( n59578 , n19047 , n34758 );
or ( n59579 , n59577 , n59578 );
and ( n59580 , n59579 , n23825 );
and ( n59581 , n22102 , n21333 );
and ( n59582 , n19047 , n34758 );
or ( n59583 , n59581 , n59582 );
and ( n59584 , n59583 , n23832 );
and ( n59585 , n45974 , n21333 );
and ( n59586 , n19047 , n34758 );
or ( n59587 , n59585 , n59586 );
and ( n59588 , n59587 , n23917 );
and ( n59589 , n19047 , n34526 );
or ( n59590 , n59572 , n59576 , n59580 , n59584 , n59588 , n59589 );
and ( n59591 , n59568 , n59590 );
and ( n59592 , n19047 , n17451 );
or ( n59593 , n59591 , n59592 );
and ( n59594 , n59593 , n23924 );
and ( n59595 , n19047 , n23926 );
or ( n59596 , n59594 , n59595 );
buf ( n59597 , n59596 );
buf ( n59598 , n59597 );
buf ( n59599 , n10613 );
buf ( n59600 , n10615 );
not ( n59601 , n24800 );
and ( n59602 , n26731 , n25222 );
and ( n59603 , n49562 , n28589 );
and ( n59604 , n26731 , n31075 );
or ( n59605 , n59603 , n59604 );
and ( n59606 , n59605 , n28594 );
and ( n59607 , n49572 , n28589 );
and ( n59608 , n26731 , n31075 );
or ( n59609 , n59607 , n59608 );
and ( n59610 , n59609 , n30269 );
and ( n59611 , n49582 , n28589 );
and ( n59612 , n26731 , n31075 );
or ( n59613 , n59611 , n59612 );
and ( n59614 , n59613 , n30982 );
and ( n59615 , n29159 , n28589 );
and ( n59616 , n26731 , n31075 );
or ( n59617 , n59615 , n59616 );
and ( n59618 , n59617 , n30989 );
and ( n59619 , n29159 , n30991 );
and ( n59620 , n49592 , n28589 );
and ( n59621 , n26731 , n31075 );
or ( n59622 , n59620 , n59621 );
and ( n59623 , n59622 , n31002 );
or ( n59624 , n59602 , n59606 , n59610 , n59614 , n59618 , n59619 , n59623 );
and ( n59625 , n59601 , n59624 );
and ( n59626 , n26731 , n24800 );
or ( n59627 , n59625 , n59626 );
and ( n59628 , n59627 , n31008 );
and ( n59629 , n25609 , n10618 );
or ( n59630 , n59628 , n59629 );
buf ( n59631 , n59630 );
buf ( n59632 , n59631 );
buf ( n59633 , n10613 );
buf ( n59634 , n10613 );
and ( n59635 , n16793 , n23924 );
and ( n59636 , n22133 , n23926 );
or ( n59637 , n59635 , n59636 );
buf ( n59638 , n59637 );
buf ( n59639 , n59638 );
not ( n59640 , n34821 );
and ( n59641 , n13299 , n14592 );
and ( n59642 , n43049 , n36350 );
and ( n59643 , n13299 , n43691 );
or ( n59644 , n59642 , n59643 );
and ( n59645 , n59644 , n14562 );
and ( n59646 , n43071 , n36350 );
and ( n59647 , n13299 , n43703 );
or ( n59648 , n59646 , n59647 );
and ( n59649 , n59648 , n14586 );
and ( n59650 , n43093 , n36345 );
and ( n59651 , n13299 , n43715 );
or ( n59652 , n59650 , n59651 );
and ( n59653 , n59652 , n14584 );
and ( n59654 , n43071 , n36345 );
and ( n59655 , n13299 , n43721 );
or ( n59656 , n59654 , n59655 );
and ( n59657 , n59656 , n37835 );
and ( n59658 , n43093 , n36345 );
and ( n59659 , n13299 , n43721 );
or ( n59660 , n59658 , n59659 );
and ( n59661 , n59660 , n37841 );
and ( n59662 , n15515 , n14564 );
and ( n59663 , n15515 , n36345 );
and ( n59664 , n13299 , n43721 );
or ( n59665 , n59663 , n59664 );
and ( n59666 , n59665 , n37847 );
or ( n59667 , n59641 , n59645 , n59649 , n59653 , n59657 , n59661 , n59662 , n59666 );
and ( n59668 , n59640 , n59667 );
and ( n59669 , n13299 , n34821 );
or ( n59670 , n59668 , n59669 );
and ( n59671 , n59670 , n16574 );
and ( n59672 , n12285 , n16576 );
or ( n59673 , n59671 , n59672 );
buf ( n59674 , n59673 );
buf ( n59675 , n59674 );
buf ( n59676 , n10615 );
buf ( n59677 , n10615 );
buf ( n59678 , n10613 );
buf ( n59679 , n10613 );
buf ( n59680 , n10613 );
buf ( n59681 , n10613 );
not ( n59682 , n24800 );
and ( n59683 , n25919 , n25222 );
and ( n59684 , n34569 , n28583 );
and ( n59685 , n25919 , n28591 );
or ( n59686 , n59684 , n59685 );
and ( n59687 , n59686 , n28594 );
and ( n59688 , n34582 , n28583 );
and ( n59689 , n25919 , n28591 );
or ( n59690 , n59688 , n59689 );
and ( n59691 , n59690 , n30269 );
and ( n59692 , n34592 , n28583 );
and ( n59693 , n25919 , n28591 );
or ( n59694 , n59692 , n59693 );
and ( n59695 , n59694 , n30982 );
and ( n59696 , n29635 , n28583 );
and ( n59697 , n25919 , n28591 );
or ( n59698 , n59696 , n59697 );
and ( n59699 , n59698 , n30989 );
and ( n59700 , n25917 , n30991 );
and ( n59701 , n34602 , n28583 );
and ( n59702 , n25919 , n28591 );
or ( n59703 , n59701 , n59702 );
and ( n59704 , n59703 , n31002 );
or ( n59705 , n59683 , n59687 , n59691 , n59695 , n59699 , n59700 , n59704 );
and ( n59706 , n59682 , n59705 );
and ( n59707 , n25919 , n24800 );
or ( n59708 , n59706 , n59707 );
and ( n59709 , n59708 , n31008 );
and ( n59710 , n25919 , n10618 );
or ( n59711 , n59709 , n59710 );
buf ( n59712 , n59711 );
buf ( n59713 , n59712 );
buf ( n59714 , n10613 );
buf ( n59715 , n10613 );
buf ( n59716 , n10615 );
buf ( n59717 , n10613 );
buf ( n59718 , n10613 );
buf ( n59719 , n10615 );
buf ( n59720 , n10613 );
buf ( n59721 , n10615 );
buf ( n59722 , n10613 );
not ( n59723 , n17451 );
and ( n59724 , n18703 , n17873 );
and ( n59725 , n40011 , n21336 );
and ( n59726 , n18703 , n42682 );
or ( n59727 , n59725 , n59726 );
and ( n59728 , n59727 , n21341 );
and ( n59729 , n40021 , n21336 );
and ( n59730 , n18703 , n42682 );
or ( n59731 , n59729 , n59730 );
and ( n59732 , n59731 , n23064 );
and ( n59733 , n40031 , n21336 );
and ( n59734 , n18703 , n42682 );
or ( n59735 , n59733 , n59734 );
and ( n59736 , n59735 , n23825 );
and ( n59737 , n22302 , n21336 );
and ( n59738 , n18703 , n42682 );
or ( n59739 , n59737 , n59738 );
and ( n59740 , n59739 , n23832 );
and ( n59741 , n22302 , n23834 );
and ( n59742 , n40041 , n21336 );
and ( n59743 , n18703 , n42682 );
or ( n59744 , n59742 , n59743 );
and ( n59745 , n59744 , n23917 );
or ( n59746 , n59724 , n59728 , n59732 , n59736 , n59740 , n59741 , n59745 );
and ( n59747 , n59723 , n59746 );
and ( n59748 , n18703 , n17451 );
or ( n59749 , n59747 , n59748 );
and ( n59750 , n59749 , n23924 );
and ( n59751 , n17960 , n23926 );
or ( n59752 , n59750 , n59751 );
buf ( n59753 , n59752 );
buf ( n59754 , n59753 );
and ( n59755 , n24341 , n31008 );
and ( n59756 , n29131 , n10618 );
or ( n59757 , n59755 , n59756 );
buf ( n59758 , n59757 );
buf ( n59759 , n59758 );
buf ( n59760 , n10615 );
and ( n59761 , n24198 , n31008 );
and ( n59762 , n29526 , n10618 );
or ( n59763 , n59761 , n59762 );
buf ( n59764 , n59763 );
buf ( n59765 , n59764 );
buf ( n59766 , n10613 );
not ( n59767 , n11333 );
and ( n59768 , n59767 , n10637 );
xor ( n59769 , n11351 , n11007 );
and ( n59770 , n59769 , n11333 );
or ( n59771 , n59768 , n59770 );
buf ( n59772 , n59771 );
buf ( n59773 , n59772 );
not ( n59774 , n34538 );
and ( n59775 , n59774 , n19356 );
and ( n59776 , n14681 , n34538 );
or ( n59777 , n59775 , n59776 );
and ( n59778 , n59777 , n23924 );
and ( n59779 , n14681 , n23926 );
or ( n59780 , n59778 , n59779 );
buf ( n59781 , n59780 );
buf ( n59782 , n59781 );
not ( n59783 , n34821 );
and ( n59784 , n13371 , n14592 );
and ( n59785 , n39404 , n36350 );
and ( n59786 , n13371 , n43691 );
or ( n59787 , n59785 , n59786 );
and ( n59788 , n59787 , n14562 );
and ( n59789 , n39423 , n36350 );
and ( n59790 , n13371 , n43703 );
or ( n59791 , n59789 , n59790 );
and ( n59792 , n59791 , n14586 );
and ( n59793 , n39442 , n36345 );
and ( n59794 , n13371 , n43715 );
or ( n59795 , n59793 , n59794 );
and ( n59796 , n59795 , n14584 );
and ( n59797 , n39423 , n36345 );
and ( n59798 , n13371 , n43721 );
or ( n59799 , n59797 , n59798 );
and ( n59800 , n59799 , n37835 );
and ( n59801 , n39442 , n36345 );
and ( n59802 , n13371 , n43721 );
or ( n59803 , n59801 , n59802 );
and ( n59804 , n59803 , n37841 );
and ( n59805 , n15647 , n14564 );
and ( n59806 , n15647 , n36345 );
and ( n59807 , n13371 , n43721 );
or ( n59808 , n59806 , n59807 );
and ( n59809 , n59808 , n37847 );
or ( n59810 , n59784 , n59788 , n59792 , n59796 , n59800 , n59804 , n59805 , n59809 );
and ( n59811 , n59783 , n59810 );
and ( n59812 , n13371 , n34821 );
or ( n59813 , n59811 , n59812 );
and ( n59814 , n59813 , n16574 );
and ( n59815 , n12303 , n16576 );
or ( n59816 , n59814 , n59815 );
buf ( n59817 , n59816 );
buf ( n59818 , n59817 );
not ( n59819 , n17451 );
and ( n59820 , n18314 , n17873 );
and ( n59821 , n34353 , n21336 );
and ( n59822 , n18314 , n42682 );
or ( n59823 , n59821 , n59822 );
and ( n59824 , n59823 , n21341 );
and ( n59825 , n34363 , n21336 );
and ( n59826 , n18314 , n42682 );
or ( n59827 , n59825 , n59826 );
and ( n59828 , n59827 , n23064 );
and ( n59829 , n34373 , n21336 );
and ( n59830 , n18314 , n42682 );
or ( n59831 , n59829 , n59830 );
and ( n59832 , n59831 , n23825 );
and ( n59833 , n21639 , n21336 );
and ( n59834 , n18314 , n42682 );
or ( n59835 , n59833 , n59834 );
and ( n59836 , n59835 , n23832 );
and ( n59837 , n21639 , n23834 );
and ( n59838 , n34383 , n21336 );
and ( n59839 , n18314 , n42682 );
or ( n59840 , n59838 , n59839 );
and ( n59841 , n59840 , n23917 );
or ( n59842 , n59820 , n59824 , n59828 , n59832 , n59836 , n59837 , n59841 );
and ( n59843 , n59819 , n59842 );
and ( n59844 , n18314 , n17451 );
or ( n59845 , n59843 , n59844 );
and ( n59846 , n59845 , n23924 );
and ( n59847 , n17875 , n23926 );
or ( n59848 , n59846 , n59847 );
buf ( n59849 , n59848 );
buf ( n59850 , n59849 );
buf ( n59851 , n10613 );
not ( n59852 , n24800 );
and ( n59853 , n50001 , n28587 );
and ( n59854 , n26159 , n39807 );
or ( n59855 , n59853 , n59854 );
and ( n59856 , n59855 , n28594 );
and ( n59857 , n50011 , n28587 );
and ( n59858 , n26159 , n39807 );
or ( n59859 , n59857 , n59858 );
and ( n59860 , n59859 , n30269 );
and ( n59861 , n50021 , n28587 );
and ( n59862 , n26159 , n39807 );
or ( n59863 , n59861 , n59862 );
and ( n59864 , n59863 , n30982 );
and ( n59865 , n29495 , n28587 );
and ( n59866 , n26159 , n39807 );
or ( n59867 , n59865 , n59866 );
and ( n59868 , n59867 , n30989 );
and ( n59869 , n50032 , n28587 );
and ( n59870 , n26159 , n39807 );
or ( n59871 , n59869 , n59870 );
and ( n59872 , n59871 , n31002 );
and ( n59873 , n26159 , n34607 );
or ( n59874 , n59856 , n59860 , n59864 , n59868 , n59872 , n59873 );
and ( n59875 , n59852 , n59874 );
and ( n59876 , n26159 , n24800 );
or ( n59877 , n59875 , n59876 );
and ( n59878 , n59877 , n31008 );
and ( n59879 , n26159 , n10618 );
or ( n59880 , n59878 , n59879 );
buf ( n59881 , n59880 );
buf ( n59882 , n59881 );
and ( n59883 , n11617 , n16574 );
and ( n59884 , n15638 , n16576 );
or ( n59885 , n59883 , n59884 );
buf ( n59886 , n59885 );
buf ( n59887 , n59886 );
buf ( n59888 , n10613 );
not ( n59889 , n34821 );
and ( n59890 , n59889 , n36311 );
and ( n59891 , n36286 , n34821 );
or ( n59892 , n59890 , n59891 );
and ( n59893 , n59892 , n16574 );
and ( n59894 , n36286 , n16576 );
or ( n59895 , n59893 , n59894 );
buf ( n59896 , n59895 );
buf ( n59897 , n59896 );
buf ( n59898 , n10613 );
buf ( n59899 , n10613 );
buf ( n59900 , n10613 );
buf ( n59901 , n10615 );
not ( n59902 , n17162 );
not ( n59903 , n17450 );
and ( n59904 , n10668 , n37947 );
not ( n59905 , n38425 );
and ( n59906 , n59905 , n38319 );
xor ( n59907 , n46213 , n46214 );
and ( n59908 , n59907 , n38425 );
or ( n59909 , n59906 , n59908 );
buf ( n59910 , n59909 );
and ( n59911 , n59910 , n19745 );
not ( n59912 , n38934 );
and ( n59913 , n59912 , n38828 );
xor ( n59914 , n46226 , n46227 );
and ( n59915 , n59914 , n38934 );
or ( n59916 , n59913 , n59915 );
buf ( n59917 , n59916 );
and ( n59918 , n59917 , n19748 );
and ( n59919 , n22160 , n21253 );
and ( n59920 , n10668 , n21255 );
or ( n59921 , n59911 , n59918 , n59919 , n59920 );
and ( n59922 , n59921 , n38980 );
or ( n59923 , n59904 , n59922 );
and ( n59924 , n59903 , n59923 );
or ( n59925 , n59924 , C0 );
and ( n59926 , n59902 , n59925 );
and ( n59927 , n59921 , n17162 );
or ( n59928 , n59926 , n59927 );
and ( n59929 , n59928 , n23924 );
not ( n59930 , n39264 );
and ( n59931 , n59930 , n39176 );
xor ( n59932 , n46250 , n46251 );
and ( n59933 , n59932 , n39264 );
or ( n59934 , n59931 , n59933 );
buf ( n59935 , n59934 );
and ( n59936 , n59935 , n23926 );
or ( n59937 , n59929 , n59936 );
buf ( n59938 , n59937 );
buf ( n59939 , n59938 );
buf ( n59940 , n10613 );
buf ( n59941 , n10613 );
not ( n59942 , n24800 );
and ( n59943 , n34656 , n28587 );
and ( n59944 , n26329 , n39807 );
or ( n59945 , n59943 , n59944 );
and ( n59946 , n59945 , n28594 );
and ( n59947 , n34674 , n28587 );
and ( n59948 , n26329 , n39807 );
or ( n59949 , n59947 , n59948 );
and ( n59950 , n59949 , n30269 );
and ( n59951 , n34692 , n28587 );
and ( n59952 , n26329 , n39807 );
or ( n59953 , n59951 , n59952 );
and ( n59954 , n59953 , n30982 );
and ( n59955 , n29395 , n28587 );
and ( n59956 , n26329 , n39807 );
or ( n59957 , n59955 , n59956 );
and ( n59958 , n59957 , n30989 );
and ( n59959 , n34714 , n28587 );
and ( n59960 , n26329 , n39807 );
or ( n59961 , n59959 , n59960 );
and ( n59962 , n59961 , n31002 );
and ( n59963 , n26329 , n34607 );
or ( n59964 , n59946 , n59950 , n59954 , n59958 , n59962 , n59963 );
and ( n59965 , n59942 , n59964 );
and ( n59966 , n26329 , n24800 );
or ( n59967 , n59965 , n59966 );
and ( n59968 , n59967 , n31008 );
and ( n59969 , n26329 , n10618 );
or ( n59970 , n59968 , n59969 );
buf ( n59971 , n59970 );
buf ( n59972 , n59971 );
buf ( n59973 , n10613 );
buf ( n59974 , n10615 );
not ( n59975 , n34804 );
and ( n59976 , n59975 , n26297 );
and ( n59977 , n14755 , n34804 );
or ( n59978 , n59976 , n59977 );
and ( n59979 , n59978 , n31008 );
and ( n59980 , n14755 , n10618 );
or ( n59981 , n59979 , n59980 );
buf ( n59982 , n59981 );
buf ( n59983 , n59982 );
and ( n59984 , n11512 , n16574 );
and ( n59985 , n15065 , n16576 );
or ( n59986 , n59984 , n59985 );
buf ( n59987 , n59986 );
buf ( n59988 , n59987 );
buf ( n59989 , n10615 );
buf ( n59990 , n10615 );
not ( n59991 , n11954 );
not ( n59992 , n12243 );
and ( n59993 , n10877 , n31187 );
not ( n59994 , n31697 );
and ( n59995 , n59994 , n31523 );
xor ( n59996 , n50357 , n50374 );
and ( n59997 , n59996 , n31697 );
or ( n59998 , n59995 , n59997 );
buf ( n59999 , n59998 );
and ( n60000 , n59999 , n14140 );
not ( n60001 , n32214 );
and ( n60002 , n60001 , n32040 );
xor ( n60003 , n50384 , n50401 );
and ( n60004 , n60003 , n32214 );
or ( n60005 , n60002 , n60004 );
buf ( n60006 , n60005 );
and ( n60007 , n60006 , n14137 );
and ( n60008 , n15667 , n14143 );
and ( n60009 , n10877 , n14141 );
or ( n60010 , n60000 , n60007 , n60008 , n60009 );
and ( n60011 , n60010 , n32236 );
or ( n60012 , n59993 , n60011 );
and ( n60013 , n59992 , n60012 );
not ( n60014 , n34038 );
and ( n60015 , n60014 , n33794 );
xor ( n60016 , n50417 , n50434 );
and ( n60017 , n60016 , n34038 );
or ( n60018 , n60015 , n60017 );
buf ( n60019 , n60018 );
and ( n60020 , n60019 , n12243 );
or ( n60021 , n60013 , n60020 );
and ( n60022 , n59991 , n60021 );
and ( n60023 , n60010 , n11954 );
or ( n60024 , n60022 , n60023 );
and ( n60025 , n60024 , n16574 );
not ( n60026 , n34327 );
and ( n60027 , n60026 , n34183 );
xor ( n60028 , n50449 , n50466 );
and ( n60029 , n60028 , n34327 );
or ( n60030 , n60027 , n60029 );
buf ( n60031 , n60030 );
and ( n60032 , n60031 , n16576 );
or ( n60033 , n60025 , n60032 );
buf ( n60034 , n60033 );
buf ( n60035 , n60034 );
buf ( n60036 , n10613 );
not ( n60037 , n34821 );
and ( n60038 , n43617 , n36345 );
and ( n60039 , n13341 , n36352 );
or ( n60040 , n60038 , n60039 );
and ( n60041 , n60040 , n14562 );
and ( n60042 , n43627 , n36345 );
and ( n60043 , n13341 , n37073 );
or ( n60044 , n60042 , n60043 );
and ( n60045 , n60044 , n14586 );
and ( n60046 , n43637 , n36350 );
and ( n60047 , n13341 , n37825 );
or ( n60048 , n60046 , n60047 );
and ( n60049 , n60048 , n14584 );
and ( n60050 , n43627 , n36350 );
and ( n60051 , n13341 , n37831 );
or ( n60052 , n60050 , n60051 );
and ( n60053 , n60052 , n37835 );
and ( n60054 , n43637 , n36350 );
and ( n60055 , n13341 , n37831 );
or ( n60056 , n60054 , n60055 );
and ( n60057 , n60056 , n37841 );
and ( n60058 , n15581 , n36350 );
and ( n60059 , n13341 , n37831 );
or ( n60060 , n60058 , n60059 );
and ( n60061 , n60060 , n37847 );
and ( n60062 , n13341 , n37849 );
or ( n60063 , n60041 , n60045 , n60049 , n60053 , n60057 , n60061 , n60062 );
and ( n60064 , n60037 , n60063 );
and ( n60065 , n13341 , n34821 );
or ( n60066 , n60064 , n60065 );
and ( n60067 , n60066 , n16574 );
and ( n60068 , n13341 , n16576 );
or ( n60069 , n60067 , n60068 );
buf ( n60070 , n60069 );
buf ( n60071 , n60070 );
not ( n60072 , n34821 );
and ( n60073 , n43688 , n36345 );
and ( n60074 , n13353 , n36352 );
or ( n60075 , n60073 , n60074 );
and ( n60076 , n60075 , n14562 );
and ( n60077 , n43700 , n36345 );
and ( n60078 , n13353 , n37073 );
or ( n60079 , n60077 , n60078 );
and ( n60080 , n60079 , n14586 );
and ( n60081 , n43712 , n36350 );
and ( n60082 , n13353 , n37825 );
or ( n60083 , n60081 , n60082 );
and ( n60084 , n60083 , n14584 );
and ( n60085 , n43700 , n36350 );
and ( n60086 , n13353 , n37831 );
or ( n60087 , n60085 , n60086 );
and ( n60088 , n60087 , n37835 );
and ( n60089 , n43712 , n36350 );
and ( n60090 , n13353 , n37831 );
or ( n60091 , n60089 , n60090 );
and ( n60092 , n60091 , n37841 );
and ( n60093 , n15603 , n36350 );
and ( n60094 , n13353 , n37831 );
or ( n60095 , n60093 , n60094 );
and ( n60096 , n60095 , n37847 );
and ( n60097 , n13353 , n37849 );
or ( n60098 , n60076 , n60080 , n60084 , n60088 , n60092 , n60096 , n60097 );
and ( n60099 , n60072 , n60098 );
and ( n60100 , n13353 , n34821 );
or ( n60101 , n60099 , n60100 );
and ( n60102 , n60101 , n16574 );
and ( n60103 , n13353 , n16576 );
or ( n60104 , n60102 , n60103 );
buf ( n60105 , n60104 );
buf ( n60106 , n60105 );
not ( n60107 , n17162 );
not ( n60108 , n17450 );
and ( n60109 , n10653 , n37947 );
not ( n60110 , n38425 );
and ( n60111 , n60110 , n38370 );
xor ( n60112 , n51306 , n51307 );
and ( n60113 , n60112 , n38425 );
or ( n60114 , n60111 , n60113 );
buf ( n60115 , n60114 );
and ( n60116 , n60115 , n19745 );
not ( n60117 , n38934 );
and ( n60118 , n60117 , n38879 );
xor ( n60119 , n51317 , n51318 );
and ( n60120 , n60119 , n38934 );
or ( n60121 , n60118 , n60120 );
buf ( n60122 , n60121 );
and ( n60123 , n60122 , n19748 );
and ( n60124 , n22100 , n21253 );
and ( n60125 , n10653 , n21255 );
or ( n60126 , n60116 , n60123 , n60124 , n60125 );
and ( n60127 , n60126 , n38980 );
or ( n60128 , n60109 , n60127 );
and ( n60129 , n60108 , n60128 );
or ( n60130 , n60129 , C0 );
and ( n60131 , n60107 , n60130 );
and ( n60132 , n60126 , n17162 );
or ( n60133 , n60131 , n60132 );
and ( n60134 , n60133 , n23924 );
not ( n60135 , n39264 );
and ( n60136 , n60135 , n39218 );
xor ( n60137 , n51339 , n51340 );
and ( n60138 , n60137 , n39264 );
or ( n60139 , n60136 , n60138 );
buf ( n60140 , n60139 );
and ( n60141 , n60140 , n23926 );
or ( n60142 , n60134 , n60141 );
buf ( n60143 , n60142 );
buf ( n60144 , n60143 );
buf ( n60145 , n10615 );
buf ( n60146 , n10615 );
buf ( n60147 , n10613 );
buf ( n60148 , n10615 );
buf ( n60149 , n10615 );
buf ( n60150 , n10615 );
buf ( n60151 , n10615 );
and ( n60152 , n11537 , n16574 );
and ( n60153 , n15110 , n16576 );
or ( n60154 , n60152 , n60153 );
buf ( n60155 , n60154 );
buf ( n60156 , n60155 );
buf ( n60157 , n10615 );
buf ( n60158 , n10615 );
not ( n60159 , n24800 );
and ( n60160 , n52160 , n28586 );
and ( n60161 , n26769 , n34573 );
or ( n60162 , n60160 , n60161 );
and ( n60163 , n60162 , n28594 );
and ( n60164 , n52170 , n28586 );
and ( n60165 , n26769 , n34573 );
or ( n60166 , n60164 , n60165 );
and ( n60167 , n60166 , n30269 );
and ( n60168 , n52180 , n28586 );
and ( n60169 , n26769 , n34573 );
or ( n60170 , n60168 , n60169 );
and ( n60171 , n60170 , n30982 );
and ( n60172 , n29146 , n28586 );
and ( n60173 , n26769 , n34573 );
or ( n60174 , n60172 , n60173 );
and ( n60175 , n60174 , n30989 );
and ( n60176 , n52191 , n28586 );
and ( n60177 , n26769 , n34573 );
or ( n60178 , n60176 , n60177 );
and ( n60179 , n60178 , n31002 );
and ( n60180 , n26769 , n34607 );
or ( n60181 , n60163 , n60167 , n60171 , n60175 , n60179 , n60180 );
and ( n60182 , n60159 , n60181 );
and ( n60183 , n26769 , n24800 );
or ( n60184 , n60182 , n60183 );
and ( n60185 , n60184 , n31008 );
and ( n60186 , n26769 , n10618 );
or ( n60187 , n60185 , n60186 );
buf ( n60188 , n60187 );
buf ( n60189 , n60188 );
buf ( n60190 , n10613 );
buf ( n60191 , n10615 );
buf ( n60192 , n10613 );
buf ( n60193 , n10613 );
buf ( n60194 , n10613 );
buf ( n60195 , n10615 );
buf ( n60196 , n10615 );
buf ( n60197 , n10615 );
not ( n60198 , n17451 );
and ( n60199 , n51973 , n21333 );
and ( n60200 , n18741 , n34758 );
or ( n60201 , n60199 , n60200 );
and ( n60202 , n60201 , n21341 );
and ( n60203 , n51983 , n21333 );
and ( n60204 , n18741 , n34758 );
or ( n60205 , n60203 , n60204 );
and ( n60206 , n60205 , n23064 );
and ( n60207 , n51993 , n21333 );
and ( n60208 , n18741 , n34758 );
or ( n60209 , n60207 , n60208 );
and ( n60210 , n60209 , n23825 );
and ( n60211 , n22282 , n21333 );
and ( n60212 , n18741 , n34758 );
or ( n60213 , n60211 , n60212 );
and ( n60214 , n60213 , n23832 );
and ( n60215 , n52004 , n21333 );
and ( n60216 , n18741 , n34758 );
or ( n60217 , n60215 , n60216 );
and ( n60218 , n60217 , n23917 );
and ( n60219 , n18741 , n34526 );
or ( n60220 , n60202 , n60206 , n60210 , n60214 , n60218 , n60219 );
and ( n60221 , n60198 , n60220 );
and ( n60222 , n18741 , n17451 );
or ( n60223 , n60221 , n60222 );
and ( n60224 , n60223 , n23924 );
and ( n60225 , n18741 , n23926 );
or ( n60226 , n60224 , n60225 );
buf ( n60227 , n60226 );
buf ( n60228 , n60227 );
buf ( n60229 , n10615 );
buf ( n60230 , n10615 );
not ( n60231 , n11954 );
not ( n60232 , n12243 );
and ( n60233 , n10925 , n31187 );
not ( n60234 , n31697 );
and ( n60235 , n60234 , n31421 );
xor ( n60236 , n50363 , n50368 );
and ( n60237 , n60236 , n31697 );
or ( n60238 , n60235 , n60237 );
buf ( n60239 , n60238 );
and ( n60240 , n60239 , n14140 );
not ( n60241 , n32214 );
and ( n60242 , n60241 , n31938 );
xor ( n60243 , n50390 , n50395 );
and ( n60244 , n60243 , n32214 );
or ( n60245 , n60242 , n60244 );
buf ( n60246 , n60245 );
and ( n60247 , n60246 , n14137 );
and ( n60248 , n15799 , n14143 );
and ( n60249 , n10925 , n14141 );
or ( n60250 , n60240 , n60247 , n60248 , n60249 );
and ( n60251 , n60250 , n32236 );
or ( n60252 , n60233 , n60251 );
and ( n60253 , n60232 , n60252 );
not ( n60254 , n34038 );
and ( n60255 , n60254 , n33650 );
xor ( n60256 , n50423 , n50428 );
and ( n60257 , n60256 , n34038 );
or ( n60258 , n60255 , n60257 );
buf ( n60259 , n60258 );
and ( n60260 , n60259 , n12243 );
or ( n60261 , n60253 , n60260 );
and ( n60262 , n60231 , n60261 );
and ( n60263 , n60250 , n11954 );
or ( n60264 , n60262 , n60263 );
and ( n60265 , n60264 , n16574 );
not ( n60266 , n34327 );
and ( n60267 , n60266 , n34099 );
xor ( n60268 , n50455 , n50460 );
and ( n60269 , n60268 , n34327 );
or ( n60270 , n60267 , n60269 );
buf ( n60271 , n60270 );
and ( n60272 , n60271 , n16576 );
or ( n60273 , n60265 , n60272 );
buf ( n60274 , n60273 );
buf ( n60275 , n60274 );
buf ( n60276 , n10615 );
not ( n60277 , n17451 );
and ( n60278 , n19147 , n17873 );
and ( n60279 , n46760 , n21330 );
and ( n60280 , n19147 , n21338 );
or ( n60281 , n60279 , n60280 );
and ( n60282 , n60281 , n21341 );
and ( n60283 , n46770 , n21330 );
and ( n60284 , n19147 , n21338 );
or ( n60285 , n60283 , n60284 );
and ( n60286 , n60285 , n23064 );
and ( n60287 , n46780 , n21330 );
and ( n60288 , n19147 , n21338 );
or ( n60289 , n60287 , n60288 );
and ( n60290 , n60289 , n23825 );
and ( n60291 , n22042 , n21330 );
and ( n60292 , n19147 , n21338 );
or ( n60293 , n60291 , n60292 );
and ( n60294 , n60293 , n23832 );
and ( n60295 , n19145 , n23834 );
and ( n60296 , n46791 , n21330 );
and ( n60297 , n19147 , n21338 );
or ( n60298 , n60296 , n60297 );
and ( n60299 , n60298 , n23917 );
or ( n60300 , n60278 , n60282 , n60286 , n60290 , n60294 , n60295 , n60299 );
and ( n60301 , n60277 , n60300 );
and ( n60302 , n19147 , n17451 );
or ( n60303 , n60301 , n60302 );
and ( n60304 , n60303 , n23924 );
and ( n60305 , n19147 , n23926 );
or ( n60306 , n60304 , n60305 );
buf ( n60307 , n60306 );
buf ( n60308 , n60307 );
not ( n60309 , n24511 );
not ( n60310 , n24799 );
buf ( n60311 , n56380 );
and ( n60312 , n60311 , n27046 );
or ( n60313 , n28506 , n28508 );
or ( n60314 , n60313 , n27049 );
and ( n60315 , n27051 , n60314 );
or ( n60316 , n60312 , n60315 );
and ( n60317 , n60316 , n28594 );
or ( n60318 , n30991 , n31002 );
or ( n60319 , n60318 , n30987 );
or ( n60320 , n60319 , n30988 );
or ( n60321 , n60320 , n30976 );
or ( n60322 , n60321 , n30977 );
or ( n60323 , n60322 , n30263 );
or ( n60324 , n60323 , n30264 );
or ( n60325 , n60324 , n30979 );
or ( n60326 , n60325 , n30266 );
or ( n60327 , n60326 , n30981 );
or ( n60328 , n60327 , n30268 );
or ( n60329 , n60328 , n25222 );
and ( n60330 , n27051 , n60329 );
or ( n60331 , n60317 , n60330 );
and ( n60332 , n60310 , n60331 );
and ( n60333 , n27051 , n24799 );
or ( n60334 , n60332 , n60333 );
and ( n60335 , n60309 , n60334 );
buf ( n60336 , n25876 );
not ( n60337 , n60336 );
buf ( n60338 , n27181 );
and ( n60339 , n60337 , n60338 );
buf ( n60340 , n60339 );
not ( n60341 , n60340 );
and ( n60342 , n60341 , n25876 );
or ( n60343 , n60342 , C0 );
buf ( n60344 , n60343 );
buf ( n60345 , n29094 );
xor ( n60346 , n60344 , n60345 );
not ( n60347 , n60346 );
not ( n60348 , n60340 );
and ( n60349 , n60348 , n27181 );
or ( n60350 , n60349 , C0 );
buf ( n60351 , n60350 );
not ( n60352 , n60351 );
buf ( n60353 , n29107 );
and ( n60354 , n60352 , n60353 );
buf ( n60355 , n27193 );
buf ( n60356 , n60355 );
not ( n60357 , n60356 );
buf ( n60358 , n29120 );
and ( n60359 , n60357 , n60358 );
buf ( n60360 , n26807 );
buf ( n60361 , n60360 );
not ( n60362 , n60361 );
buf ( n60363 , n29133 );
and ( n60364 , n60362 , n60363 );
buf ( n60365 , n26773 );
buf ( n60366 , n60365 );
not ( n60367 , n60366 );
buf ( n60368 , n29146 );
and ( n60369 , n60367 , n60368 );
buf ( n60370 , n26739 );
buf ( n60371 , n60370 );
not ( n60372 , n60371 );
buf ( n60373 , n29159 );
and ( n60374 , n60372 , n60373 );
buf ( n60375 , n26705 );
buf ( n60376 , n60375 );
not ( n60377 , n60376 );
buf ( n60378 , n29172 );
and ( n60379 , n60377 , n60378 );
buf ( n60380 , n26671 );
buf ( n60381 , n60380 );
not ( n60382 , n60381 );
buf ( n60383 , n29185 );
and ( n60384 , n60382 , n60383 );
buf ( n60385 , n26637 );
buf ( n60386 , n60385 );
not ( n60387 , n60386 );
buf ( n60388 , n29198 );
and ( n60389 , n60387 , n60388 );
buf ( n60390 , n26603 );
buf ( n60391 , n60390 );
not ( n60392 , n60391 );
buf ( n60393 , n29211 );
and ( n60394 , n60392 , n60393 );
buf ( n60395 , n26569 );
buf ( n60396 , n60395 );
not ( n60397 , n60396 );
buf ( n60398 , n29224 );
and ( n60399 , n60397 , n60398 );
buf ( n60400 , n26535 );
buf ( n60401 , n60400 );
not ( n60402 , n60401 );
buf ( n60403 , n29237 );
and ( n60404 , n60402 , n60403 );
buf ( n60405 , n26501 );
buf ( n60406 , n60405 );
not ( n60407 , n60406 );
buf ( n60408 , n29295 );
and ( n60409 , n60407 , n60408 );
buf ( n60410 , n26467 );
buf ( n60411 , n60410 );
not ( n60412 , n60411 );
buf ( n60413 , n29315 );
and ( n60414 , n60412 , n60413 );
buf ( n60415 , n26433 );
buf ( n60416 , n60415 );
not ( n60417 , n60416 );
buf ( n60418 , n29335 );
and ( n60419 , n60417 , n60418 );
buf ( n60420 , n26399 );
buf ( n60421 , n60420 );
not ( n60422 , n60421 );
buf ( n60423 , n29355 );
and ( n60424 , n60422 , n60423 );
buf ( n60425 , n26365 );
buf ( n60426 , n60425 );
not ( n60427 , n60426 );
buf ( n60428 , n29375 );
and ( n60429 , n60427 , n60428 );
buf ( n60430 , n26331 );
buf ( n60431 , n60430 );
not ( n60432 , n60431 );
buf ( n60433 , n29395 );
and ( n60434 , n60432 , n60433 );
buf ( n60435 , n26297 );
buf ( n60436 , n60435 );
not ( n60437 , n60436 );
buf ( n60438 , n29415 );
and ( n60439 , n60437 , n60438 );
buf ( n60440 , n26263 );
buf ( n60441 , n60440 );
not ( n60442 , n60441 );
buf ( n60443 , n29435 );
and ( n60444 , n60442 , n60443 );
buf ( n60445 , n26229 );
buf ( n60446 , n60445 );
not ( n60447 , n60446 );
buf ( n60448 , n29455 );
and ( n60449 , n60447 , n60448 );
buf ( n60450 , n26195 );
buf ( n60451 , n60450 );
not ( n60452 , n60451 );
buf ( n60453 , n29475 );
and ( n60454 , n60452 , n60453 );
buf ( n60455 , n26161 );
buf ( n60456 , n60455 );
not ( n60457 , n60456 );
buf ( n60458 , n29495 );
and ( n60459 , n60457 , n60458 );
buf ( n60460 , n26127 );
buf ( n60461 , n60460 );
not ( n60462 , n60461 );
buf ( n60463 , n29515 );
and ( n60464 , n60462 , n60463 );
buf ( n60465 , n26093 );
buf ( n60466 , n60465 );
not ( n60467 , n60466 );
buf ( n60468 , n29535 );
and ( n60469 , n60467 , n60468 );
buf ( n60470 , n26059 );
buf ( n60471 , n60470 );
not ( n60472 , n60471 );
buf ( n60473 , n29555 );
and ( n60474 , n60472 , n60473 );
buf ( n60475 , n26025 );
buf ( n60476 , n60475 );
not ( n60477 , n60476 );
buf ( n60478 , n29575 );
and ( n60479 , n60477 , n60478 );
buf ( n60480 , n25991 );
buf ( n60481 , n60480 );
not ( n60482 , n60481 );
buf ( n60483 , n29595 );
and ( n60484 , n60482 , n60483 );
buf ( n60485 , n25958 );
buf ( n60486 , n60485 );
not ( n60487 , n60486 );
buf ( n60488 , n29615 );
and ( n60489 , n60487 , n60488 );
buf ( n60490 , n25925 );
buf ( n60491 , n60490 );
not ( n60492 , n60491 );
buf ( n60493 , n29635 );
and ( n60494 , n60492 , n60493 );
buf ( n60495 , n25894 );
buf ( n60496 , n60495 );
not ( n60497 , n60496 );
buf ( n60498 , n29655 );
and ( n60499 , n60497 , n60498 );
buf ( n60500 , n25863 );
buf ( n60501 , n60500 );
not ( n60502 , n60501 );
buf ( n60503 , n28892 );
and ( n60504 , n60502 , n60503 );
xnor ( n60505 , n60496 , n60498 );
and ( n60506 , n60504 , n60505 );
or ( n60507 , n60499 , n60506 );
xnor ( n60508 , n60491 , n60493 );
and ( n60509 , n60507 , n60508 );
or ( n60510 , n60494 , n60509 );
xnor ( n60511 , n60486 , n60488 );
and ( n60512 , n60510 , n60511 );
or ( n60513 , n60489 , n60512 );
xnor ( n60514 , n60481 , n60483 );
and ( n60515 , n60513 , n60514 );
or ( n60516 , n60484 , n60515 );
xnor ( n60517 , n60476 , n60478 );
and ( n60518 , n60516 , n60517 );
or ( n60519 , n60479 , n60518 );
xnor ( n60520 , n60471 , n60473 );
and ( n60521 , n60519 , n60520 );
or ( n60522 , n60474 , n60521 );
xnor ( n60523 , n60466 , n60468 );
and ( n60524 , n60522 , n60523 );
or ( n60525 , n60469 , n60524 );
xnor ( n60526 , n60461 , n60463 );
and ( n60527 , n60525 , n60526 );
or ( n60528 , n60464 , n60527 );
xnor ( n60529 , n60456 , n60458 );
and ( n60530 , n60528 , n60529 );
or ( n60531 , n60459 , n60530 );
xnor ( n60532 , n60451 , n60453 );
and ( n60533 , n60531 , n60532 );
or ( n60534 , n60454 , n60533 );
xnor ( n60535 , n60446 , n60448 );
and ( n60536 , n60534 , n60535 );
or ( n60537 , n60449 , n60536 );
xnor ( n60538 , n60441 , n60443 );
and ( n60539 , n60537 , n60538 );
or ( n60540 , n60444 , n60539 );
xnor ( n60541 , n60436 , n60438 );
and ( n60542 , n60540 , n60541 );
or ( n60543 , n60439 , n60542 );
xnor ( n60544 , n60431 , n60433 );
and ( n60545 , n60543 , n60544 );
or ( n60546 , n60434 , n60545 );
xnor ( n60547 , n60426 , n60428 );
and ( n60548 , n60546 , n60547 );
or ( n60549 , n60429 , n60548 );
xnor ( n60550 , n60421 , n60423 );
and ( n60551 , n60549 , n60550 );
or ( n60552 , n60424 , n60551 );
xnor ( n60553 , n60416 , n60418 );
and ( n60554 , n60552 , n60553 );
or ( n60555 , n60419 , n60554 );
xnor ( n60556 , n60411 , n60413 );
and ( n60557 , n60555 , n60556 );
or ( n60558 , n60414 , n60557 );
xnor ( n60559 , n60406 , n60408 );
and ( n60560 , n60558 , n60559 );
or ( n60561 , n60409 , n60560 );
xnor ( n60562 , n60401 , n60403 );
and ( n60563 , n60561 , n60562 );
or ( n60564 , n60404 , n60563 );
xnor ( n60565 , n60396 , n60398 );
and ( n60566 , n60564 , n60565 );
or ( n60567 , n60399 , n60566 );
xnor ( n60568 , n60391 , n60393 );
and ( n60569 , n60567 , n60568 );
or ( n60570 , n60394 , n60569 );
xnor ( n60571 , n60386 , n60388 );
and ( n60572 , n60570 , n60571 );
or ( n60573 , n60389 , n60572 );
xnor ( n60574 , n60381 , n60383 );
and ( n60575 , n60573 , n60574 );
or ( n60576 , n60384 , n60575 );
xnor ( n60577 , n60376 , n60378 );
and ( n60578 , n60576 , n60577 );
or ( n60579 , n60379 , n60578 );
xnor ( n60580 , n60371 , n60373 );
and ( n60581 , n60579 , n60580 );
or ( n60582 , n60374 , n60581 );
xnor ( n60583 , n60366 , n60368 );
and ( n60584 , n60582 , n60583 );
or ( n60585 , n60369 , n60584 );
xnor ( n60586 , n60361 , n60363 );
and ( n60587 , n60585 , n60586 );
or ( n60588 , n60364 , n60587 );
xnor ( n60589 , n60356 , n60358 );
and ( n60590 , n60588 , n60589 );
or ( n60591 , n60359 , n60590 );
xnor ( n60592 , n60351 , n60353 );
and ( n60593 , n60591 , n60592 );
or ( n60594 , n60354 , n60593 );
and ( n60595 , n60347 , n60594 );
not ( n60596 , n60345 );
and ( n60597 , n60596 , n60344 );
and ( n60598 , n60597 , n60346 );
or ( n60599 , n60595 , n60598 );
buf ( n60600 , n60599 );
not ( n60601 , n60600 );
or ( n60602 , n60601 , n27051 );
and ( n60603 , n60602 , n25221 );
or ( n60604 , n60600 , n27051 );
and ( n60605 , n60604 , n25219 );
buf ( n60606 , n25876 );
buf ( n60607 , n29094 );
xor ( n60608 , n60606 , n60607 );
not ( n60609 , n60608 );
buf ( n60610 , n29107 );
not ( n60611 , n60610 );
buf ( n60612 , n27181 );
and ( n60613 , n60611 , n60612 );
buf ( n60614 , n29120 );
not ( n60615 , n60614 );
buf ( n60616 , n27193 );
and ( n60617 , n60615 , n60616 );
buf ( n60618 , n29133 );
not ( n60619 , n60618 );
buf ( n60620 , n26807 );
and ( n60621 , n60619 , n60620 );
buf ( n60622 , n29146 );
not ( n60623 , n60622 );
buf ( n60624 , n26773 );
and ( n60625 , n60623 , n60624 );
buf ( n60626 , n29159 );
not ( n60627 , n60626 );
buf ( n60628 , n26739 );
and ( n60629 , n60627 , n60628 );
buf ( n60630 , n29172 );
not ( n60631 , n60630 );
buf ( n60632 , n26705 );
and ( n60633 , n60631 , n60632 );
buf ( n60634 , n29185 );
not ( n60635 , n60634 );
buf ( n60636 , n26671 );
and ( n60637 , n60635 , n60636 );
buf ( n60638 , n29198 );
not ( n60639 , n60638 );
buf ( n60640 , n26637 );
and ( n60641 , n60639 , n60640 );
buf ( n60642 , n29211 );
not ( n60643 , n60642 );
buf ( n60644 , n26603 );
and ( n60645 , n60643 , n60644 );
buf ( n60646 , n29224 );
not ( n60647 , n60646 );
buf ( n60648 , n26569 );
and ( n60649 , n60647 , n60648 );
buf ( n60650 , n29237 );
not ( n60651 , n60650 );
buf ( n60652 , n26535 );
and ( n60653 , n60651 , n60652 );
buf ( n60654 , n29295 );
not ( n60655 , n60654 );
buf ( n60656 , n26501 );
and ( n60657 , n60655 , n60656 );
buf ( n60658 , n29315 );
not ( n60659 , n60658 );
buf ( n60660 , n26467 );
and ( n60661 , n60659 , n60660 );
buf ( n60662 , n29335 );
not ( n60663 , n60662 );
buf ( n60664 , n26433 );
and ( n60665 , n60663 , n60664 );
buf ( n60666 , n29355 );
not ( n60667 , n60666 );
buf ( n60668 , n26399 );
and ( n60669 , n60667 , n60668 );
buf ( n60670 , n29375 );
not ( n60671 , n60670 );
buf ( n60672 , n26365 );
and ( n60673 , n60671 , n60672 );
buf ( n60674 , n29395 );
not ( n60675 , n60674 );
buf ( n60676 , n26331 );
and ( n60677 , n60675 , n60676 );
buf ( n60678 , n29415 );
not ( n60679 , n60678 );
buf ( n60680 , n26297 );
and ( n60681 , n60679 , n60680 );
buf ( n60682 , n29435 );
not ( n60683 , n60682 );
buf ( n60684 , n26263 );
and ( n60685 , n60683 , n60684 );
buf ( n60686 , n29455 );
not ( n60687 , n60686 );
buf ( n60688 , n26229 );
and ( n60689 , n60687 , n60688 );
buf ( n60690 , n29475 );
not ( n60691 , n60690 );
buf ( n60692 , n26195 );
and ( n60693 , n60691 , n60692 );
buf ( n60694 , n29495 );
not ( n60695 , n60694 );
buf ( n60696 , n26161 );
and ( n60697 , n60695 , n60696 );
buf ( n60698 , n29515 );
not ( n60699 , n60698 );
buf ( n60700 , n26127 );
and ( n60701 , n60699 , n60700 );
buf ( n60702 , n29535 );
not ( n60703 , n60702 );
buf ( n60704 , n26093 );
and ( n60705 , n60703 , n60704 );
buf ( n60706 , n29555 );
not ( n60707 , n60706 );
buf ( n60708 , n26059 );
and ( n60709 , n60707 , n60708 );
buf ( n60710 , n29575 );
not ( n60711 , n60710 );
buf ( n60712 , n26025 );
and ( n60713 , n60711 , n60712 );
buf ( n60714 , n29595 );
not ( n60715 , n60714 );
buf ( n60716 , n25991 );
and ( n60717 , n60715 , n60716 );
buf ( n60718 , n29615 );
not ( n60719 , n60718 );
buf ( n60720 , n25958 );
and ( n60721 , n60719 , n60720 );
buf ( n60722 , n29635 );
not ( n60723 , n60722 );
buf ( n60724 , n25925 );
and ( n60725 , n60723 , n60724 );
buf ( n60726 , n29655 );
not ( n60727 , n60726 );
buf ( n60728 , n25894 );
and ( n60729 , n60727 , n60728 );
buf ( n60730 , n28892 );
not ( n60731 , n60730 );
buf ( n60732 , n25863 );
and ( n60733 , n60731 , n60732 );
xnor ( n60734 , n60728 , n60726 );
and ( n60735 , n60733 , n60734 );
or ( n60736 , n60729 , n60735 );
xnor ( n60737 , n60724 , n60722 );
and ( n60738 , n60736 , n60737 );
or ( n60739 , n60725 , n60738 );
xnor ( n60740 , n60720 , n60718 );
and ( n60741 , n60739 , n60740 );
or ( n60742 , n60721 , n60741 );
xnor ( n60743 , n60716 , n60714 );
and ( n60744 , n60742 , n60743 );
or ( n60745 , n60717 , n60744 );
xnor ( n60746 , n60712 , n60710 );
and ( n60747 , n60745 , n60746 );
or ( n60748 , n60713 , n60747 );
xnor ( n60749 , n60708 , n60706 );
and ( n60750 , n60748 , n60749 );
or ( n60751 , n60709 , n60750 );
xnor ( n60752 , n60704 , n60702 );
and ( n60753 , n60751 , n60752 );
or ( n60754 , n60705 , n60753 );
xnor ( n60755 , n60700 , n60698 );
and ( n60756 , n60754 , n60755 );
or ( n60757 , n60701 , n60756 );
xnor ( n60758 , n60696 , n60694 );
and ( n60759 , n60757 , n60758 );
or ( n60760 , n60697 , n60759 );
xnor ( n60761 , n60692 , n60690 );
and ( n60762 , n60760 , n60761 );
or ( n60763 , n60693 , n60762 );
xnor ( n60764 , n60688 , n60686 );
and ( n60765 , n60763 , n60764 );
or ( n60766 , n60689 , n60765 );
xnor ( n60767 , n60684 , n60682 );
and ( n60768 , n60766 , n60767 );
or ( n60769 , n60685 , n60768 );
xnor ( n60770 , n60680 , n60678 );
and ( n60771 , n60769 , n60770 );
or ( n60772 , n60681 , n60771 );
xnor ( n60773 , n60676 , n60674 );
and ( n60774 , n60772 , n60773 );
or ( n60775 , n60677 , n60774 );
xnor ( n60776 , n60672 , n60670 );
and ( n60777 , n60775 , n60776 );
or ( n60778 , n60673 , n60777 );
xnor ( n60779 , n60668 , n60666 );
and ( n60780 , n60778 , n60779 );
or ( n60781 , n60669 , n60780 );
xnor ( n60782 , n60664 , n60662 );
and ( n60783 , n60781 , n60782 );
or ( n60784 , n60665 , n60783 );
xnor ( n60785 , n60660 , n60658 );
and ( n60786 , n60784 , n60785 );
or ( n60787 , n60661 , n60786 );
xnor ( n60788 , n60656 , n60654 );
and ( n60789 , n60787 , n60788 );
or ( n60790 , n60657 , n60789 );
xnor ( n60791 , n60652 , n60650 );
and ( n60792 , n60790 , n60791 );
or ( n60793 , n60653 , n60792 );
xnor ( n60794 , n60648 , n60646 );
and ( n60795 , n60793 , n60794 );
or ( n60796 , n60649 , n60795 );
xnor ( n60797 , n60644 , n60642 );
and ( n60798 , n60796 , n60797 );
or ( n60799 , n60645 , n60798 );
xnor ( n60800 , n60640 , n60638 );
and ( n60801 , n60799 , n60800 );
or ( n60802 , n60641 , n60801 );
xnor ( n60803 , n60636 , n60634 );
and ( n60804 , n60802 , n60803 );
or ( n60805 , n60637 , n60804 );
xnor ( n60806 , n60632 , n60630 );
and ( n60807 , n60805 , n60806 );
or ( n60808 , n60633 , n60807 );
xnor ( n60809 , n60628 , n60626 );
and ( n60810 , n60808 , n60809 );
or ( n60811 , n60629 , n60810 );
xnor ( n60812 , n60624 , n60622 );
and ( n60813 , n60811 , n60812 );
or ( n60814 , n60625 , n60813 );
xnor ( n60815 , n60620 , n60618 );
and ( n60816 , n60814 , n60815 );
or ( n60817 , n60621 , n60816 );
xnor ( n60818 , n60616 , n60614 );
and ( n60819 , n60817 , n60818 );
or ( n60820 , n60617 , n60819 );
xnor ( n60821 , n60612 , n60610 );
and ( n60822 , n60820 , n60821 );
or ( n60823 , n60613 , n60822 );
and ( n60824 , n60609 , n60823 );
not ( n60825 , n60606 );
and ( n60826 , n60825 , n60607 );
and ( n60827 , n60826 , n60608 );
or ( n60828 , n60824 , n60827 );
buf ( n60829 , n60828 );
or ( n60830 , n60829 , n27051 );
and ( n60831 , n60830 , n25217 );
not ( n60832 , n60829 );
or ( n60833 , n60832 , n27051 );
and ( n60834 , n60833 , n28594 );
buf ( n60835 , n25876 );
buf ( n60836 , n29094 );
xor ( n60837 , n60835 , n60836 );
buf ( n60838 , n27181 );
buf ( n60839 , n29107 );
xor ( n60840 , n60838 , n60839 );
or ( n60841 , n60837 , n60840 );
buf ( n60842 , n27193 );
buf ( n60843 , n29120 );
xor ( n60844 , n60842 , n60843 );
or ( n60845 , n60841 , n60844 );
buf ( n60846 , n26807 );
buf ( n60847 , n29133 );
xor ( n60848 , n60846 , n60847 );
or ( n60849 , n60845 , n60848 );
buf ( n60850 , n26773 );
buf ( n60851 , n29146 );
xor ( n60852 , n60850 , n60851 );
or ( n60853 , n60849 , n60852 );
buf ( n60854 , n26739 );
buf ( n60855 , n29159 );
xor ( n60856 , n60854 , n60855 );
or ( n60857 , n60853 , n60856 );
buf ( n60858 , n26705 );
buf ( n60859 , n29172 );
xor ( n60860 , n60858 , n60859 );
or ( n60861 , n60857 , n60860 );
buf ( n60862 , n26671 );
buf ( n60863 , n29185 );
xor ( n60864 , n60862 , n60863 );
or ( n60865 , n60861 , n60864 );
buf ( n60866 , n26637 );
buf ( n60867 , n29198 );
xor ( n60868 , n60866 , n60867 );
or ( n60869 , n60865 , n60868 );
buf ( n60870 , n26603 );
buf ( n60871 , n29211 );
xor ( n60872 , n60870 , n60871 );
or ( n60873 , n60869 , n60872 );
buf ( n60874 , n26569 );
buf ( n60875 , n29224 );
xor ( n60876 , n60874 , n60875 );
or ( n60877 , n60873 , n60876 );
buf ( n60878 , n26535 );
buf ( n60879 , n29237 );
xor ( n60880 , n60878 , n60879 );
or ( n60881 , n60877 , n60880 );
buf ( n60882 , n26501 );
buf ( n60883 , n29295 );
xor ( n60884 , n60882 , n60883 );
or ( n60885 , n60881 , n60884 );
buf ( n60886 , n26467 );
buf ( n60887 , n29315 );
xor ( n60888 , n60886 , n60887 );
or ( n60889 , n60885 , n60888 );
buf ( n60890 , n26433 );
buf ( n60891 , n29335 );
xor ( n60892 , n60890 , n60891 );
or ( n60893 , n60889 , n60892 );
buf ( n60894 , n26399 );
buf ( n60895 , n29355 );
xor ( n60896 , n60894 , n60895 );
or ( n60897 , n60893 , n60896 );
buf ( n60898 , n26365 );
buf ( n60899 , n29375 );
xor ( n60900 , n60898 , n60899 );
or ( n60901 , n60897 , n60900 );
buf ( n60902 , n26331 );
buf ( n60903 , n29395 );
xor ( n60904 , n60902 , n60903 );
or ( n60905 , n60901 , n60904 );
buf ( n60906 , n26297 );
buf ( n60907 , n29415 );
xor ( n60908 , n60906 , n60907 );
or ( n60909 , n60905 , n60908 );
buf ( n60910 , n26263 );
buf ( n60911 , n29435 );
xor ( n60912 , n60910 , n60911 );
or ( n60913 , n60909 , n60912 );
buf ( n60914 , n26229 );
buf ( n60915 , n29455 );
xor ( n60916 , n60914 , n60915 );
or ( n60917 , n60913 , n60916 );
buf ( n60918 , n26195 );
buf ( n60919 , n29475 );
xor ( n60920 , n60918 , n60919 );
or ( n60921 , n60917 , n60920 );
buf ( n60922 , n26161 );
buf ( n60923 , n29495 );
xor ( n60924 , n60922 , n60923 );
or ( n60925 , n60921 , n60924 );
buf ( n60926 , n26127 );
buf ( n60927 , n29515 );
xor ( n60928 , n60926 , n60927 );
or ( n60929 , n60925 , n60928 );
buf ( n60930 , n26093 );
buf ( n60931 , n29535 );
xor ( n60932 , n60930 , n60931 );
or ( n60933 , n60929 , n60932 );
buf ( n60934 , n26059 );
buf ( n60935 , n29555 );
xor ( n60936 , n60934 , n60935 );
or ( n60937 , n60933 , n60936 );
buf ( n60938 , n26025 );
buf ( n60939 , n29575 );
xor ( n60940 , n60938 , n60939 );
or ( n60941 , n60937 , n60940 );
buf ( n60942 , n25991 );
buf ( n60943 , n29595 );
xor ( n60944 , n60942 , n60943 );
or ( n60945 , n60941 , n60944 );
buf ( n60946 , n25958 );
buf ( n60947 , n29615 );
xor ( n60948 , n60946 , n60947 );
or ( n60949 , n60945 , n60948 );
buf ( n60950 , n25925 );
buf ( n60951 , n29635 );
xor ( n60952 , n60950 , n60951 );
or ( n60953 , n60949 , n60952 );
buf ( n60954 , n25894 );
buf ( n60955 , n29655 );
xor ( n60956 , n60954 , n60955 );
or ( n60957 , n60953 , n60956 );
buf ( n60958 , n25863 );
buf ( n60959 , n28892 );
xor ( n60960 , n60958 , n60959 );
or ( n60961 , n60957 , n60960 );
not ( n60962 , n60961 );
buf ( n60963 , n60962 );
not ( n60964 , n60963 );
or ( n60965 , n60964 , n27051 );
and ( n60966 , n60965 , n30268 );
or ( n60967 , n60963 , n27051 );
and ( n60968 , n60967 , n30981 );
buf ( n60969 , n25876 );
buf ( n60970 , n29094 );
xor ( n60971 , n60969 , n60970 );
not ( n60972 , n60971 );
buf ( n60973 , n27181 );
not ( n60974 , n60973 );
buf ( n60975 , n29107 );
and ( n60976 , n60974 , n60975 );
buf ( n60977 , n27193 );
not ( n60978 , n60977 );
buf ( n60979 , n29120 );
nand ( n60980 , n60978 , n60979 );
buf ( n60981 , n26807 );
not ( n60982 , n60981 );
buf ( n60983 , n29133 );
nand ( n60984 , n60982 , n60983 );
buf ( n60985 , n26773 );
not ( n60986 , n60985 );
buf ( n60987 , n29146 );
and ( n60988 , n60986 , n60987 );
buf ( n60989 , n26739 );
not ( n60990 , n60989 );
buf ( n60991 , n29159 );
and ( n60992 , n60990 , n60991 );
buf ( n60993 , n26705 );
not ( n60994 , n60993 );
buf ( n60995 , n29172 );
and ( n60996 , n60994 , n60995 );
buf ( n60997 , n26671 );
not ( n60998 , n60997 );
buf ( n60999 , n29185 );
and ( n61000 , n60998 , n60999 );
buf ( n61001 , n26637 );
not ( n61002 , n61001 );
buf ( n61003 , n29198 );
and ( n61004 , n61002 , n61003 );
buf ( n61005 , n26603 );
not ( n61006 , n61005 );
buf ( n61007 , n29211 );
and ( n61008 , n61006 , n61007 );
buf ( n61009 , n26569 );
not ( n61010 , n61009 );
buf ( n61011 , n29224 );
and ( n61012 , n61010 , n61011 );
buf ( n61013 , n26535 );
not ( n61014 , n61013 );
buf ( n61015 , n29237 );
and ( n61016 , n61014 , n61015 );
buf ( n61017 , n26501 );
not ( n61018 , n61017 );
buf ( n61019 , n29295 );
and ( n61020 , n61018 , n61019 );
buf ( n61021 , n26467 );
not ( n61022 , n61021 );
buf ( n61023 , n29315 );
and ( n61024 , n61022 , n61023 );
buf ( n61025 , n26433 );
not ( n61026 , n61025 );
buf ( n61027 , n29335 );
and ( n61028 , n61026 , n61027 );
buf ( n61029 , n26399 );
not ( n61030 , n61029 );
buf ( n61031 , n29355 );
and ( n61032 , n61030 , n61031 );
buf ( n61033 , n26365 );
not ( n61034 , n61033 );
buf ( n61035 , n29375 );
and ( n61036 , n61034 , n61035 );
buf ( n61037 , n26331 );
not ( n61038 , n61037 );
buf ( n61039 , n29395 );
and ( n61040 , n61038 , n61039 );
buf ( n61041 , n26297 );
not ( n61042 , n61041 );
buf ( n61043 , n29415 );
and ( n61044 , n61042 , n61043 );
buf ( n61045 , n26263 );
not ( n61046 , n61045 );
buf ( n61047 , n29435 );
and ( n61048 , n61046 , n61047 );
buf ( n61049 , n26229 );
not ( n61050 , n61049 );
buf ( n61051 , n29455 );
and ( n61052 , n61050 , n61051 );
buf ( n61053 , n26195 );
not ( n61054 , n61053 );
buf ( n61055 , n29475 );
and ( n61056 , n61054 , n61055 );
buf ( n61057 , n26161 );
not ( n61058 , n61057 );
buf ( n61059 , n29495 );
and ( n61060 , n61058 , n61059 );
buf ( n61061 , n26127 );
not ( n61062 , n61061 );
buf ( n61063 , n29515 );
and ( n61064 , n61062 , n61063 );
buf ( n61065 , n26093 );
not ( n61066 , n61065 );
buf ( n61067 , n29535 );
and ( n61068 , n61066 , n61067 );
buf ( n61069 , n26059 );
not ( n61070 , n61069 );
buf ( n61071 , n29555 );
and ( n61072 , n61070 , n61071 );
buf ( n61073 , n26025 );
not ( n61074 , n61073 );
buf ( n61075 , n29575 );
and ( n61076 , n61074 , n61075 );
buf ( n61077 , n25991 );
not ( n61078 , n61077 );
buf ( n61079 , n29595 );
and ( n61080 , n61078 , n61079 );
buf ( n61081 , n25958 );
not ( n61082 , n61081 );
buf ( n61083 , n29615 );
and ( n61084 , n61082 , n61083 );
buf ( n61085 , n25925 );
not ( n61086 , n61085 );
buf ( n61087 , n29635 );
and ( n61088 , n61086 , n61087 );
buf ( n61089 , n25894 );
not ( n61090 , n61089 );
buf ( n61091 , n29655 );
and ( n61092 , n61090 , n61091 );
buf ( n61093 , n25863 );
not ( n61094 , n61093 );
buf ( n61095 , n28892 );
and ( n61096 , n61094 , n61095 );
xnor ( n61097 , n61089 , n61091 );
and ( n61098 , n61096 , n61097 );
or ( n61099 , n61092 , n61098 );
xnor ( n61100 , n61085 , n61087 );
and ( n61101 , n61099 , n61100 );
or ( n61102 , n61088 , n61101 );
xnor ( n61103 , n61081 , n61083 );
and ( n61104 , n61102 , n61103 );
or ( n61105 , n61084 , n61104 );
xnor ( n61106 , n61077 , n61079 );
and ( n61107 , n61105 , n61106 );
or ( n61108 , n61080 , n61107 );
xnor ( n61109 , n61073 , n61075 );
and ( n61110 , n61108 , n61109 );
or ( n61111 , n61076 , n61110 );
xnor ( n61112 , n61069 , n61071 );
and ( n61113 , n61111 , n61112 );
or ( n61114 , n61072 , n61113 );
xnor ( n61115 , n61065 , n61067 );
and ( n61116 , n61114 , n61115 );
or ( n61117 , n61068 , n61116 );
xnor ( n61118 , n61061 , n61063 );
and ( n61119 , n61117 , n61118 );
or ( n61120 , n61064 , n61119 );
xnor ( n61121 , n61057 , n61059 );
and ( n61122 , n61120 , n61121 );
or ( n61123 , n61060 , n61122 );
xnor ( n61124 , n61053 , n61055 );
and ( n61125 , n61123 , n61124 );
or ( n61126 , n61056 , n61125 );
xnor ( n61127 , n61049 , n61051 );
and ( n61128 , n61126 , n61127 );
or ( n61129 , n61052 , n61128 );
xnor ( n61130 , n61045 , n61047 );
and ( n61131 , n61129 , n61130 );
or ( n61132 , n61048 , n61131 );
xnor ( n61133 , n61041 , n61043 );
and ( n61134 , n61132 , n61133 );
or ( n61135 , n61044 , n61134 );
xnor ( n61136 , n61037 , n61039 );
and ( n61137 , n61135 , n61136 );
or ( n61138 , n61040 , n61137 );
xnor ( n61139 , n61033 , n61035 );
and ( n61140 , n61138 , n61139 );
or ( n61141 , n61036 , n61140 );
xnor ( n61142 , n61029 , n61031 );
and ( n61143 , n61141 , n61142 );
or ( n61144 , n61032 , n61143 );
xnor ( n61145 , n61025 , n61027 );
and ( n61146 , n61144 , n61145 );
or ( n61147 , n61028 , n61146 );
xnor ( n61148 , n61021 , n61023 );
and ( n61149 , n61147 , n61148 );
or ( n61150 , n61024 , n61149 );
xnor ( n61151 , n61017 , n61019 );
and ( n61152 , n61150 , n61151 );
or ( n61153 , n61020 , n61152 );
xnor ( n61154 , n61013 , n61015 );
and ( n61155 , n61153 , n61154 );
or ( n61156 , n61016 , n61155 );
xnor ( n61157 , n61009 , n61011 );
and ( n61158 , n61156 , n61157 );
or ( n61159 , n61012 , n61158 );
xnor ( n61160 , n61005 , n61007 );
and ( n61161 , n61159 , n61160 );
or ( n61162 , n61008 , n61161 );
xnor ( n61163 , n61001 , n61003 );
and ( n61164 , n61162 , n61163 );
or ( n61165 , n61004 , n61164 );
xnor ( n61166 , n60997 , n60999 );
and ( n61167 , n61165 , n61166 );
or ( n61168 , n61000 , n61167 );
xnor ( n61169 , n60993 , n60995 );
and ( n61170 , n61168 , n61169 );
or ( n61171 , n60996 , n61170 );
xnor ( n61172 , n60989 , n60991 );
and ( n61173 , n61171 , n61172 );
or ( n61174 , n60992 , n61173 );
xnor ( n61175 , n60985 , n60987 );
and ( n61176 , n61174 , n61175 );
or ( n61177 , n60988 , n61176 );
xnor ( n61178 , n60981 , n60983 );
and ( n61179 , n61177 , n61178 );
or ( n61180 , n60984 , n61179 );
xnor ( n61181 , n60977 , n60979 );
and ( n61182 , n61180 , n61181 );
or ( n61183 , n60980 , n61182 );
xnor ( n61184 , n60973 , n60975 );
and ( n61185 , n61183 , n61184 );
or ( n61186 , n60976 , n61185 );
and ( n61187 , n60972 , n61186 );
not ( n61188 , n60970 );
and ( n61189 , n61188 , n60969 );
and ( n61190 , n61189 , n60971 );
or ( n61191 , n61187 , n61190 );
buf ( n61192 , n61191 );
not ( n61193 , n61192 );
or ( n61194 , n61193 , n27051 );
and ( n61195 , n61194 , n30266 );
or ( n61196 , n61192 , n27051 );
and ( n61197 , n61196 , n30979 );
and ( n61198 , n60601 , n30264 );
and ( n61199 , n60600 , n30263 );
and ( n61200 , n60829 , n30977 );
and ( n61201 , n60832 , n30976 );
and ( n61202 , n60964 , n30988 );
and ( n61203 , n60963 , n30987 );
and ( n61204 , n61193 , n30991 );
and ( n61205 , n61192 , n31002 );
or ( n61206 , n60603 , n60605 , n60831 , n60834 , n60966 , n60968 , n61195 , n61197 , n61198 , n61199 , n61200 , n61201 , n61202 , n61203 , n61204 , n61205 );
and ( n61207 , n61206 , n24511 );
or ( n61208 , n60335 , n61207 );
and ( n61209 , n61208 , n31008 );
and ( n61210 , n27051 , n10618 );
or ( n61211 , n61209 , n61210 );
buf ( n61212 , n61211 );
buf ( n61213 , n61212 );
buf ( n61214 , n10613 );
not ( n61215 , n11954 );
not ( n61216 , n12243 );
and ( n61217 , n10805 , n31187 );
not ( n61218 , n31697 );
and ( n61219 , n61218 , n31676 );
xor ( n61220 , n56878 , n56891 );
and ( n61221 , n61220 , n31697 );
or ( n61222 , n61219 , n61221 );
buf ( n61223 , n61222 );
and ( n61224 , n61223 , n14140 );
not ( n61225 , n32214 );
and ( n61226 , n61225 , n32193 );
xor ( n61227 , n56901 , n56914 );
and ( n61228 , n61227 , n32214 );
or ( n61229 , n61226 , n61228 );
buf ( n61230 , n61229 );
and ( n61231 , n61230 , n14137 );
and ( n61232 , n15469 , n14143 );
and ( n61233 , n10805 , n14141 );
or ( n61234 , n61224 , n61231 , n61232 , n61233 );
and ( n61235 , n61234 , n32236 );
or ( n61236 , n61217 , n61235 );
and ( n61237 , n61216 , n61236 );
not ( n61238 , n34038 );
and ( n61239 , n61238 , n34010 );
xor ( n61240 , n56930 , n56943 );
and ( n61241 , n61240 , n34038 );
or ( n61242 , n61239 , n61241 );
buf ( n61243 , n61242 );
and ( n61244 , n61243 , n12243 );
or ( n61245 , n61237 , n61244 );
and ( n61246 , n61215 , n61245 );
and ( n61247 , n61234 , n11954 );
or ( n61248 , n61246 , n61247 );
and ( n61249 , n61248 , n16574 );
not ( n61250 , n34327 );
and ( n61251 , n61250 , n34309 );
xor ( n61252 , n56958 , n56971 );
and ( n61253 , n61252 , n34327 );
or ( n61254 , n61251 , n61253 );
buf ( n61255 , n61254 );
and ( n61256 , n61255 , n16576 );
or ( n61257 , n61249 , n61256 );
buf ( n61258 , n61257 );
buf ( n61259 , n61258 );
buf ( n61260 , n10613 );
buf ( n61261 , n10613 );
buf ( n61262 , n10615 );
not ( n61263 , n24800 );
and ( n61264 , n26665 , n25222 );
and ( n61265 , n48044 , n28583 );
and ( n61266 , n26665 , n28591 );
or ( n61267 , n61265 , n61266 );
and ( n61268 , n61267 , n28594 );
and ( n61269 , n48054 , n28583 );
and ( n61270 , n26665 , n28591 );
or ( n61271 , n61269 , n61270 );
and ( n61272 , n61271 , n30269 );
and ( n61273 , n48064 , n28583 );
and ( n61274 , n26665 , n28591 );
or ( n61275 , n61273 , n61274 );
and ( n61276 , n61275 , n30982 );
and ( n61277 , n29185 , n28583 );
and ( n61278 , n26665 , n28591 );
or ( n61279 , n61277 , n61278 );
and ( n61280 , n61279 , n30989 );
and ( n61281 , n26663 , n30991 );
and ( n61282 , n48075 , n28583 );
and ( n61283 , n26665 , n28591 );
or ( n61284 , n61282 , n61283 );
and ( n61285 , n61284 , n31002 );
or ( n61286 , n61264 , n61268 , n61272 , n61276 , n61280 , n61281 , n61285 );
and ( n61287 , n61263 , n61286 );
and ( n61288 , n26665 , n24800 );
or ( n61289 , n61287 , n61288 );
and ( n61290 , n61289 , n31008 );
and ( n61291 , n26665 , n10618 );
or ( n61292 , n61290 , n61291 );
buf ( n61293 , n61292 );
buf ( n61294 , n61293 );
buf ( n61295 , n10613 );
not ( n61296 , n17451 );
and ( n61297 , n18538 , n17873 );
and ( n61298 , n34754 , n21336 );
and ( n61299 , n18538 , n42682 );
or ( n61300 , n61298 , n61299 );
and ( n61301 , n61300 , n21341 );
and ( n61302 , n34767 , n21336 );
and ( n61303 , n18538 , n42682 );
or ( n61304 , n61302 , n61303 );
and ( n61305 , n61304 , n23064 );
and ( n61306 , n34777 , n21336 );
and ( n61307 , n18538 , n42682 );
or ( n61308 , n61306 , n61307 );
and ( n61309 , n61308 , n23825 );
and ( n61310 , n22402 , n21336 );
and ( n61311 , n18538 , n42682 );
or ( n61312 , n61310 , n61311 );
and ( n61313 , n61312 , n23832 );
and ( n61314 , n22402 , n23834 );
and ( n61315 , n34787 , n21336 );
and ( n61316 , n18538 , n42682 );
or ( n61317 , n61315 , n61316 );
and ( n61318 , n61317 , n23917 );
or ( n61319 , n61297 , n61301 , n61305 , n61309 , n61313 , n61314 , n61318 );
and ( n61320 , n61296 , n61319 );
and ( n61321 , n18538 , n17451 );
or ( n61322 , n61320 , n61321 );
and ( n61323 , n61322 , n23924 );
and ( n61324 , n17885 , n23926 );
or ( n61325 , n61323 , n61324 );
buf ( n61326 , n61325 );
buf ( n61327 , n61326 );
not ( n61328 , n17451 );
and ( n61329 , n42969 , n21333 );
and ( n61330 , n18877 , n34758 );
or ( n61331 , n61329 , n61330 );
and ( n61332 , n61331 , n21341 );
and ( n61333 , n42979 , n21333 );
and ( n61334 , n18877 , n34758 );
or ( n61335 , n61333 , n61334 );
and ( n61336 , n61335 , n23064 );
and ( n61337 , n42989 , n21333 );
and ( n61338 , n18877 , n34758 );
or ( n61339 , n61337 , n61338 );
and ( n61340 , n61339 , n23825 );
and ( n61341 , n22202 , n21333 );
and ( n61342 , n18877 , n34758 );
or ( n61343 , n61341 , n61342 );
and ( n61344 , n61343 , n23832 );
and ( n61345 , n42999 , n21333 );
and ( n61346 , n18877 , n34758 );
or ( n61347 , n61345 , n61346 );
and ( n61348 , n61347 , n23917 );
and ( n61349 , n18877 , n34526 );
or ( n61350 , n61332 , n61336 , n61340 , n61344 , n61348 , n61349 );
and ( n61351 , n61328 , n61350 );
and ( n61352 , n18877 , n17451 );
or ( n61353 , n61351 , n61352 );
and ( n61354 , n61353 , n23924 );
and ( n61355 , n18877 , n23926 );
or ( n61356 , n61354 , n61355 );
buf ( n61357 , n61356 );
buf ( n61358 , n61357 );
buf ( n61359 , n10613 );
not ( n61360 , n34821 );
and ( n61361 , n55616 , n36347 );
and ( n61362 , n14607 , n39408 );
or ( n61363 , n61361 , n61362 );
and ( n61364 , n61363 , n14562 );
and ( n61365 , n55625 , n36348 );
and ( n61366 , n14607 , n39427 );
or ( n61367 , n61365 , n61366 );
and ( n61368 , n61367 , n14586 );
and ( n61369 , n55634 , n36347 );
and ( n61370 , n14607 , n39446 );
or ( n61371 , n61369 , n61370 );
and ( n61372 , n61371 , n14584 );
and ( n61373 , n55625 , n36348 );
and ( n61374 , n14607 , n39453 );
or ( n61375 , n61373 , n61374 );
and ( n61376 , n61375 , n37835 );
and ( n61377 , n55634 , n36348 );
and ( n61378 , n14607 , n39453 );
or ( n61379 , n61377 , n61378 );
and ( n61380 , n61379 , n37841 );
and ( n61381 , n14952 , n36348 );
and ( n61382 , n14607 , n39453 );
or ( n61383 , n61381 , n61382 );
and ( n61384 , n61383 , n37847 );
and ( n61385 , n14607 , n37849 );
or ( n61386 , n61364 , n61368 , n61372 , n61376 , n61380 , n61384 , n61385 );
and ( n61387 , n61360 , n61386 );
and ( n61388 , n14607 , n34821 );
or ( n61389 , n61387 , n61388 );
and ( n61390 , n61389 , n16574 );
and ( n61391 , n14607 , n16576 );
or ( n61392 , n61390 , n61391 );
buf ( n61393 , n61392 );
buf ( n61394 , n61393 );
buf ( n61395 , n10615 );
buf ( n61396 , n10615 );
buf ( n61397 , n10613 );
buf ( n61398 , n10613 );
buf ( n61399 , n10613 );
not ( n61400 , n17451 );
and ( n61401 , n19452 , n17873 );
and ( n61402 , n45354 , n21330 );
and ( n61403 , n19452 , n21338 );
or ( n61404 , n61402 , n61403 );
and ( n61405 , n61404 , n21341 );
and ( n61406 , n45364 , n21330 );
and ( n61407 , n19452 , n21338 );
or ( n61408 , n61406 , n61407 );
and ( n61409 , n61408 , n23064 );
and ( n61410 , n45374 , n21330 );
and ( n61411 , n19452 , n21338 );
or ( n61412 , n61410 , n61411 );
and ( n61413 , n61412 , n23825 );
and ( n61414 , n21880 , n21330 );
and ( n61415 , n19452 , n21338 );
or ( n61416 , n61414 , n61415 );
and ( n61417 , n61416 , n23832 );
and ( n61418 , n19450 , n23834 );
and ( n61419 , n45384 , n21330 );
and ( n61420 , n19452 , n21338 );
or ( n61421 , n61419 , n61420 );
and ( n61422 , n61421 , n23917 );
or ( n61423 , n61401 , n61405 , n61409 , n61413 , n61417 , n61418 , n61422 );
and ( n61424 , n61400 , n61423 );
and ( n61425 , n19452 , n17451 );
or ( n61426 , n61424 , n61425 );
and ( n61427 , n61426 , n23924 );
and ( n61428 , n19452 , n23926 );
or ( n61429 , n61427 , n61428 );
buf ( n61430 , n61429 );
buf ( n61431 , n61430 );
not ( n61432 , n17451 );
and ( n61433 , n19249 , n17873 );
and ( n61434 , n47430 , n21330 );
and ( n61435 , n19249 , n21338 );
or ( n61436 , n61434 , n61435 );
and ( n61437 , n61436 , n21341 );
and ( n61438 , n47440 , n21330 );
and ( n61439 , n19249 , n21338 );
or ( n61440 , n61438 , n61439 );
and ( n61441 , n61440 , n23064 );
and ( n61442 , n47450 , n21330 );
and ( n61443 , n19249 , n21338 );
or ( n61444 , n61442 , n61443 );
and ( n61445 , n61444 , n23825 );
and ( n61446 , n21958 , n21330 );
and ( n61447 , n19249 , n21338 );
or ( n61448 , n61446 , n61447 );
and ( n61449 , n61448 , n23832 );
and ( n61450 , n19247 , n23834 );
and ( n61451 , n47461 , n21330 );
and ( n61452 , n19249 , n21338 );
or ( n61453 , n61451 , n61452 );
and ( n61454 , n61453 , n23917 );
or ( n61455 , n61433 , n61437 , n61441 , n61445 , n61449 , n61450 , n61454 );
and ( n61456 , n61432 , n61455 );
and ( n61457 , n19249 , n17451 );
or ( n61458 , n61456 , n61457 );
and ( n61459 , n61458 , n23924 );
and ( n61460 , n19249 , n23926 );
or ( n61461 , n61459 , n61460 );
buf ( n61462 , n61461 );
buf ( n61463 , n61462 );
buf ( n61464 , n10615 );
buf ( n61465 , n10613 );
buf ( n61466 , n10615 );
buf ( n61467 , n10613 );
buf ( n61468 , n10615 );
buf ( n61469 , n10615 );
buf ( n61470 , n10615 );
not ( n61471 , n34821 );
and ( n61472 , n47213 , n36345 );
and ( n61473 , n13147 , n36352 );
or ( n61474 , n61472 , n61473 );
and ( n61475 , n61474 , n14562 );
and ( n61476 , n13147 , n37073 );
or ( n61477 , C0 , n61476 );
and ( n61478 , n61477 , n14586 );
and ( n61479 , n13147 , n37825 );
or ( n61480 , C0 , n61479 );
and ( n61481 , n61480 , n14584 );
and ( n61482 , n13147 , n37831 );
or ( n61483 , C0 , n61482 );
and ( n61484 , n61483 , n37835 );
and ( n61485 , n13147 , n37831 );
or ( n61486 , C0 , n61485 );
and ( n61487 , n61486 , n37841 );
and ( n61488 , n14934 , n36350 );
and ( n61489 , n13147 , n37831 );
or ( n61490 , n61488 , n61489 );
and ( n61491 , n61490 , n37847 );
and ( n61492 , n13147 , n37849 );
or ( n61493 , n61475 , n61478 , n61481 , n61484 , n61487 , n61491 , n61492 );
and ( n61494 , n61471 , n61493 );
and ( n61495 , n13147 , n34821 );
or ( n61496 , n61494 , n61495 );
and ( n61497 , n61496 , n16574 );
and ( n61498 , n13147 , n16576 );
or ( n61499 , n61497 , n61498 );
buf ( n61500 , n61499 );
buf ( n61501 , n61500 );
buf ( n61502 , n10615 );
buf ( n61503 , n10613 );
buf ( n61504 , n10613 );
not ( n61505 , n11954 );
not ( n61506 , n12243 );
and ( n61507 , n10845 , n31187 );
not ( n61508 , n31697 );
and ( n61509 , n61508 , n31591 );
xor ( n61510 , n56883 , n56886 );
and ( n61511 , n61510 , n31697 );
or ( n61512 , n61509 , n61511 );
buf ( n61513 , n61512 );
and ( n61514 , n61513 , n14140 );
not ( n61515 , n32214 );
and ( n61516 , n61515 , n32108 );
xor ( n61517 , n56906 , n56909 );
and ( n61518 , n61517 , n32214 );
or ( n61519 , n61516 , n61518 );
buf ( n61520 , n61519 );
and ( n61521 , n61520 , n14137 );
and ( n61522 , n15579 , n14143 );
and ( n61523 , n10845 , n14141 );
or ( n61524 , n61514 , n61521 , n61522 , n61523 );
and ( n61525 , n61524 , n32236 );
or ( n61526 , n61507 , n61525 );
and ( n61527 , n61506 , n61526 );
not ( n61528 , n34038 );
and ( n61529 , n61528 , n33890 );
xor ( n61530 , n56935 , n56938 );
and ( n61531 , n61530 , n34038 );
or ( n61532 , n61529 , n61531 );
buf ( n61533 , n61532 );
and ( n61534 , n61533 , n12243 );
or ( n61535 , n61527 , n61534 );
and ( n61536 , n61505 , n61535 );
and ( n61537 , n61524 , n11954 );
or ( n61538 , n61536 , n61537 );
and ( n61539 , n61538 , n16574 );
not ( n61540 , n34327 );
and ( n61541 , n61540 , n34239 );
xor ( n61542 , n56963 , n56966 );
and ( n61543 , n61542 , n34327 );
or ( n61544 , n61541 , n61543 );
buf ( n61545 , n61544 );
and ( n61546 , n61545 , n16576 );
or ( n61547 , n61539 , n61546 );
buf ( n61548 , n61547 );
buf ( n61549 , n61548 );
buf ( n61550 , n10613 );
buf ( n61551 , n10613 );
buf ( n61552 , n10615 );
not ( n61553 , n34538 );
and ( n61554 , n61553 , n18546 );
and ( n61555 , n14825 , n34538 );
or ( n61556 , n61554 , n61555 );
and ( n61557 , n61556 , n23924 );
and ( n61558 , n14825 , n23926 );
or ( n61559 , n61557 , n61558 );
buf ( n61560 , n61559 );
buf ( n61561 , n61560 );
buf ( n61562 , n10613 );
buf ( n61563 , n10613 );
not ( n61564 , n24800 );
and ( n61565 , n43420 , n28586 );
and ( n61566 , n26701 , n34573 );
or ( n61567 , n61565 , n61566 );
and ( n61568 , n61567 , n28594 );
and ( n61569 , n43436 , n28586 );
and ( n61570 , n26701 , n34573 );
or ( n61571 , n61569 , n61570 );
and ( n61572 , n61571 , n30269 );
and ( n61573 , n43452 , n28586 );
and ( n61574 , n26701 , n34573 );
or ( n61575 , n61573 , n61574 );
and ( n61576 , n61575 , n30982 );
and ( n61577 , n29172 , n28586 );
and ( n61578 , n26701 , n34573 );
or ( n61579 , n61577 , n61578 );
and ( n61580 , n61579 , n30989 );
and ( n61581 , n43471 , n28586 );
and ( n61582 , n26701 , n34573 );
or ( n61583 , n61581 , n61582 );
and ( n61584 , n61583 , n31002 );
and ( n61585 , n26701 , n34607 );
or ( n61586 , n61568 , n61572 , n61576 , n61580 , n61584 , n61585 );
and ( n61587 , n61564 , n61586 );
and ( n61588 , n26701 , n24800 );
or ( n61589 , n61587 , n61588 );
and ( n61590 , n61589 , n31008 );
and ( n61591 , n26701 , n10618 );
or ( n61592 , n61590 , n61591 );
buf ( n61593 , n61592 );
buf ( n61594 , n61593 );
not ( n61595 , n17451 );
and ( n61596 , n19011 , n17873 );
and ( n61597 , n58841 , n21330 );
and ( n61598 , n19011 , n21338 );
or ( n61599 , n61597 , n61598 );
and ( n61600 , n61599 , n21341 );
and ( n61601 , n58851 , n21330 );
and ( n61602 , n19011 , n21338 );
or ( n61603 , n61601 , n61602 );
and ( n61604 , n61603 , n23064 );
and ( n61605 , n58861 , n21330 );
and ( n61606 , n19011 , n21338 );
or ( n61607 , n61605 , n61606 );
and ( n61608 , n61607 , n23825 );
and ( n61609 , n22122 , n21330 );
and ( n61610 , n19011 , n21338 );
or ( n61611 , n61609 , n61610 );
and ( n61612 , n61611 , n23832 );
and ( n61613 , n19009 , n23834 );
and ( n61614 , n58872 , n21330 );
and ( n61615 , n19011 , n21338 );
or ( n61616 , n61614 , n61615 );
and ( n61617 , n61616 , n23917 );
or ( n61618 , n61596 , n61600 , n61604 , n61608 , n61612 , n61613 , n61617 );
and ( n61619 , n61595 , n61618 );
and ( n61620 , n19011 , n17451 );
or ( n61621 , n61619 , n61620 );
and ( n61622 , n61621 , n23924 );
and ( n61623 , n19011 , n23926 );
or ( n61624 , n61622 , n61623 );
buf ( n61625 , n61624 );
buf ( n61626 , n61625 );
not ( n61627 , n24800 );
and ( n61628 , n26563 , n25222 );
and ( n61629 , n45874 , n28583 );
and ( n61630 , n26563 , n28591 );
or ( n61631 , n61629 , n61630 );
and ( n61632 , n61631 , n28594 );
and ( n61633 , n45884 , n28583 );
and ( n61634 , n26563 , n28591 );
or ( n61635 , n61633 , n61634 );
and ( n61636 , n61635 , n30269 );
and ( n61637 , n45894 , n28583 );
and ( n61638 , n26563 , n28591 );
or ( n61639 , n61637 , n61638 );
and ( n61640 , n61639 , n30982 );
and ( n61641 , n29224 , n28583 );
and ( n61642 , n26563 , n28591 );
or ( n61643 , n61641 , n61642 );
and ( n61644 , n61643 , n30989 );
and ( n61645 , n26561 , n30991 );
and ( n61646 , n45905 , n28583 );
and ( n61647 , n26563 , n28591 );
or ( n61648 , n61646 , n61647 );
and ( n61649 , n61648 , n31002 );
or ( n61650 , n61628 , n61632 , n61636 , n61640 , n61644 , n61645 , n61649 );
and ( n61651 , n61627 , n61650 );
and ( n61652 , n26563 , n24800 );
or ( n61653 , n61651 , n61652 );
and ( n61654 , n61653 , n31008 );
and ( n61655 , n26563 , n10618 );
or ( n61656 , n61654 , n61655 );
buf ( n61657 , n61656 );
buf ( n61658 , n61657 );
not ( n61659 , n24511 );
not ( n61660 , n24799 );
and ( n61661 , n10685 , n40154 );
not ( n61662 , n40632 );
and ( n61663 , n61662 , n40475 );
xor ( n61664 , n40640 , n40660 );
and ( n61665 , n61664 , n40632 );
or ( n61666 , n61663 , n61665 );
buf ( n61667 , n61666 );
and ( n61668 , n61667 , n27046 );
not ( n61669 , n41147 );
and ( n61670 , n61669 , n40990 );
xor ( n61671 , n41155 , n41175 );
and ( n61672 , n61671 , n41147 );
or ( n61673 , n61670 , n61672 );
buf ( n61674 , n61673 );
and ( n61675 , n61674 , n27049 );
and ( n61676 , n29473 , n28506 );
and ( n61677 , n10685 , n28508 );
or ( n61678 , n61668 , n61675 , n61676 , n61677 );
and ( n61679 , n61678 , n41199 );
or ( n61680 , n61661 , n61679 );
and ( n61681 , n61660 , n61680 );
xor ( n61682 , n41596 , n41604 );
xor ( n61683 , n61682 , n41791 );
buf ( n61684 , n61683 );
and ( n61685 , n61684 , n27046 );
xor ( n61686 , n42168 , n42169 );
xor ( n61687 , n61686 , n42287 );
buf ( n61688 , n61687 );
and ( n61689 , n61688 , n27049 );
and ( n61690 , n29473 , n42306 );
or ( n61691 , n61685 , n61689 , n61690 );
buf ( n61692 , n61691 );
and ( n61693 , C1 , n61692 );
or ( n61694 , n61693 , C0 );
buf ( n61695 , n61694 );
not ( n61696 , n61695 );
buf ( n61697 , n61696 );
buf ( n61698 , n61697 );
not ( n61699 , n61698 );
and ( n61700 , C1 , n61699 );
or ( n61701 , n61700 , C0 );
buf ( n61702 , n61701 );
and ( n61703 , n61702 , n24799 );
or ( n61704 , n61681 , n61703 );
and ( n61705 , n61659 , n61704 );
and ( n61706 , n61678 , n24511 );
or ( n61707 , n61705 , n61706 );
and ( n61708 , n61707 , n31008 );
not ( n61709 , n42601 );
and ( n61710 , n61709 , n42471 );
xor ( n61711 , n42609 , n42629 );
and ( n61712 , n61711 , n42601 );
or ( n61713 , n61710 , n61712 );
buf ( n61714 , n61713 );
and ( n61715 , n61714 , n10618 );
or ( n61716 , n61708 , n61715 );
buf ( n61717 , n61716 );
buf ( n61718 , n61717 );
buf ( n61719 , n10613 );
and ( n61720 , n24078 , n31008 );
and ( n61721 , n29209 , n10618 );
or ( n61722 , n61720 , n61721 );
buf ( n61723 , n61722 );
buf ( n61724 , n61723 );
not ( n61725 , n24800 );
and ( n61726 , n47500 , n28587 );
and ( n61727 , n26499 , n39807 );
or ( n61728 , n61726 , n61727 );
and ( n61729 , n61728 , n28594 );
and ( n61730 , n47510 , n28587 );
and ( n61731 , n26499 , n39807 );
or ( n61732 , n61730 , n61731 );
and ( n61733 , n61732 , n30269 );
and ( n61734 , n47520 , n28587 );
and ( n61735 , n26499 , n39807 );
or ( n61736 , n61734 , n61735 );
and ( n61737 , n61736 , n30982 );
and ( n61738 , n29295 , n28587 );
and ( n61739 , n26499 , n39807 );
or ( n61740 , n61738 , n61739 );
and ( n61741 , n61740 , n30989 );
and ( n61742 , n47531 , n28587 );
and ( n61743 , n26499 , n39807 );
or ( n61744 , n61742 , n61743 );
and ( n61745 , n61744 , n31002 );
and ( n61746 , n26499 , n34607 );
or ( n61747 , n61729 , n61733 , n61737 , n61741 , n61745 , n61746 );
and ( n61748 , n61725 , n61747 );
and ( n61749 , n26499 , n24800 );
or ( n61750 , n61748 , n61749 );
and ( n61751 , n61750 , n31008 );
and ( n61752 , n26499 , n10618 );
or ( n61753 , n61751 , n61752 );
buf ( n61754 , n61753 );
buf ( n61755 , n61754 );
buf ( n61756 , n10613 );
buf ( n61757 , n10613 );
buf ( n61758 , n10615 );
buf ( n61759 , n10615 );
buf ( n61760 , n10615 );
buf ( n61761 , n10615 );
buf ( n61762 , n10615 );
not ( n61763 , n12243 );
or ( n61764 , n11954 , n61763 );
not ( n61765 , n61764 );
and ( n61766 , n12243 , n61765 );
and ( n61767 , n61766 , n16574 );
buf ( n61768 , n61767 );
buf ( n61769 , n61768 );
not ( n61770 , n11333 );
and ( n61771 , n61770 , n11244 );
xor ( n61772 , n11337 , n11365 );
and ( n61773 , n61772 , n11333 );
or ( n61774 , n61771 , n61773 );
buf ( n61775 , n61774 );
buf ( n61776 , n61775 );
buf ( n61777 , n10613 );
buf ( n61778 , n10613 );
buf ( n61779 , n10613 );
buf ( n61780 , n10613 );
buf ( n61781 , n10613 );
buf ( n61782 , n10613 );
buf ( n61783 , n10613 );
not ( n61784 , n34821 );
and ( n61785 , n13179 , n14592 );
and ( n61786 , n46418 , n36350 );
and ( n61787 , n13179 , n43691 );
or ( n61788 , n61786 , n61787 );
and ( n61789 , n61788 , n14562 );
and ( n61790 , n46436 , n36350 );
and ( n61791 , n13179 , n43703 );
or ( n61792 , n61790 , n61791 );
and ( n61793 , n61792 , n14586 );
and ( n61794 , n46454 , n36345 );
and ( n61795 , n13179 , n43715 );
or ( n61796 , n61794 , n61795 );
and ( n61797 , n61796 , n14584 );
and ( n61798 , n46436 , n36345 );
and ( n61799 , n13179 , n43721 );
or ( n61800 , n61798 , n61799 );
and ( n61801 , n61800 , n37835 );
and ( n61802 , n46454 , n36345 );
and ( n61803 , n13179 , n43721 );
or ( n61804 , n61802 , n61803 );
and ( n61805 , n61804 , n37841 );
and ( n61806 , n15022 , n14564 );
and ( n61807 , n15022 , n36345 );
and ( n61808 , n13179 , n43721 );
or ( n61809 , n61807 , n61808 );
and ( n61810 , n61809 , n37847 );
or ( n61811 , n61785 , n61789 , n61793 , n61797 , n61801 , n61805 , n61806 , n61810 );
and ( n61812 , n61784 , n61811 );
and ( n61813 , n13179 , n34821 );
or ( n61814 , n61812 , n61813 );
and ( n61815 , n61814 , n16574 );
and ( n61816 , n12255 , n16576 );
or ( n61817 , n61815 , n61816 );
buf ( n61818 , n61817 );
buf ( n61819 , n61818 );
buf ( n61820 , n10613 );
not ( n61821 , n34804 );
and ( n61822 , n61821 , n26365 );
and ( n61823 , n14743 , n34804 );
or ( n61824 , n61822 , n61823 );
and ( n61825 , n61824 , n31008 );
and ( n61826 , n14743 , n10618 );
or ( n61827 , n61825 , n61826 );
buf ( n61828 , n61827 );
buf ( n61829 , n61828 );
buf ( n61830 , n10613 );
buf ( n61831 , n10613 );
buf ( n61832 , n10613 );
buf ( n61833 , n10613 );
not ( n61834 , n24511 );
not ( n61835 , n24799 );
and ( n61836 , n10675 , n40154 );
not ( n61837 , n40632 );
and ( n61838 , n61837 , n40509 );
xor ( n61839 , n40638 , n40662 );
and ( n61840 , n61839 , n40632 );
or ( n61841 , n61838 , n61840 );
buf ( n61842 , n61841 );
and ( n61843 , n61842 , n27046 );
not ( n61844 , n41147 );
and ( n61845 , n61844 , n41024 );
xor ( n61846 , n41153 , n41177 );
and ( n61847 , n61846 , n41147 );
or ( n61848 , n61845 , n61847 );
buf ( n61849 , n61848 );
and ( n61850 , n61849 , n27049 );
and ( n61851 , n29433 , n28506 );
and ( n61852 , n10675 , n28508 );
or ( n61853 , n61843 , n61850 , n61851 , n61852 );
and ( n61854 , n61853 , n41199 );
or ( n61855 , n61836 , n61854 );
and ( n61856 , n61835 , n61855 );
xor ( n61857 , n41564 , n41572 );
xor ( n61858 , n61857 , n41797 );
buf ( n61859 , n61858 );
and ( n61860 , n61859 , n27046 );
xor ( n61861 , n42150 , n42151 );
xor ( n61862 , n61861 , n42293 );
buf ( n61863 , n61862 );
and ( n61864 , n61863 , n27049 );
and ( n61865 , n29433 , n42306 );
or ( n61866 , n61860 , n61864 , n61865 );
buf ( n61867 , n61866 );
and ( n61868 , C1 , n61867 );
or ( n61869 , n61868 , C0 );
buf ( n61870 , n61869 );
not ( n61871 , n61870 );
buf ( n61872 , n61871 );
buf ( n61873 , n61872 );
not ( n61874 , n61873 );
and ( n61875 , C1 , n61874 );
or ( n61876 , n61875 , C0 );
buf ( n61877 , n61876 );
and ( n61878 , n61877 , n24799 );
or ( n61879 , n61856 , n61878 );
and ( n61880 , n61834 , n61879 );
and ( n61881 , n61853 , n24511 );
or ( n61882 , n61880 , n61881 );
and ( n61883 , n61882 , n31008 );
not ( n61884 , n42601 );
and ( n61885 , n61884 , n42499 );
xor ( n61886 , n42607 , n42631 );
and ( n61887 , n61886 , n42601 );
or ( n61888 , n61885 , n61887 );
buf ( n61889 , n61888 );
and ( n61890 , n61889 , n10618 );
or ( n61891 , n61883 , n61890 );
buf ( n61892 , n61891 );
buf ( n61893 , n61892 );
not ( n61894 , n34821 );
and ( n61895 , n13229 , n14592 );
and ( n61896 , n45746 , n36348 );
and ( n61897 , n13229 , n43530 );
or ( n61898 , n61896 , n61897 );
and ( n61899 , n61898 , n14562 );
and ( n61900 , n45762 , n36347 );
and ( n61901 , n13229 , n43543 );
or ( n61902 , n61900 , n61901 );
and ( n61903 , n61902 , n14586 );
and ( n61904 , n45778 , n36348 );
and ( n61905 , n13229 , n43556 );
or ( n61906 , n61904 , n61905 );
and ( n61907 , n61906 , n14584 );
and ( n61908 , n45762 , n36347 );
and ( n61909 , n13229 , n43563 );
or ( n61910 , n61908 , n61909 );
and ( n61911 , n61910 , n37835 );
and ( n61912 , n45778 , n36347 );
and ( n61913 , n13229 , n43563 );
or ( n61914 , n61912 , n61913 );
and ( n61915 , n61914 , n37841 );
and ( n61916 , n13227 , n14564 );
and ( n61917 , n15082 , n36347 );
and ( n61918 , n13229 , n43563 );
or ( n61919 , n61917 , n61918 );
and ( n61920 , n61919 , n37847 );
or ( n61921 , n61895 , n61899 , n61903 , n61907 , n61911 , n61915 , n61916 , n61920 );
and ( n61922 , n61894 , n61921 );
and ( n61923 , n13229 , n34821 );
or ( n61924 , n61922 , n61923 );
and ( n61925 , n61924 , n16574 );
and ( n61926 , n13229 , n16576 );
or ( n61927 , n61925 , n61926 );
buf ( n61928 , n61927 );
buf ( n61929 , n61928 );
buf ( n61930 , n10615 );
not ( n61931 , n24800 );
and ( n61932 , n26119 , n25222 );
and ( n61933 , n49846 , n28589 );
and ( n61934 , n26119 , n31075 );
or ( n61935 , n61933 , n61934 );
and ( n61936 , n61935 , n28594 );
and ( n61937 , n49856 , n28589 );
and ( n61938 , n26119 , n31075 );
or ( n61939 , n61937 , n61938 );
and ( n61940 , n61939 , n30269 );
and ( n61941 , n49866 , n28589 );
and ( n61942 , n26119 , n31075 );
or ( n61943 , n61941 , n61942 );
and ( n61944 , n61943 , n30982 );
and ( n61945 , n29515 , n28589 );
and ( n61946 , n26119 , n31075 );
or ( n61947 , n61945 , n61946 );
and ( n61948 , n61947 , n30989 );
and ( n61949 , n29515 , n30991 );
and ( n61950 , n49876 , n28589 );
and ( n61951 , n26119 , n31075 );
or ( n61952 , n61950 , n61951 );
and ( n61953 , n61952 , n31002 );
or ( n61954 , n61932 , n61936 , n61940 , n61944 , n61948 , n61949 , n61953 );
and ( n61955 , n61931 , n61954 );
and ( n61956 , n26119 , n24800 );
or ( n61957 , n61955 , n61956 );
and ( n61958 , n61957 , n31008 );
and ( n61959 , n25339 , n10618 );
or ( n61960 , n61958 , n61959 );
buf ( n61961 , n61960 );
buf ( n61962 , n61961 );
not ( n61963 , n24800 );
and ( n61964 , n48044 , n28587 );
and ( n61965 , n26669 , n39807 );
or ( n61966 , n61964 , n61965 );
and ( n61967 , n61966 , n28594 );
and ( n61968 , n48054 , n28587 );
and ( n61969 , n26669 , n39807 );
or ( n61970 , n61968 , n61969 );
and ( n61971 , n61970 , n30269 );
and ( n61972 , n48064 , n28587 );
and ( n61973 , n26669 , n39807 );
or ( n61974 , n61972 , n61973 );
and ( n61975 , n61974 , n30982 );
and ( n61976 , n29185 , n28587 );
and ( n61977 , n26669 , n39807 );
or ( n61978 , n61976 , n61977 );
and ( n61979 , n61978 , n30989 );
and ( n61980 , n48075 , n28587 );
and ( n61981 , n26669 , n39807 );
or ( n61982 , n61980 , n61981 );
and ( n61983 , n61982 , n31002 );
and ( n61984 , n26669 , n34607 );
or ( n61985 , n61967 , n61971 , n61975 , n61979 , n61983 , n61984 );
and ( n61986 , n61963 , n61985 );
and ( n61987 , n26669 , n24800 );
or ( n61988 , n61986 , n61987 );
and ( n61989 , n61988 , n31008 );
and ( n61990 , n26669 , n10618 );
or ( n61991 , n61989 , n61990 );
buf ( n61992 , n61991 );
buf ( n61993 , n61992 );
buf ( n61994 , n10615 );
not ( n61995 , n34821 );
and ( n61996 , n14605 , n14592 );
and ( n61997 , n55616 , n36348 );
and ( n61998 , n14605 , n43530 );
or ( n61999 , n61997 , n61998 );
and ( n62000 , n61999 , n14562 );
and ( n62001 , n55625 , n36347 );
and ( n62002 , n14605 , n43543 );
or ( n62003 , n62001 , n62002 );
and ( n62004 , n62003 , n14586 );
and ( n62005 , n55634 , n36348 );
and ( n62006 , n14605 , n43556 );
or ( n62007 , n62005 , n62006 );
and ( n62008 , n62007 , n14584 );
and ( n62009 , n55625 , n36347 );
and ( n62010 , n14605 , n43563 );
or ( n62011 , n62009 , n62010 );
and ( n62012 , n62011 , n37835 );
and ( n62013 , n55634 , n36347 );
and ( n62014 , n14605 , n43563 );
or ( n62015 , n62013 , n62014 );
and ( n62016 , n62015 , n37841 );
and ( n62017 , n14603 , n14564 );
and ( n62018 , n14952 , n36347 );
and ( n62019 , n14605 , n43563 );
or ( n62020 , n62018 , n62019 );
and ( n62021 , n62020 , n37847 );
or ( n62022 , n61996 , n62000 , n62004 , n62008 , n62012 , n62016 , n62017 , n62021 );
and ( n62023 , n61995 , n62022 );
and ( n62024 , n14605 , n34821 );
or ( n62025 , n62023 , n62024 );
and ( n62026 , n62025 , n16574 );
and ( n62027 , n14605 , n16576 );
or ( n62028 , n62026 , n62027 );
buf ( n62029 , n62028 );
buf ( n62030 , n62029 );
buf ( n62031 , n10613 );
buf ( n62032 , n10615 );
buf ( n62033 , n10613 );
buf ( n62034 , n10615 );
buf ( n62035 , n10615 );
not ( n62036 , n17451 );
and ( n62037 , n34353 , n21334 );
and ( n62038 , n18511 , n34492 );
or ( n62039 , n62037 , n62038 );
and ( n62040 , n62039 , n21341 );
and ( n62041 , n34363 , n21334 );
and ( n62042 , n18511 , n34492 );
or ( n62043 , n62041 , n62042 );
and ( n62044 , n62043 , n23064 );
and ( n62045 , n34373 , n21334 );
and ( n62046 , n18511 , n34492 );
or ( n62047 , n62045 , n62046 );
and ( n62048 , n62047 , n23825 );
and ( n62049 , n21639 , n21334 );
and ( n62050 , n18511 , n34492 );
or ( n62051 , n62049 , n62050 );
and ( n62052 , n62051 , n23832 );
and ( n62053 , n34383 , n21334 );
and ( n62054 , n18511 , n34492 );
or ( n62055 , n62053 , n62054 );
and ( n62056 , n62055 , n23917 );
and ( n62057 , n18511 , n34526 );
or ( n62058 , n62040 , n62044 , n62048 , n62052 , n62056 , n62057 );
and ( n62059 , n62036 , n62058 );
and ( n62060 , n18511 , n17451 );
or ( n62061 , n62059 , n62060 );
and ( n62062 , n62061 , n23924 );
and ( n62063 , n18511 , n23926 );
or ( n62064 , n62062 , n62063 );
buf ( n62065 , n62064 );
buf ( n62066 , n62065 );
buf ( n62067 , n10615 );
buf ( n62068 , n10615 );
buf ( n62069 , n10615 );
buf ( n62070 , n10615 );
buf ( n62071 , n10613 );
buf ( n62072 , n10613 );
not ( n62073 , n24800 );
and ( n62074 , n26221 , n25222 );
and ( n62075 , n53614 , n28589 );
and ( n62076 , n26221 , n31075 );
or ( n62077 , n62075 , n62076 );
and ( n62078 , n62077 , n28594 );
and ( n62079 , n53624 , n28589 );
and ( n62080 , n26221 , n31075 );
or ( n62081 , n62079 , n62080 );
and ( n62082 , n62081 , n30269 );
and ( n62083 , n53634 , n28589 );
and ( n62084 , n26221 , n31075 );
or ( n62085 , n62083 , n62084 );
and ( n62086 , n62085 , n30982 );
and ( n62087 , n29455 , n28589 );
and ( n62088 , n26221 , n31075 );
or ( n62089 , n62087 , n62088 );
and ( n62090 , n62089 , n30989 );
and ( n62091 , n29455 , n30991 );
and ( n62092 , n53645 , n28589 );
and ( n62093 , n26221 , n31075 );
or ( n62094 , n62092 , n62093 );
and ( n62095 , n62094 , n31002 );
or ( n62096 , n62074 , n62078 , n62082 , n62086 , n62090 , n62091 , n62095 );
and ( n62097 , n62073 , n62096 );
and ( n62098 , n26221 , n24800 );
or ( n62099 , n62097 , n62098 );
and ( n62100 , n62099 , n31008 );
and ( n62101 , n25384 , n10618 );
or ( n62102 , n62100 , n62101 );
buf ( n62103 , n62102 );
buf ( n62104 , n62103 );
buf ( n62105 , n10613 );
buf ( n62106 , n10613 );
buf ( n62107 , n10613 );
not ( n62108 , n34821 );
and ( n62109 , n53772 , n36347 );
and ( n62110 , n13510 , n39408 );
or ( n62111 , n62109 , n62110 );
and ( n62112 , n62111 , n14562 );
and ( n62113 , n53782 , n36348 );
and ( n62114 , n13510 , n39427 );
or ( n62115 , n62113 , n62114 );
and ( n62116 , n62115 , n14586 );
and ( n62117 , n53792 , n36347 );
and ( n62118 , n13510 , n39446 );
or ( n62119 , n62117 , n62118 );
and ( n62120 , n62119 , n14584 );
and ( n62121 , n53782 , n36348 );
and ( n62122 , n13510 , n39453 );
or ( n62123 , n62121 , n62122 );
and ( n62124 , n62123 , n37835 );
and ( n62125 , n53792 , n36348 );
and ( n62126 , n13510 , n39453 );
or ( n62127 , n62125 , n62126 );
and ( n62128 , n62127 , n37841 );
and ( n62129 , n15866 , n36348 );
and ( n62130 , n13510 , n39453 );
or ( n62131 , n62129 , n62130 );
and ( n62132 , n62131 , n37847 );
and ( n62133 , n13510 , n37849 );
or ( n62134 , n62112 , n62116 , n62120 , n62124 , n62128 , n62132 , n62133 );
and ( n62135 , n62108 , n62134 );
and ( n62136 , n13510 , n34821 );
or ( n62137 , n62135 , n62136 );
and ( n62138 , n62137 , n16574 );
and ( n62139 , n13510 , n16576 );
or ( n62140 , n62138 , n62139 );
buf ( n62141 , n62140 );
buf ( n62142 , n62141 );
buf ( n62143 , n10613 );
buf ( n62144 , n10615 );
buf ( n62145 , n10615 );
not ( n62146 , n34821 );
and ( n62147 , n13349 , n14592 );
and ( n62148 , n43688 , n36348 );
and ( n62149 , n13349 , n43530 );
or ( n62150 , n62148 , n62149 );
and ( n62151 , n62150 , n14562 );
and ( n62152 , n43700 , n36347 );
and ( n62153 , n13349 , n43543 );
or ( n62154 , n62152 , n62153 );
and ( n62155 , n62154 , n14586 );
and ( n62156 , n43712 , n36348 );
and ( n62157 , n13349 , n43556 );
or ( n62158 , n62156 , n62157 );
and ( n62159 , n62158 , n14584 );
and ( n62160 , n43700 , n36347 );
and ( n62161 , n13349 , n43563 );
or ( n62162 , n62160 , n62161 );
and ( n62163 , n62162 , n37835 );
and ( n62164 , n43712 , n36347 );
and ( n62165 , n13349 , n43563 );
or ( n62166 , n62164 , n62165 );
and ( n62167 , n62166 , n37841 );
and ( n62168 , n13347 , n14564 );
and ( n62169 , n15603 , n36347 );
and ( n62170 , n13349 , n43563 );
or ( n62171 , n62169 , n62170 );
and ( n62172 , n62171 , n37847 );
or ( n62173 , n62147 , n62151 , n62155 , n62159 , n62163 , n62167 , n62168 , n62172 );
and ( n62174 , n62146 , n62173 );
and ( n62175 , n13349 , n34821 );
or ( n62176 , n62174 , n62175 );
and ( n62177 , n62176 , n16574 );
and ( n62178 , n13349 , n16576 );
or ( n62179 , n62177 , n62178 );
buf ( n62180 , n62179 );
buf ( n62181 , n62180 );
buf ( n62182 , n10613 );
not ( n62183 , n24800 );
and ( n62184 , n26631 , n25222 );
and ( n62185 , n54833 , n28583 );
and ( n62186 , n26631 , n28591 );
or ( n62187 , n62185 , n62186 );
and ( n62188 , n62187 , n28594 );
and ( n62189 , n54843 , n28583 );
and ( n62190 , n26631 , n28591 );
or ( n62191 , n62189 , n62190 );
and ( n62192 , n62191 , n30269 );
and ( n62193 , n54853 , n28583 );
and ( n62194 , n26631 , n28591 );
or ( n62195 , n62193 , n62194 );
and ( n62196 , n62195 , n30982 );
and ( n62197 , n29198 , n28583 );
and ( n62198 , n26631 , n28591 );
or ( n62199 , n62197 , n62198 );
and ( n62200 , n62199 , n30989 );
and ( n62201 , n26629 , n30991 );
and ( n62202 , n54863 , n28583 );
and ( n62203 , n26631 , n28591 );
or ( n62204 , n62202 , n62203 );
and ( n62205 , n62204 , n31002 );
or ( n62206 , n62184 , n62188 , n62192 , n62196 , n62200 , n62201 , n62205 );
and ( n62207 , n62183 , n62206 );
and ( n62208 , n26631 , n24800 );
or ( n62209 , n62207 , n62208 );
and ( n62210 , n62209 , n31008 );
and ( n62211 , n26631 , n10618 );
or ( n62212 , n62210 , n62211 );
buf ( n62213 , n62212 );
buf ( n62214 , n62213 );
not ( n62215 , n17451 );
and ( n62216 , n19179 , n17873 );
and ( n62217 , n46077 , n21336 );
and ( n62218 , n19179 , n42682 );
or ( n62219 , n62217 , n62218 );
and ( n62220 , n62219 , n21341 );
and ( n62221 , n46087 , n21336 );
and ( n62222 , n19179 , n42682 );
or ( n62223 , n62221 , n62222 );
and ( n62224 , n62223 , n23064 );
and ( n62225 , n46097 , n21336 );
and ( n62226 , n19179 , n42682 );
or ( n62227 , n62225 , n62226 );
and ( n62228 , n62227 , n23825 );
and ( n62229 , n21984 , n21336 );
and ( n62230 , n19179 , n42682 );
or ( n62231 , n62229 , n62230 );
and ( n62232 , n62231 , n23832 );
and ( n62233 , n21984 , n23834 );
and ( n62234 , n46108 , n21336 );
and ( n62235 , n19179 , n42682 );
or ( n62236 , n62234 , n62235 );
and ( n62237 , n62236 , n23917 );
or ( n62238 , n62216 , n62220 , n62224 , n62228 , n62232 , n62233 , n62237 );
and ( n62239 , n62215 , n62238 );
and ( n62240 , n19179 , n17451 );
or ( n62241 , n62239 , n62240 );
and ( n62242 , n62241 , n23924 );
and ( n62243 , n18170 , n23926 );
or ( n62244 , n62242 , n62243 );
buf ( n62245 , n62244 );
buf ( n62246 , n62245 );
not ( n62247 , n17451 );
and ( n62248 , n39576 , n21333 );
and ( n62249 , n19319 , n34758 );
or ( n62250 , n62248 , n62249 );
and ( n62251 , n62250 , n21341 );
and ( n62252 , n39586 , n21333 );
and ( n62253 , n19319 , n34758 );
or ( n62254 , n62252 , n62253 );
and ( n62255 , n62254 , n23064 );
and ( n62256 , n39596 , n21333 );
and ( n62257 , n19319 , n34758 );
or ( n62258 , n62256 , n62257 );
and ( n62259 , n62258 , n23825 );
and ( n62260 , n21932 , n21333 );
and ( n62261 , n19319 , n34758 );
or ( n62262 , n62260 , n62261 );
and ( n62263 , n62262 , n23832 );
and ( n62264 , n39606 , n21333 );
and ( n62265 , n19319 , n34758 );
or ( n62266 , n62264 , n62265 );
and ( n62267 , n62266 , n23917 );
and ( n62268 , n19319 , n34526 );
or ( n62269 , n62251 , n62255 , n62259 , n62263 , n62267 , n62268 );
and ( n62270 , n62247 , n62269 );
and ( n62271 , n19319 , n17451 );
or ( n62272 , n62270 , n62271 );
and ( n62273 , n62272 , n23924 );
and ( n62274 , n19319 , n23926 );
or ( n62275 , n62273 , n62274 );
buf ( n62276 , n62275 );
buf ( n62277 , n62276 );
buf ( n62278 , n10613 );
not ( n62279 , n17451 );
and ( n62280 , n18637 , n17873 );
and ( n62281 , n47363 , n21330 );
and ( n62282 , n18637 , n21338 );
or ( n62283 , n62281 , n62282 );
and ( n62284 , n62283 , n21341 );
and ( n62285 , n47373 , n21330 );
and ( n62286 , n18637 , n21338 );
or ( n62287 , n62285 , n62286 );
and ( n62288 , n62287 , n23064 );
and ( n62289 , n47383 , n21330 );
and ( n62290 , n18637 , n21338 );
or ( n62291 , n62289 , n62290 );
and ( n62292 , n62291 , n23825 );
and ( n62293 , n22342 , n21330 );
and ( n62294 , n18637 , n21338 );
or ( n62295 , n62293 , n62294 );
and ( n62296 , n62295 , n23832 );
and ( n62297 , n18635 , n23834 );
and ( n62298 , n47394 , n21330 );
and ( n62299 , n18637 , n21338 );
or ( n62300 , n62298 , n62299 );
and ( n62301 , n62300 , n23917 );
or ( n62302 , n62280 , n62284 , n62288 , n62292 , n62296 , n62297 , n62301 );
and ( n62303 , n62279 , n62302 );
and ( n62304 , n18637 , n17451 );
or ( n62305 , n62303 , n62304 );
and ( n62306 , n62305 , n23924 );
and ( n62307 , n18637 , n23926 );
or ( n62308 , n62306 , n62307 );
buf ( n62309 , n62308 );
buf ( n62310 , n62309 );
buf ( n62311 , n10613 );
not ( n62312 , n17451 );
and ( n62313 , n47430 , n21334 );
and ( n62314 , n19253 , n34492 );
or ( n62315 , n62313 , n62314 );
and ( n62316 , n62315 , n21341 );
and ( n62317 , n47440 , n21334 );
and ( n62318 , n19253 , n34492 );
or ( n62319 , n62317 , n62318 );
and ( n62320 , n62319 , n23064 );
and ( n62321 , n47450 , n21334 );
and ( n62322 , n19253 , n34492 );
or ( n62323 , n62321 , n62322 );
and ( n62324 , n62323 , n23825 );
and ( n62325 , n21958 , n21334 );
and ( n62326 , n19253 , n34492 );
or ( n62327 , n62325 , n62326 );
and ( n62328 , n62327 , n23832 );
and ( n62329 , n47461 , n21334 );
and ( n62330 , n19253 , n34492 );
or ( n62331 , n62329 , n62330 );
and ( n62332 , n62331 , n23917 );
and ( n62333 , n19253 , n34526 );
or ( n62334 , n62316 , n62320 , n62324 , n62328 , n62332 , n62333 );
and ( n62335 , n62312 , n62334 );
and ( n62336 , n19253 , n17451 );
or ( n62337 , n62335 , n62336 );
and ( n62338 , n62337 , n23924 );
and ( n62339 , n19253 , n23926 );
or ( n62340 , n62338 , n62339 );
buf ( n62341 , n62340 );
buf ( n62342 , n62341 );
buf ( n62343 , n10615 );
buf ( n62344 , n10615 );
not ( n62345 , n34821 );
and ( n62346 , n46418 , n36347 );
and ( n62347 , n13183 , n39408 );
or ( n62348 , n62346 , n62347 );
and ( n62349 , n62348 , n14562 );
and ( n62350 , n46436 , n36348 );
and ( n62351 , n13183 , n39427 );
or ( n62352 , n62350 , n62351 );
and ( n62353 , n62352 , n14586 );
and ( n62354 , n46454 , n36347 );
and ( n62355 , n13183 , n39446 );
or ( n62356 , n62354 , n62355 );
and ( n62357 , n62356 , n14584 );
and ( n62358 , n46436 , n36348 );
and ( n62359 , n13183 , n39453 );
or ( n62360 , n62358 , n62359 );
and ( n62361 , n62360 , n37835 );
and ( n62362 , n46454 , n36348 );
and ( n62363 , n13183 , n39453 );
or ( n62364 , n62362 , n62363 );
and ( n62365 , n62364 , n37841 );
and ( n62366 , n15022 , n36348 );
and ( n62367 , n13183 , n39453 );
or ( n62368 , n62366 , n62367 );
and ( n62369 , n62368 , n37847 );
and ( n62370 , n13183 , n37849 );
or ( n62371 , n62349 , n62353 , n62357 , n62361 , n62365 , n62369 , n62370 );
and ( n62372 , n62345 , n62371 );
and ( n62373 , n13183 , n34821 );
or ( n62374 , n62372 , n62373 );
and ( n62375 , n62374 , n16574 );
and ( n62376 , n13183 , n16576 );
or ( n62377 , n62375 , n62376 );
buf ( n62378 , n62377 );
buf ( n62379 , n62378 );
not ( n62380 , n34821 );
and ( n62381 , n13203 , n14592 );
and ( n62382 , n47932 , n36350 );
and ( n62383 , n13203 , n43691 );
or ( n62384 , n62382 , n62383 );
and ( n62385 , n62384 , n14562 );
and ( n62386 , n47942 , n36350 );
and ( n62387 , n13203 , n43703 );
or ( n62388 , n62386 , n62387 );
and ( n62389 , n62388 , n14586 );
and ( n62390 , n47952 , n36345 );
and ( n62391 , n13203 , n43715 );
or ( n62392 , n62390 , n62391 );
and ( n62393 , n62392 , n14584 );
and ( n62394 , n47942 , n36345 );
and ( n62395 , n13203 , n43721 );
or ( n62396 , n62394 , n62395 );
and ( n62397 , n62396 , n37835 );
and ( n62398 , n47952 , n36345 );
and ( n62399 , n13203 , n43721 );
or ( n62400 , n62398 , n62399 );
and ( n62401 , n62400 , n37841 );
and ( n62402 , n15052 , n14564 );
and ( n62403 , n15052 , n36345 );
and ( n62404 , n13203 , n43721 );
or ( n62405 , n62403 , n62404 );
and ( n62406 , n62405 , n37847 );
or ( n62407 , n62381 , n62385 , n62389 , n62393 , n62397 , n62401 , n62402 , n62406 );
and ( n62408 , n62380 , n62407 );
and ( n62409 , n13203 , n34821 );
or ( n62410 , n62408 , n62409 );
and ( n62411 , n62410 , n16574 );
and ( n62412 , n12261 , n16576 );
or ( n62413 , n62411 , n62412 );
buf ( n62414 , n62413 );
buf ( n62415 , n62414 );
not ( n62416 , n24800 );
and ( n62417 , n26597 , n25222 );
and ( n62418 , n42864 , n28583 );
and ( n62419 , n26597 , n28591 );
or ( n62420 , n62418 , n62419 );
and ( n62421 , n62420 , n28594 );
and ( n62422 , n42884 , n28583 );
and ( n62423 , n26597 , n28591 );
or ( n62424 , n62422 , n62423 );
and ( n62425 , n62424 , n30269 );
and ( n62426 , n42904 , n28583 );
and ( n62427 , n26597 , n28591 );
or ( n62428 , n62426 , n62427 );
and ( n62429 , n62428 , n30982 );
and ( n62430 , n29211 , n28583 );
and ( n62431 , n26597 , n28591 );
or ( n62432 , n62430 , n62431 );
and ( n62433 , n62432 , n30989 );
and ( n62434 , n26595 , n30991 );
and ( n62435 , n42929 , n28583 );
and ( n62436 , n26597 , n28591 );
or ( n62437 , n62435 , n62436 );
and ( n62438 , n62437 , n31002 );
or ( n62439 , n62417 , n62421 , n62425 , n62429 , n62433 , n62434 , n62438 );
and ( n62440 , n62416 , n62439 );
and ( n62441 , n26597 , n24800 );
or ( n62442 , n62440 , n62441 );
and ( n62443 , n62442 , n31008 );
and ( n62444 , n26597 , n10618 );
or ( n62445 , n62443 , n62444 );
buf ( n62446 , n62445 );
buf ( n62447 , n62446 );
not ( n62448 , n24800 );
and ( n62449 , n26357 , n25222 );
and ( n62450 , n51562 , n28589 );
and ( n62451 , n26357 , n31075 );
or ( n62452 , n62450 , n62451 );
and ( n62453 , n62452 , n28594 );
and ( n62454 , n51572 , n28589 );
and ( n62455 , n26357 , n31075 );
or ( n62456 , n62454 , n62455 );
and ( n62457 , n62456 , n30269 );
and ( n62458 , n51582 , n28589 );
and ( n62459 , n26357 , n31075 );
or ( n62460 , n62458 , n62459 );
and ( n62461 , n62460 , n30982 );
and ( n62462 , n29375 , n28589 );
and ( n62463 , n26357 , n31075 );
or ( n62464 , n62462 , n62463 );
and ( n62465 , n62464 , n30989 );
and ( n62466 , n29375 , n30991 );
or ( n62467 , n51592 , n28589 );
and ( n62468 , n26357 , n31075 );
or ( n62469 , n62467 , n62468 );
and ( n62470 , n62469 , n31002 );
or ( n62471 , n62449 , n62453 , n62457 , n62461 , n62465 , n62466 , n62470 );
and ( n62472 , n62448 , n62471 );
and ( n62473 , n26357 , n24800 );
or ( n62474 , n62472 , n62473 );
and ( n62475 , n62474 , n31008 );
and ( n62476 , n25444 , n10618 );
or ( n62477 , n62475 , n62476 );
buf ( n62478 , n62477 );
buf ( n62479 , n62478 );
buf ( n62480 , n10613 );
buf ( n62481 , n10615 );
buf ( n62482 , n10613 );
buf ( n62483 , n10615 );
buf ( n62484 , n10613 );
buf ( n62485 , n10615 );
buf ( n62486 , n10615 );
buf ( n62487 , n10613 );
buf ( n62488 , n10613 );
buf ( n62489 , n10615 );
buf ( n62490 , n10613 );
buf ( n62491 , n10613 );
not ( n62492 , n24800 );
and ( n62493 , n26427 , n25222 );
and ( n62494 , n39662 , n28583 );
and ( n62495 , n26427 , n28591 );
or ( n62496 , n62494 , n62495 );
and ( n62497 , n62496 , n28594 );
and ( n62498 , n39678 , n28583 );
and ( n62499 , n26427 , n28591 );
or ( n62500 , n62498 , n62499 );
and ( n62501 , n62500 , n30269 );
and ( n62502 , n39694 , n28583 );
and ( n62503 , n26427 , n28591 );
or ( n62504 , n62502 , n62503 );
and ( n62505 , n62504 , n30982 );
and ( n62506 , n29335 , n28583 );
and ( n62507 , n26427 , n28591 );
or ( n62508 , n62506 , n62507 );
and ( n62509 , n62508 , n30989 );
and ( n62510 , n26425 , n30991 );
and ( n62511 , n39713 , n28583 );
and ( n62512 , n26427 , n28591 );
or ( n62513 , n62511 , n62512 );
and ( n62514 , n62513 , n31002 );
or ( n62515 , n62493 , n62497 , n62501 , n62505 , n62509 , n62510 , n62514 );
and ( n62516 , n62492 , n62515 );
and ( n62517 , n26427 , n24800 );
or ( n62518 , n62516 , n62517 );
and ( n62519 , n62518 , n31008 );
and ( n62520 , n26427 , n10618 );
or ( n62521 , n62519 , n62520 );
buf ( n62522 , n62521 );
buf ( n62523 , n62522 );
not ( n62524 , n24800 );
and ( n62525 , n26325 , n25222 );
and ( n62526 , n34656 , n28583 );
and ( n62527 , n26325 , n28591 );
or ( n62528 , n62526 , n62527 );
and ( n62529 , n62528 , n28594 );
and ( n62530 , n34674 , n28583 );
and ( n62531 , n26325 , n28591 );
or ( n62532 , n62530 , n62531 );
and ( n62533 , n62532 , n30269 );
and ( n62534 , n34692 , n28583 );
and ( n62535 , n26325 , n28591 );
or ( n62536 , n62534 , n62535 );
and ( n62537 , n62536 , n30982 );
and ( n62538 , n29395 , n28583 );
and ( n62539 , n26325 , n28591 );
or ( n62540 , n62538 , n62539 );
and ( n62541 , n62540 , n30989 );
and ( n62542 , n26323 , n30991 );
and ( n62543 , n34714 , n28583 );
and ( n62544 , n26325 , n28591 );
or ( n62545 , n62543 , n62544 );
and ( n62546 , n62545 , n31002 );
or ( n62547 , n62525 , n62529 , n62533 , n62537 , n62541 , n62542 , n62546 );
and ( n62548 , n62524 , n62547 );
and ( n62549 , n26325 , n24800 );
or ( n62550 , n62548 , n62549 );
and ( n62551 , n62550 , n31008 );
and ( n62552 , n26325 , n10618 );
or ( n62553 , n62551 , n62552 );
buf ( n62554 , n62553 );
buf ( n62555 , n62554 );
buf ( n62556 , n10615 );
buf ( n62557 , n10615 );
buf ( n62558 , n10613 );
buf ( n62559 , n10613 );
buf ( n62560 , n10615 );
buf ( n62561 , n10615 );
not ( n62562 , n17451 );
and ( n62563 , n18602 , n17873 );
and ( n62564 , n48952 , n21336 );
and ( n62565 , n18602 , n42682 );
or ( n62566 , n62564 , n62565 );
and ( n62567 , n62566 , n21341 );
and ( n62568 , n48962 , n21336 );
and ( n62569 , n18602 , n42682 );
or ( n62570 , n62568 , n62569 );
and ( n62571 , n62570 , n23064 );
and ( n62572 , n48972 , n21336 );
and ( n62573 , n18602 , n42682 );
or ( n62574 , n62572 , n62573 );
and ( n62575 , n62574 , n23825 );
and ( n62576 , n22362 , n21336 );
and ( n62577 , n18602 , n42682 );
or ( n62578 , n62576 , n62577 );
and ( n62579 , n62578 , n23832 );
and ( n62580 , n22362 , n23834 );
and ( n62581 , n48982 , n21336 );
and ( n62582 , n18602 , n42682 );
or ( n62583 , n62581 , n62582 );
and ( n62584 , n62583 , n23917 );
or ( n62585 , n62563 , n62567 , n62571 , n62575 , n62579 , n62580 , n62584 );
and ( n62586 , n62562 , n62585 );
and ( n62587 , n18602 , n17451 );
or ( n62588 , n62586 , n62587 );
and ( n62589 , n62588 , n23924 );
and ( n62590 , n17915 , n23926 );
or ( n62591 , n62589 , n62590 );
buf ( n62592 , n62591 );
buf ( n62593 , n62592 );
and ( n62594 , n24238 , n31008 );
and ( n62595 , n29626 , n10618 );
or ( n62596 , n62594 , n62595 );
buf ( n62597 , n62596 );
buf ( n62598 , n62597 );
buf ( n62599 , n10613 );
buf ( n62600 , n10613 );
buf ( n62601 , n10615 );
and ( n62602 , n17008 , n23924 );
and ( n62603 , n21904 , n23926 );
or ( n62604 , n62602 , n62603 );
buf ( n62605 , n62604 );
buf ( n62606 , n62605 );
buf ( n62607 , n10615 );
buf ( n62608 , n10613 );
buf ( n62609 , n10613 );
buf ( n62610 , n10615 );
not ( n62611 , n24800 );
and ( n62612 , n45874 , n28587 );
and ( n62613 , n26567 , n39807 );
or ( n62614 , n62612 , n62613 );
and ( n62615 , n62614 , n28594 );
and ( n62616 , n45884 , n28587 );
and ( n62617 , n26567 , n39807 );
or ( n62618 , n62616 , n62617 );
and ( n62619 , n62618 , n30269 );
and ( n62620 , n45894 , n28587 );
and ( n62621 , n26567 , n39807 );
or ( n62622 , n62620 , n62621 );
and ( n62623 , n62622 , n30982 );
and ( n62624 , n29224 , n28587 );
and ( n62625 , n26567 , n39807 );
or ( n62626 , n62624 , n62625 );
and ( n62627 , n62626 , n30989 );
and ( n62628 , n45905 , n28587 );
and ( n62629 , n26567 , n39807 );
or ( n62630 , n62628 , n62629 );
and ( n62631 , n62630 , n31002 );
and ( n62632 , n26567 , n34607 );
or ( n62633 , n62615 , n62619 , n62623 , n62627 , n62631 , n62632 );
and ( n62634 , n62611 , n62633 );
and ( n62635 , n26567 , n24800 );
or ( n62636 , n62634 , n62635 );
and ( n62637 , n62636 , n31008 );
and ( n62638 , n26567 , n10618 );
or ( n62639 , n62637 , n62638 );
buf ( n62640 , n62639 );
buf ( n62641 , n62640 );
buf ( n62642 , n10615 );
buf ( n62643 , n10613 );
not ( n62644 , n17451 );
and ( n62645 , n19111 , n17873 );
and ( n62646 , n39499 , n21336 );
and ( n62647 , n19111 , n42682 );
or ( n62648 , n62646 , n62647 );
and ( n62649 , n62648 , n21341 );
and ( n62650 , n39509 , n21336 );
and ( n62651 , n19111 , n42682 );
or ( n62652 , n62650 , n62651 );
and ( n62653 , n62652 , n23064 );
and ( n62654 , n39519 , n21336 );
and ( n62655 , n19111 , n42682 );
or ( n62656 , n62654 , n62655 );
and ( n62657 , n62656 , n23825 );
and ( n62658 , n22062 , n21336 );
and ( n62659 , n19111 , n42682 );
or ( n62660 , n62658 , n62659 );
and ( n62661 , n62660 , n23832 );
and ( n62662 , n22062 , n23834 );
and ( n62663 , n39529 , n21336 );
and ( n62664 , n19111 , n42682 );
or ( n62665 , n62663 , n62664 );
and ( n62666 , n62665 , n23917 );
or ( n62667 , n62645 , n62649 , n62653 , n62657 , n62661 , n62662 , n62666 );
and ( n62668 , n62644 , n62667 );
and ( n62669 , n19111 , n17451 );
or ( n62670 , n62668 , n62669 );
and ( n62671 , n62670 , n23924 );
and ( n62672 , n18140 , n23926 );
or ( n62673 , n62671 , n62672 );
buf ( n62674 , n62673 );
buf ( n62675 , n62674 );
buf ( n62676 , n10613 );
buf ( n62677 , n10615 );
buf ( n62678 , n10613 );
buf ( n62679 , n10613 );
not ( n62680 , n24511 );
not ( n62681 , n24799 );
and ( n62682 , n10705 , n40154 );
not ( n62683 , n40632 );
and ( n62684 , n62683 , n40407 );
xor ( n62685 , n40644 , n40656 );
and ( n62686 , n62685 , n40632 );
or ( n62687 , n62684 , n62686 );
buf ( n62688 , n62687 );
and ( n62689 , n62688 , n27046 );
not ( n62690 , n41147 );
and ( n62691 , n62690 , n40922 );
xor ( n62692 , n41159 , n41171 );
and ( n62693 , n62692 , n41147 );
or ( n62694 , n62691 , n62693 );
buf ( n62695 , n62694 );
and ( n62696 , n62695 , n27049 );
and ( n62697 , n29553 , n28506 );
and ( n62698 , n10705 , n28508 );
or ( n62699 , n62689 , n62696 , n62697 , n62698 );
and ( n62700 , n62699 , n41199 );
or ( n62701 , n62682 , n62700 );
and ( n62702 , n62681 , n62701 );
xor ( n62703 , n41660 , n41668 );
xor ( n62704 , n62703 , n41779 );
buf ( n62705 , n62704 );
and ( n62706 , n62705 , n27046 );
xor ( n62707 , n42204 , n42205 );
xor ( n62708 , n62707 , n42275 );
buf ( n62709 , n62708 );
and ( n62710 , n62709 , n27049 );
and ( n62711 , n29553 , n42306 );
or ( n62712 , n62706 , n62710 , n62711 );
buf ( n62713 , n62712 );
and ( n62714 , C1 , n62713 );
or ( n62715 , n62714 , C0 );
buf ( n62716 , n62715 );
not ( n62717 , n62716 );
buf ( n62718 , n62717 );
buf ( n62719 , n62718 );
not ( n62720 , n62719 );
and ( n62721 , C1 , n62720 );
or ( n62722 , n62721 , C0 );
buf ( n62723 , n62722 );
and ( n62724 , n62723 , n24799 );
or ( n62725 , n62702 , n62724 );
and ( n62726 , n62680 , n62725 );
and ( n62727 , n62699 , n24511 );
or ( n62728 , n62726 , n62727 );
and ( n62729 , n62728 , n31008 );
not ( n62730 , n42601 );
and ( n62731 , n62730 , n42415 );
xor ( n62732 , n42613 , n42625 );
and ( n62733 , n62732 , n42601 );
or ( n62734 , n62731 , n62733 );
buf ( n62735 , n62734 );
and ( n62736 , n62735 , n10618 );
or ( n62737 , n62729 , n62736 );
buf ( n62738 , n62737 );
buf ( n62739 , n62738 );
buf ( n62740 , n10615 );
not ( n62741 , n34821 );
and ( n62742 , n57357 , n36345 );
and ( n62743 , n13257 , n36352 );
or ( n62744 , n62742 , n62743 );
and ( n62745 , n62744 , n14562 );
and ( n62746 , n57367 , n36345 );
and ( n62747 , n13257 , n37073 );
or ( n62748 , n62746 , n62747 );
and ( n62749 , n62748 , n14586 );
and ( n62750 , n57377 , n36350 );
and ( n62751 , n13257 , n37825 );
or ( n62752 , n62750 , n62751 );
and ( n62753 , n62752 , n14584 );
and ( n62754 , n57367 , n36350 );
and ( n62755 , n13257 , n37831 );
or ( n62756 , n62754 , n62755 );
and ( n62757 , n62756 , n37835 );
and ( n62758 , n57377 , n36350 );
and ( n62759 , n13257 , n37831 );
or ( n62760 , n62758 , n62759 );
and ( n62761 , n62760 , n37841 );
and ( n62762 , n15112 , n36350 );
and ( n62763 , n13257 , n37831 );
or ( n62764 , n62762 , n62763 );
and ( n62765 , n62764 , n37847 );
and ( n62766 , n13257 , n37849 );
or ( n62767 , n62745 , n62749 , n62753 , n62757 , n62761 , n62765 , n62766 );
and ( n62768 , n62741 , n62767 );
and ( n62769 , n13257 , n34821 );
or ( n62770 , n62768 , n62769 );
and ( n62771 , n62770 , n16574 );
and ( n62772 , n13257 , n16576 );
or ( n62773 , n62771 , n62772 );
buf ( n62774 , n62773 );
buf ( n62775 , n62774 );
buf ( n62776 , n10613 );
buf ( n62777 , n10615 );
buf ( n62778 , n10615 );
buf ( n62779 , n10613 );
not ( n62780 , n17162 );
not ( n62781 , n17450 );
and ( n62782 , n10718 , n37947 );
not ( n62783 , n38425 );
and ( n62784 , n62783 , n38149 );
xor ( n62785 , n38437 , n38443 );
and ( n62786 , n62785 , n38425 );
or ( n62787 , n62784 , n62786 );
buf ( n62788 , n62787 );
and ( n62789 , n62788 , n19745 );
not ( n62790 , n38934 );
and ( n62791 , n62790 , n38658 );
xor ( n62792 , n38946 , n38952 );
and ( n62793 , n62792 , n38934 );
or ( n62794 , n62791 , n62793 );
buf ( n62795 , n62794 );
and ( n62796 , n62795 , n19748 );
and ( n62797 , n22360 , n21253 );
and ( n62798 , n10718 , n21255 );
or ( n62799 , n62789 , n62796 , n62797 , n62798 );
and ( n62800 , n62799 , n38980 );
or ( n62801 , n62782 , n62800 );
and ( n62802 , n62781 , n62801 );
or ( n62803 , n62802 , C0 );
and ( n62804 , n62780 , n62803 );
and ( n62805 , n62799 , n17162 );
or ( n62806 , n62804 , n62805 );
and ( n62807 , n62806 , n23924 );
not ( n62808 , n39264 );
and ( n62809 , n62808 , n39036 );
xor ( n62810 , n39276 , n39282 );
and ( n62811 , n62810 , n39264 );
or ( n62812 , n62809 , n62811 );
buf ( n62813 , n62812 );
and ( n62814 , n62813 , n23926 );
or ( n62815 , n62807 , n62814 );
buf ( n62816 , n62815 );
buf ( n62817 , n62816 );
not ( n62818 , n17451 );
and ( n62819 , n58841 , n21334 );
and ( n62820 , n19015 , n34492 );
or ( n62821 , n62819 , n62820 );
and ( n62822 , n62821 , n21341 );
and ( n62823 , n58851 , n21334 );
and ( n62824 , n19015 , n34492 );
or ( n62825 , n62823 , n62824 );
and ( n62826 , n62825 , n23064 );
and ( n62827 , n58861 , n21334 );
and ( n62828 , n19015 , n34492 );
or ( n62829 , n62827 , n62828 );
and ( n62830 , n62829 , n23825 );
and ( n62831 , n22122 , n21334 );
and ( n62832 , n19015 , n34492 );
or ( n62833 , n62831 , n62832 );
and ( n62834 , n62833 , n23832 );
and ( n62835 , n58872 , n21334 );
and ( n62836 , n19015 , n34492 );
or ( n62837 , n62835 , n62836 );
and ( n62838 , n62837 , n23917 );
and ( n62839 , n19015 , n34526 );
or ( n62840 , n62822 , n62826 , n62830 , n62834 , n62838 , n62839 );
and ( n62841 , n62818 , n62840 );
and ( n62842 , n19015 , n17451 );
or ( n62843 , n62841 , n62842 );
and ( n62844 , n62843 , n23924 );
and ( n62845 , n19015 , n23926 );
or ( n62846 , n62844 , n62845 );
buf ( n62847 , n62846 );
buf ( n62848 , n62847 );
buf ( n62849 , n10613 );
buf ( n62850 , n10613 );
buf ( n62851 , n10613 );
buf ( n62852 , n10615 );
buf ( n62853 , n10615 );
not ( n62854 , n34804 );
and ( n62855 , n62854 , n26059 );
and ( n62856 , n14797 , n34804 );
or ( n62857 , n62855 , n62856 );
and ( n62858 , n62857 , n31008 );
and ( n62859 , n14797 , n10618 );
or ( n62860 , n62858 , n62859 );
buf ( n62861 , n62860 );
buf ( n62862 , n62861 );
not ( n62863 , n11333 );
and ( n62864 , n62863 , n11142 );
xnor ( n62865 , n11343 , n11359 );
and ( n62866 , n62865 , n11333 );
or ( n62867 , n62864 , n62866 );
buf ( n62868 , n62867 );
buf ( n62869 , n62868 );
buf ( n62870 , n10615 );
not ( n62871 , n11954 );
not ( n62872 , n12243 );
and ( n62873 , n10813 , n31187 );
not ( n62874 , n31697 );
and ( n62875 , n62874 , n31659 );
xor ( n62876 , n56879 , n56890 );
and ( n62877 , n62876 , n31697 );
or ( n62878 , n62875 , n62877 );
buf ( n62879 , n62878 );
and ( n62880 , n62879 , n14140 );
not ( n62881 , n32214 );
and ( n62882 , n62881 , n32176 );
xor ( n62883 , n56902 , n56913 );
and ( n62884 , n62883 , n32214 );
or ( n62885 , n62882 , n62884 );
buf ( n62886 , n62885 );
and ( n62887 , n62886 , n14137 );
and ( n62888 , n15491 , n14143 );
and ( n62889 , n10813 , n14141 );
or ( n62890 , n62880 , n62887 , n62888 , n62889 );
and ( n62891 , n62890 , n32236 );
or ( n62892 , n62873 , n62891 );
and ( n62893 , n62872 , n62892 );
not ( n62894 , n34038 );
and ( n62895 , n62894 , n33986 );
xor ( n62896 , n56931 , n56942 );
and ( n62897 , n62896 , n34038 );
or ( n62898 , n62895 , n62897 );
buf ( n62899 , n62898 );
and ( n62900 , n62899 , n12243 );
or ( n62901 , n62893 , n62900 );
and ( n62902 , n62871 , n62901 );
and ( n62903 , n62890 , n11954 );
or ( n62904 , n62902 , n62903 );
and ( n62905 , n62904 , n16574 );
not ( n62906 , n34327 );
and ( n62907 , n62906 , n34295 );
xor ( n62908 , n56959 , n56970 );
and ( n62909 , n62908 , n34327 );
or ( n62910 , n62907 , n62909 );
buf ( n62911 , n62910 );
and ( n62912 , n62911 , n16576 );
or ( n62913 , n62905 , n62912 );
buf ( n62914 , n62913 );
buf ( n62915 , n62914 );
buf ( n62916 , n10613 );
buf ( n62917 , n10615 );
not ( n62918 , n11954 );
not ( n62919 , n12243 );
and ( n62920 , n10885 , n31187 );
not ( n62921 , n31697 );
and ( n62922 , n62921 , n31506 );
xor ( n62923 , n50358 , n50373 );
and ( n62924 , n62923 , n31697 );
or ( n62925 , n62922 , n62924 );
buf ( n62926 , n62925 );
and ( n62927 , n62926 , n14140 );
not ( n62928 , n32214 );
and ( n62929 , n62928 , n32023 );
xor ( n62930 , n50385 , n50400 );
and ( n62931 , n62930 , n32214 );
or ( n62932 , n62929 , n62931 );
buf ( n62933 , n62932 );
and ( n62934 , n62933 , n14137 );
and ( n62935 , n15689 , n14143 );
and ( n62936 , n10885 , n14141 );
or ( n62937 , n62927 , n62934 , n62935 , n62936 );
and ( n62938 , n62937 , n32236 );
or ( n62939 , n62920 , n62938 );
and ( n62940 , n62919 , n62939 );
not ( n62941 , n34038 );
and ( n62942 , n62941 , n33770 );
xor ( n62943 , n50418 , n50433 );
and ( n62944 , n62943 , n34038 );
or ( n62945 , n62942 , n62944 );
buf ( n62946 , n62945 );
and ( n62947 , n62946 , n12243 );
or ( n62948 , n62940 , n62947 );
and ( n62949 , n62918 , n62948 );
and ( n62950 , n62937 , n11954 );
or ( n62951 , n62949 , n62950 );
and ( n62952 , n62951 , n16574 );
not ( n62953 , n34327 );
and ( n62954 , n62953 , n34169 );
xor ( n62955 , n50450 , n50465 );
and ( n62956 , n62955 , n34327 );
or ( n62957 , n62954 , n62956 );
buf ( n62958 , n62957 );
and ( n62959 , n62958 , n16576 );
or ( n62960 , n62952 , n62959 );
buf ( n62961 , n62960 );
buf ( n62962 , n62961 );
buf ( n62963 , n10613 );
buf ( n62964 , n10613 );
buf ( n62965 , n10613 );
buf ( n62966 , n10613 );
buf ( n62967 , n10613 );
buf ( n62968 , n10613 );
buf ( n62969 , n10615 );
not ( n62970 , n17451 );
and ( n62971 , n45354 , n21334 );
and ( n62972 , n19456 , n34492 );
or ( n62973 , n62971 , n62972 );
and ( n62974 , n62973 , n21341 );
and ( n62975 , n45364 , n21334 );
and ( n62976 , n19456 , n34492 );
or ( n62977 , n62975 , n62976 );
and ( n62978 , n62977 , n23064 );
and ( n62979 , n45374 , n21334 );
and ( n62980 , n19456 , n34492 );
or ( n62981 , n62979 , n62980 );
and ( n62982 , n62981 , n23825 );
and ( n62983 , n21880 , n21334 );
and ( n62984 , n19456 , n34492 );
or ( n62985 , n62983 , n62984 );
and ( n62986 , n62985 , n23832 );
and ( n62987 , n45384 , n21334 );
and ( n62988 , n19456 , n34492 );
or ( n62989 , n62987 , n62988 );
and ( n62990 , n62989 , n23917 );
and ( n62991 , n19456 , n34526 );
or ( n62992 , n62974 , n62978 , n62982 , n62986 , n62990 , n62991 );
and ( n62993 , n62970 , n62992 );
and ( n62994 , n19456 , n17451 );
or ( n62995 , n62993 , n62994 );
and ( n62996 , n62995 , n23924 );
and ( n62997 , n19456 , n23926 );
or ( n62998 , n62996 , n62997 );
buf ( n62999 , n62998 );
buf ( n63000 , n62999 );
buf ( n63001 , n10613 );
buf ( n63002 , n10615 );
buf ( n63003 , n10613 );
buf ( n63004 , n10615 );
buf ( n63005 , n10615 );
buf ( n63006 , n10613 );
buf ( n63007 , n10613 );
not ( n63008 , n11954 );
not ( n63009 , n12243 );
and ( n63010 , n10837 , n31187 );
not ( n63011 , n31697 );
and ( n63012 , n63011 , n31608 );
xor ( n63013 , n56882 , n56887 );
and ( n63014 , n63013 , n31697 );
or ( n63015 , n63012 , n63014 );
buf ( n63016 , n63015 );
and ( n63017 , n63016 , n14140 );
not ( n63018 , n32214 );
and ( n63019 , n63018 , n32125 );
xor ( n63020 , n56905 , n56910 );
and ( n63021 , n63020 , n32214 );
or ( n63022 , n63019 , n63021 );
buf ( n63023 , n63022 );
and ( n63024 , n63023 , n14137 );
and ( n63025 , n15557 , n14143 );
and ( n63026 , n10837 , n14141 );
or ( n63027 , n63017 , n63024 , n63025 , n63026 );
and ( n63028 , n63027 , n32236 );
or ( n63029 , n63010 , n63028 );
and ( n63030 , n63009 , n63029 );
not ( n63031 , n34038 );
and ( n63032 , n63031 , n33914 );
xor ( n63033 , n56934 , n56939 );
and ( n63034 , n63033 , n34038 );
or ( n63035 , n63032 , n63034 );
buf ( n63036 , n63035 );
and ( n63037 , n63036 , n12243 );
or ( n63038 , n63030 , n63037 );
and ( n63039 , n63008 , n63038 );
and ( n63040 , n63027 , n11954 );
or ( n63041 , n63039 , n63040 );
and ( n63042 , n63041 , n16574 );
not ( n63043 , n34327 );
and ( n63044 , n63043 , n34253 );
xor ( n63045 , n56962 , n56967 );
and ( n63046 , n63045 , n34327 );
or ( n63047 , n63044 , n63046 );
buf ( n63048 , n63047 );
and ( n63049 , n63048 , n16576 );
or ( n63050 , n63042 , n63049 );
buf ( n63051 , n63050 );
buf ( n63052 , n63051 );
buf ( n63053 , n10613 );
buf ( n63054 , n10615 );
not ( n63055 , n34804 );
and ( n63056 , n63055 , n26195 );
and ( n63057 , n14773 , n34804 );
or ( n63058 , n63056 , n63057 );
and ( n63059 , n63058 , n31008 );
and ( n63060 , n14773 , n10618 );
or ( n63061 , n63059 , n63060 );
buf ( n63062 , n63061 );
buf ( n63063 , n63062 );
not ( n63064 , n24511 );
not ( n63065 , n24799 );
and ( n63066 , n10645 , n40154 );
not ( n63067 , n40632 );
and ( n63068 , n63067 , n40611 );
xor ( n63069 , n43752 , n43757 );
and ( n63070 , n63069 , n40632 );
or ( n63071 , n63068 , n63070 );
buf ( n63072 , n63071 );
and ( n63073 , n63072 , n27046 );
not ( n63074 , n41147 );
and ( n63075 , n63074 , n41126 );
xor ( n63076 , n43767 , n43772 );
and ( n63077 , n63076 , n41147 );
or ( n63078 , n63075 , n63077 );
buf ( n63079 , n63078 );
and ( n63080 , n63079 , n27049 );
and ( n63081 , n29313 , n28506 );
and ( n63082 , n10645 , n28508 );
or ( n63083 , n63073 , n63080 , n63081 , n63082 );
and ( n63084 , n63083 , n41199 );
or ( n63085 , n63066 , n63084 );
and ( n63086 , n63065 , n63085 );
xor ( n63087 , n43815 , n43823 );
xor ( n63088 , n63087 , n43866 );
buf ( n63089 , n63088 );
and ( n63090 , n63089 , n27046 );
xor ( n63091 , n43896 , n43897 );
xor ( n63092 , n63091 , n43926 );
buf ( n63093 , n63092 );
and ( n63094 , n63093 , n27049 );
and ( n63095 , n29313 , n42306 );
or ( n63096 , n63090 , n63094 , n63095 );
buf ( n63097 , n63096 );
and ( n63098 , C1 , n63097 );
or ( n63099 , n63098 , C0 );
buf ( n63100 , n63099 );
not ( n63101 , n63100 );
buf ( n63102 , n63101 );
buf ( n63103 , n63102 );
not ( n63104 , n63103 );
and ( n63105 , C1 , n63104 );
or ( n63106 , n63105 , C0 );
buf ( n63107 , n63106 );
and ( n63108 , n63107 , n24799 );
or ( n63109 , n63086 , n63108 );
and ( n63110 , n63064 , n63109 );
and ( n63111 , n63083 , n24511 );
or ( n63112 , n63110 , n63111 );
and ( n63113 , n63112 , n31008 );
not ( n63114 , n42601 );
and ( n63115 , n63114 , n42583 );
xor ( n63116 , n43955 , n43960 );
and ( n63117 , n63116 , n42601 );
or ( n63118 , n63115 , n63117 );
buf ( n63119 , n63118 );
and ( n63120 , n63119 , n10618 );
or ( n63121 , n63113 , n63120 );
buf ( n63122 , n63121 );
buf ( n63123 , n63122 );
buf ( n63124 , n10615 );
not ( n63125 , n34821 );
and ( n63126 , n13169 , n14592 );
and ( n63127 , n49057 , n36348 );
and ( n63128 , n13169 , n43530 );
or ( n63129 , n63127 , n63128 );
and ( n63130 , n63129 , n14562 );
and ( n63131 , n49067 , n36347 );
and ( n63132 , n13169 , n43543 );
or ( n63133 , n63131 , n63132 );
and ( n63134 , n63133 , n14586 );
and ( n63135 , n49077 , n36348 );
and ( n63136 , n13169 , n43556 );
or ( n63137 , n63135 , n63136 );
and ( n63138 , n63137 , n14584 );
and ( n63139 , n49067 , n36347 );
and ( n63140 , n13169 , n43563 );
or ( n63141 , n63139 , n63140 );
and ( n63142 , n63141 , n37835 );
and ( n63143 , n49077 , n36347 );
and ( n63144 , n13169 , n43563 );
or ( n63145 , n63143 , n63144 );
and ( n63146 , n63145 , n37841 );
and ( n63147 , n13167 , n14564 );
and ( n63148 , n15007 , n36347 );
and ( n63149 , n13169 , n43563 );
or ( n63150 , n63148 , n63149 );
and ( n63151 , n63150 , n37847 );
or ( n63152 , n63126 , n63130 , n63134 , n63138 , n63142 , n63146 , n63147 , n63151 );
and ( n63153 , n63125 , n63152 );
and ( n63154 , n13169 , n34821 );
or ( n63155 , n63153 , n63154 );
and ( n63156 , n63155 , n16574 );
and ( n63157 , n13169 , n16576 );
or ( n63158 , n63156 , n63157 );
buf ( n63159 , n63158 );
buf ( n63160 , n63159 );
buf ( n63161 , n10613 );
not ( n63162 , n11954 );
not ( n63163 , n12243 );
and ( n63164 , n10917 , n31187 );
not ( n63165 , n31697 );
and ( n63166 , n63165 , n31438 );
xor ( n63167 , n50362 , n50369 );
and ( n63168 , n63167 , n31697 );
or ( n63169 , n63166 , n63168 );
buf ( n63170 , n63169 );
and ( n63171 , n63170 , n14140 );
not ( n63172 , n32214 );
and ( n63173 , n63172 , n31955 );
xor ( n63174 , n50389 , n50396 );
and ( n63175 , n63174 , n32214 );
or ( n63176 , n63173 , n63175 );
buf ( n63177 , n63176 );
and ( n63178 , n63177 , n14137 );
and ( n63179 , n15777 , n14143 );
and ( n63180 , n10917 , n14141 );
or ( n63181 , n63171 , n63178 , n63179 , n63180 );
and ( n63182 , n63181 , n32236 );
or ( n63183 , n63164 , n63182 );
and ( n63184 , n63163 , n63183 );
not ( n63185 , n34038 );
and ( n63186 , n63185 , n33674 );
xor ( n63187 , n50422 , n50429 );
and ( n63188 , n63187 , n34038 );
or ( n63189 , n63186 , n63188 );
buf ( n63190 , n63189 );
and ( n63191 , n63190 , n12243 );
or ( n63192 , n63184 , n63191 );
and ( n63193 , n63162 , n63192 );
and ( n63194 , n63181 , n11954 );
or ( n63195 , n63193 , n63194 );
and ( n63196 , n63195 , n16574 );
not ( n63197 , n34327 );
and ( n63198 , n63197 , n34113 );
xor ( n63199 , n50454 , n50461 );
and ( n63200 , n63199 , n34327 );
or ( n63201 , n63198 , n63200 );
buf ( n63202 , n63201 );
and ( n63203 , n63202 , n16576 );
or ( n63204 , n63196 , n63203 );
buf ( n63205 , n63204 );
buf ( n63206 , n63205 );
buf ( n63207 , n10613 );
buf ( n63208 , n10613 );
buf ( n63209 , n10613 );
buf ( n63210 , n10613 );
not ( n63211 , n34821 );
and ( n63212 , n13241 , n14592 );
and ( n63213 , n53712 , n36348 );
and ( n63214 , n13241 , n43530 );
or ( n63215 , n63213 , n63214 );
and ( n63216 , n63215 , n14562 );
and ( n63217 , n53722 , n36347 );
and ( n63218 , n13241 , n43543 );
or ( n63219 , n63217 , n63218 );
and ( n63220 , n63219 , n14586 );
and ( n63221 , n53732 , n36348 );
and ( n63222 , n13241 , n43556 );
or ( n63223 , n63221 , n63222 );
and ( n63224 , n63223 , n14584 );
and ( n63225 , n53722 , n36347 );
and ( n63226 , n13241 , n43563 );
or ( n63227 , n63225 , n63226 );
and ( n63228 , n63227 , n37835 );
and ( n63229 , n53732 , n36347 );
and ( n63230 , n13241 , n43563 );
or ( n63231 , n63229 , n63230 );
and ( n63232 , n63231 , n37841 );
and ( n63233 , n13239 , n14564 );
and ( n63234 , n15097 , n36347 );
and ( n63235 , n13241 , n43563 );
or ( n63236 , n63234 , n63235 );
and ( n63237 , n63236 , n37847 );
or ( n63238 , n63212 , n63216 , n63220 , n63224 , n63228 , n63232 , n63233 , n63237 );
and ( n63239 , n63211 , n63238 );
and ( n63240 , n13241 , n34821 );
or ( n63241 , n63239 , n63240 );
and ( n63242 , n63241 , n16574 );
and ( n63243 , n13241 , n16576 );
or ( n63244 , n63242 , n63243 );
buf ( n63245 , n63244 );
buf ( n63246 , n63245 );
not ( n63247 , n11333 );
and ( n63248 , n63247 , n11023 );
xor ( n63249 , n11350 , n11352 );
and ( n63250 , n63249 , n11333 );
or ( n63251 , n63248 , n63250 );
buf ( n63252 , n63251 );
buf ( n63253 , n63252 );
buf ( n63254 , n10613 );
buf ( n63255 , n10615 );
buf ( n63256 , n10615 );
buf ( n63257 , n10615 );
buf ( n63258 , n10613 );
buf ( n63259 , n10615 );
not ( n63260 , n17451 );
and ( n63261 , n18807 , n17873 );
nand ( n63262 , n46858 , n21330 );
and ( n63263 , n18807 , n21338 );
or ( n63264 , n63262 , n63263 );
and ( n63265 , n63264 , n21341 );
and ( n63266 , n46868 , n21330 );
and ( n63267 , n18807 , n21338 );
or ( n63268 , n63266 , n63267 );
and ( n63269 , n63268 , n23064 );
and ( n63270 , n46878 , n21330 );
and ( n63271 , n18807 , n21338 );
or ( n63272 , n63270 , n63271 );
and ( n63273 , n63272 , n23825 );
and ( n63274 , n22242 , n21330 );
and ( n63275 , n18807 , n21338 );
or ( n63276 , n63274 , n63275 );
and ( n63277 , n63276 , n23832 );
and ( n63278 , n18805 , n23834 );
and ( n63279 , n46888 , n21330 );
and ( n63280 , n18807 , n21338 );
or ( n63281 , n63279 , n63280 );
and ( n63282 , n63281 , n23917 );
or ( n63283 , n63261 , n63265 , n63269 , n63273 , n63277 , n63278 , n63282 );
and ( n63284 , n63260 , n63283 );
and ( n63285 , n18807 , n17451 );
or ( n63286 , n63284 , n63285 );
and ( n63287 , n63286 , n23924 );
and ( n63288 , n18807 , n23926 );
or ( n63289 , n63287 , n63288 );
buf ( n63290 , n63289 );
buf ( n63291 , n63290 );
buf ( n63292 , n10615 );
buf ( n63293 , n10613 );
not ( n63294 , n17451 );
and ( n63295 , n43338 , n21333 );
and ( n63296 , n18911 , n34758 );
or ( n63297 , n63295 , n63296 );
and ( n63298 , n63297 , n21341 );
and ( n63299 , n43348 , n21333 );
and ( n63300 , n18911 , n34758 );
or ( n63301 , n63299 , n63300 );
and ( n63302 , n63301 , n23064 );
and ( n63303 , n43358 , n21333 );
and ( n63304 , n18911 , n34758 );
or ( n63305 , n63303 , n63304 );
and ( n63306 , n63305 , n23825 );
and ( n63307 , n22182 , n21333 );
and ( n63308 , n18911 , n34758 );
or ( n63309 , n63307 , n63308 );
and ( n63310 , n63309 , n23832 );
and ( n63311 , n43368 , n21333 );
and ( n63312 , n18911 , n34758 );
or ( n63313 , n63311 , n63312 );
and ( n63314 , n63313 , n23917 );
and ( n63315 , n18911 , n34526 );
or ( n63316 , n63298 , n63302 , n63306 , n63310 , n63314 , n63315 );
and ( n63317 , n63294 , n63316 );
and ( n63318 , n18911 , n17451 );
or ( n63319 , n63317 , n63318 );
and ( n63320 , n63319 , n23924 );
and ( n63321 , n18911 , n23926 );
or ( n63322 , n63320 , n63321 );
buf ( n63323 , n63322 );
buf ( n63324 , n63323 );
buf ( n63325 , n10613 );
buf ( n63326 , n10613 );
buf ( n63327 , n10613 );
not ( n63328 , n34538 );
and ( n63329 , n63328 , n19017 );
and ( n63330 , n14741 , n34538 );
or ( n63331 , n63329 , n63330 );
and ( n63332 , n63331 , n23924 );
and ( n63333 , n14741 , n23926 );
or ( n63334 , n63332 , n63333 );
buf ( n63335 , n63334 );
buf ( n63336 , n63335 );
not ( n63337 , n34538 );
and ( n63338 , n63337 , n18711 );
and ( n63339 , n14795 , n34538 );
or ( n63340 , n63338 , n63339 );
and ( n63341 , n63340 , n23924 );
and ( n63342 , n14795 , n23926 );
or ( n63343 , n63341 , n63342 );
buf ( n63344 , n63343 );
buf ( n63345 , n63344 );
buf ( n63346 , n10615 );
buf ( n63347 , n10615 );
not ( n63348 , n17451 );
and ( n63349 , n39326 , n21333 );
and ( n63350 , n19081 , n34758 );
or ( n63351 , n63349 , n63350 );
and ( n63352 , n63351 , n21341 );
and ( n63353 , n39336 , n21333 );
and ( n63354 , n19081 , n34758 );
or ( n63355 , n63353 , n63354 );
and ( n63356 , n63355 , n23064 );
and ( n63357 , n39346 , n21333 );
and ( n63358 , n19081 , n34758 );
or ( n63359 , n63357 , n63358 );
and ( n63360 , n63359 , n23825 );
and ( n63361 , n22082 , n21333 );
and ( n63362 , n19081 , n34758 );
or ( n63363 , n63361 , n63362 );
and ( n63364 , n63363 , n23832 );
and ( n63365 , n39356 , n21333 );
and ( n63366 , n19081 , n34758 );
or ( n63367 , n63365 , n63366 );
and ( n63368 , n63367 , n23917 );
and ( n63369 , n19081 , n34526 );
or ( n63370 , n63352 , n63356 , n63360 , n63364 , n63368 , n63369 );
and ( n63371 , n63348 , n63370 );
and ( n63372 , n19081 , n17451 );
or ( n63373 , n63371 , n63372 );
and ( n63374 , n63373 , n23924 );
and ( n63375 , n19081 , n23926 );
or ( n63376 , n63374 , n63375 );
buf ( n63377 , n63376 );
buf ( n63378 , n63377 );
buf ( n63379 , n10615 );
buf ( n63380 , n10615 );
buf ( n63381 , n10613 );
buf ( n63382 , n10613 );
not ( n63383 , n24800 );
and ( n63384 , n26629 , n25222 );
and ( n63385 , n54833 , n28589 );
and ( n63386 , n26629 , n31075 );
or ( n63387 , n63385 , n63386 );
and ( n63388 , n63387 , n28594 );
and ( n63389 , n54843 , n28589 );
and ( n63390 , n26629 , n31075 );
or ( n63391 , n63389 , n63390 );
and ( n63392 , n63391 , n30269 );
and ( n63393 , n54853 , n28589 );
and ( n63394 , n26629 , n31075 );
or ( n63395 , n63393 , n63394 );
and ( n63396 , n63395 , n30982 );
and ( n63397 , n29198 , n28589 );
and ( n63398 , n26629 , n31075 );
or ( n63399 , n63397 , n63398 );
and ( n63400 , n63399 , n30989 );
and ( n63401 , n29198 , n30991 );
and ( n63402 , n54863 , n28589 );
and ( n63403 , n26629 , n31075 );
or ( n63404 , n63402 , n63403 );
and ( n63405 , n63404 , n31002 );
or ( n63406 , n63384 , n63388 , n63392 , n63396 , n63400 , n63401 , n63405 );
and ( n63407 , n63383 , n63406 );
and ( n63408 , n26629 , n24800 );
or ( n63409 , n63407 , n63408 );
and ( n63410 , n63409 , n31008 );
and ( n63411 , n25564 , n10618 );
or ( n63412 , n63410 , n63411 );
buf ( n63413 , n63412 );
buf ( n63414 , n63413 );
buf ( n63415 , n10613 );
not ( n63416 , n34821 );
and ( n63417 , n55549 , n36347 );
and ( n63418 , n13158 , n39408 );
or ( n63419 , n63417 , n63418 );
and ( n63420 , n63419 , n14562 );
and ( n63421 , n55559 , n36348 );
and ( n63422 , n13158 , n39427 );
or ( n63423 , n63421 , n63422 );
and ( n63424 , n63423 , n14586 );
and ( n63425 , n55569 , n36347 );
and ( n63426 , n13158 , n39446 );
or ( n63427 , n63425 , n63426 );
and ( n63428 , n63427 , n14584 );
and ( n63429 , n55559 , n36348 );
and ( n63430 , n13158 , n39453 );
or ( n63431 , n63429 , n63430 );
and ( n63432 , n63431 , n37835 );
and ( n63433 , n55569 , n36348 );
and ( n63434 , n13158 , n39453 );
or ( n63435 , n63433 , n63434 );
and ( n63436 , n63435 , n37841 );
and ( n63437 , n14992 , n36348 );
and ( n63438 , n13158 , n39453 );
or ( n63439 , n63437 , n63438 );
and ( n63440 , n63439 , n37847 );
and ( n63441 , n13158 , n37849 );
or ( n63442 , n63420 , n63424 , n63428 , n63432 , n63436 , n63440 , n63441 );
and ( n63443 , n63416 , n63442 );
and ( n63444 , n13158 , n34821 );
or ( n63445 , n63443 , n63444 );
and ( n63446 , n63445 , n16574 );
and ( n63447 , n13158 , n16576 );
or ( n63448 , n63446 , n63447 );
buf ( n63449 , n63448 );
buf ( n63450 , n63449 );
buf ( n63451 , n10613 );
buf ( n63452 , n10615 );
not ( n63453 , n34538 );
and ( n63454 , n63453 , n19221 );
and ( n63455 , n14705 , n34538 );
or ( n63456 , n63454 , n63455 );
and ( n63457 , n63456 , n23924 );
and ( n63458 , n14705 , n23926 );
or ( n63459 , n63457 , n63458 );
buf ( n63460 , n63459 );
buf ( n63461 , n63460 );
not ( n63462 , n34821 );
and ( n63463 , n45165 , n36345 );
and ( n63464 , n13269 , n36352 );
or ( n63465 , n63463 , n63464 );
and ( n63466 , n63465 , n14562 );
and ( n63467 , n45181 , n36345 );
and ( n63468 , n13269 , n37073 );
or ( n63469 , n63467 , n63468 );
and ( n63470 , n63469 , n14586 );
and ( n63471 , n45197 , n36350 );
and ( n63472 , n13269 , n37825 );
or ( n63473 , n63471 , n63472 );
and ( n63474 , n63473 , n14584 );
and ( n63475 , n45181 , n36350 );
and ( n63476 , n13269 , n37831 );
or ( n63477 , n63475 , n63476 );
and ( n63478 , n63477 , n37835 );
and ( n63479 , n45197 , n36350 );
and ( n63480 , n13269 , n37831 );
or ( n63481 , n63479 , n63480 );
and ( n63482 , n63481 , n37841 );
and ( n63483 , n15449 , n36350 );
and ( n63484 , n13269 , n37831 );
or ( n63485 , n63483 , n63484 );
and ( n63486 , n63485 , n37847 );
and ( n63487 , n13269 , n37849 );
or ( n63488 , n63466 , n63470 , n63474 , n63478 , n63482 , n63486 , n63487 );
and ( n63489 , n63462 , n63488 );
and ( n63490 , n13269 , n34821 );
or ( n63491 , n63489 , n63490 );
and ( n63492 , n63491 , n16574 );
and ( n63493 , n13269 , n16576 );
or ( n63494 , n63492 , n63493 );
buf ( n63495 , n63494 );
buf ( n63496 , n63495 );
not ( n63497 , n34804 );
and ( n63498 , n63497 , n25958 );
and ( n63499 , n14815 , n34804 );
or ( n63500 , n63498 , n63499 );
and ( n63501 , n63500 , n31008 );
and ( n63502 , n14815 , n10618 );
or ( n63503 , n63501 , n63502 );
buf ( n63504 , n63503 );
buf ( n63505 , n63504 );
not ( n63506 , n34538 );
and ( n63507 , n63506 , n18779 );
and ( n63508 , n14783 , n34538 );
or ( n63509 , n63507 , n63508 );
and ( n63510 , n63509 , n23924 );
and ( n63511 , n14783 , n23926 );
or ( n63512 , n63510 , n63511 );
buf ( n63513 , n63512 );
buf ( n63514 , n63513 );
buf ( n63515 , n10615 );
and ( n63516 , n24182 , n31008 );
and ( n63517 , n29486 , n10618 );
or ( n63518 , n63516 , n63517 );
buf ( n63519 , n63518 );
buf ( n63520 , n63519 );
buf ( n63521 , n10613 );
not ( n63522 , n17162 );
not ( n63523 , n17450 );
and ( n63524 , n10643 , n37947 );
not ( n63525 , n38425 );
and ( n63526 , n63525 , n38404 );
xor ( n63527 , n52275 , n52276 );
and ( n63528 , n63527 , n38425 );
or ( n63529 , n63526 , n63528 );
buf ( n63530 , n63529 );
and ( n63531 , n63530 , n19745 );
not ( n63532 , n38934 );
and ( n63533 , n63532 , n38913 );
xor ( n63534 , n52286 , n52287 );
and ( n63535 , n63534 , n38934 );
or ( n63536 , n63533 , n63535 );
buf ( n63537 , n63536 );
and ( n63538 , n63537 , n19748 );
and ( n63539 , n22060 , n21253 );
and ( n63540 , n10643 , n21255 );
or ( n63541 , n63531 , n63538 , n63539 , n63540 );
and ( n63542 , n63541 , n38980 );
or ( n63543 , n63524 , n63542 );
and ( n63544 , n63523 , n63543 );
or ( n63545 , n63544 , C0 );
and ( n63546 , n63522 , n63545 );
and ( n63547 , n63541 , n17162 );
or ( n63548 , n63546 , n63547 );
and ( n63549 , n63548 , n23924 );
not ( n63550 , n39264 );
and ( n63551 , n63550 , n39246 );
xor ( n63552 , n52308 , n52309 );
and ( n63553 , n63552 , n39264 );
or ( n63554 , n63551 , n63553 );
buf ( n63555 , n63554 );
and ( n63556 , n63555 , n23926 );
or ( n63557 , n63549 , n63556 );
buf ( n63558 , n63557 );
buf ( n63559 , n63558 );
not ( n63560 , n34538 );
and ( n63561 , n63560 , n18577 );
and ( n63562 , n14819 , n34538 );
or ( n63563 , n63561 , n63562 );
and ( n63564 , n63563 , n23924 );
and ( n63565 , n14819 , n23926 );
or ( n63566 , n63564 , n63565 );
buf ( n63567 , n63566 );
buf ( n63568 , n63567 );
buf ( n63569 , n10615 );
buf ( n63570 , n10615 );
buf ( n63571 , n10615 );
not ( n63572 , n34821 );
and ( n63573 , n59483 , n36347 );
and ( n63574 , n13435 , n39408 );
or ( n63575 , n63573 , n63574 );
and ( n63576 , n63575 , n14562 );
and ( n63577 , n59493 , n36348 );
and ( n63578 , n13435 , n39427 );
or ( n63579 , n63577 , n63578 );
and ( n63580 , n63579 , n14586 );
and ( n63581 , n59503 , n36347 );
and ( n63582 , n13435 , n39446 );
or ( n63583 , n63581 , n63582 );
and ( n63584 , n63583 , n14584 );
and ( n63585 , n59493 , n36348 );
and ( n63586 , n13435 , n39453 );
or ( n63587 , n63585 , n63586 );
and ( n63588 , n63587 , n37835 );
and ( n63589 , n59503 , n36348 );
and ( n63590 , n13435 , n39453 );
or ( n63591 , n63589 , n63590 );
and ( n63592 , n63591 , n37841 );
and ( n63593 , n15757 , n36348 );
and ( n63594 , n13435 , n39453 );
or ( n63595 , n63593 , n63594 );
and ( n63596 , n63595 , n37847 );
and ( n63597 , n13435 , n37849 );
or ( n63598 , n63576 , n63580 , n63584 , n63588 , n63592 , n63596 , n63597 );
and ( n63599 , n63572 , n63598 );
and ( n63600 , n13435 , n34821 );
or ( n63601 , n63599 , n63600 );
and ( n63602 , n63601 , n16574 );
and ( n63603 , n13435 , n16576 );
or ( n63604 , n63602 , n63603 );
buf ( n63605 , n63604 );
buf ( n63606 , n63605 );
not ( n63607 , n34821 );
and ( n63608 , n13431 , n14592 );
and ( n63609 , n59483 , n36350 );
and ( n63610 , n13431 , n43691 );
or ( n63611 , n63609 , n63610 );
and ( n63612 , n63611 , n14562 );
and ( n63613 , n59493 , n36350 );
and ( n63614 , n13431 , n43703 );
or ( n63615 , n63613 , n63614 );
and ( n63616 , n63615 , n14586 );
and ( n63617 , n59503 , n36345 );
and ( n63618 , n13431 , n43715 );
or ( n63619 , n63617 , n63618 );
and ( n63620 , n63619 , n14584 );
and ( n63621 , n59493 , n36345 );
and ( n63622 , n13431 , n43721 );
or ( n63623 , n63621 , n63622 );
and ( n63624 , n63623 , n37835 );
and ( n63625 , n59503 , n36345 );
and ( n63626 , n13431 , n43721 );
or ( n63627 , n63625 , n63626 );
and ( n63628 , n63627 , n37841 );
and ( n63629 , n15757 , n14564 );
and ( n63630 , n15757 , n36345 );
and ( n63631 , n13431 , n43721 );
or ( n63632 , n63630 , n63631 );
and ( n63633 , n63632 , n37847 );
or ( n63634 , n63608 , n63612 , n63616 , n63620 , n63624 , n63628 , n63629 , n63633 );
and ( n63635 , n63607 , n63634 );
and ( n63636 , n13431 , n34821 );
or ( n63637 , n63635 , n63636 );
and ( n63638 , n63637 , n16574 );
and ( n63639 , n12318 , n16576 );
or ( n63640 , n63638 , n63639 );
buf ( n63641 , n63640 );
buf ( n63642 , n63641 );
buf ( n63643 , n10613 );
not ( n63644 , n17451 );
and ( n63645 , n18604 , n17873 );
and ( n63646 , n48952 , n21330 );
and ( n63647 , n18604 , n21338 );
or ( n63648 , n63646 , n63647 );
and ( n63649 , n63648 , n21341 );
and ( n63650 , n48962 , n21330 );
and ( n63651 , n18604 , n21338 );
or ( n63652 , n63650 , n63651 );
and ( n63653 , n63652 , n23064 );
and ( n63654 , n48972 , n21330 );
and ( n63655 , n18604 , n21338 );
or ( n63656 , n63654 , n63655 );
and ( n63657 , n63656 , n23825 );
and ( n63658 , n22362 , n21330 );
and ( n63659 , n18604 , n21338 );
or ( n63660 , n63658 , n63659 );
and ( n63661 , n63660 , n23832 );
and ( n63662 , n18602 , n23834 );
and ( n63663 , n48982 , n21330 );
and ( n63664 , n18604 , n21338 );
or ( n63665 , n63663 , n63664 );
and ( n63666 , n63665 , n23917 );
or ( n63667 , n63645 , n63649 , n63653 , n63657 , n63661 , n63662 , n63666 );
and ( n63668 , n63644 , n63667 );
and ( n63669 , n18604 , n17451 );
or ( n63670 , n63668 , n63669 );
and ( n63671 , n63670 , n23924 );
and ( n63672 , n18604 , n23926 );
or ( n63673 , n63671 , n63672 );
buf ( n63674 , n63673 );
buf ( n63675 , n63674 );
buf ( n63676 , n10615 );
buf ( n63677 , n10615 );
buf ( n63678 , n10615 );
buf ( n63679 , n10615 );
buf ( n63680 , n10615 );
buf ( n63681 , n10613 );
not ( n63682 , n34821 );
and ( n63683 , n13253 , n14592 );
and ( n63684 , n57357 , n36348 );
and ( n63685 , n13253 , n43530 );
or ( n63686 , n63684 , n63685 );
and ( n63687 , n63686 , n14562 );
and ( n63688 , n57367 , n36347 );
and ( n63689 , n13253 , n43543 );
or ( n63690 , n63688 , n63689 );
and ( n63691 , n63690 , n14586 );
and ( n63692 , n57377 , n36348 );
and ( n63693 , n13253 , n43556 );
or ( n63694 , n63692 , n63693 );
and ( n63695 , n63694 , n14584 );
and ( n63696 , n57367 , n36347 );
and ( n63697 , n13253 , n43563 );
or ( n63698 , n63696 , n63697 );
and ( n63699 , n63698 , n37835 );
and ( n63700 , n57377 , n36347 );
and ( n63701 , n13253 , n43563 );
or ( n63702 , n63700 , n63701 );
and ( n63703 , n63702 , n37841 );
and ( n63704 , n13251 , n14564 );
and ( n63705 , n15112 , n36347 );
and ( n63706 , n13253 , n43563 );
or ( n63707 , n63705 , n63706 );
and ( n63708 , n63707 , n37847 );
or ( n63709 , n63683 , n63687 , n63691 , n63695 , n63699 , n63703 , n63704 , n63708 );
and ( n63710 , n63682 , n63709 );
and ( n63711 , n13253 , n34821 );
or ( n63712 , n63710 , n63711 );
and ( n63713 , n63712 , n16574 );
and ( n63714 , n13253 , n16576 );
or ( n63715 , n63713 , n63714 );
buf ( n63716 , n63715 );
buf ( n63717 , n63716 );
buf ( n63718 , n10615 );
buf ( n63719 , n10613 );
not ( n63720 , n34538 );
and ( n63721 , n63720 , n19289 );
and ( n63722 , n14693 , n34538 );
or ( n63723 , n63721 , n63722 );
and ( n63724 , n63723 , n23924 );
and ( n63725 , n14693 , n23926 );
or ( n63726 , n63724 , n63725 );
buf ( n63727 , n63726 );
buf ( n63728 , n63727 );
buf ( n63729 , n10615 );
buf ( n63730 , n10615 );
buf ( n63731 , n10613 );
buf ( n63732 , n10613 );
buf ( n63733 , n10615 );
buf ( n63734 , n10615 );
not ( n63735 , n11954 );
not ( n63736 , n12243 );
and ( n63737 , n10821 , n31187 );
not ( n63738 , n31697 );
and ( n63739 , n63738 , n31642 );
xor ( n63740 , n56880 , n56889 );
and ( n63741 , n63740 , n31697 );
or ( n63742 , n63739 , n63741 );
buf ( n63743 , n63742 );
and ( n63744 , n63743 , n14140 );
not ( n63745 , n32214 );
and ( n63746 , n63745 , n32159 );
xor ( n63747 , n56903 , n56912 );
and ( n63748 , n63747 , n32214 );
or ( n63749 , n63746 , n63748 );
buf ( n63750 , n63749 );
and ( n63751 , n63750 , n14137 );
and ( n63752 , n15513 , n14143 );
and ( n63753 , n10821 , n14141 );
or ( n63754 , n63744 , n63751 , n63752 , n63753 );
and ( n63755 , n63754 , n32236 );
or ( n63756 , n63737 , n63755 );
and ( n63757 , n63736 , n63756 );
not ( n63758 , n34038 );
and ( n63759 , n63758 , n33962 );
xor ( n63760 , n56932 , n56941 );
and ( n63761 , n63760 , n34038 );
or ( n63762 , n63759 , n63761 );
buf ( n63763 , n63762 );
and ( n63764 , n63763 , n12243 );
or ( n63765 , n63757 , n63764 );
and ( n63766 , n63735 , n63765 );
and ( n63767 , n63754 , n11954 );
or ( n63768 , n63766 , n63767 );
and ( n63769 , n63768 , n16574 );
not ( n63770 , n34327 );
and ( n63771 , n63770 , n34281 );
xor ( n63772 , n56960 , n56969 );
and ( n63773 , n63772 , n34327 );
or ( n63774 , n63771 , n63773 );
buf ( n63775 , n63774 );
and ( n63776 , n63775 , n16576 );
or ( n63777 , n63769 , n63776 );
buf ( n63778 , n63777 );
buf ( n63779 , n63778 );
not ( n63780 , n17451 );
and ( n63781 , n52940 , n21333 );
and ( n63782 , n18523 , n34758 );
or ( n63783 , n63781 , n63782 );
and ( n63784 , n63783 , n21341 );
and ( n63785 , n18523 , n34758 );
buf ( n63786 , n63785 );
and ( n63787 , n63786 , n23064 );
and ( n63788 , n18523 , n34758 );
buf ( n63789 , n63788 );
and ( n63790 , n63789 , n23825 );
and ( n63791 , n21841 , n21333 );
and ( n63792 , n18523 , n34758 );
or ( n63793 , n63791 , n63792 );
and ( n63794 , n63793 , n23832 );
and ( n63795 , n52959 , n21333 );
and ( n63796 , n18523 , n34758 );
or ( n63797 , n63795 , n63796 );
and ( n63798 , n63797 , n23917 );
and ( n63799 , n18523 , n34526 );
or ( n63800 , n63784 , n63787 , n63790 , n63794 , n63798 , n63799 );
and ( n63801 , n63780 , n63800 );
and ( n63802 , n18523 , n17451 );
or ( n63803 , n63801 , n63802 );
and ( n63804 , n63803 , n23924 );
and ( n63805 , n18523 , n23926 );
or ( n63806 , n63804 , n63805 );
buf ( n63807 , n63806 );
buf ( n63808 , n63807 );
buf ( n63809 , n10613 );
not ( n63810 , n11954 );
not ( n63811 , n12243 );
and ( n63812 , n10829 , n31187 );
not ( n63813 , n31697 );
and ( n63814 , n63813 , n31625 );
xor ( n63815 , n56881 , n56888 );
and ( n63816 , n63815 , n31697 );
or ( n63817 , n63814 , n63816 );
buf ( n63818 , n63817 );
and ( n63819 , n63818 , n14140 );
not ( n63820 , n32214 );
and ( n63821 , n63820 , n32142 );
xor ( n63822 , n56904 , n56911 );
and ( n63823 , n63822 , n32214 );
or ( n63824 , n63821 , n63823 );
buf ( n63825 , n63824 );
and ( n63826 , n63825 , n14137 );
and ( n63827 , n15535 , n14143 );
and ( n63828 , n10829 , n14141 );
or ( n63829 , n63819 , n63826 , n63827 , n63828 );
and ( n63830 , n63829 , n32236 );
or ( n63831 , n63812 , n63830 );
and ( n63832 , n63811 , n63831 );
not ( n63833 , n34038 );
and ( n63834 , n63833 , n33938 );
xor ( n63835 , n56933 , n56940 );
and ( n63836 , n63835 , n34038 );
or ( n63837 , n63834 , n63836 );
buf ( n63838 , n63837 );
and ( n63839 , n63838 , n12243 );
or ( n63840 , n63832 , n63839 );
and ( n63841 , n63810 , n63840 );
and ( n63842 , n63829 , n11954 );
or ( n63843 , n63841 , n63842 );
and ( n63844 , n63843 , n16574 );
not ( n63845 , n34327 );
and ( n63846 , n63845 , n34267 );
xor ( n63847 , n56961 , n56968 );
and ( n63848 , n63847 , n34327 );
or ( n63849 , n63846 , n63848 );
buf ( n63850 , n63849 );
and ( n63851 , n63850 , n16576 );
or ( n63852 , n63844 , n63851 );
buf ( n63853 , n63852 );
buf ( n63854 , n63853 );
buf ( n63855 , n10613 );
buf ( n63856 , n10613 );
not ( n63857 , n24800 );
and ( n63858 , n31072 , n28587 );
and ( n63859 , n26193 , n39807 );
or ( n63860 , n63858 , n63859 );
and ( n63861 , n63860 , n28594 );
and ( n63862 , n31102 , n28587 );
and ( n63863 , n26193 , n39807 );
or ( n63864 , n63862 , n63863 );
and ( n63865 , n63864 , n30269 );
and ( n63866 , n31130 , n28587 );
and ( n63867 , n26193 , n39807 );
or ( n63868 , n63866 , n63867 );
and ( n63869 , n63868 , n30982 );
and ( n63870 , n29475 , n28587 );
and ( n63871 , n26193 , n39807 );
or ( n63872 , n63870 , n63871 );
and ( n63873 , n63872 , n30989 );
and ( n63874 , n31168 , n28587 );
and ( n63875 , n26193 , n39807 );
or ( n63876 , n63874 , n63875 );
and ( n63877 , n63876 , n31002 );
and ( n63878 , n26193 , n34607 );
or ( n63879 , n63861 , n63865 , n63869 , n63873 , n63877 , n63878 );
and ( n63880 , n63857 , n63879 );
and ( n63881 , n26193 , n24800 );
or ( n63882 , n63880 , n63881 );
and ( n63883 , n63882 , n31008 );
and ( n63884 , n26193 , n10618 );
or ( n63885 , n63883 , n63884 );
buf ( n63886 , n63885 );
buf ( n63887 , n63886 );
not ( n63888 , n24800 );
and ( n63889 , n45549 , n28586 );
and ( n63890 , n25987 , n34573 );
or ( n63891 , n63889 , n63890 );
and ( n63892 , n63891 , n28594 );
and ( n63893 , n45559 , n28586 );
and ( n63894 , n25987 , n34573 );
or ( n63895 , n63893 , n63894 );
and ( n63896 , n63895 , n30269 );
and ( n63897 , n45569 , n28586 );
and ( n63898 , n25987 , n34573 );
or ( n63899 , n63897 , n63898 );
and ( n63900 , n63899 , n30982 );
and ( n63901 , n29595 , n28586 );
and ( n63902 , n25987 , n34573 );
or ( n63903 , n63901 , n63902 );
and ( n63904 , n63903 , n30989 );
and ( n63905 , n45580 , n28586 );
and ( n63906 , n25987 , n34573 );
or ( n63907 , n63905 , n63906 );
and ( n63908 , n63907 , n31002 );
and ( n63909 , n25987 , n34607 );
or ( n63910 , n63892 , n63896 , n63900 , n63904 , n63908 , n63909 );
and ( n63911 , n63888 , n63910 );
and ( n63912 , n25987 , n24800 );
or ( n63913 , n63911 , n63912 );
and ( n63914 , n63913 , n31008 );
and ( n63915 , n25987 , n10618 );
or ( n63916 , n63914 , n63915 );
buf ( n63917 , n63916 );
buf ( n63918 , n63917 );
buf ( n63919 , n10613 );
not ( n63920 , n34821 );
and ( n63921 , n13289 , n14592 );
and ( n63922 , n51156 , n36348 );
and ( n63923 , n13289 , n43530 );
or ( n63924 , n63922 , n63923 );
and ( n63925 , n63924 , n14562 );
and ( n63926 , n51166 , n36347 );
and ( n63927 , n13289 , n43543 );
or ( n63928 , n63926 , n63927 );
and ( n63929 , n63928 , n14586 );
and ( n63930 , n51176 , n36348 );
and ( n63931 , n13289 , n43556 );
or ( n63932 , n63930 , n63931 );
and ( n63933 , n63932 , n14584 );
and ( n63934 , n51166 , n36347 );
and ( n63935 , n13289 , n43563 );
or ( n63936 , n63934 , n63935 );
and ( n63937 , n63936 , n37835 );
and ( n63938 , n51176 , n36347 );
and ( n63939 , n13289 , n43563 );
or ( n63940 , n63938 , n63939 );
and ( n63941 , n63940 , n37841 );
and ( n63942 , n13287 , n14564 );
and ( n63943 , n15493 , n36347 );
and ( n63944 , n13289 , n43563 );
or ( n63945 , n63943 , n63944 );
and ( n63946 , n63945 , n37847 );
or ( n63947 , n63921 , n63925 , n63929 , n63933 , n63937 , n63941 , n63942 , n63946 );
or ( n63948 , n63920 , n63947 );
or ( n63949 , n13289 , n34821 );
or ( n63950 , n63948 , n63949 );
and ( n63951 , n63950 , n16574 );
and ( n63952 , n13289 , n16576 );
or ( n63953 , n63951 , n63952 );
buf ( n63954 , n63953 );
buf ( n63955 , n63954 );
buf ( n63956 , n10615 );
not ( n63957 , n17451 );
and ( n63958 , n46858 , n21334 );
and ( n63959 , n18811 , n34492 );
or ( n63960 , n63958 , n63959 );
and ( n63961 , n63960 , n21341 );
and ( n63962 , n46868 , n21334 );
and ( n63963 , n18811 , n34492 );
or ( n63964 , n63962 , n63963 );
and ( n63965 , n63964 , n23064 );
and ( n63966 , n46878 , n21334 );
and ( n63967 , n18811 , n34492 );
or ( n63968 , n63966 , n63967 );
and ( n63969 , n63968 , n23825 );
and ( n63970 , n22242 , n21334 );
and ( n63971 , n18811 , n34492 );
or ( n63972 , n63970 , n63971 );
and ( n63973 , n63972 , n23832 );
and ( n63974 , n46888 , n21334 );
and ( n63975 , n18811 , n34492 );
or ( n63976 , n63974 , n63975 );
and ( n63977 , n63976 , n23917 );
and ( n63978 , n18811 , n34526 );
or ( n63979 , n63961 , n63965 , n63969 , n63973 , n63977 , n63978 );
and ( n63980 , n63957 , n63979 );
and ( n63981 , n18811 , n17451 );
or ( n63982 , n63980 , n63981 );
and ( n63983 , n63982 , n23924 );
and ( n63984 , n18811 , n23926 );
or ( n63985 , n63983 , n63984 );
buf ( n63986 , n63985 );
buf ( n63987 , n63986 );
buf ( n63988 , n10613 );
buf ( n63989 , n10615 );
and ( n63990 , n16900 , n23924 );
and ( n63991 , n21351 , n23926 );
or ( n63992 , n63990 , n63991 );
buf ( n63993 , n63992 );
buf ( n63994 , n63993 );
not ( n63995 , n34821 );
and ( n63996 , n36271 , n36347 );
and ( n63997 , n13411 , n39408 );
or ( n63998 , n63996 , n63997 );
and ( n63999 , n63998 , n14562 );
and ( n64000 , n37069 , n36348 );
and ( n64001 , n13411 , n39427 );
or ( n64002 , n64000 , n64001 );
and ( n64003 , n64002 , n14586 );
and ( n64004 , n37822 , n36347 );
and ( n64005 , n13411 , n39446 );
or ( n64006 , n64004 , n64005 );
and ( n64007 , n64006 , n14584 );
and ( n64008 , n37069 , n36348 );
and ( n64009 , n13411 , n39453 );
or ( n64010 , n64008 , n64009 );
and ( n64011 , n64010 , n37835 );
and ( n64012 , n37822 , n36348 );
and ( n64013 , n13411 , n39453 );
or ( n64014 , n64012 , n64013 );
and ( n64015 , n64014 , n37841 );
and ( n64016 , n15713 , n36348 );
and ( n64017 , n13411 , n39453 );
or ( n64018 , n64016 , n64017 );
and ( n64019 , n64018 , n37847 );
and ( n64020 , n13411 , n37849 );
or ( n64021 , n63999 , n64003 , n64007 , n64011 , n64015 , n64019 , n64020 );
and ( n64022 , n63995 , n64021 );
and ( n64023 , n13411 , n34821 );
or ( n64024 , n64022 , n64023 );
and ( n64025 , n64024 , n16574 );
and ( n64026 , n13411 , n16576 );
or ( n64027 , n64025 , n64026 );
buf ( n64028 , n64027 );
buf ( n64029 , n64028 );
and ( n64030 , n11665 , n16574 );
and ( n64031 , n15770 , n16576 );
or ( n64032 , n64030 , n64031 );
buf ( n64033 , n64032 );
buf ( n64034 , n64033 );
buf ( n64035 , n10615 );
not ( n64036 , n34821 );
and ( n64037 , n55549 , n36345 );
and ( n64038 , n13160 , n36352 );
or ( n64039 , n64037 , n64038 );
and ( n64040 , n64039 , n14562 );
and ( n64041 , n55559 , n36345 );
and ( n64042 , n13160 , n37073 );
or ( n64043 , n64041 , n64042 );
and ( n64044 , n64043 , n14586 );
and ( n64045 , n55569 , n36350 );
and ( n64046 , n13160 , n37825 );
or ( n64047 , n64045 , n64046 );
and ( n64048 , n64047 , n14584 );
and ( n64049 , n55559 , n36350 );
and ( n64050 , n13160 , n37831 );
or ( n64051 , n64049 , n64050 );
and ( n64052 , n64051 , n37835 );
and ( n64053 , n55569 , n36350 );
and ( n64054 , n13160 , n37831 );
or ( n64055 , n64053 , n64054 );
and ( n64056 , n64055 , n37841 );
and ( n64057 , n14992 , n36350 );
and ( n64058 , n13160 , n37831 );
or ( n64059 , n64057 , n64058 );
and ( n64060 , n64059 , n37847 );
and ( n64061 , n13160 , n37849 );
or ( n64062 , n64040 , n64044 , n64048 , n64052 , n64056 , n64060 , n64061 );
and ( n64063 , n64036 , n64062 );
and ( n64064 , n13160 , n34821 );
or ( n64065 , n64063 , n64064 );
and ( n64066 , n64065 , n16574 );
and ( n64067 , n13160 , n16576 );
or ( n64068 , n64066 , n64067 );
buf ( n64069 , n64068 );
buf ( n64070 , n64069 );
not ( n64071 , n34821 );
and ( n64072 , n13215 , n14592 );
and ( n64073 , n57550 , n36350 );
and ( n64074 , n13215 , n43691 );
or ( n64075 , n64073 , n64074 );
and ( n64076 , n64075 , n14562 );
and ( n64077 , n57560 , n36350 );
and ( n64078 , n13215 , n43703 );
or ( n64079 , n64077 , n64078 );
and ( n64080 , n64079 , n14586 );
and ( n64081 , n57570 , n36345 );
and ( n64082 , n13215 , n43715 );
or ( n64083 , n64081 , n64082 );
and ( n64084 , n64083 , n14584 );
and ( n64085 , n57560 , n36345 );
and ( n64086 , n13215 , n43721 );
or ( n64087 , n64085 , n64086 );
and ( n64088 , n64087 , n37835 );
and ( n64089 , n57570 , n36345 );
and ( n64090 , n13215 , n43721 );
or ( n64091 , n64089 , n64090 );
and ( n64092 , n64091 , n37841 );
and ( n64093 , n15067 , n14564 );
and ( n64094 , n15067 , n36345 );
and ( n64095 , n13215 , n43721 );
or ( n64096 , n64094 , n64095 );
and ( n64097 , n64096 , n37847 );
or ( n64098 , n64072 , n64076 , n64080 , n64084 , n64088 , n64092 , n64093 , n64097 );
and ( n64099 , n64071 , n64098 );
and ( n64100 , n13215 , n34821 );
or ( n64101 , n64099 , n64100 );
and ( n64102 , n64101 , n16574 );
and ( n64103 , n12264 , n16576 );
or ( n64104 , n64102 , n64103 );
buf ( n64105 , n64104 );
buf ( n64106 , n64105 );
buf ( n64107 , n10615 );
buf ( n64108 , n10615 );
buf ( n64109 , n10615 );
buf ( n64110 , n10613 );
buf ( n64111 , n10615 );
not ( n64112 , n24800 );
and ( n64113 , n56393 , n28586 );
and ( n64114 , n27177 , n34573 );
or ( n64115 , n64113 , n64114 );
and ( n64116 , n64115 , n28594 );
and ( n64117 , n56402 , n28586 );
and ( n64118 , n27177 , n34573 );
or ( n64119 , n64117 , n64118 );
and ( n64120 , n64119 , n30269 );
and ( n64121 , n56411 , n28586 );
and ( n64122 , n27177 , n34573 );
or ( n64123 , n64121 , n64122 );
and ( n64124 , n64123 , n30982 );
and ( n64125 , n29107 , n28586 );
and ( n64126 , n27177 , n34573 );
or ( n64127 , n64125 , n64126 );
and ( n64128 , n64127 , n30989 );
and ( n64129 , n56421 , n28586 );
and ( n64130 , n27177 , n34573 );
or ( n64131 , n64129 , n64130 );
and ( n64132 , n64131 , n31002 );
and ( n64133 , n27177 , n34607 );
or ( n64134 , n64116 , n64120 , n64124 , n64128 , n64132 , n64133 );
and ( n64135 , n64112 , n64134 );
and ( n64136 , n27177 , n24800 );
or ( n64137 , n64135 , n64136 );
and ( n64138 , n64137 , n31008 );
and ( n64139 , n27177 , n10618 );
or ( n64140 , n64138 , n64139 );
buf ( n64141 , n64140 );
buf ( n64142 , n64141 );
buf ( n64143 , n10615 );
buf ( n64144 , n10615 );
buf ( n64145 , n10615 );
not ( n64146 , n17162 );
not ( n64147 , n17450 );
and ( n64148 , n10703 , n37947 );
not ( n64149 , n38425 );
and ( n64150 , n64149 , n38200 );
xor ( n64151 , n38434 , n38446 );
and ( n64152 , n64151 , n38425 );
xor ( n64153 , n64150 , n64152 );
not ( n64154 , n64153 );
and ( n64155 , n64154 , n19745 );
not ( n64156 , n38934 );
and ( n64157 , n64156 , n38709 );
xor ( n64158 , n38943 , n38955 );
and ( n64159 , n64158 , n38934 );
or ( n64160 , n64157 , n64159 );
buf ( n64161 , n64160 );
and ( n64162 , n64161 , n19748 );
and ( n64163 , n22300 , n21253 );
and ( n64164 , n10703 , n21255 );
or ( n64165 , n64155 , n64162 , n64163 , n64164 );
and ( n64166 , n64165 , n38980 );
or ( n64167 , n64148 , n64166 );
and ( n64168 , n64147 , n64167 );
or ( n64169 , n64168 , C0 );
and ( n64170 , n64146 , n64169 );
and ( n64171 , n64165 , n17162 );
or ( n64172 , n64170 , n64171 );
and ( n64173 , n64172 , n23924 );
not ( n64174 , n39264 );
and ( n64175 , n64174 , n39078 );
xor ( n64176 , n39273 , n39285 );
and ( n64177 , n64176 , n39264 );
or ( n64178 , n64175 , n64177 );
buf ( n64179 , n64178 );
and ( n64180 , n64179 , n23926 );
or ( n64181 , n64173 , n64180 );
buf ( n64182 , n64181 );
buf ( n64183 , n64182 );
buf ( n64184 , n10615 );
buf ( n64185 , n10615 );
buf ( n64186 , n10613 );
buf ( n64187 , n10613 );
buf ( n64188 , n10613 );
buf ( n64189 , n10613 );
buf ( n64190 , n10615 );
buf ( n64191 , n10613 );
buf ( n64192 , n10613 );
and ( n64193 , n24357 , n31008 );
and ( n64194 , n29157 , n10618 );
or ( n64195 , n64193 , n64194 );
buf ( n64196 , n64195 );
buf ( n64197 , n64196 );
not ( n64198 , n11954 );
not ( n64199 , n12243 );
and ( n64200 , n10893 , n31187 );
not ( n64201 , n31697 );
and ( n64202 , n64201 , n31489 );
xor ( n64203 , n50359 , n50372 );
and ( n64204 , n64203 , n31697 );
or ( n64205 , n64202 , n64204 );
buf ( n64206 , n64205 );
and ( n64207 , n64206 , n14140 );
not ( n64208 , n32214 );
and ( n64209 , n64208 , n32006 );
xor ( n64210 , n50386 , n50399 );
and ( n64211 , n64210 , n32214 );
or ( n64212 , n64209 , n64211 );
buf ( n64213 , n64212 );
and ( n64214 , n64213 , n14137 );
and ( n64215 , n15711 , n14143 );
and ( n64216 , n10893 , n14141 );
or ( n64217 , n64207 , n64214 , n64215 , n64216 );
and ( n64218 , n64217 , n32236 );
or ( n64219 , n64200 , n64218 );
and ( n64220 , n64199 , n64219 );
not ( n64221 , n34038 );
and ( n64222 , n64221 , n33746 );
xor ( n64223 , n50419 , n50432 );
and ( n64224 , n64223 , n34038 );
or ( n64225 , n64222 , n64224 );
buf ( n64226 , n64225 );
and ( n64227 , n64226 , n12243 );
or ( n64228 , n64220 , n64227 );
and ( n64229 , n64198 , n64228 );
and ( n64230 , n64217 , n11954 );
or ( n64231 , n64229 , n64230 );
and ( n64232 , n64231 , n16574 );
not ( n64233 , n34327 );
and ( n64234 , n64233 , n34155 );
xor ( n64235 , n50451 , n50464 );
and ( n64236 , n64235 , n34327 );
or ( n64237 , n64234 , n64236 );
buf ( n64238 , n64237 );
and ( n64239 , n64238 , n16576 );
or ( n64240 , n64232 , n64239 );
buf ( n64241 , n64240 );
buf ( n64242 , n64241 );
not ( n64243 , n34821 );
and ( n64244 , n13433 , n14592 );
and ( n64245 , n59483 , n36348 );
and ( n64246 , n13433 , n43530 );
or ( n64247 , n64245 , n64246 );
and ( n64248 , n64247 , n14562 );
and ( n64249 , n59493 , n36347 );
and ( n64250 , n13433 , n43543 );
or ( n64251 , n64249 , n64250 );
and ( n64252 , n64251 , n14586 );
and ( n64253 , n59503 , n36348 );
and ( n64254 , n13433 , n43556 );
or ( n64255 , n64253 , n64254 );
and ( n64256 , n64255 , n14584 );
and ( n64257 , n59493 , n36347 );
and ( n64258 , n13433 , n43563 );
or ( n64259 , n64257 , n64258 );
and ( n64260 , n64259 , n37835 );
and ( n64261 , n59503 , n36347 );
and ( n64262 , n13433 , n43563 );
or ( n64263 , n64261 , n64262 );
and ( n64264 , n64263 , n37841 );
and ( n64265 , n13431 , n14564 );
and ( n64266 , n15757 , n36347 );
and ( n64267 , n13433 , n43563 );
or ( n64268 , n64266 , n64267 );
and ( n64269 , n64268 , n37847 );
or ( n64270 , n64244 , n64248 , n64252 , n64256 , n64260 , n64264 , n64265 , n64269 );
and ( n64271 , n64243 , n64270 );
and ( n64272 , n13433 , n34821 );
or ( n64273 , n64271 , n64272 );
and ( n64274 , n64273 , n16574 );
and ( n64275 , n13433 , n16576 );
or ( n64276 , n64274 , n64275 );
buf ( n64277 , n64276 );
buf ( n64278 , n64277 );
buf ( n64279 , n10613 );
not ( n64280 , n24800 );
and ( n64281 , n26017 , n25222 );
and ( n64282 , n39803 , n28589 );
and ( n64283 , n26017 , n31075 );
or ( n64284 , n64282 , n64283 );
and ( n64285 , n64284 , n28594 );
and ( n64286 , n39816 , n28589 );
and ( n64287 , n26017 , n31075 );
or ( n64288 , n64286 , n64287 );
and ( n64289 , n64288 , n30269 );
and ( n64290 , n39826 , n28589 );
and ( n64291 , n26017 , n31075 );
or ( n64292 , n64290 , n64291 );
and ( n64293 , n64292 , n30982 );
and ( n64294 , n29575 , n28589 );
and ( n64295 , n26017 , n31075 );
or ( n64296 , n64294 , n64295 );
and ( n64297 , n64296 , n30989 );
and ( n64298 , n29575 , n30991 );
and ( n64299 , n39836 , n28589 );
and ( n64300 , n26017 , n31075 );
or ( n64301 , n64299 , n64300 );
and ( n64302 , n64301 , n31002 );
or ( n64303 , n64281 , n64285 , n64289 , n64293 , n64297 , n64298 , n64302 );
and ( n64304 , n64280 , n64303 );
and ( n64305 , n26017 , n24800 );
or ( n64306 , n64304 , n64305 );
and ( n64307 , n64306 , n31008 );
and ( n64308 , n25294 , n10618 );
or ( n64309 , n64307 , n64308 );
buf ( n64310 , n64309 );
buf ( n64311 , n64310 );
not ( n64312 , n34821 );
and ( n64313 , n13359 , n14592 );
and ( n64314 , n45647 , n36350 );
and ( n64315 , n13359 , n43691 );
or ( n64316 , n64314 , n64315 );
and ( n64317 , n64316 , n14562 );
and ( n64318 , n45657 , n36350 );
and ( n64319 , n13359 , n43703 );
or ( n64320 , n64318 , n64319 );
and ( n64321 , n64320 , n14586 );
and ( n64322 , n45667 , n36345 );
and ( n64323 , n13359 , n43715 );
or ( n64324 , n64322 , n64323 );
and ( n64325 , n64324 , n14584 );
and ( n64326 , n45657 , n36345 );
and ( n64327 , n13359 , n43721 );
or ( n64328 , n64326 , n64327 );
and ( n64329 , n64328 , n37835 );
and ( n64330 , n45667 , n36345 );
and ( n64331 , n13359 , n43721 );
or ( n64332 , n64330 , n64331 );
and ( n64333 , n64332 , n37841 );
and ( n64334 , n15625 , n14564 );
and ( n64335 , n15625 , n36345 );
and ( n64336 , n13359 , n43721 );
or ( n64337 , n64335 , n64336 );
and ( n64338 , n64337 , n37847 );
or ( n64339 , n64313 , n64317 , n64321 , n64325 , n64329 , n64333 , n64334 , n64338 );
and ( n64340 , n64312 , n64339 );
and ( n64341 , n13359 , n34821 );
or ( n64342 , n64340 , n64341 );
and ( n64343 , n64342 , n16574 );
and ( n64344 , n12300 , n16576 );
or ( n64345 , n64343 , n64344 );
buf ( n64346 , n64345 );
buf ( n64347 , n64346 );
not ( n64348 , n17451 );
and ( n64349 , n58841 , n21333 );
and ( n64350 , n19013 , n34758 );
or ( n64351 , n64349 , n64350 );
and ( n64352 , n64351 , n21341 );
and ( n64353 , n58851 , n21333 );
and ( n64354 , n19013 , n34758 );
or ( n64355 , n64353 , n64354 );
and ( n64356 , n64355 , n23064 );
and ( n64357 , n58861 , n21333 );
and ( n64358 , n19013 , n34758 );
or ( n64359 , n64357 , n64358 );
and ( n64360 , n64359 , n23825 );
and ( n64361 , n22122 , n21333 );
and ( n64362 , n19013 , n34758 );
or ( n64363 , n64361 , n64362 );
and ( n64364 , n64363 , n23832 );
and ( n64365 , n58872 , n21333 );
and ( n64366 , n19013 , n34758 );
or ( n64367 , n64365 , n64366 );
and ( n64368 , n64367 , n23917 );
and ( n64369 , n19013 , n34526 );
or ( n64370 , n64352 , n64356 , n64360 , n64364 , n64368 , n64369 );
and ( n64371 , n64348 , n64370 );
and ( n64372 , n19013 , n17451 );
or ( n64373 , n64371 , n64372 );
and ( n64374 , n64373 , n23924 );
and ( n64375 , n19013 , n23926 );
or ( n64376 , n64374 , n64375 );
buf ( n64377 , n64376 );
buf ( n64378 , n64377 );
buf ( n64379 , n10613 );
buf ( n64380 , n10613 );
buf ( n64381 , n10615 );
buf ( n64382 , n10615 );
not ( n64383 , n11954 );
not ( n64384 , n12243 );
and ( n64385 , n10909 , n31187 );
not ( n64386 , n31697 );
and ( n64387 , n64386 , n31455 );
xor ( n64388 , n50361 , n50370 );
and ( n64389 , n64388 , n31697 );
or ( n64390 , n64387 , n64389 );
buf ( n64391 , n64390 );
and ( n64392 , n64391 , n14140 );
not ( n64393 , n32214 );
and ( n64394 , n64393 , n31972 );
xor ( n64395 , n50388 , n50397 );
and ( n64396 , n64395 , n32214 );
or ( n64397 , n64394 , n64396 );
buf ( n64398 , n64397 );
and ( n64399 , n64398 , n14137 );
and ( n64400 , n15755 , n14143 );
and ( n64401 , n10909 , n14141 );
or ( n64402 , n64392 , n64399 , n64400 , n64401 );
and ( n64403 , n64402 , n32236 );
or ( n64404 , n64385 , n64403 );
and ( n64405 , n64384 , n64404 );
not ( n64406 , n34038 );
and ( n64407 , n64406 , n33698 );
xor ( n64408 , n50421 , n50430 );
and ( n64409 , n64408 , n34038 );
or ( n64410 , n64407 , n64409 );
buf ( n64411 , n64410 );
and ( n64412 , n64411 , n12243 );
or ( n64413 , n64405 , n64412 );
and ( n64414 , n64383 , n64413 );
and ( n64415 , n64402 , n11954 );
or ( n64416 , n64414 , n64415 );
and ( n64417 , n64416 , n16574 );
not ( n64418 , n34327 );
and ( n64419 , n64418 , n34127 );
xor ( n64420 , n50453 , n50462 );
and ( n64421 , n64420 , n34327 );
or ( n64422 , n64419 , n64421 );
buf ( n64423 , n64422 );
and ( n64424 , n64423 , n16576 );
or ( n64425 , n64417 , n64424 );
buf ( n64426 , n64425 );
buf ( n64427 , n64426 );
buf ( n64428 , n10615 );
buf ( n64429 , n10613 );
buf ( n64430 , n10615 );
not ( n64431 , n17451 );
and ( n64432 , n47363 , n21334 );
and ( n64433 , n18641 , n34492 );
or ( n64434 , n64432 , n64433 );
and ( n64435 , n64434 , n21341 );
and ( n64436 , n47373 , n21334 );
and ( n64437 , n18641 , n34492 );
or ( n64438 , n64436 , n64437 );
and ( n64439 , n64438 , n23064 );
and ( n64440 , n47383 , n21334 );
and ( n64441 , n18641 , n34492 );
or ( n64442 , n64440 , n64441 );
and ( n64443 , n64442 , n23825 );
and ( n64444 , n22342 , n21334 );
and ( n64445 , n18641 , n34492 );
or ( n64446 , n64444 , n64445 );
and ( n64447 , n64446 , n23832 );
and ( n64448 , n47394 , n21334 );
and ( n64449 , n18641 , n34492 );
or ( n64450 , n64448 , n64449 );
and ( n64451 , n64450 , n23917 );
and ( n64452 , n18641 , n34526 );
or ( n64453 , n64435 , n64439 , n64443 , n64447 , n64451 , n64452 );
and ( n64454 , n64431 , n64453 );
and ( n64455 , n18641 , n17451 );
or ( n64456 , n64454 , n64455 );
and ( n64457 , n64456 , n23924 );
and ( n64458 , n18641 , n23926 );
or ( n64459 , n64457 , n64458 );
buf ( n64460 , n64459 );
buf ( n64461 , n64460 );
and ( n64462 , n11569 , n16574 );
and ( n64463 , n15506 , n16576 );
or ( n64464 , n64462 , n64463 );
buf ( n64465 , n64464 );
buf ( n64466 , n64465 );
buf ( n64467 , n10613 );
buf ( n64468 , n10615 );
not ( n64469 , n24800 );
and ( n64470 , n26765 , n25222 );
and ( n64471 , n52160 , n28589 );
and ( n64472 , n26765 , n31075 );
or ( n64473 , n64471 , n64472 );
and ( n64474 , n64473 , n28594 );
and ( n64475 , n52170 , n28589 );
and ( n64476 , n26765 , n31075 );
or ( n64477 , n64475 , n64476 );
and ( n64478 , n64477 , n30269 );
and ( n64479 , n52180 , n28589 );
and ( n64480 , n26765 , n31075 );
or ( n64481 , n64479 , n64480 );
and ( n64482 , n64481 , n30982 );
and ( n64483 , n29146 , n28589 );
and ( n64484 , n26765 , n31075 );
or ( n64485 , n64483 , n64484 );
and ( n64486 , n64485 , n30989 );
and ( n64487 , n29146 , n30991 );
and ( n64488 , n52191 , n28589 );
and ( n64489 , n26765 , n31075 );
or ( n64490 , n64488 , n64489 );
and ( n64491 , n64490 , n31002 );
or ( n64492 , n64470 , n64474 , n64478 , n64482 , n64486 , n64487 , n64491 );
and ( n64493 , n64469 , n64492 );
and ( n64494 , n26765 , n24800 );
or ( n64495 , n64493 , n64494 );
and ( n64496 , n64495 , n31008 );
and ( n64497 , n25624 , n10618 );
or ( n64498 , n64496 , n64497 );
buf ( n64499 , n64498 );
buf ( n64500 , n64499 );
buf ( n64501 , n10615 );
buf ( n64502 , n10615 );
buf ( n64503 , n10615 );
not ( n64504 , n17451 );
and ( n64505 , n42746 , n21333 );
and ( n64506 , n18945 , n34758 );
or ( n64507 , n64505 , n64506 );
and ( n64508 , n64507 , n21341 );
and ( n64509 , n42756 , n21333 );
and ( n64510 , n18945 , n34758 );
or ( n64511 , n64509 , n64510 );
and ( n64512 , n64511 , n23064 );
and ( n64513 , n42766 , n21333 );
and ( n64514 , n18945 , n34758 );
or ( n64515 , n64513 , n64514 );
and ( n64516 , n64515 , n23825 );
and ( n64517 , n22162 , n21333 );
and ( n64518 , n18945 , n34758 );
or ( n64519 , n64517 , n64518 );
and ( n64520 , n64519 , n23832 );
and ( n64521 , n42776 , n21333 );
and ( n64522 , n18945 , n34758 );
or ( n64523 , n64521 , n64522 );
and ( n64524 , n64523 , n23917 );
and ( n64525 , n18945 , n34526 );
or ( n64526 , n64508 , n64512 , n64516 , n64520 , n64524 , n64525 );
and ( n64527 , n64504 , n64526 );
and ( n64528 , n18945 , n17451 );
or ( n64529 , n64527 , n64528 );
and ( n64530 , n64529 , n23924 );
and ( n64531 , n18945 , n23926 );
or ( n64532 , n64530 , n64531 );
buf ( n64533 , n64532 );
buf ( n64534 , n64533 );
buf ( n64535 , n10613 );
not ( n64536 , n24800 );
and ( n64537 , n27187 , n25222 );
and ( n64538 , n55800 , n28583 );
and ( n64539 , n27187 , n28591 );
or ( n64540 , n64538 , n64539 );
and ( n64541 , n64540 , n28594 );
and ( n64542 , n55812 , n28583 );
and ( n64543 , n27187 , n28591 );
or ( n64544 , n64542 , n64543 );
and ( n64545 , n64544 , n30269 );
and ( n64546 , n55824 , n28583 );
and ( n64547 , n27187 , n28591 );
or ( n64548 , n64546 , n64547 );
and ( n64549 , n64548 , n30982 );
and ( n64550 , n29120 , n28583 );
and ( n64551 , n27187 , n28591 );
or ( n64552 , n64550 , n64551 );
and ( n64553 , n64552 , n30989 );
and ( n64554 , n27185 , n30991 );
and ( n64555 , n55834 , n28583 );
and ( n64556 , n27187 , n28591 );
or ( n64557 , n64555 , n64556 );
and ( n64558 , n64557 , n31002 );
or ( n64559 , n64537 , n64541 , n64545 , n64549 , n64553 , n64554 , n64558 );
and ( n64560 , n64536 , n64559 );
and ( n64561 , n27187 , n24800 );
or ( n64562 , n64560 , n64561 );
and ( n64563 , n64562 , n31008 );
and ( n64564 , n27187 , n10618 );
or ( n64565 , n64563 , n64564 );
buf ( n64566 , n64565 );
buf ( n64567 , n64566 );
buf ( n64568 , n10615 );
not ( n64569 , n34821 );
and ( n64570 , n57550 , n36347 );
and ( n64571 , n13219 , n39408 );
or ( n64572 , n64570 , n64571 );
and ( n64573 , n64572 , n14562 );
and ( n64574 , n57560 , n36348 );
and ( n64575 , n13219 , n39427 );
or ( n64576 , n64574 , n64575 );
and ( n64577 , n64576 , n14586 );
and ( n64578 , n57570 , n36347 );
and ( n64579 , n13219 , n39446 );
or ( n64580 , n64578 , n64579 );
and ( n64581 , n64580 , n14584 );
and ( n64582 , n57560 , n36348 );
and ( n64583 , n13219 , n39453 );
or ( n64584 , n64582 , n64583 );
and ( n64585 , n64584 , n37835 );
and ( n64586 , n57570 , n36348 );
and ( n64587 , n13219 , n39453 );
or ( n64588 , n64586 , n64587 );
and ( n64589 , n64588 , n37841 );
and ( n64590 , n15067 , n36348 );
and ( n64591 , n13219 , n39453 );
or ( n64592 , n64590 , n64591 );
and ( n64593 , n64592 , n37847 );
and ( n64594 , n13219 , n37849 );
or ( n64595 , n64573 , n64577 , n64581 , n64585 , n64589 , n64593 , n64594 );
and ( n64596 , n64569 , n64595 );
and ( n64597 , n13219 , n34821 );
or ( n64598 , n64596 , n64597 );
and ( n64599 , n64598 , n16574 );
and ( n64600 , n13219 , n16576 );
or ( n64601 , n64599 , n64600 );
buf ( n64602 , n64601 );
buf ( n64603 , n64602 );
buf ( n64604 , n10613 );
buf ( n64605 , n10615 );
buf ( n64606 , n10615 );
and ( n64607 , n24373 , n31008 );
and ( n64608 , n29183 , n10618 );
or ( n64609 , n64607 , n64608 );
buf ( n64610 , n64609 );
buf ( n64611 , n64610 );
buf ( n64612 , n10613 );
buf ( n64613 , n10613 );
buf ( n64614 , n10615 );
not ( n64615 , n24800 );
and ( n64616 , n27175 , n25222 );
and ( n64617 , n56393 , n28583 );
and ( n64618 , n27175 , n28591 );
or ( n64619 , n64617 , n64618 );
and ( n64620 , n64619 , n28594 );
and ( n64621 , n56402 , n28583 );
and ( n64622 , n27175 , n28591 );
or ( n64623 , n64621 , n64622 );
and ( n64624 , n64623 , n30269 );
and ( n64625 , n56411 , n28583 );
and ( n64626 , n27175 , n28591 );
or ( n64627 , n64625 , n64626 );
and ( n64628 , n64627 , n30982 );
and ( n64629 , n29107 , n28583 );
and ( n64630 , n27175 , n28591 );
or ( n64631 , n64629 , n64630 );
and ( n64632 , n64631 , n30989 );
and ( n64633 , n27173 , n30991 );
and ( n64634 , n56421 , n28583 );
and ( n64635 , n27175 , n28591 );
or ( n64636 , n64634 , n64635 );
and ( n64637 , n64636 , n31002 );
or ( n64638 , n64616 , n64620 , n64624 , n64628 , n64632 , n64633 , n64637 );
and ( n64639 , n64615 , n64638 );
and ( n64640 , n27175 , n24800 );
or ( n64641 , n64639 , n64640 );
and ( n64642 , n64641 , n31008 );
and ( n64643 , n27175 , n10618 );
or ( n64644 , n64642 , n64643 );
buf ( n64645 , n64644 );
buf ( n64646 , n64645 );
buf ( n64647 , n10613 );
not ( n64648 , n34538 );
and ( n64649 , n64648 , n20496 );
and ( n64650 , n14657 , n34538 );
or ( n64651 , n64649 , n64650 );
and ( n64652 , n64651 , n23924 );
and ( n64653 , n14657 , n23926 );
or ( n64654 , n64652 , n64653 );
buf ( n64655 , n64654 );
buf ( n64656 , n64655 );
buf ( n64657 , n10613 );
buf ( n64658 , n10615 );
buf ( n64659 , n10615 );
buf ( n64660 , n10613 );
not ( n64661 , n11954 );
not ( n64662 , n12243 );
and ( n64663 , n10901 , n31187 );
not ( n64664 , n31697 );
and ( n64665 , n64664 , n31472 );
xor ( n64666 , n50360 , n50371 );
and ( n64667 , n64666 , n31697 );
or ( n64668 , n64665 , n64667 );
buf ( n64669 , n64668 );
and ( n64670 , n64669 , n14140 );
not ( n64671 , n32214 );
and ( n64672 , n64671 , n31989 );
xor ( n64673 , n50387 , n50398 );
and ( n64674 , n64673 , n32214 );
or ( n64675 , n64672 , n64674 );
buf ( n64676 , n64675 );
and ( n64677 , n64676 , n14137 );
and ( n64678 , n15733 , n14143 );
and ( n64679 , n10901 , n14141 );
or ( n64680 , n64670 , n64677 , n64678 , n64679 );
and ( n64681 , n64680 , n32236 );
or ( n64682 , n64663 , n64681 );
and ( n64683 , n64662 , n64682 );
not ( n64684 , n34038 );
and ( n64685 , n64684 , n33722 );
xor ( n64686 , n50420 , n50431 );
and ( n64687 , n64686 , n34038 );
or ( n64688 , n64685 , n64687 );
buf ( n64689 , n64688 );
and ( n64690 , n64689 , n12243 );
or ( n64691 , n64683 , n64690 );
and ( n64692 , n64661 , n64691 );
and ( n64693 , n64680 , n11954 );
or ( n64694 , n64692 , n64693 );
and ( n64695 , n64694 , n16574 );
not ( n64696 , n34327 );
and ( n64697 , n64696 , n34141 );
xor ( n64698 , n50452 , n50463 );
and ( n64699 , n64698 , n34327 );
or ( n64700 , n64697 , n64699 );
buf ( n64701 , n64700 );
and ( n64702 , n64701 , n16576 );
or ( n64703 , n64695 , n64702 );
buf ( n64704 , n64703 );
buf ( n64705 , n64704 );
buf ( n64706 , n10613 );
buf ( n64707 , n10615 );
not ( n64708 , n17451 );
and ( n64709 , n49126 , n21333 );
and ( n64710 , n18979 , n34758 );
or ( n64711 , n64709 , n64710 );
and ( n64712 , n64711 , n21341 );
and ( n64713 , n49136 , n21333 );
and ( n64714 , n18979 , n34758 );
or ( n64715 , n64713 , n64714 );
and ( n64716 , n64715 , n23064 );
and ( n64717 , n49146 , n21333 );
and ( n64718 , n18979 , n34758 );
or ( n64719 , n64717 , n64718 );
and ( n64720 , n64719 , n23825 );
and ( n64721 , n22142 , n21333 );
and ( n64722 , n18979 , n34758 );
or ( n64723 , n64721 , n64722 );
and ( n64724 , n64723 , n23832 );
and ( n64725 , n49157 , n21333 );
and ( n64726 , n18979 , n34758 );
or ( n64727 , n64725 , n64726 );
and ( n64728 , n64727 , n23917 );
and ( n64729 , n18979 , n34526 );
or ( n64730 , n64712 , n64716 , n64720 , n64724 , n64728 , n64729 );
and ( n64731 , n64708 , n64730 );
and ( n64732 , n18979 , n17451 );
or ( n64733 , n64731 , n64732 );
and ( n64734 , n64733 , n23924 );
and ( n64735 , n18979 , n23926 );
or ( n64736 , n64734 , n64735 );
buf ( n64737 , n64736 );
buf ( n64738 , n64737 );
buf ( n64739 , n10615 );
buf ( n64740 , n10613 );
buf ( n64741 , n10615 );
and ( n64742 , n24102 , n31008 );
and ( n64743 , n29248 , n10618 );
or ( n64744 , n64742 , n64743 );
buf ( n64745 , n64744 );
buf ( n64746 , n64745 );
buf ( n64747 , n10613 );
buf ( n64748 , n10613 );
buf ( n64749 , n10615 );
buf ( n64750 , n10613 );
buf ( n64751 , n10613 );
not ( n64752 , n34804 );
and ( n64753 , n64752 , n25894 );
and ( n64754 , n14827 , n34804 );
or ( n64755 , n64753 , n64754 );
and ( n64756 , n64755 , n31008 );
and ( n64757 , n14827 , n10618 );
or ( n64758 , n64756 , n64757 );
buf ( n64759 , n64758 );
buf ( n64760 , n64759 );
buf ( n64761 , n10613 );
not ( n64762 , n17451 );
and ( n64763 , n49126 , n21334 );
and ( n64764 , n18981 , n34492 );
or ( n64765 , n64763 , n64764 );
and ( n64766 , n64765 , n21341 );
and ( n64767 , n49136 , n21334 );
and ( n64768 , n18981 , n34492 );
or ( n64769 , n64767 , n64768 );
and ( n64770 , n64769 , n23064 );
and ( n64771 , n49146 , n21334 );
and ( n64772 , n18981 , n34492 );
or ( n64773 , n64771 , n64772 );
and ( n64774 , n64773 , n23825 );
and ( n64775 , n22142 , n21334 );
and ( n64776 , n18981 , n34492 );
or ( n64777 , n64775 , n64776 );
and ( n64778 , n64777 , n23832 );
and ( n64779 , n49157 , n21334 );
and ( n64780 , n18981 , n34492 );
or ( n64781 , n64779 , n64780 );
and ( n64782 , n64781 , n23917 );
and ( n64783 , n18981 , n34526 );
or ( n64784 , n64766 , n64770 , n64774 , n64778 , n64782 , n64783 );
and ( n64785 , n64762 , n64784 );
and ( n64786 , n18981 , n17451 );
or ( n64787 , n64785 , n64786 );
and ( n64788 , n64787 , n23924 );
and ( n64789 , n18981 , n23926 );
or ( n64790 , n64788 , n64789 );
buf ( n64791 , n64790 );
buf ( n64792 , n64791 );
buf ( n64793 , n10615 );
not ( n64794 , n17451 );
and ( n64795 , n46760 , n21334 );
and ( n64796 , n19151 , n34492 );
or ( n64797 , n64795 , n64796 );
and ( n64798 , n64797 , n21341 );
and ( n64799 , n46770 , n21334 );
and ( n64800 , n19151 , n34492 );
or ( n64801 , n64799 , n64800 );
and ( n64802 , n64801 , n23064 );
and ( n64803 , n46780 , n21334 );
and ( n64804 , n19151 , n34492 );
or ( n64805 , n64803 , n64804 );
and ( n64806 , n64805 , n23825 );
and ( n64807 , n22042 , n21334 );
and ( n64808 , n19151 , n34492 );
or ( n64809 , n64807 , n64808 );
and ( n64810 , n64809 , n23832 );
and ( n64811 , n46791 , n21334 );
and ( n64812 , n19151 , n34492 );
or ( n64813 , n64811 , n64812 );
and ( n64814 , n64813 , n23917 );
and ( n64815 , n19151 , n34526 );
or ( n64816 , n64798 , n64802 , n64806 , n64810 , n64814 , n64815 );
and ( n64817 , n64794 , n64816 );
and ( n64818 , n19151 , n17451 );
or ( n64819 , n64817 , n64818 );
and ( n64820 , n64819 , n23924 );
and ( n64821 , n19151 , n23926 );
or ( n64822 , n64820 , n64821 );
buf ( n64823 , n64822 );
buf ( n64824 , n64823 );
buf ( n64825 , n10613 );
buf ( n64826 , n10615 );
buf ( n64827 , n10615 );
and ( n64828 , n24230 , n31008 );
and ( n64829 , n29606 , n10618 );
or ( n64830 , n64828 , n64829 );
buf ( n64831 , n64830 );
buf ( n64832 , n64831 );
not ( n64833 , n17451 );
and ( n64834 , n18839 , n17873 );
and ( n64835 , n34488 , n21336 );
and ( n64836 , n18839 , n42682 );
or ( n64837 , n64835 , n64836 );
and ( n64838 , n64837 , n21341 );
and ( n64839 , n34501 , n21336 );
and ( n64840 , n18839 , n42682 );
or ( n64841 , n64839 , n64840 );
and ( n64842 , n64841 , n23064 );
and ( n64843 , n34511 , n21336 );
and ( n64844 , n18839 , n42682 );
or ( n64845 , n64843 , n64844 );
and ( n64846 , n64845 , n23825 );
and ( n64847 , n22222 , n21336 );
and ( n64848 , n18839 , n42682 );
or ( n64849 , n64847 , n64848 );
and ( n64850 , n64849 , n23832 );
and ( n64851 , n22222 , n23834 );
and ( n64852 , n34521 , n21336 );
and ( n64853 , n18839 , n42682 );
or ( n64854 , n64852 , n64853 );
and ( n64855 , n64854 , n23917 );
or ( n64856 , n64834 , n64838 , n64842 , n64846 , n64850 , n64851 , n64855 );
and ( n64857 , n64833 , n64856 );
and ( n64858 , n18839 , n17451 );
or ( n64859 , n64857 , n64858 );
and ( n64860 , n64859 , n23924 );
and ( n64861 , n18020 , n23926 );
or ( n64862 , n64860 , n64861 );
buf ( n64863 , n64862 );
buf ( n64864 , n64863 );
buf ( n64865 , n10615 );
not ( n64866 , n17451 );
and ( n64867 , n18737 , n17873 );
and ( n64868 , n51973 , n21336 );
and ( n64869 , n18737 , n42682 );
or ( n64870 , n64868 , n64869 );
and ( n64871 , n64870 , n21341 );
and ( n64872 , n51983 , n21336 );
and ( n64873 , n18737 , n42682 );
or ( n64874 , n64872 , n64873 );
and ( n64875 , n64874 , n23064 );
and ( n64876 , n51993 , n21336 );
and ( n64877 , n18737 , n42682 );
or ( n64878 , n64876 , n64877 );
and ( n64879 , n64878 , n23825 );
and ( n64880 , n22282 , n21336 );
and ( n64881 , n18737 , n42682 );
or ( n64882 , n64880 , n64881 );
and ( n64883 , n64882 , n23832 );
and ( n64884 , n22282 , n23834 );
and ( n64885 , n52004 , n21336 );
and ( n64886 , n18737 , n42682 );
or ( n64887 , n64885 , n64886 );
and ( n64888 , n64887 , n23917 );
or ( n64889 , n64867 , n64871 , n64875 , n64879 , n64883 , n64884 , n64888 );
and ( n64890 , n64866 , n64889 );
and ( n64891 , n18737 , n17451 );
or ( n64892 , n64890 , n64891 );
and ( n64893 , n64892 , n23924 );
and ( n64894 , n17975 , n23926 );
or ( n64895 , n64893 , n64894 );
buf ( n64896 , n64895 );
buf ( n64897 , n64896 );
buf ( n64898 , n10615 );
and ( C0 , n10618 , n10617 );
or ( C1 , n10618 , n10617 );
endmodule

