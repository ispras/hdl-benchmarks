//NOTE: no-implementation module stub

module SREG16MC (
    input wire DSPCLK,
    input wire MMR_web,
    input wire SCTL_we_PSET,
    input wire [15:0] DMD_SCTL,
    output reg [15:0] SCTL,
    input wire RST
);

endmodule
