// IWLS benchmark module "sbc" printed on Wed May 29 21:45:28 2002
module sbc(ACKl, BUS_Inactive, GRANTi, LastRQSTi, SBCResetPCC, PCCReq, PCCReqCode0, PCCReqCode1, PCCReqCode2, PCCReqCode3, PCCConfirm, RQSTi, SingleStep, STARTi, TM0i, TM1i, VACKl, VTM0i, VSACKi, ACKi, RESETi, SlotSpace_Id_Match, PCCSawReset, CoherencyState1i, CoherencyState2i, NuBusActive, PCCAck, PCCsync, STARTo, Tag_Match, TM1l, VTM0l, VTM1l, PCCAckCode, VACKi, physrecXXXXstate0, physrecXXXXstate1, wdcntXXXXstate1, wdcntXXXXstate2, wdcntXXXXstate3, physrecXXXXNextState0, physrecXXXXNextState1, wdcntXXXXNextState1, wdcntXXXXNextState2, wdcntXXXXNextState3, masterXXXXArb_active, masterXXXXEn_ABufo, masterXXXXEn_PDBufi, masterXXXXL_PDBufi, masterXXXXEn_VDBufi, masterXXXXEn_PDBufo, masterXXXXL_DBufo_if_TM0, masterXXXXRQSTo, masterXXXXSBC_WriteCache, nubusXXXXNuBusActive, nubusXXXXL_PABufi, resetXXXXSBCResetPCC, resetXXXXReset, slaveXXXXL_VABufi, slaveXXXXSBCReq, slaveXXXXSBCReqCode0, slaveXXXXSBCReqCode1, slaveXXXXSBCReqCode2, slaveXXXXSnoopAddrFromProc, slaveXXXXSnoopVTag_W, slaveXXXXSnoopState_W, slaveXXXXGenerateNextState, slaveXXXXSnoopVTagState_R, virmachXXXXEn_VDBufo, virmachXXXXSBCsetDirty, virmachXXXXSBCCacheRelease, virmachXXXXSBCConfigure, wdcntXXXXwd_cnt0, wdcntXXXXwd_cnt1, wdcntXXXXwd_cnt2, encodemuxXXXXMX_AD_8, nextstateXXXXCoherencyState2o, orXXXXACKo, orXXXXEn_CNTL, orXXXXRESETo, orXXXXTM0o, orXXXXTM1o, orXXXXEn_START, orXXXXSBCAck, orXXXXSBCAckCodelatch, orXXXXSBCAckCode0, orXXXXSBCAckCode1, orXXXXSBCAckCode2, orXXXXSBCAckCode3, orXXXXSTARTo, orXXXXEn_VCNTL, orXXXXVSACKo, orXXXXVACKo, orXXXXVTM0o, orXXXXVTM1o, orXXXXL_DBufo);
input
  PCCsync,
  wdcntXXXXstate1,
  wdcntXXXXstate2,
  wdcntXXXXstate3,
  SlotSpace_Id_Match,
  CoherencyState1i,
  CoherencyState2i,
  NuBusActive,
  Tag_Match,
  physrecXXXXstate0,
  physrecXXXXstate1,
  PCCReqCode0,
  PCCReqCode1,
  PCCReqCode2,
  PCCReqCode3,
  RESETi,
  PCCAckCode,
  PCCAck,
  GRANTi,
  STARTi,
  STARTo,
  RQSTi,
  ACKi,
  ACKl,
  TM0i,
  PCCReq,
  TM1i,
  TM1l,
  SingleStep,
  BUS_Inactive,
  SBCResetPCC,
  VACKi,
  VACKl,
  PCCConfirm,
  VTM0i,
  VTM0l,
  VTM1l,
  VSACKi,
  PCCSawReset,
  LastRQSTi;
output
  orXXXXVSACKo,
  orXXXXL_DBufo,
  orXXXXACKo,
  orXXXXEn_VCNTL,
  orXXXXEn_CNTL,
  virmachXXXXSBCConfigure,
  masterXXXXRQSTo,
  orXXXXRESETo,
  orXXXXSBCAckCodelatch,
  masterXXXXEn_ABufo,
  slaveXXXXSnoopAddrFromProc,
  virmachXXXXSBCCacheRelease,
  physrecXXXXNextState0,
  physrecXXXXNextState1,
  orXXXXSTARTo,
  slaveXXXXSnoopVTagState_R,
  encodemuxXXXXMX_AD_8,
  masterXXXXL_PDBufi,
  resetXXXXReset,
  slaveXXXXGenerateNextState,
  resetXXXXSBCResetPCC,
  masterXXXXL_DBufo_if_TM0,
  slaveXXXXSBCReqCode0,
  slaveXXXXSBCReqCode1,
  slaveXXXXSBCReqCode2,
  orXXXXTM1o,
  orXXXXTM0o,
  masterXXXXArb_active,
  masterXXXXEn_PDBufi,
  nubusXXXXL_PABufi,
  masterXXXXEn_PDBufo,
  orXXXXVTM1o,
  orXXXXVTM0o,
  virmachXXXXEn_VDBufo,
  slaveXXXXL_VABufi,
  masterXXXXEn_VDBufi,
  slaveXXXXSBCReq,
  orXXXXSBCAckCode0,
  orXXXXSBCAckCode1,
  orXXXXSBCAckCode2,
  orXXXXSBCAckCode3,
  wdcntXXXXwd_cnt0,
  wdcntXXXXwd_cnt1,
  wdcntXXXXwd_cnt2,
  nubusXXXXNuBusActive,
  orXXXXEn_START,
  orXXXXSBCAck,
  slaveXXXXSnoopState_W,
  slaveXXXXSnoopVTag_W,
  nextstateXXXXCoherencyState2o,
  orXXXXVACKo,
  masterXXXXSBC_WriteCache,
  wdcntXXXXNextState1,
  wdcntXXXXNextState2,
  wdcntXXXXNextState3,
  virmachXXXXSBCsetDirty;
reg
  masterXXXXstate0,
  masterXXXXstate1,
  masterXXXXstate2,
  masterXXXXstate3,
  V_transmit_begin,
  wdcntXXXXstate0,
  P_receive_begin,
  UpdateDone,
  UpdateReq,
  virmachXXXXstate0,
  virmachXXXXstate1,
  resetXXXXstate0,
  resetXXXXstate1,
  resetXXXXstate2,
  wd_cnt_test,
  Reset_wd_cnt,
  Set_ex_wd_cnt1,
  Intr_req,
  Intr_done,
  Gen_Reset,
  Incr_wd_cnt,
  slaveXXXXstate0,
  slaveXXXXstate1,
  slaveXXXXstate2,
  nubusXXXXstate0,
  nubusXXXXstate1,
  P_receive_cancel;
wire
  \[145] ,
  \[15247] ,
  \[146] ,
  \[147] ,
  \[10061] ,
  \[14676]* ,
  \[14883] ,
  \[14862]* ,
  masterXXXXACKo,
  \[150] ,
  \[151] ,
  \[14529] ,
  \[152] ,
  \[14911] ,
  \[154] ,
  \[155] ,
  \[14627] ,
  \[156] ,
  \[14627]* ,
  \{nubusXXXXNuBusActive} ,
  \[157] ,
  \[14816] ,
  \[158] ,
  \[159] ,
  \[14531] ,
  \[15452] ,
  \{physrecXXXXNextState1} ,
  \{resetXXXXSBCResetPCC} ,
  \[15030]* ,
  \[10750]_inv ,
  \{orXXXXReset_wd_cnt_x} ,
  \[160] ,
  \[15169] ,
  \[161] ,
  \[162] ,
  \{orXXXXSBCAckCode1} ,
  \{orXXXXSBCAckCode2} ,
  \{virmachXXXXNextState1} ,
  \{slaveXXXXL_VABufi} ,
  \{orXXXXSBCAckCode3} ,
  \[165] ,
  \[14535] ,
  \[166] ,
  \[14928] ,
  \[10653] ,
  \[14984]* ,
  \[84] ,
  \{virmachXXXXNextState0} ,
  \[169] ,
  \[85] ,
  \{orXXXXSBCAckCode0} ,
  \{orXXXXTM1o} ,
  \[86] ,
  \[87] ,
  \[15074] ,
  \[14797]* ,
  \[88] ,
  \[14443] ,
  \[89] ,
  \{masterXXXXSBC_WriteCache} ,
  \{masterXXXXUpdateReq} ,
  \{orXXXXACKo} ,
  \[173] ,
  \[90] ,
  \[91] ,
  \[176] ,
  \[92] ,
  \[177] ,
  \[93] ,
  \{orXXXXEn_CNTL} ,
  \[178] ,
  \[10703]_inv* ,
  \[94] ,
  \[179] ,
  \[95] ,
  \[96] ,
  \{orXXXXVTM0o} ,
  \[97] ,
  \[98] ,
  \[100] ,
  \[99] ,
  \[101] ,
  \[2536] ,
  \{orXXXXIncr_wd_cnt} ,
  \{slaveXXXXNextState1} ,
  \[102] ,
  \{slaveXXXXNextState2} ,
  \[103] ,
  \{orXXXXEn_VCNTL} ,
  \[104] ,
  \{slaveXXXXNextState0} ,
  \[105] ,
  \[106] ,
  \[107] ,
  \[108] ,
  \[202] ,
  \[15017] ,
  \[109] ,
  \[15190] ,
  \[203] ,
  \[1048] ,
  \[15192] ,
  \{orXXXXVSACKo} ,
  \[14654] ,
  \[14467] ,
  \[206] ,
  \[207] ,
  \[14469] ,
  \[208] ,
  \[14852] ,
  \{orXXXXEn_START} ,
  \[209] ,
  \[111] ,
  \[15198] ,
  \{slaveXXXXSBCReq} ,
  \{masterXXXXNextState1} ,
  \[14902]* ,
  \[112] ,
  \[14567] ,
  \{masterXXXXNextState2} ,
  \[15021] ,
  \[14661] ,
  \[113] ,
  \{masterXXXXNextState3} ,
  \[10748]_inv ,
  \[114] ,
  \[191] ,
  \[2836] ,
  \{wdcntXXXXwd_cnt_test} ,
  \[116] ,
  \[193] ,
  \[210] ,
  \{nubusXXXXL_PABufi} ,
  \{resetXXXXNextState1} ,
  \[15676] ,
  \[117] ,
  \[15219] ,
  \[211] ,
  \{orXXXXRESETo} ,
  \{slaveXXXXSBCReqCode0} ,
  \{resetXXXXNextState2} ,
  \[212] ,
  \{masterXXXXNextState0} ,
  \{virmachXXXXSBCConfigure} ,
  \[119] ,
  \[213] ,
  \[214] ,
  \[10889]_inv ,
  \{slaveXXXXSBCReqCode1} ,
  \[15030] ,
  \[120] ,
  \[121] ,
  masterXXXXVSACKo,
  \[122] ,
  \[14764] ,
  \[123] ,
  \[124] ,
  \[15228] ,
  \{orXXXXSBCAck} ,
  \[125] ,
  \[126] ,
  \[128] ,
  \[129] ,
  \[15223] ,
  \{nubusXXXXNextState0} ,
  \[14676] ,
  \{orXXXXL_DBufo} ,
  \[10507]_inv ,
  \{nubusXXXXNextState1} ,
  \[130] ,
  \[10749]_inv ,
  \[131] ,
  \[15041] ,
  \[14681] ,
  \[133] ,
  \[134] ,
  \[135] ,
  \[136] ,
  \{slaveXXXXSnoopState_W} ,
  \[137] ,
  \[138] ,
  \[14417] ,
  \[139] ,
  \[14857]* ,
  \{orXXXXVACKo} ,
  \[15334] ,
  \{orXXXXSBCAckCodelatch} ,
  \[140] ,
  \[14976] ,
  \[141] ,
  \[14902] ,
  \[142] ,
  \[143] ,
  \[144] ;
assign
  orXXXXVSACKo = \{orXXXXVSACKo} ,
  \[145]  = masterXXXXstate2 & ~STARTi,
  \[15247]  = ~\[10889]_inv  & (~masterXXXXstate3 & (masterXXXXstate2 & ~ACKl)),
  \[146]  = ~\[128]  & GRANTi,
  \[147]  = VSACKi | ~VTM0i,
  \[10061]  = (~\[193]  & \[169] ) | ((~\[193]  & ~CoherencyState2i) | (\[144]  & ~slaveXXXXstate1)),
  \[14676]*  = ~\[14676] ,
  \[14883]  = (\[209]  & (~nubusXXXXstate0 & SlotSpace_Id_Match)) | (\[207]  & ~Intr_done),
  orXXXXL_DBufo = \{orXXXXL_DBufo} ,
  orXXXXACKo = \{orXXXXACKo} ,
  \[14862]*  = \[15041]  | \[15219] ,
  orXXXXEn_VCNTL = \{orXXXXEn_VCNTL} ,
  masterXXXXACKo = 0,
  \[150]  = (~\[114]  & VSACKi) | (masterXXXXstate1 & ~ACKl),
  \[151]  = \[10507]_inv  | PCCReqCode2,
  \[14529]  = (\[134]  & (~masterXXXXstate0 & ~SBCResetPCC)) | ((\[15223]  & (STARTi & ~SBCResetPCC)) | \[161] ),
  \[152]  = ~VTM0l | STARTo,
  \[14911]  = (\[140]  & (~P_receive_cancel & (~physrecXXXXstate0 & ~TM1i))) | ((\[140]  & (~P_receive_cancel & (~physrecXXXXstate0 & ~TM0i))) | (\[140]  & (~wd_cnt_test & ~physrecXXXXstate0))),
  \[154]  = ~nubusXXXXstate1 | STARTi,
  \[155]  = (\[141]  & \[10749]_inv ) | (~\[138]  & ~PCCConfirm),
  \[14627]  = (\[137]  & \[121] ) | (\[137]  & ~\[14911] ),
  orXXXXEn_CNTL = \{orXXXXEn_CNTL} ,
  \[156]  = ~\[10889]_inv  & ACKl,
  \[14627]*  = ~\[14627] ,
  \{nubusXXXXNuBusActive}  = (\[112]  & (\[2536]  & ~Intr_done)) | ((\[158]  & ~\[2536] ) | \[209] ),
  \[157]  = ~masterXXXXstate1 & ~SBCResetPCC,
  \[14816]  = (\[156]  & (\[145]  & ~masterXXXXstate3)) | (\[135]  & (masterXXXXstate1 & ACKl)),
  \[158]  = \[124]  & nubusXXXXstate0,
  virmachXXXXSBCConfigure = \{virmachXXXXSBCConfigure} ,
  \[159]  = ~\[143]  & (~\[131]  & (\[113]  & (~masterXXXXstate0 & (~RQSTi & ~SBCResetPCC)))),
  \[14531]  = (~\[141]  & (~\[128]  & ~SBCResetPCC)) | ((\[179]  & \[134] ) | (~\[10889]_inv  & \[15223] )),
  \[15452]  = \[208]  & ~virmachXXXXstate1,
  \{physrecXXXXNextState1}  = (\[117]  & (P_receive_begin & physrecXXXXstate0)) | ((\[210]  & wd_cnt_test) | ((\[160]  & ~P_receive_cancel) | (\[160]  & physrecXXXXstate0))),
  masterXXXXRQSTo = \[14531] ,
  orXXXXRESETo = \{orXXXXRESETo} ,
  \{resetXXXXSBCResetPCC}  = (resetXXXXstate1 & ~PCCSawReset) | (resetXXXXstate2 | (resetXXXXstate0 | RESETi)),
  orXXXXSBCAckCodelatch = \{orXXXXSBCAckCodelatch} ,
  \[15030]*  = ~\[15030] ,
  \[10750]_inv  = \[193]  | (\[125]  | (~slaveXXXXstate2 | ~Tag_Match)),
  \{orXXXXReset_wd_cnt_x}  = (\[10507]_inv  & \[14443] ) | ((\[10507]_inv  & PCCReqCode1) | ((\[14764]  & ~slaveXXXXstate0) | (~\[151]  | \[15017] ))),
  \[160]  = \[117]  & ~ACKi,
  \[15169]  = \[15452]  & wd_cnt_test,
  \[161]  = \[146]  & ~SBCResetPCC,
  \[162]  = \[112]  & ~slaveXXXXstate0,
  masterXXXXEn_ABufo = \[14535] ,
  \{orXXXXSBCAckCode1}  = (\[123]  & (ACKi & ~TM0i)) | ((\[140]  & ~wd_cnt_test) | ((\[140]  & physrecXXXXstate0) | ((\[14816]  & ~TM0i) | ((\[14911]  & TM1i) | (\[14911]  & TM0i))))),
  \{orXXXXSBCAckCode2}  = (\[123]  & (~\[14928]  & (~TM1i & TM0i))) | ((ACKi & (TM1i & (~TM0i & ~SBCResetPCC))) | ((~\[141]  & (\[14469]  & PCCReqCode2)) | ((\[141]  & (\[14469]  & PCCConfirm)) | ((\[14816]  & (~TM1i & TM0i)) | ((~\[15676]  & (resetXXXXstate2 & ~resetXXXXstate1)) | ((\[140]  & ~wd_cnt_test) | ((\[140]  & physrecXXXXstate0) | ((\[1048]  & \[14469] ) | ((\[14911]  & ~TM0i) | (\{orXXXXSBCAckCode1}  & TM1i)))))))))),
  \{virmachXXXXNextState1}  = (P_receive_cancel & (~virmachXXXXstate1 & (~virmachXXXXstate0 & ~SBCResetPCC))) | ((\[208]  & (virmachXXXXstate1 & ~VACKi)) | (\[15192]  & ~PCCAck)),
  \{slaveXXXXL_VABufi}  = (\[213]  & (\[136]  & (~Intr_req & (slaveXXXXstate0 & ~VSACKi)))) | ((\[136]  & (~Intr_req & (ACKi & (~VSACKi & STARTi)))) | ((\[129]  & (~slaveXXXXstate0 & (ACKi & STARTi))) | ((\[120]  & (~slaveXXXXstate2 & (~slaveXXXXstate0 & ACKi))) | ((\[213]  & (\[129]  & ~slaveXXXXstate0)) | ((\[136]  & (~slaveXXXXstate0 & ACKi)) | RESETi))))),
  \{orXXXXSBCAckCode3}  = (resetXXXXstate2 & ~RESETi) | ~\[14627] ,
  \[165]  = ~Incr_wd_cnt | ~wdcntXXXXstate3,
  \[14535]  = ~\[130]  & (~\[10749]_inv  & ~SBCResetPCC),
  \[166]  = PCCReqCode2 | PCCReqCode0,
  \[14928]  = (\[210]  & wd_cnt_test) | (\[123]  & ~ACKi),
  \[10653]  = (\[145]  & (masterXXXXstate0 & (~LastRQSTi & ACKl))) | ((masterXXXXstate1 & (masterXXXXstate0 & (~LastRQSTi & ACKl))) | (~\[130]  & masterXXXXstate2)),
  \[14984]*  = (\[142]  & (~Incr_wd_cnt & wdcntXXXXstate3)) | ((\[142]  & (wdcntXXXXstate0 & wdcntXXXXstate3)) | (\[14797]*  & (wdcntXXXXstate3 & wdcntXXXXstate2))),
  \[84]  = \{masterXXXXNextState0} ,
  \{virmachXXXXNextState0}  = (~\[15192]  & \{virmachXXXXNextState1} ) | ((\[15192]  & ~\{virmachXXXXNextState1} ) | \[214] ),
  \[169]  = ~TM1l | ~CoherencyState1i,
  \[85]  = \{masterXXXXNextState1} ,
  \{orXXXXSBCAckCode0}  = \[14469]  | \[14911] ,
  \{orXXXXTM1o}  = (\[151]  & ~PCCReqCode1) | (~\[191]  | (~\[14862]*  | PCCReqCode0)),
  \[86]  = \{masterXXXXNextState2} ,
  slaveXXXXSnoopAddrFromProc = \[14681] ,
  virmachXXXXSBCCacheRelease = \[15169] ,
  \[87]  = \{masterXXXXNextState3} ,
  physrecXXXXNextState0 = \[14928] ,
  physrecXXXXNextState1 = \{physrecXXXXNextState1} ,
  \[15074]  = (masterXXXXstate3 & (~masterXXXXstate1 & ~SingleStep)) | (\[143]  & ~masterXXXXstate1),
  \[14797]*  = (~\[165]  & (\[142]  & ~wdcntXXXXstate2)) | ((\[165]  & (\[142]  & wdcntXXXXstate2)) | (\[142]  & (wdcntXXXXstate2 & wdcntXXXXstate1))),
  \[88]  = \{nubusXXXXNextState0} ,
  orXXXXSTARTo = \[14567] ,
  \[14443]  = \[151]  & PCCReqCode0,
  \[89]  = \{nubusXXXXNextState1} ,
  \{masterXXXXSBC_WriteCache}  = (masterXXXXstate2 & (VSACKi & ~ACKl)) | ((\[145]  & ~ACKl) | (\[135]  | \[14902] )),
  \{masterXXXXUpdateReq}  = (\[157]  & (~UpdateDone & ~masterXXXXstate0)) | (masterXXXXVSACKo | ~PCCReqCode1),
  \{orXXXXACKo}  = 1,
  \[173]  = masterXXXXstate2 | RQSTi,
  \[90]  = \{slaveXXXXNextState0} ,
  \[91]  = \{slaveXXXXNextState1} ,
  \[176]  = ~VTM1l & ~TM1l,
  \[92]  = \{slaveXXXXNextState2} ,
  \[177]  = \[135]  & ~ACKl,
  \[93]  = \[14976] ,
  \{orXXXXEn_CNTL}  = (\[133]  & (\[124]  & ~SlotSpace_Id_Match)) | ((\[158]  & \[133] ) | (~\[14661]  & ~SBCResetPCC)),
  \[178]  = \[139]  & \[129] ,
  \[10703]_inv*  = (\[177]  & (\[147]  & ~\[131] )) | ((\[177]  & \[126] ) | (\[177]  & masterXXXXstate1)),
  \[94]  = \{resetXXXXNextState1} ,
  \[179]  = \[10889]_inv  & ~SBCResetPCC,
  \[95]  = \{resetXXXXNextState2} ,
  slaveXXXXSnoopVTagState_R = \[14764] ,
  \[96]  = \{virmachXXXXNextState0} ,
  \{orXXXXVTM0o}  = (\[15452]  & ~wd_cnt_test) | ((\[15452]  & ~PCCAckCode) | (masterXXXXVSACKo | \[14852] )),
  \[97]  = \{virmachXXXXNextState1} ,
  \[98]  = \[15030]* ,
  \[100]  = \[14883] ,
  \[99]  = \[14627]* ,
  \[101]  = \[15190] ,
  \[2536]  = (\[211]  & STARTi) | (~\[154]  & nubusXXXXstate0),
  \{orXXXXIncr_wd_cnt}  = (~V_transmit_begin & (VTM0i & ~SBCResetPCC)) | ((\[210]  & ~\[14928] ) | ((\[15247]  & TM0i) | ((\[15247]  & STARTi) | \[214] ))),
  \{slaveXXXXNextState1}  = (\[120]  & (slaveXXXXstate2 & (PCCsync & (~RESETi & ACKi)))) | ((~\[125]  & (\[120]  & (~\[14764]  & PCCsync))) | ((~slaveXXXXstate2 & (TM1l & (~RESETi & ACKi))) | ((~slaveXXXXstate2 & (~RESETi & (ACKi & ~STARTi))) | ((~\[125]  & (\[10061]  & ~\[14764] )) | ((\[14764]  & (slaveXXXXstate0 & TM1l)) | ((\[14764]  & ~STARTi) | slaveXXXXstate1)))))),
  \[102]  = \{masterXXXXUpdateReq} ,
  \{slaveXXXXNextState2}  = (\[144]  & (~\[125]  & (slaveXXXXstate2 & ~slaveXXXXstate1))) | ((\[136]  & (\[112]  & (~Intr_req & NuBusActive))) | ((\[162]  & (~\[120]  & slaveXXXXstate2)) | ((\[162]  & (slaveXXXXstate2 & PCCsync)) | ((\[136]  & (~\[125]  & VSACKi)) | ((~\[206]  & ~RESETi) | ((\[178]  & ~\[14764] ) | ((\[162]  & \[136] ) | ((\[139]  & \[136] ) | (\[14764]  & ~PCCsync))))))))),
  \[103]  = \[14681] ,
  \{orXXXXEn_VCNTL}  = (~\[131]  & (~\[10749]_inv  & (~RQSTi & ~SBCResetPCC))) | ((\[212]  & (VSACKi & STARTi)) | ((~\[138]  & (PCCConfirm & ~SBCResetPCC)) | ((\[177]  & masterXXXXstate2) | (\[15192]  | (\[15452]  | \[14852] ))))),
  \[104]  = \{orXXXXReset_wd_cnt_x} ,
  \{slaveXXXXNextState0}  = (~\[125]  & (slaveXXXXstate1 & VSACKi)) | ((\[178]  & VTM0l) | ((~\[125]  & \[10061] ) | (~\[125]  & ~slaveXXXXstate2))),
  encodemuxXXXXMX_AD_8 = \[15198] ,
  masterXXXXL_PDBufi = \[10703]_inv* ,
  \[105]  = \[14467] ,
  resetXXXXReset = \[15676] ,
  \[106]  = \{orXXXXIncr_wd_cnt} ,
  \[107]  = \{wdcntXXXXwd_cnt_test} ,
  \[108]  = \[14443] ,
  \[202]  = 0,
  \[15017]  = \[145]  & (\[135]  & (VSACKi & VTM0i)),
  \[109]  = \[15017] ,
  \[15190]  = (\[206]  & slaveXXXXstate0) | (\[206]  & RESETi),
  \[203]  = ~Gen_Reset | (resetXXXXstate1 | resetXXXXstate0),
  \[1048]  = (~\[131]  & (\[113]  & (~masterXXXXstate0 & (SingleStep & PCCReq)))) | ((~\[131]  & (\[113]  & (~masterXXXXstate0 & (RQSTi & PCCReq)))) | (~\[10748]_inv  & PCCReqCode1)),
  \[15192]  = (V_transmit_begin & (~P_receive_cancel & (~virmachXXXXstate0 & ~SBCResetPCC))) | (virmachXXXXstate1 & (~virmachXXXXstate0 & ~SBCResetPCC)),
  slaveXXXXGenerateNextState = \[14676]* ,
  \{orXXXXVSACKo}  = (\[176]  & (\[10061]  & (\[15190]  & (VTM0l & (Tag_Match & ~RESETi))))) | ((~\[144]  & (\[10061]  & (\[15190]  & (~CoherencyState2i & ~RESETi)))) | ((\[15190]  & (~slaveXXXXstate2 & ~RESETi)) | (\[214]  | (\[15192]  | (masterXXXXVSACKo | (\[15334]  | \[14764] )))))),
  \[14654]  = (\[136]  & (\[124]  & (Intr_req & (slaveXXXXstate0 & (~PCCsync & (NuBusActive & ~VSACKi)))))) | (\[162]  & (slaveXXXXstate2 & ~slaveXXXXstate1)),
  \[14467]  = (\[10507]_inv  & (PCCReqCode2 & PCCReqCode0)) | ((~\[166]  & \[10507]_inv ) | ((~\[166]  & PCCReqCode1) | (~\[113]  & PCCReqCode0))),
  \[206]  = slaveXXXXstate2 | (~slaveXXXXstate1 | ~PCCAck),
  \[207]  = \[158]  & ~nubusXXXXstate1,
  \[14469]  = (~\[137]  & (masterXXXXstate3 & PCCReqCode2)) | ((\[155]  & ~SBCResetPCC) | ((~\[137]  & PCCReqCode0) | (\[1048]  & ~SBCResetPCC))),
  \[208]  = virmachXXXXstate0 & ~SBCResetPCC,
  \[14852]  = ~\[10750]_inv  & (~TM1l & CoherencyState2i),
  \{orXXXXEn_START}  = (\[117]  & (~\[14911]  & ~LastRQSTi)) | ((~\{physrecXXXXNextState1}  & (~ACKi & ~SBCResetPCC)) | ((physrecXXXXstate0 & (~SBCResetPCC & ~LastRQSTi)) | ((~\[14661]  & ~SBCResetPCC) | ((\{physrecXXXXNextState1}  & P_receive_begin) | ((\{physrecXXXXNextState1}  & ~physrecXXXXstate0) | \[15247] ))))),
  \[209]  = ~\[133]  & \[124] ,
  resetXXXXSBCResetPCC = \{resetXXXXSBCResetPCC} ,
  \[111]  = \[14852] ,
  \[15198]  = \[116]  & (~PCCReqCode3 & ~PCCReqCode2),
  \{slaveXXXXSBCReq}  = ~\[14676]  | \[14654] ,
  \{masterXXXXNextState1}  = (~\[143]  & (~\[121]  & (~\[15074]  & ~SBCResetPCC))) | ((~\[143]  & (~\[121]  & (~masterXXXXstate2 & ~SBCResetPCC))) | ((~\[143]  & (~\[15074]  & (RQSTi & ~SBCResetPCC))) | ((~\[143]  & (~masterXXXXstate2 & (RQSTi & ~SBCResetPCC))) | ((~\[114]  & (VSACKi & (~SBCResetPCC & GRANTi))) | ((\[161]  & \[10749]_inv ) | ((\[161]  & ~PCCConfirm) | ((\[161]  & ~BUS_Inactive) | ~\[14902] ))))))),
  \[14902]*  = ~\[14902] ,
  \[112]  = ~RESETi & ~ACKi,
  \[14567]  = (\[159]  & ~SingleStep) | (\[141]  & ~SBCResetPCC),
  \{masterXXXXNextState2}  = (\[159]  & (\[15074]  & \[15198] )) | ((\[159]  & (\[15074]  & ~PCCReqCode0)) | ((masterXXXXstate3 & (masterXXXXstate1 & ~SBCResetPCC)) | ((\[157]  & ~UpdateDone) | (~\[147]  | (~\[10889]_inv  | masterXXXXstate2))))),
  \[15021]  = \[146]  & (~VSACKi & BUS_Inactive),
  \[14661]  = (~\[121]  & (~\[10653]  & (~\[10748]_inv  & BUS_Inactive))) | ((\[131]  & (~\[10653]  & BUS_Inactive)) | (\[146]  & ~\[10653] )),
  \[113]  = ~PCCReqCode2 | ~PCCReqCode1,
  \{masterXXXXNextState3}  = (\[179]  & (\[157]  & (\[121]  & (~\[119]  & (PCCReqCode3 & PCCReq))))) | ((\[179]  & (\[157]  & (~\[15074]  & (masterXXXXstate3 & ~RQSTi)))) | ((\[179]  & (\[157]  & (masterXXXXstate3 & (~RQSTi & ~PCCReq)))) | ((\[157]  & (~\[119]  & (~RQSTi & (PCCReqCode2 & PCCReqCode0)))) | ((\[157]  & (~\[119]  & (~RQSTi & (PCCReqCode1 & ~PCCReqCode0)))) | ((~\[157]  & (\[119]  & (masterXXXXstate3 & ~SBCResetPCC))) | ((\[157]  & (\[156]  & (VSACKi & ~LastRQSTi))) | ((\[156]  & (\[10653]  & (VSACKi & ~VACKl))) | ((\[156]  & (masterXXXXstate2 & (~VSACKi & ~LastRQSTi))) | ((\[141]  & (\[14529]  & (~PCCReqCode2 & ~PCCReqCode1))) | ((\[141]  & (\[14529]  & (PCCReqCode2 & PCCReqCode0))) | ((\[141]  & (\[14529]  & (PCCReqCode1 & ~PCCReqCode0))) | ((~\[119]  & (~\[10889]_inv  & (~\[14816]  & ~\[15041] ))) | ((\[179]  & (\[10653]  & ~RQSTi)) | ((\[159]  & (~PCCReqCode2 & ~PCCReqCode1)) | ((\[141]  & (\[14529]  & ~PCCConfirm)) | ((\[141]  & (\[14529]  & PCCReqCode3)) | ((\[141]  & (\[14529]  & ~PCCReq)) | ((~\[119]  & (~\[10889]_inv  & ~VTM0i)) | ((~\[119]  & (\[14816]  & VSACKi)) | ((\[119]  & (\[14529]  & ~masterXXXXstate2)) | ((\[177]  & \[126] ) | ((\[10653]  & \[14816] ) | (\[15041]  & ~RQSTi))))))))))))))))))))))),
  \[10748]_inv  = masterXXXXstate2 | (masterXXXXstate1 | (masterXXXXstate0 | (~PCCReqCode3 | ~PCCReq))),
  \[114]  = masterXXXXstate3 | ~masterXXXXstate1,
  masterXXXXL_DBufo_if_TM0 = \[15247] ,
  \[191]  = ~\[10507]_inv  | \[14467] ,
  \[2836]  = (\[157]  & (UpdateDone & (masterXXXXstate2 & ~masterXXXXstate0))) | ((resetXXXXstate2 & ~RESETi) | \[14816] ),
  slaveXXXXSBCReqCode0 = \{slaveXXXXSBCReqCode0} ,
  slaveXXXXSBCReqCode1 = \{slaveXXXXSBCReqCode1} ,
  \{wdcntXXXXwd_cnt_test}  = (\[14857]*  & (\[14797]*  & (~Incr_wd_cnt & wdcntXXXXstate3))) | ((\[14857]*  & (\[14797]*  & (Incr_wd_cnt & wdcntXXXXstate2))) | ~\[15030] ),
  slaveXXXXSBCReqCode2 = \[14654] ,
  \[116]  = PCCReqCode1 | ~PCCReqCode0,
  \[193]  = slaveXXXXstate1 | ~VTM0l,
  \[210]  = \[160]  & TM0i,
  orXXXXTM1o = \{orXXXXTM1o} ,
  \{nubusXXXXL_PABufi}  = (\[213]  & \[211] ) | ((\[2536]  & ACKi) | (~Intr_done | ~RESETi)),
  \{resetXXXXNextState1}  = (\{resetXXXXSBCResetPCC}  & (~PCCSawReset & ~RESETi)) | \[15676] ,
  \[15676]  = RESETi & resetXXXXstate2,
  \[117]  = physrecXXXXstate1 & ~SBCResetPCC,
  \[15219]  = \[207]  & Intr_done,
  \[211]  = ~nubusXXXXstate1 & ~nubusXXXXstate0,
  orXXXXTM0o = \[14862]* ,
  \{orXXXXRESETo}  = (\[211]  & (~\[122]  & (ACKi & ~STARTi))) | ((~\[122]  & (nubusXXXXstate1 & (nubusXXXXstate0 & STARTi))) | ((\[139]  & (~nubusXXXXstate1 & nubusXXXXstate0)) | ~\[14627] )),
  \{slaveXXXXSBCReqCode0}  = (\[14852]  & ~\{slaveXXXXSBCReqCode1} ) | (\{slaveXXXXSBCReqCode1}  & TM1l),
  \{resetXXXXNextState2}  = (\[203]  & RESETi) | \[15676] ,
  masterXXXXArb_active = \[14529] ,
  \[212]  = ~\[131]  & ~\[10889]_inv ,
  \{masterXXXXNextState0}  = (\[138]  & (~\[15223]  & (SBCResetPCC & GRANTi))) | ((\[138]  & (STARTi & (SBCResetPCC & GRANTi))) | ((\[15021]  & (~\[15223]  & (~PCCConfirm & SBCResetPCC))) | ((\[15021]  & (STARTi & (~PCCConfirm & SBCResetPCC))) | ((~\[147]  & (\[135]  & masterXXXXstate2)) | ((\[145]  & (\[135]  & VSACKi)) | ((\[128]  & (~\[15223]  & SBCResetPCC)) | ((\[128]  & (STARTi & SBCResetPCC)) | ((\[114]  & (~\[10889]_inv  & VACKl)) | ((\[212]  & ~\[15041] ) | ((\[159]  & ~SingleStep) | ((\[150]  & ~\[10889]_inv ) | ((~\[15041]  & \[10703]_inv* ) | \[15247] )))))))))))),
  \{virmachXXXXSBCConfigure}  = (~\[15192]  & ~PCCAck) | \[15452] ,
  masterXXXXEn_PDBufi = \[10703]_inv* ,
  nubusXXXXL_PABufi = \{nubusXXXXL_PABufi} ,
  masterXXXXEn_PDBufo = \[15247] ,
  \[119]  = ~masterXXXXstate3 | masterXXXXstate2,
  \[213]  = ~ACKi & ~STARTi,
  \[214]  = ~\[15169]  & \[15452] ,
  \[10889]_inv  = ~masterXXXXstate0 | SBCResetPCC,
  orXXXXVTM1o = \[14417] ,
  orXXXXVTM0o = \{orXXXXVTM0o} ,
  virmachXXXXEn_VDBufo = \[15452] ,
  slaveXXXXL_VABufi = \{slaveXXXXL_VABufi} ,
  \{slaveXXXXSBCReqCode1}  = (\[176]  & (~\[10750]_inv  & ~CoherencyState1i)) | ((~\[169]  & (~\[10750]_inv  & ~CoherencyState2i)) | (\[14852]  & ~VTM1l)),
  \[15030]  = (~Set_ex_wd_cnt1 & ~SBCResetPCC) | ((~wdcntXXXXstate0 & SBCResetPCC) | ((wdcntXXXXstate3 & SBCResetPCC) | ((wdcntXXXXstate2 & SBCResetPCC) | ((wdcntXXXXstate1 & ~SBCResetPCC) | ~Reset_wd_cnt)))),
  masterXXXXEn_VDBufi = \[14902]* ,
  \[120]  = Intr_req | SlotSpace_Id_Match,
  \[121]  = \[116]  | PCCReqCode2,
  masterXXXXVSACKo = ~\[14443]  | PCCReqCode2,
  \[122]  = Intr_done | RESETi,
  \[14764]  = (\[178]  & ~\[152] ) | (\[129]  & ~\[125] ),
  \[123]  = (\[117]  & P_receive_cancel) | (physrecXXXXstate0 & ~SBCResetPCC),
  slaveXXXXSBCReq = \{slaveXXXXSBCReq} ,
  \[124]  = \[112]  & ~STARTi,
  \[15228]  = \[208]  & (virmachXXXXstate1 & (VACKi & VTM0i)),
  \{orXXXXSBCAck}  = 1,
  \[125]  = ~slaveXXXXstate0 | RESETi,
  \[126]  = (\[145]  & ~VSACKi) | (VSACKi & STARTi),
  \[128]  = \[114]  | ~masterXXXXstate2,
  \[129]  = ~slaveXXXXstate2 & ~slaveXXXXstate1,
  \[15223]  = ~masterXXXXstate3 & (~masterXXXXstate2 & (~masterXXXXstate1 & masterXXXXstate0)),
  orXXXXSBCAckCode0 = \{orXXXXSBCAckCode0} ,
  orXXXXSBCAckCode1 = \{orXXXXSBCAckCode1} ,
  orXXXXSBCAckCode2 = \{orXXXXSBCAckCode2} ,
  orXXXXSBCAckCode3 = \{orXXXXSBCAckCode3} ,
  wdcntXXXXwd_cnt0 = \[14984]* ,
  wdcntXXXXwd_cnt1 = \[14797]* ,
  wdcntXXXXwd_cnt2 = \[14857]* ,
  nubusXXXXNuBusActive = \{nubusXXXXNuBusActive} ,
  orXXXXEn_START = \{orXXXXEn_START} ,
  \{nubusXXXXNextState0}  = (\[139]  & (~nubusXXXXstate0 & ~TM1i)) | (\[209]  | \[207] ),
  \[14676]  = (~\[14852]  & (~\{slaveXXXXSBCReqCode1}  & ~CoherencyState1i)) | ((TM1l & CoherencyState2i) | \[10750]_inv ),
  orXXXXSBCAck = \{orXXXXSBCAck} ,
  \{orXXXXL_DBufo}  = (\[191]  & ~\[14443] ) | ((~\[15192]  & ~PCCAck) | (\{virmachXXXXSBCConfigure}  & ~\[15169] )),
  slaveXXXXSnoopState_W = \{slaveXXXXSnoopState_W} ,
  \[10507]_inv  = \[143]  | (\[130]  | (SingleStep | SBCResetPCC)),
  \{nubusXXXXNextState1}  = (\[154]  & (\[122]  & (~\[2536]  & ~ACKi))) | (\[122]  & (~\[2536]  & (SlotSpace_Id_Match & ~ACKi))),
  \[130]  = ~masterXXXXstate3 | masterXXXXstate0,
  \[10749]_inv  = \[143]  | (~\[113]  | SingleStep),
  \[131]  = \[119]  | masterXXXXstate1,
  slaveXXXXSnoopVTag_W = \[14681] ,
  \[15041]  = \[212]  & (~VSACKi & ~SingleStep),
  \[14681]  = (\[129]  & (\[112]  & (~\[14764]  & (UpdateReq & VTM0l)))) | ((\[129]  & (\[124]  & (~\[14764]  & UpdateReq))) | (\[162]  & (\[136]  & UpdateReq))),
  \[133]  = Intr_done | ~nubusXXXXstate1,
  \[134]  = (~\[173]  & ~\[15074] ) | (~\[119]  & masterXXXXstate1),
  \[135]  = ~\[10889]_inv  & masterXXXXstate3,
  \[136]  = slaveXXXXstate2 & slaveXXXXstate1,
  \{slaveXXXXSnoopState_W}  = ~\[14676]  | \[14681] ,
  \[137]  = \[10748]_inv  | SBCResetPCC,
  \[138]  = \[10749]_inv  | ~\[15021] ,
  nextstateXXXXCoherencyState2o = \[15334] ,
  orXXXXVACKo = \{orXXXXVACKo} ,
  \[14417]  = \[14443]  & PCCReqCode1,
  \[139]  = \[112]  & STARTi,
  \[14857]*  = (\[142]  & (~\[14797]*  & wdcntXXXXstate2)) | (\[142]  & wdcntXXXXstate1),
  \{orXXXXVACKo}  = \[15041]  | \[15169] ,
  \[15334]  = \[176]  & CoherencyState2i,
  \{orXXXXSBCAckCodelatch}  = (~physrecXXXXstate1 & (ACKi & ~SBCResetPCC)) | ((~physrecXXXXstate0 & (ACKi & ~SBCResetPCC)) | (\[15041]  | (\[2836]  | \[14469] ))),
  \[140]  = \[117]  & ACKi,
  \[14976]  = ~\[203]  & (~resetXXXXstate2 & RESETi),
  masterXXXXSBC_WriteCache = \{masterXXXXSBC_WriteCache} ,
  \[141]  = \[15021]  & ~SingleStep,
  \[14902]  = \[10889]_inv ,
  wdcntXXXXNextState1 = \[14857]* ,
  wdcntXXXXNextState2 = \[14797]* ,
  \[142]  = Reset_wd_cnt & SBCResetPCC,
  wdcntXXXXNextState3 = \[14984]* ,
  \[143]  = PCCReqCode3 | ~PCCReq,
  virmachXXXXSBCsetDirty = \[15228] ,
  \[144]  = (\[176]  & ~CoherencyState2i) | ((~CoherencyState2i & ~CoherencyState1i) | ~Tag_Match);
always begin
  masterXXXXstate0 = \[84] ;
  masterXXXXstate1 = \[85] ;
  masterXXXXstate2 = \[86] ;
  masterXXXXstate3 = \[87] ;
  V_transmit_begin = \[111] ;
  wdcntXXXXstate0 = \[98] ;
  P_receive_begin = \[108] ;
  UpdateDone = \[103] ;
  UpdateReq = \[102] ;
  virmachXXXXstate0 = \[96] ;
  virmachXXXXstate1 = \[97] ;
  resetXXXXstate0 = \[93] ;
  resetXXXXstate1 = \[94] ;
  resetXXXXstate2 = \[95] ;
  wd_cnt_test = \[107] ;
  Reset_wd_cnt = \[104] ;
  Set_ex_wd_cnt1 = \[105] ;
  Intr_req = \[100] ;
  Intr_done = \[101] ;
  Gen_Reset = \[99] ;
  Incr_wd_cnt = \[106] ;
  slaveXXXXstate0 = \[90] ;
  slaveXXXXstate1 = \[91] ;
  slaveXXXXstate2 = \[92] ;
  nubusXXXXstate0 = \[88] ;
  nubusXXXXstate1 = \[89] ;
  P_receive_cancel = \[109] ;
end
initial begin
  masterXXXXstate0 = 0;
  masterXXXXstate1 = 0;
  masterXXXXstate2 = 0;
  masterXXXXstate3 = 0;
  V_transmit_begin = 0;
  wdcntXXXXstate0 = 0;
  P_receive_begin = 0;
  UpdateDone = 0;
  UpdateReq = 0;
  virmachXXXXstate0 = 0;
  virmachXXXXstate1 = 0;
  resetXXXXstate0 = 0;
  resetXXXXstate1 = 0;
  resetXXXXstate2 = 0;
  wd_cnt_test = 0;
  Reset_wd_cnt = 0;
  Set_ex_wd_cnt1 = 0;
  Intr_req = 0;
  Intr_done = 0;
  Gen_Reset = 0;
  Incr_wd_cnt = 0;
  slaveXXXXstate0 = 0;
  slaveXXXXstate1 = 0;
  slaveXXXXstate2 = 0;
  nubusXXXXstate0 = 0;
  nubusXXXXstate1 = 0;
  P_receive_cancel = 0;
end
endmodule

