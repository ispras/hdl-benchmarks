module test ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , 
 n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , 
 n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , 
 n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , 
 n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , 
 n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , 
 n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , 
 n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , 
 n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , 
 n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , 
 n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , 
 n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , 
 n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , 
 n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , 
 n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , 
 n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , 
 n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , 
 n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , 
 n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , 
 n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , 
 n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , 
 n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , 
 n221 , n222 , n223 , n224 , n225 , n226 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , 
 n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , 
 n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , 
 n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , 
 n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , 
 n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , 
 n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , 
 n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , 
 n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , 
 n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 ;
output n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , 
 n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , 
 n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , 
 n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , 
 n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , 
 n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , 
 n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , 
 n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , 
 n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , 
 n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , 
 n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , 
 n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , 
 n220 , n221 , n222 , n223 , n224 , n225 , n226 ;
wire n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , 
 n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , 
 n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , 
 n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , 
 n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , 
 n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , 
 n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , 
 n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , 
 n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , 
 n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , 
 n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , 
 n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , 
 n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , 
 n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , 
 n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , 
 n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , 
 n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , 
 n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , 
 n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , 
 n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , 
 n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , 
 n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , 
 n675 , n676 , n677 , n678 , n679 , n680 , n29489 , n29490 , n29491 , n29492 , 
 n29493 , n29494 , n29495 , n29496 , n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , 
 n29503 , n29504 , n29505 , n29506 , n29507 , n29508 , n29509 , n29510 , n29511 , n29512 , 
 n29513 , n29514 , n29515 , n29516 , n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , 
 n29523 , n29524 , n29525 , n29526 , n29527 , n29528 , n29529 , n29530 , n29531 , n29532 , 
 n29533 , n29534 , n29535 , n29536 , n29537 , n29538 , n29539 , n29540 , n29541 , n29542 , 
 n29543 , n29544 , n29545 , n29546 , n29547 , n29548 , n29549 , n29550 , n29551 , n29552 , 
 n29553 , n29554 , n29555 , n29556 , n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , 
 n29563 , n29564 , n29565 , n29566 , n29567 , n29568 , n29569 , n29570 , n29571 , n29572 , 
 n29573 , n29574 , n29575 , n29576 , n29577 , n29578 , n29579 , n29580 , n29581 , n29582 , 
 n29583 , n29584 , n29585 , n29586 , n29587 , n29588 , n29589 , n29590 , n29591 , n29592 , 
 n29593 , n29594 , n29595 , n29596 , n29597 , n29598 , n29599 , n29600 , n29601 , n29602 , 
 n29603 , n29604 , n29605 , n29606 , n29607 , n29608 , n29609 , n29610 , n29611 , n29612 , 
 n29613 , n29614 , n29615 , n29616 , n29617 , n29618 , n29619 , n29620 , n29621 , n29622 , 
 n29623 , n29624 , n29625 , n29626 , n29627 , n29628 , n29629 , n29630 , n29631 , n29632 , 
 n29633 , n29634 , n29635 , n29636 , n29637 , n29638 , n29639 , n29640 , n29641 , n29642 , 
 n29643 , n29644 , n29645 , n29646 , n29647 , n29648 , n29649 , n29650 , n29651 , n29652 , 
 n29653 , n29654 , n29655 , n29656 , n29657 , n29658 , n29659 , n29660 , n29661 , n29662 , 
 n29663 , n29664 , n29665 , n29666 , n29667 , n29668 , n29669 , n29670 , n29671 , n29672 , 
 n29673 , n29674 , n29675 , n29676 , n29677 , n29678 , n29679 , n29680 , n29681 , n29682 , 
 n29683 , n29684 , n29685 , n29686 , n29687 , n29688 , n29689 , n29690 , n29691 , n29692 , 
 n29693 , n29694 , n29695 , n29696 , n29697 , n29698 , n29699 , n29700 , n29701 , n29702 , 
 n29703 , n29704 , n29705 , n29706 , n29707 , n29708 , n29709 , n29710 , n29711 , n29712 , 
 n29713 , n29714 , n29715 , n29716 , n29717 , n29718 , n29719 , n29720 , n29721 , n29722 , 
 n29723 , n29724 , n29725 , n29726 , n29727 , n29728 , n29729 , n29730 , n29731 , n29732 , 
 n29733 , n29734 , n29735 , n29736 , n29737 , n29738 , n29739 , n29740 , n29741 , n29742 , 
 n29743 , n29744 , n29745 , n29746 , n29747 , n29748 , n29749 , n29750 , n29751 , n29752 , 
 n29753 , n29754 , n29755 , n29756 , n29757 , n29758 , n29759 , n29760 , n29761 , n29762 , 
 n29763 , n29764 , n29765 , n684 , n29767 , n686 , n687 , n29770 , n689 , n690 , 
 n691 , n692 , n693 , n29776 , n695 , n696 , n697 , n698 , n699 , n700 , 
 n701 , n29784 , n703 , n29786 , n705 , n706 , n707 , n708 , n709 , n29792 , 
 n711 , n712 , n29795 , n714 , n29797 , n716 , n717 , n718 , n29801 , n720 , 
 n29803 , n722 , n723 , n724 , n725 , n29808 , n727 , n29810 , n729 , n730 , 
 n731 , n732 , n733 , n734 , n29817 , n736 , n29819 , n29820 , n29821 , n743 , 
 n29823 , n29824 , n29825 , n29826 , n29827 , n29828 , n29829 , n751 , n752 , n753 , 
 n754 , n758 , n29835 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , 
 n770 , n29844 , n29845 , n29846 , n774 , n775 , n776 , n777 , n778 , n782 , 
 n29853 , n784 , n29855 , n786 , n787 , n29858 , n789 , n790 , n791 , n792 , 
 n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n29871 , n802 , 
 n29873 , n804 , n29875 , n806 , n29877 , n29878 , n809 , n29880 , n814 , n29882 , 
 n29883 , n817 , n818 , n819 , n820 , n29888 , n822 , n823 , n824 , n825 , 
 n29893 , n827 , n828 , n829 , n29897 , n831 , n29899 , n29900 , n834 , n835 , 
 n29903 , n29904 , n29905 , n842 , n29907 , n844 , n845 , n846 , n847 , n29912 , 
 n849 , n29914 , n851 , n852 , n29917 , n854 , n855 , n29920 , n857 , n858 , 
 n29923 , n860 , n29925 , n29926 , n863 , n29928 , n868 , n29930 , n29931 , n871 , 
 n29933 , n29934 , n29935 , n875 , n876 , n29938 , n878 , n29940 , n29941 , n29942 , 
 n29943 , n883 , n29945 , n29946 , n886 , n887 , n888 , n29950 , n890 , n891 , 
 n892 , n893 , n894 , n895 , n896 , n897 , n29959 , n899 , n900 , n901 , 
 n902 , n903 , n904 , n29966 , n29967 , n907 , n908 , n909 , n910 , n914 , 
 n29973 , n29974 , n917 , n29976 , n919 , n29978 , n29979 , n922 , n923 , n924 , 
 n925 , n29984 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , 
 n29993 , n936 , n29995 , n29996 , n939 , n29998 , n941 , n942 , n943 , n944 , 
 n945 , n30004 , n950 , n30006 , n952 , n30008 , n954 , n955 , n956 , n957 , 
 n30013 , n959 , n30015 , n961 , n30017 , n963 , n964 , n30020 , n30021 , n967 , 
 n30023 , n969 , n970 , n971 , n30027 , n973 , n974 , n30030 , n976 , n30032 , 
 n30033 , n30034 , n980 , n30036 , n30037 , n30038 , n30039 , n30040 , n986 , n30042 , 
 n30043 , n989 , n30045 , n994 , n30047 , n996 , n30049 , n998 , n999 , n1000 , 
 n1001 , n1002 , n1003 , n1004 , n30057 , n1006 , n30059 , n1008 , n1009 , n30062 , 
 n30063 , n1012 , n30065 , n30066 , n1015 , n30068 , n30069 , n30070 , n1019 , n30072 , 
 n1024 , n1025 , n30075 , n1027 , n1028 , n1029 , n1030 , n1031 , n30081 , n1033 , 
 n1034 , n1035 , n1036 , n1037 , n30087 , n1039 , n30089 , n1041 , n30091 , n1043 , 
 n30093 , n1045 , n1046 , n30096 , n30097 , n1049 , n30099 , n30100 , n1052 , n30102 , 
 n30103 , n1055 , n1056 , n30106 , n30107 , n1059 , n30109 , n30110 , n1062 , n30112 , 
 n30113 , n1065 , n30115 , n1067 , n1068 , n1069 , n30119 , n30120 , n1072 , n30122 , 
 n30123 , n30124 , n1076 , n30126 , n30127 , n30128 , n1080 , n30130 , n1085 , n30132 , 
 n1087 , n1088 , n30135 , n30136 , n1091 , n30138 , n30139 , n1094 , n30141 , n30142 , 
 n1097 , n1098 , n30145 , n30146 , n1101 , n30148 , n30149 , n1104 , n30151 , n30152 , 
 n1107 , n30154 , n30155 , n1110 , n30157 , n30158 , n1113 , n30160 , n30161 , n1116 , 
 n30163 , n1118 , n30165 , n1120 , n1121 , n30168 , n30169 , n1127 , n30171 , n30172 , 
 n1130 , n30174 , n1132 , n1133 , n30177 , n30178 , n30179 , n30180 , n1138 , n30182 , 
 n1140 , n30184 , n1142 , n30186 , n1144 , n1145 , n30189 , n1147 , n30191 , n1149 , 
 n30193 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n30202 , 
 n1160 , n30204 , n30205 , n1163 , n1164 , n1165 , n30209 , n30210 , n1168 , n30212 , 
 n1170 , n30214 , n30215 , n1173 , n1174 , n1175 , n30219 , n1177 , n1178 , n1179 , 
 n30223 , n1181 , n1182 , n1183 , n1187 , n30228 , n1189 , n1190 , n1191 , n30232 , 
 n30233 , n1194 , n30235 , n1196 , n30237 , n1198 , n1199 , n1200 , n1201 , n1202 , 
 n1203 , n1204 , n30245 , n30246 , n1207 , n30248 , n30249 , n1210 , n30251 , n30252 , 
 n1213 , n1214 , n30255 , n30256 , n30257 , n30258 , n30259 , n1223 , n30261 , n30262 , 
 n30263 , n30264 , n30265 , n1229 , n1230 , n30268 , n1232 , n30270 , n1234 , n1235 , 
 n30273 , n30274 , n30275 , n1239 , n30277 , n30278 , n1242 , n30280 , n30281 , n30282 , 
 n1246 , n30284 , n30285 , n1249 , n30287 , n30288 , n1252 , n1253 , n1254 , n1255 , 
 n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , 
 n1266 , n1267 , n30305 , n1269 , n1270 , n1271 , n1272 , n30310 , n1274 , n30312 , 
 n1276 , n1277 , n30315 , n1279 , n30317 , n1281 , n30319 , n1283 , n30321 , n30322 , 
 n1286 , n1287 , n1288 , n30326 , n30327 , n1291 , n30329 , n30330 , n30331 , n1295 , 
 n1296 , n1297 , n30335 , n30336 , n1300 , n1301 , n1302 , n30340 , n1304 , n1305 , 
 n1309 , n30344 , n30345 , n1312 , n1313 , n30348 , n30349 , n1316 , n1317 , n1318 , 
 n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n30359 , n30360 , n1327 , n1328 , 
 n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n30369 , n30370 , n1337 , n30372 , 
 n1342 , n30374 , n1344 , n1345 , n30377 , n30378 , n30379 , n30380 , n30381 , n1351 , 
 n30383 , n30384 , n1354 , n1355 , n30387 , n1357 , n1358 , n1359 , n1360 , n1361 , 
 n1362 , n1363 , n1364 , n1365 , n1366 , n30398 , n1368 , n1369 , n30401 , n30402 , 
 n1372 , n30404 , n30405 , n1375 , n30407 , n30408 , n1378 , n30410 , n1380 , n30412 , 
 n30413 , n1383 , n1384 , n1385 , n30417 , n30418 , n1388 , n1389 , n1390 , n30422 , 
 n1392 , n1393 , n1394 , n30426 , n30427 , n30428 , n1398 , n30430 , n30431 , n1401 , 
 n1402 , n1403 , n1404 , n1405 , n1409 , n30438 , n1411 , n1412 , n1413 , n1414 , 
 n1415 , n30444 , n30445 , n1418 , n30447 , n1420 , n1421 , n1422 , n1423 , n1424 , 
 n30453 , n1426 , n30455 , n1428 , n1429 , n30458 , n30459 , n1432 , n30461 , n30462 , 
 n1435 , n30464 , n30465 , n30466 , n1439 , n30468 , n1441 , n1442 , n1443 , n1444 , 
 n1445 , n1446 , n1447 , n1448 , n1449 , n30478 , n1451 , n1452 , n1453 , n30482 , 
 n30483 , n1459 , n1460 , n1461 , n30487 , n1463 , n1464 , n1465 , n1466 , n1467 , 
 n30493 , n1469 , n1470 , n1471 , n1472 , n1473 , n30499 , n1475 , n30501 , n1477 , 
 n1478 , n30504 , n1480 , n1481 , n1482 , n1483 , n1484 , n30510 , n1486 , n1487 , 
 n1488 , n30514 , n30515 , n1491 , n30517 , n30518 , n1494 , n30520 , n30521 , n30522 , 
 n1498 , n30524 , n30525 , n1501 , n30527 , n30528 , n1504 , n30530 , n1506 , n30532 , 
 n1508 , n1509 , n30535 , n30536 , n1512 , n30538 , n30539 , n1515 , n30541 , n30542 , 
 n1518 , n1519 , n30545 , n30546 , n1522 , n30548 , n30549 , n30550 , n30551 , n30552 , 
 n30553 , n30554 , n1530 , n30556 , n1532 , n30558 , n30559 , n30560 , n30561 , n1537 , 
 n30563 , n1539 , n30565 , n30566 , n1542 , n30568 , n30569 , n1545 , n30571 , n1547 , 
 n1548 , n1549 , n1550 , n30576 , n1552 , n30578 , n1554 , n1555 , n30581 , n30582 , 
 n1558 , n30584 , n30585 , n1561 , n30587 , n30588 , n1564 , n30590 , n30591 , n1567 , 
 n1568 , n30594 , n1573 , n30596 , n30597 , n1576 , n30599 , n30600 , n30601 , n1580 , 
 n30603 , n1582 , n1583 , n30606 , n1585 , n30608 , n1587 , n1588 , n30611 , n30612 , 
 n1591 , n30614 , n30615 , n1594 , n30617 , n30618 , n30619 , n1598 , n30621 , n30622 , 
 n1604 , n30624 , n30625 , n1607 , n1608 , n30628 , n30629 , n1611 , n1612 , n1613 , 
 n30633 , n1615 , n1616 , n1617 , n30637 , n1619 , n1620 , n1621 , n1622 , n1623 , 
 n1624 , n1625 , n30645 , n1627 , n30647 , n30648 , n30649 , n30650 , n30651 , n1633 , 
 n30653 , n1635 , n1636 , n30656 , n1638 , n30658 , n1640 , n1641 , n30661 , n30662 , 
 n1644 , n30664 , n30665 , n1647 , n30667 , n1649 , n30669 , n1651 , n30671 , n30672 , 
 n30673 , n30674 , n1656 , n30676 , n1658 , n1659 , n30679 , n1661 , n30681 , n1663 , 
 n1664 , n30684 , n30685 , n1667 , n30687 , n30688 , n1670 , n30690 , n30691 , n30692 , 
 n1677 , n30694 , n30695 , n1680 , n30697 , n30698 , n1683 , n30700 , n1685 , n30702 , 
 n30703 , n1688 , n30705 , n1690 , n30707 , n30708 , n30709 , n30710 , n1695 , n30712 , 
 n1697 , n30714 , n30715 , n1700 , n30717 , n30718 , n30719 , n1704 , n30721 , n1706 , 
 n1707 , n30724 , n1709 , n30726 , n1711 , n1712 , n30729 , n30730 , n1715 , n30732 , 
 n30733 , n1718 , n30735 , n30736 , n30737 , n1722 , n30739 , n30740 , n1725 , n30742 , 
 n30743 , n1728 , n30745 , n1730 , n1731 , n1732 , n1733 , n30750 , n30751 , n30752 , 
 n30753 , n1741 , n1742 , n30756 , n30757 , n1745 , n30759 , n30760 , n1748 , n30762 , 
 n1750 , n1751 , n30765 , n30766 , n30767 , n1755 , n30769 , n1757 , n1758 , n1759 , 
 n30773 , n1761 , n30775 , n1763 , n1764 , n30778 , n30779 , n1767 , n30781 , n30782 , 
 n1770 , n30784 , n1772 , n1773 , n1774 , n30788 , n1776 , n30790 , n1778 , n30792 , 
 n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , 
 n1790 , n30804 , n1792 , n1793 , n1794 , n1795 , n1796 , n30810 , n1798 , n1799 , 
 n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , 
 n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n30830 , n1818 , n1819 , 
 n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n30839 , n30840 , n30841 , n1829 , 
 n30843 , n1831 , n30845 , n30846 , n30847 , n30848 , n1836 , n30850 , n30851 , n30852 , 
 n1840 , n30854 , n30855 , n1843 , n30857 , n1845 , n1846 , n1847 , n30861 , n1849 , 
 n1850 , n30864 , n30865 , n1853 , n30867 , n30868 , n30869 , n1857 , n30871 , n30872 , 
 n1860 , n30874 , n30875 , n1863 , n30877 , n1865 , n30879 , n1870 , n30881 , n30882 , 
 n1873 , n30884 , n30885 , n30886 , n1877 , n30888 , n30889 , n1880 , n1881 , n30892 , 
 n1883 , n1884 , n1885 , n30896 , n30897 , n1888 , n30899 , n30900 , n1891 , n30902 , 
 n1893 , n30904 , n30905 , n1896 , n30907 , n1898 , n30909 , n30910 , n30911 , n30912 , 
 n1906 , n1907 , n1908 , n1909 , n30917 , n1911 , n30919 , n1913 , n1914 , n1915 , 
 n30923 , n1917 , n30925 , n1919 , n30927 , n1921 , n1922 , n1923 , n1924 , n30932 , 
 n30933 , n30934 , n1928 , n30936 , n30937 , n1931 , n30939 , n1933 , n1934 , n1935 , 
 n30943 , n30944 , n1938 , n30946 , n30947 , n1941 , n30949 , n1943 , n1944 , n30952 , 
 n1946 , n30954 , n1948 , n1949 , n30957 , n30958 , n1952 , n30960 , n30961 , n1955 , 
 n30963 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , 
 n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n30982 , 
 n30983 , n30984 , n30985 , n30986 , n30987 , n1981 , n30989 , n1983 , n30991 , n30992 , 
 n1986 , n30994 , n30995 , n30996 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , 
 n1999 , n2000 , n2001 , n31006 , n2003 , n2004 , n31009 , n2006 , n31011 , n31012 , 
 n31013 , n31014 , n2011 , n31016 , n31017 , n2014 , n31019 , n31020 , n2017 , n31022 , 
 n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , 
 n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , 
 n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n31049 , n2046 , n31051 , n2048 , 
 n2049 , n31054 , n2051 , n31056 , n2053 , n31058 , n31059 , n2056 , n31061 , n2058 , 
 n31063 , n2063 , n31065 , n2065 , n31067 , n2067 , n2068 , n31070 , n31071 , n31072 , 
 n2072 , n31074 , n31075 , n2075 , n31077 , n31078 , n2078 , n31080 , n2080 , n2081 , 
 n31083 , n31084 , n2084 , n31086 , n2086 , n31088 , n2088 , n31090 , n2090 , n2091 , 
 n2092 , n31094 , n31095 , n2095 , n31097 , n31098 , n2098 , n31100 , n2100 , n2101 , 
 n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n31112 , 
 n31113 , n2113 , n31115 , n2115 , n31117 , n31118 , n31119 , n31120 , n2120 , n31122 , 
 n31123 , n31124 , n2124 , n31126 , n2126 , n2127 , n2128 , n2129 , n2130 , n31132 , 
 n31133 , n2133 , n31135 , n31136 , n31137 , n2137 , n31139 , n2139 , n2140 , n2141 , 
 n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n31151 , n2151 , 
 n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n31159 , n2159 , n2160 , n31162 , 
 n2162 , n31164 , n31165 , n2165 , n2166 , n31168 , n31169 , n31170 , n2170 , n31172 , 
 n31173 , n2173 , n31175 , n31176 , n2176 , n31178 , n31179 , n31180 , n2180 , n31182 , 
 n2182 , n31184 , n31185 , n31186 , n31187 , n2187 , n31189 , n31190 , n2190 , n31192 , 
 n31193 , n2193 , n31195 , n31196 , n2196 , n31198 , n31199 , n2199 , n31201 , n31202 , 
 n2202 , n2206 , n31205 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n31212 , 
 n2215 , n2216 , n31215 , n31216 , n2219 , n31218 , n31219 , n2222 , n31221 , n2224 , 
 n31223 , n31224 , n2227 , n31226 , n31227 , n2230 , n31229 , n2232 , n2233 , n2234 , 
 n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n31241 , n2247 , 
 n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , 
 n2258 , n2259 , n2260 , n2261 , n2262 , n31258 , n31259 , n2265 , n31261 , n2267 , 
 n2268 , n2269 , n2270 , n2271 , n31267 , n31268 , n31269 , n2275 , n31271 , n31272 , 
 n31273 , n2279 , n31275 , n31276 , n2282 , n31278 , n2284 , n31280 , n31281 , n31282 , 
 n2288 , n31284 , n2290 , n31286 , n31287 , n31288 , n31289 , n2295 , n31291 , n31292 , 
 n2298 , n31294 , n31295 , n2301 , n2302 , n31298 , n31299 , n2305 , n31301 , n31302 , 
 n2308 , n2309 , n2310 , n2311 , n31307 , n31308 , n2314 , n31310 , n2316 , n31312 , 
 n2318 , n2319 , n31315 , n31316 , n31317 , n2323 , n31319 , n31320 , n2326 , n31322 , 
 n31323 , n2329 , n31325 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , 
 n31333 , n2339 , n31335 , n2341 , n2342 , n31338 , n31339 , n31340 , n2346 , n31342 , 
 n31343 , n2349 , n31345 , n31346 , n2352 , n31348 , n2354 , n2355 , n2356 , n2357 , 
 n2358 , n31354 , n2360 , n31356 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , 
 n2368 , n31364 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n31372 , 
 n2378 , n31374 , n2380 , n2381 , n31377 , n31378 , n2384 , n31380 , n31381 , n31382 , 
 n2388 , n31384 , n31385 , n2391 , n31387 , n31388 , n31389 , n31390 , n2396 , n31392 , 
 n31393 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n31400 , n2409 , n2410 , 
 n2411 , n2412 , n31405 , n2414 , n2415 , n31408 , n31409 , n31410 , n2419 , n31412 , 
 n31413 , n2422 , n31415 , n31416 , n2425 , n31418 , n31419 , n2428 , n31421 , n2430 , 
 n31423 , n2432 , n2433 , n31426 , n31427 , n31428 , n2437 , n31430 , n31431 , n2440 , 
 n31433 , n31434 , n2443 , n31436 , n31437 , n2446 , n31439 , n2448 , n2449 , n2450 , 
 n2451 , n2452 , n2453 , n31446 , n2455 , n31448 , n2457 , n2458 , n31451 , n31452 , 
 n31453 , n2462 , n31455 , n31456 , n2465 , n31458 , n31459 , n2468 , n31461 , n31462 , 
 n31463 , n31464 , n2473 , n31466 , n2475 , n31468 , n31469 , n31470 , n2479 , n31472 , 
 n2481 , n2482 , n2483 , n2484 , n31477 , n31478 , n31479 , n31480 , n31481 , n31482 , 
 n2491 , n31484 , n2493 , n2494 , n31487 , n2496 , n2497 , n2498 , n2499 , n2500 , 
 n31493 , n31494 , n2503 , n31496 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , 
 n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , 
 n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n31519 , n2528 , n31521 , n2530 , 
 n2531 , n31524 , n31525 , n2534 , n31527 , n31528 , n31529 , n2538 , n31531 , n31532 , 
 n2541 , n31534 , n31535 , n31536 , n2545 , n31538 , n2547 , n2548 , n31541 , n31542 , 
 n31543 , n2552 , n31545 , n31546 , n2555 , n31548 , n31549 , n2558 , n31551 , n31552 , 
 n2561 , n2562 , n2563 , n2564 , n2565 , n31558 , n2567 , n31560 , n31561 , n2573 , 
 n31563 , n2575 , n31565 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n31572 , 
 n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n31581 , n31582 , 
 n2594 , n31584 , n31585 , n2597 , n31587 , n2599 , n2600 , n31590 , n31591 , n31592 , 
 n2604 , n31594 , n31595 , n2607 , n31597 , n31598 , n2610 , n31600 , n2612 , n31602 , 
 n2614 , n31604 , n2616 , n2617 , n31607 , n31608 , n31609 , n2621 , n31611 , n31612 , 
 n2624 , n31614 , n31615 , n2627 , n31617 , n2629 , n2630 , n2631 , n2632 , n2633 , 
 n2634 , n31624 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , 
 n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n31640 , n2652 , n2653 , 
 n2654 , n2655 , n31645 , n31646 , n2658 , n31648 , n31649 , n2661 , n2662 , n2663 , 
 n2664 , n2665 , n2666 , n2667 , n2668 , n31658 , n2670 , n31660 , n31661 , n2673 , 
 n2674 , n31664 , n2676 , n31666 , n2678 , n31668 , n31669 , n2681 , n31671 , n31672 , 
 n31673 , n2685 , n31675 , n2687 , n2688 , n31678 , n31679 , n31680 , n2692 , n31682 , 
 n31683 , n2695 , n31685 , n31686 , n2698 , n31688 , n31689 , n2701 , n31691 , n31692 , 
 n2704 , n31694 , n2706 , n31696 , n31697 , n31698 , n31699 , n2711 , n31701 , n31702 , 
 n31703 , n2715 , n31705 , n31706 , n31707 , n2719 , n31709 , n2721 , n2722 , n31712 , 
 n2724 , n31714 , n2726 , n31716 , n31717 , n2729 , n31719 , n31720 , n2732 , n31722 , 
 n31723 , n2738 , n31725 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , 
 n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n31739 , n2754 , n31741 , n2756 , 
 n31743 , n2758 , n2759 , n2760 , n31747 , n31748 , n2763 , n31750 , n31751 , n2766 , 
 n31753 , n31754 , n2769 , n31756 , n2771 , n2772 , n31759 , n2774 , n31761 , n2776 , 
 n31763 , n31764 , n2779 , n31766 , n2781 , n2782 , n31769 , n2784 , n31771 , n2786 , 
 n2787 , n31774 , n31775 , n31776 , n2791 , n31778 , n31779 , n2794 , n31781 , n31782 , 
 n2797 , n31784 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , 
 n2807 , n2808 , n2809 , n2810 , n2811 , n31798 , n2813 , n2814 , n2815 , n2816 , 
 n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n31811 , n31812 , 
 n31813 , n2828 , n31815 , n2830 , n31817 , n31818 , n31819 , n31820 , n2835 , n31822 , 
 n31823 , n31824 , n2839 , n31826 , n31827 , n2842 , n31829 , n31830 , n2845 , n2846 , 
 n31833 , n2848 , n31835 , n31836 , n2851 , n31838 , n2853 , n31840 , n31841 , n31842 , 
 n2857 , n2858 , n31845 , n31846 , n2861 , n31848 , n31849 , n2864 , n31851 , n2866 , 
 n31853 , n31854 , n31855 , n2870 , n2871 , n31858 , n31859 , n31860 , n2875 , n2876 , 
 n31863 , n31864 , n2879 , n31866 , n2881 , n31868 , n31869 , n31870 , n2885 , n31872 , 
 n2887 , n31874 , n31875 , n31876 , n2894 , n2895 , n31879 , n31880 , n2898 , n31882 , 
 n31883 , n2901 , n2902 , n2903 , n31887 , n2905 , n31889 , n2907 , n2908 , n2909 , 
 n2910 , n2911 , n31895 , n2913 , n31897 , n31898 , n2916 , n2917 , n2918 , n31902 , 
 n31903 , n31904 , n2922 , n31906 , n2924 , n31908 , n31909 , n31910 , n2928 , n2929 , 
 n31913 , n31914 , n2932 , n2933 , n31917 , n31918 , n2936 , n2937 , n2938 , n31922 , 
 n31923 , n31924 , n31925 , n31926 , n2944 , n31928 , n2946 , n31930 , n31931 , n31932 , 
 n31933 , n2951 , n31935 , n31936 , n31937 , n2955 , n31939 , n31940 , n2958 , n31942 , 
 n31943 , n2961 , n2962 , n31946 , n31947 , n31948 , n31949 , n31950 , n2968 , n2969 , 
 n31953 , n31954 , n2972 , n2973 , n31957 , n31958 , n31959 , n2977 , n2978 , n31962 , 
 n31963 , n2981 , n31965 , n31966 , n2984 , n2985 , n31969 , n2987 , n2988 , n31972 , 
 n31973 , n2991 , n31975 , n31976 , n2994 , n31978 , n31979 , n2997 , n31981 , n31982 , 
 n3000 , n3001 , n31985 , n31986 , n3004 , n31988 , n31989 , n31990 , n3008 , n31992 , 
 n3010 , n3011 , n31995 , n31996 , n3014 , n3015 , n31999 , n32000 , n3018 , n32002 , 
 n3020 , n32004 , n32005 , n32006 , n3024 , n32008 , n32009 , n3027 , n3028 , n32012 , 
 n3030 , n3031 , n32015 , n32016 , n3034 , n3035 , n32019 , n32020 , n3041 , n32022 , 
 n32023 , n3044 , n3045 , n32026 , n32027 , n3048 , n32029 , n32030 , n32031 , n3052 , 
 n32033 , n32034 , n3055 , n3056 , n32037 , n32038 , n3059 , n3060 , n32041 , n32042 , 
 n3063 , n3064 , n32045 , n32046 , n3067 , n32048 , n3069 , n32050 , n32051 , n3072 , 
 n32053 , n32054 , n32055 , n3076 , n32057 , n3078 , n32059 , n32060 , n32061 , n3082 , 
 n3083 , n32064 , n32065 , n3086 , n3087 , n32068 , n32069 , n32070 , n3091 , n32072 , 
 n3093 , n32074 , n32075 , n32076 , n3097 , n3098 , n32079 , n32080 , n3101 , n3102 , 
 n32083 , n32084 , n32085 , n32086 , n32087 , n3108 , n32089 , n3110 , n32091 , n32092 , 
 n32093 , n3114 , n3115 , n32096 , n3117 , n3118 , n32099 , n32100 , n3121 , n32102 , 
 n32103 , n3124 , n3125 , n32106 , n3127 , n3128 , n3129 , n32110 , n3131 , n32112 , 
 n32113 , n3134 , n3135 , n3136 , n32117 , n3138 , n3139 , n3140 , n3141 , n3142 , 
 n3143 , n32124 , n32125 , n3146 , n32127 , n32128 , n3149 , n3150 , n32131 , n3152 , 
 n3153 , n3154 , n32135 , n3156 , n32137 , n32138 , n3159 , n32140 , n32141 , n3162 , 
 n32143 , n32144 , n32145 , n3166 , n3167 , n32148 , n3169 , n3170 , n32151 , n32152 , 
 n3176 , n3177 , n32155 , n3179 , n3180 , n3181 , n3182 , n3183 , n32161 , n3185 , 
 n32163 , n3187 , n32165 , n32166 , n32167 , n3191 , n32169 , n3193 , n32171 , n3195 , 
 n32173 , n32174 , n3198 , n3199 , n32177 , n3201 , n3202 , n32180 , n32181 , n3205 , 
 n32183 , n32184 , n3208 , n3209 , n32187 , n3211 , n3212 , n32190 , n32191 , n32192 , 
 n3216 , n3217 , n32195 , n3219 , n32197 , n32198 , n3222 , n32200 , n32201 , n32202 , 
 n3226 , n32204 , n32205 , n3229 , n3230 , n32208 , n32209 , n3233 , n3234 , n32212 , 
 n3236 , n32214 , n3238 , n3239 , n32217 , n3241 , n3242 , n3243 , n3244 , n3245 , 
 n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , 
 n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , 
 n3266 , n3267 , n3268 , n32246 , n32247 , n32248 , n3272 , n32250 , n32251 , n3275 , 
 n3276 , n32254 , n32255 , n3279 , n32257 , n32258 , n32259 , n3283 , n32261 , n32262 , 
 n3286 , n3287 , n32265 , n32266 , n3290 , n3291 , n32269 , n32270 , n32271 , n32272 , 
 n32273 , n3297 , n32275 , n32276 , n3303 , n3304 , n32279 , n32280 , n3307 , n32282 , 
 n32283 , n3310 , n32285 , n32286 , n3313 , n3314 , n32289 , n32290 , n32291 , n3318 , 
 n3319 , n32294 , n32295 , n3322 , n32297 , n32298 , n3325 , n32300 , n32301 , n32302 , 
 n3329 , n32304 , n32305 , n32306 , n3333 , n32308 , n32309 , n3336 , n32311 , n3338 , 
 n32313 , n32314 , n32315 , n3342 , n32317 , n32318 , n3345 , n32320 , n32321 , n3348 , 
 n32323 , n32324 , n3351 , n3352 , n3353 , n32328 , n32329 , n32330 , n32331 , n32332 , 
 n3359 , n3360 , n3361 , n32336 , n32337 , n3364 , n32339 , n32340 , n3367 , n3368 , 
 n32343 , n3370 , n32345 , n32346 , n32347 , n3374 , n32349 , n32350 , n3377 , n32352 , 
 n32353 , n3380 , n3381 , n32356 , n3383 , n3384 , n3385 , n3386 , n3387 , n32362 , 
 n32363 , n32364 , n3391 , n3392 , n32367 , n3394 , n3395 , n32370 , n32371 , n3398 , 
 n32373 , n32374 , n3401 , n3402 , n32377 , n3404 , n3405 , n3406 , n3407 , n3408 , 
 n3409 , n32384 , n3411 , n32386 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , 
 n3422 , n32394 , n32395 , n32396 , n32397 , n32398 , n3428 , n32400 , n32401 , n3431 , 
 n3432 , n32404 , n32405 , n3435 , n32407 , n32408 , n3438 , n3439 , n32411 , n32412 , 
 n3442 , n32414 , n32415 , n3445 , n32417 , n32418 , n3448 , n3449 , n32421 , n3451 , 
 n3452 , n3453 , n32425 , n3455 , n3456 , n3457 , n32429 , n3459 , n3460 , n3461 , 
 n3462 , n3463 , n3464 , n3465 , n3466 , n32438 , n3468 , n3469 , n3470 , n3471 , 
 n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , 
 n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , 
 n3492 , n3493 , n32465 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , 
 n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , 
 n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n32489 , n3522 , n3523 , n3524 , 
 n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , 
 n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , 
 n3545 , n32514 , n32515 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , 
 n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n32529 , n3562 , n3563 , n32532 , 
 n3565 , n3566 , n32535 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , 
 n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , 
 n3585 , n3586 , n3587 , n3588 , n3589 , n32558 , n32559 , n32560 , n3593 , n32562 , 
 n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , 
 n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n32580 , n3616 , n3617 , 
 n3618 , n3619 , n3620 , n3621 , n3622 , n32588 , n32589 , n3625 , n32591 , n32592 , 
 n3628 , n3629 , n32595 , n32596 , n32597 , n3633 , n32599 , n32600 , n3636 , n3637 , 
 n32603 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , 
 n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n32619 , n32620 , n32621 , n32622 , 
 n3658 , n32624 , n32625 , n3661 , n32627 , n32628 , n3664 , n32630 , n3666 , n3667 , 
 n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , 
 n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n32652 , 
 n32653 , n32654 , n3690 , n32656 , n32657 , n3693 , n32659 , n32660 , n32661 , n3697 , 
 n32663 , n32664 , n3703 , n3704 , n32667 , n3706 , n3707 , n3708 , n3709 , n3710 , 
 n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , 
 n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , 
 n3731 , n3732 , n3733 , n32696 , n32697 , n3736 , n32699 , n32700 , n32701 , n3740 , 
 n32703 , n32704 , n32705 , n3744 , n3745 , n32708 , n32709 , n3748 , n32711 , n32712 , 
 n3751 , n3752 , n32715 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , 
 n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , 
 n3771 , n32734 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , 
 n3784 , n3785 , n3786 , n3787 , n32747 , n3789 , n3790 , n3791 , n3792 , n3793 , 
 n3794 , n3795 , n3796 , n32756 , n32757 , n32758 , n3800 , n32760 , n3802 , n3803 , 
 n3804 , n3805 , n3806 , n32766 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , 
 n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , 
 n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , 
 n3834 , n3835 , n3836 , n3837 , n32797 , n3842 , n3843 , n3844 , n3845 , n3846 , 
 n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , 
 n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , 
 n32823 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , 
 n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , 
 n3887 , n3888 , n3889 , n3890 , n3891 , n32848 , n3896 , n3897 , n3898 , n3899 , 
 n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , 
 n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n32870 , n3918 , n3919 , 
 n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , 
 n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n32891 , n3942 , 
 n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , 
 n3953 , n3954 , n3955 , n3956 , n32907 , n3958 , n3959 , n3960 , n3961 , n3962 , 
 n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n32922 , 
 n3976 , n32924 , n3978 , n32926 , n3980 , n3981 , n3982 , n32930 , n32931 , n3985 , 
 n32933 , n3987 , n32935 , n3989 , n3990 , n3991 , n3992 , n32940 , n3994 , n3995 , 
 n3996 , n3997 , n3998 , n32946 , n32947 , n32948 , n32949 , n32950 , n32951 , n4005 , 
 n4006 , n32954 , n32955 , n4009 , n32957 , n32958 , n32959 , n4013 , n32961 , n32962 , 
 n4016 , n4017 , n32965 , n32966 , n4020 , n4021 , n32969 , n32970 , n32971 , n32972 , 
 n4026 , n32974 , n4028 , n4029 , n4030 , n32978 , n32979 , n4033 , n32981 , n4035 , 
 n32983 , n4037 , n32985 , n4039 , n4040 , n32988 , n32989 , n32990 , n4044 , n4045 , 
 n32993 , n4047 , n4048 , n32996 , n32997 , n4051 , n32999 , n33000 , n33001 , n4055 , 
 n33003 , n33004 , n4058 , n33006 , n33007 , n4061 , n33009 , n33010 , n4064 , n4065 , 
 n33013 , n4067 , n4068 , n33016 , n33017 , n33018 , n4072 , n4073 , n33021 , n33022 , 
 n33023 , n33024 , n4078 , n33026 , n4080 , n33028 , n33029 , n33030 , n33031 , n4085 , 
 n33033 , n33034 , n33035 , n4089 , n33037 , n33038 , n4092 , n33040 , n4094 , n33042 , 
 n33043 , n4097 , n33045 , n33046 , n33047 , n4101 , n4102 , n33050 , n4104 , n4105 , 
 n33053 , n33054 , n4108 , n4109 , n33057 , n4111 , n4112 , n4113 , n33061 , n4115 , 
 n33063 , n33064 , n33065 , n33066 , n4120 , n33068 , n33069 , n33070 , n4124 , n4125 , 
 n33073 , n4127 , n4128 , n33076 , n33077 , n4131 , n4132 , n33080 , n33081 , n33082 , 
 n33083 , n33084 , n33085 , n33086 , n33087 , n33088 , n33089 , n33090 , n33091 , n33092 , 
 n4146 , n33094 , n33095 , n4149 , n33097 , n33098 , n33099 , n4153 , n4154 , n33102 , 
 n4156 , n4157 , n33105 , n33106 , n4160 , n4161 , n33109 , n33110 , n4164 , n33112 , 
 n33113 , n4170 , n33115 , n33116 , n4173 , n33118 , n33119 , n33120 , n4180 , n33122 , 
 n33123 , n33124 , n4184 , n33126 , n33127 , n33128 , n33129 , n33130 , n4190 , n33132 , 
 n4192 , n4193 , n33135 , n33136 , n4196 , n4197 , n33139 , n33140 , n4200 , n33142 , 
 n33143 , n4203 , n33145 , n33146 , n4206 , n33148 , n33149 , n33150 , n4210 , n33152 , 
 n33153 , n4213 , n4214 , n33156 , n4216 , n4217 , n4218 , n4219 , n4220 , n33162 , 
 n4222 , n4223 , n4224 , n4225 , n33167 , n4227 , n4228 , n4229 , n33171 , n33172 , 
 n4232 , n33174 , n33175 , n4235 , n33177 , n33178 , n33179 , n4239 , n4240 , n4241 , 
 n4242 , n4243 , n4244 , n33186 , n4249 , n33188 , n33189 , n4252 , n4253 , n4254 , 
 n33193 , n4259 , n4260 , n33196 , n33197 , n33198 , n33199 , n4265 , n33201 , n4267 , 
 n4268 , n4269 , n4270 , n4271 , n4272 , n33208 , n4274 , n4275 , n4276 , n33212 , 
 n4278 , n33214 , n4280 , n4281 , n4282 , n4283 , n4284 , n33220 , n4286 , n33222 , 
 n33223 , n4289 , n33225 , n33226 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , 
 n33233 , n4299 , n4300 , n33236 , n4302 , n33238 , n4304 , n4305 , n33241 , n33242 , 
 n4308 , n33244 , n33245 , n4311 , n33247 , n33248 , n4314 , n4315 , n4316 , n33252 , 
 n33253 , n4319 , n33255 , n4321 , n33257 , n4323 , n4324 , n33260 , n33261 , n4327 , 
 n33263 , n33264 , n33265 , n33266 , n33267 , n4333 , n33269 , n4335 , n33271 , n33272 , 
 n4341 , n33274 , n33275 , n4344 , n33277 , n33278 , n4347 , n4348 , n33281 , n33282 , 
 n4354 , n33284 , n4356 , n33286 , n4358 , n4359 , n33289 , n33290 , n33291 , n4363 , 
 n33293 , n33294 , n4366 , n33296 , n33297 , n4369 , n33299 , n33300 , n4372 , n4373 , 
 n4374 , n33304 , n33305 , n4377 , n33307 , n33308 , n4380 , n33310 , n33311 , n33312 , 
 n4384 , n4385 , n33315 , n33316 , n4388 , n4389 , n4390 , n4391 , n4392 , n33322 , 
 n33323 , n4395 , n4396 , n4397 , n33327 , n33328 , n4400 , n33330 , n4402 , n33332 , 
 n4404 , n4405 , n33335 , n33336 , n33337 , n4409 , n33339 , n33340 , n33341 , n33342 , 
 n33343 , n4415 , n33345 , n33346 , n33347 , n4419 , n33349 , n4421 , n33351 , n33352 , 
 n33353 , n33354 , n4426 , n33356 , n33357 , n4429 , n33359 , n33360 , n33361 , n33362 , 
 n33363 , n4435 , n4436 , n4437 , n4438 , n4439 , n33369 , n33370 , n33371 , n33372 , 
 n33373 , n33374 , n4449 , n4450 , n33377 , n4452 , n33379 , n33380 , n33381 , n33382 , 
 n33383 , n33384 , n4462 , n4463 , n4464 , n4465 , n4466 , n33390 , n4468 , n33392 , 
 n33393 , n4471 , n33395 , n33396 , n33397 , n4475 , n33399 , n33400 , n4478 , n33402 , 
 n33403 , n33404 , n33405 , n33406 , n4484 , n4485 , n4486 , n4487 , n33411 , n33412 , 
 n33413 , n4491 , n33415 , n33416 , n4494 , n33418 , n4496 , n33420 , n4498 , n33422 , 
 n33423 , n4501 , n33425 , n33426 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , 
 n4510 , n4511 , n4512 , n33436 , n4514 , n33438 , n33439 , n4517 , n4518 , n4519 , 
 n33443 , n33444 , n33445 , n4523 , n33447 , n33448 , n4526 , n33450 , n33451 , n4529 , 
 n33453 , n33454 , n4532 , n33456 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , 
 n4540 , n4541 , n4542 , n4543 , n4544 , n33468 , n33469 , n33470 , n33471 , n4549 , 
 n4550 , n4551 , n4552 , n4553 , n4554 , n33478 , n4559 , n33480 , n4561 , n33482 , 
 n4563 , n4564 , n4565 , n33486 , n33487 , n4571 , n4572 , n4573 , n4574 , n4575 , 
 n33493 , n4577 , n4578 , n4579 , n4580 , n4581 , n33499 , n4583 , n4584 , n4585 , 
 n33503 , n33504 , n4588 , n4589 , n4590 , n33508 , n4592 , n4593 , n4594 , n33512 , 
 n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , 
 n4606 , n33524 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , 
 n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , 
 n4626 , n33544 , n33545 , n4629 , n33547 , n4631 , n33549 , n33550 , n4634 , n33552 , 
 n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n33560 , n33561 , n33562 , 
 n33563 , n4647 , n33565 , n33566 , n33567 , n4651 , n33569 , n33570 , n33571 , n4655 , 
 n33573 , n4657 , n33575 , n4659 , n33577 , n33578 , n4662 , n33580 , n4664 , n33582 , 
 n33583 , n4667 , n33585 , n33586 , n33587 , n33588 , n33589 , n4673 , n33591 , n4675 , 
 n33593 , n33594 , n4681 , n33596 , n33597 , n4684 , n33599 , n4689 , n4690 , n4691 , 
 n33603 , n33604 , n4694 , n33606 , n33607 , n33608 , n4698 , n33610 , n4700 , n4701 , 
 n33613 , n4703 , n33615 , n4705 , n33617 , n33618 , n4708 , n33620 , n33621 , n33622 , 
 n33623 , n4713 , n33625 , n4715 , n4716 , n4717 , n4718 , n4719 , n33631 , n4721 , 
 n33633 , n33634 , n4724 , n33636 , n33637 , n33638 , n4728 , n33640 , n4730 , n4731 , 
 n33643 , n33644 , n33645 , n4735 , n33647 , n33648 , n4738 , n33650 , n33651 , n4741 , 
 n33653 , n33654 , n4744 , n4745 , n4746 , n33658 , n4748 , n4749 , n4750 , n4751 , 
 n4752 , n33664 , n4754 , n33666 , n4756 , n33668 , n4758 , n4759 , n33671 , n4761 , 
 n33673 , n4763 , n33675 , n4765 , n4766 , n33678 , n4768 , n33680 , n33681 , n4771 , 
 n4772 , n4773 , n4774 , n33686 , n33687 , n33688 , n4778 , n33690 , n33691 , n4781 , 
 n4782 , n4783 , n4784 , n4785 , n33697 , n4787 , n33699 , n4789 , n4790 , n4791 , 
 n4792 , n4793 , n33705 , n4795 , n4796 , n33708 , n33709 , n33710 , n4800 , n4801 , 
 n4802 , n4803 , n4804 , n4805 , n33717 , n4810 , n33719 , n33720 , n4813 , n33722 , 
 n4818 , n4819 , n33725 , n4821 , n33727 , n4823 , n33729 , n33730 , n33731 , n4827 , 
 n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , 
 n4838 , n4839 , n4840 , n33746 , n4842 , n33748 , n4844 , n33750 , n4846 , n4847 , 
 n4848 , n4849 , n4850 , n4851 , n4852 , n33758 , n33759 , n4855 , n33761 , n33762 , 
 n4858 , n33764 , n33765 , n4861 , n33767 , n4863 , n4864 , n33770 , n4866 , n4867 , 
 n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n33782 , 
 n4878 , n33784 , n33785 , n33786 , n33787 , n4883 , n4884 , n33790 , n33791 , n4887 , 
 n33793 , n33794 , n33795 , n33796 , n33797 , n33798 , n4894 , n33800 , n4896 , n4897 , 
 n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , 
 n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , 
 n4918 , n33824 , n4920 , n33826 , n4922 , n4923 , n33829 , n4925 , n33831 , n4927 , 
 n4928 , n4929 , n4930 , n4931 , n33837 , n4933 , n33839 , n33840 , n33841 , n33842 , 
 n33843 , n33844 , n4940 , n33846 , n4942 , n4943 , n4944 , n33850 , n4949 , n33852 , 
 n4951 , n4952 , n33855 , n4957 , n33857 , n4959 , n4960 , n33860 , n4962 , n4963 , 
 n4964 , n4965 , n4966 , n33866 , n4968 , n4969 , n33869 , n33870 , n4972 , n33872 , 
 n33873 , n4975 , n33875 , n33876 , n33877 , n4979 , n33879 , n33880 , n4982 , n33882 , 
 n33883 , n33884 , n4986 , n33886 , n4988 , n33888 , n33889 , n4991 , n4992 , n4993 , 
 n4994 , n4995 , n33895 , n33896 , n4998 , n33898 , n33899 , n5001 , n5002 , n5003 , 
 n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , 
 n5014 , n33914 , n5016 , n5017 , n5018 , n5019 , n33919 , n33920 , n33921 , n5023 , 
 n5024 , n33924 , n5026 , n33926 , n33927 , n33928 , n5030 , n33930 , n33931 , n33932 , 
 n5034 , n33934 , n5036 , n33936 , n33937 , n5039 , n33939 , n33940 , n5042 , n33942 , 
 n33943 , n5045 , n33945 , n5047 , n33947 , n5049 , n5050 , n5051 , n5052 , n5053 , 
 n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n33962 , 
 n33963 , n5065 , n33965 , n5067 , n5068 , n5069 , n33969 , n5071 , n33971 , n33972 , 
 n5074 , n5075 , n33975 , n33976 , n5078 , n5079 , n33979 , n33980 , n5082 , n5083 , 
 n5084 , n33984 , n33985 , n33986 , n5088 , n5089 , n5090 , n5091 , n33991 , n33992 , 
 n33993 , n33994 , n33995 , n5100 , n5101 , n33998 , n5106 , n34000 , n5108 , n34002 , 
 n5110 , n34004 , n34005 , n5113 , n34007 , n34008 , n5116 , n34010 , n34011 , n5119 , 
 n34013 , n34014 , n34015 , n5123 , n5124 , n34018 , n5126 , n34020 , n34021 , n5129 , 
 n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n34029 , n5137 , n34031 , n34032 , 
 n5140 , n34034 , n34035 , n5143 , n5144 , n34038 , n5146 , n5147 , n34041 , n34042 , 
 n5150 , n5151 , n34045 , n5153 , n34047 , n5155 , n5156 , n34050 , n34051 , n5159 , 
 n34053 , n34054 , n5162 , n34056 , n34057 , n34058 , n5166 , n34060 , n34061 , n5169 , 
 n34063 , n34064 , n5172 , n34066 , n5174 , n34068 , n5176 , n5177 , n34071 , n5179 , 
 n34073 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n34081 , n5189 , 
 n34083 , n34084 , n5192 , n34086 , n34087 , n5195 , n34089 , n5197 , n34091 , n5199 , 
 n5200 , n34094 , n34095 , n5203 , n34097 , n34098 , n5206 , n34100 , n5208 , n5209 , 
 n34103 , n5211 , n34105 , n5213 , n5214 , n34108 , n5216 , n34110 , n5218 , n34112 , 
 n5220 , n34114 , n5222 , n5223 , n34117 , n5225 , n5226 , n34120 , n5228 , n34122 , 
 n34123 , n34124 , n5232 , n34126 , n34127 , n5235 , n34129 , n5237 , n5238 , n5239 , 
 n5240 , n5241 , n5242 , n5243 , n34137 , n34138 , n34139 , n34140 , n5248 , n5249 , 
 n34143 , n34144 , n5252 , n34146 , n34147 , n34148 , n34149 , n34150 , n34151 , n5265 , 
 n34153 , n5267 , n5268 , n34156 , n5270 , n34158 , n5272 , n5273 , n5274 , n34162 , 
 n34163 , n5277 , n34165 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , 
 n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , 
 n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n34189 , n5303 , n5304 , n5305 , 
 n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n34200 , n5314 , n34202 , 
 n5316 , n34204 , n34205 , n34206 , n5320 , n5321 , n5322 , n5323 , n5324 , n34212 , 
 n5326 , n34214 , n5328 , n34216 , n5330 , n34218 , n5332 , n5333 , n5334 , n5335 , 
 n5336 , n5337 , n5338 , n34226 , n34227 , n5341 , n34229 , n5343 , n5344 , n5345 , 
 n34233 , n34234 , n5348 , n34236 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , 
 n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n34249 , n34250 , n5364 , n34252 , 
 n34253 , n34254 , n5368 , n34256 , n34257 , n5371 , n5372 , n34260 , n34261 , n5375 , 
 n5376 , n34264 , n34265 , n5379 , n5380 , n5381 , n5382 , n34270 , n34271 , n5385 , 
 n5386 , n34274 , n5388 , n34276 , n34277 , n5391 , n5392 , n34280 , n5394 , n5395 , 
 n5396 , n5397 , n34285 , n5399 , n34287 , n5401 , n34289 , n5403 , n34291 , n5405 , 
 n5406 , n34294 , n34295 , n5409 , n34297 , n34298 , n5412 , n34300 , n34301 , n34302 , 
 n5416 , n34304 , n34305 , n5419 , n34307 , n34308 , n34309 , n34310 , n34311 , n5428 , 
 n5429 , n34314 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , 
 n5442 , n5443 , n34325 , n34326 , n5446 , n34328 , n5448 , n34330 , n5450 , n5451 , 
 n5452 , n5453 , n5454 , n5455 , n5456 , n34338 , n5458 , n34340 , n34341 , n34342 , 
 n5462 , n34344 , n5464 , n34346 , n5466 , n5467 , n34349 , n34350 , n5470 , n34352 , 
 n34353 , n5473 , n34355 , n34356 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , 
 n5482 , n34364 , n5484 , n34366 , n34367 , n5487 , n34369 , n5489 , n5490 , n34372 , 
 n5492 , n34374 , n5494 , n5495 , n34377 , n34378 , n5498 , n34380 , n34381 , n34382 , 
 n34383 , n34384 , n34385 , n5505 , n34387 , n34388 , n5508 , n34390 , n5510 , n34392 , 
 n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , 
 n5522 , n5523 , n34405 , n5525 , n34407 , n34408 , n5528 , n5529 , n5530 , n5531 , 
 n5532 , n34414 , n34415 , n5535 , n34417 , n5537 , n5538 , n5539 , n5540 , n5541 , 
 n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , 
 n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , 
 n5562 , n5563 , n5564 , n34446 , n34447 , n5567 , n5568 , n5569 , n5570 , n34452 , 
 n34453 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , 
 n5582 , n34464 , n34465 , n34466 , n5586 , n5587 , n34469 , n5589 , n34471 , n34472 , 
 n34473 , n5596 , n34475 , n34476 , n34477 , n5603 , n5604 , n34480 , n5606 , n5607 , 
 n34483 , n34484 , n5610 , n5611 , n34487 , n34488 , n5614 , n5615 , n5616 , n5617 , 
 n5618 , n34494 , n34495 , n5621 , n34497 , n34498 , n5624 , n5625 , n34501 , n34502 , 
 n34503 , n5629 , n34505 , n5631 , n5632 , n34508 , n5634 , n5635 , n5636 , n34512 , 
 n34513 , n5639 , n34515 , n34516 , n34517 , n5643 , n5644 , n34520 , n5646 , n5647 , 
 n34523 , n34524 , n5650 , n5651 , n34527 , n34528 , n34529 , n34530 , n5656 , n34532 , 
 n34533 , n34534 , n5660 , n34536 , n34537 , n5663 , n5664 , n34540 , n34541 , n5667 , 
 n5668 , n34544 , n5670 , n34546 , n5672 , n34548 , n5674 , n5675 , n34551 , n34552 , 
 n5678 , n5679 , n34555 , n5681 , n34557 , n34558 , n5684 , n5685 , n34561 , n34562 , 
 n34563 , n5689 , n34565 , n34566 , n5692 , n34568 , n34569 , n34570 , n34571 , n34572 , 
 n5698 , n34574 , n5700 , n34576 , n34577 , n34578 , n34579 , n5705 , n34581 , n34582 , 
 n34583 , n5709 , n34585 , n34586 , n5712 , n34588 , n34589 , n5715 , n5716 , n5717 , 
 n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n34599 , n5725 , n34601 , n5727 , 
 n5728 , n5729 , n5730 , n34606 , n5732 , n5733 , n34609 , n5735 , n34611 , n34612 , 
 n34613 , n5739 , n34615 , n5741 , n5742 , n5743 , n5744 , n34620 , n34621 , n5747 , 
 n5748 , n34624 , n34625 , n34626 , n5755 , n34628 , n34629 , n5761 , n5762 , n5763 , 
 n5764 , n5765 , n5766 , n34636 , n5768 , n5769 , n5770 , n5771 , n5772 , n34642 , 
 n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , 
 n34653 , n5785 , n5786 , n34656 , n34657 , n5789 , n5790 , n5791 , n5792 , n5793 , 
 n34663 , n5795 , n5796 , n5797 , n34667 , n5799 , n5800 , n5801 , n5802 , n5803 , 
 n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , 
 n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , 
 n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , 
 n5834 , n5835 , n5836 , n5837 , n34707 , n5839 , n5840 , n5841 , n5842 , n5843 , 
 n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n34720 , n5852 , n5853 , 
 n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , 
 n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , 
 n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , 
 n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n34762 , 
 n34763 , n34764 , n5896 , n34766 , n34767 , n5899 , n5900 , n34770 , n34771 , n5903 , 
 n34773 , n34774 , n34775 , n5907 , n34777 , n5909 , n34779 , n34780 , n34781 , n5913 , 
 n5914 , n34784 , n34785 , n34786 , n34787 , n34788 , n34789 , n34790 , n34791 , n34792 , 
 n34793 , n5928 , n34795 , n34796 , n34797 , n34798 , n5936 , n34800 , n34801 , n34802 , 
 n5940 , n34804 , n34805 , n5943 , n34807 , n5945 , n34809 , n34810 , n34811 , n5949 , 
 n34813 , n34814 , n5952 , n5953 , n34817 , n34818 , n5956 , n34820 , n34821 , n34822 , 
 n5960 , n5961 , n34825 , n5963 , n5964 , n34828 , n34829 , n5967 , n5968 , n34832 , 
 n5970 , n5971 , n34835 , n34836 , n34837 , n34838 , n5976 , n5977 , n34841 , n5979 , 
 n5980 , n34844 , n34845 , n5983 , n34847 , n34848 , n34849 , n5987 , n5988 , n5989 , 
 n5990 , n34854 , n34855 , n5993 , n5994 , n34858 , n34859 , n5997 , n34861 , n34862 , 
 n6000 , n6001 , n34865 , n34866 , n6004 , n6005 , n34869 , n34870 , n6008 , n6009 , 
 n6010 , n34874 , n34875 , n6013 , n34877 , n6015 , n6016 , n34880 , n6018 , n6019 , 
 n34883 , n34884 , n34885 , n6023 , n34887 , n34888 , n6026 , n6027 , n34891 , n34892 , 
 n6030 , n6031 , n34895 , n34896 , n6034 , n6035 , n6036 , n34900 , n34901 , n34902 , 
 n34903 , n6041 , n6042 , n34906 , n6044 , n6045 , n34909 , n34910 , n6048 , n34912 , 
 n34913 , n34914 , n6052 , n34916 , n34917 , n6055 , n6056 , n34920 , n34921 , n34922 , 
 n34923 , n6061 , n34925 , n6063 , n6064 , n6065 , n6066 , n34930 , n6068 , n6069 , 
 n34933 , n34934 , n6072 , n34936 , n34937 , n34938 , n6076 , n34940 , n34941 , n6079 , 
 n6080 , n34944 , n34945 , n34946 , n34947 , n6088 , n34949 , n6093 , n6094 , n34952 , 
 n6096 , n6097 , n34955 , n34956 , n6100 , n34958 , n6102 , n6103 , n6104 , n6105 , 
 n6106 , n6107 , n34965 , n34966 , n34967 , n34968 , n6112 , n34970 , n34971 , n34972 , 
 n6116 , n34974 , n6118 , n34976 , n6120 , n6121 , n34979 , n34980 , n6124 , n34982 , 
 n34983 , n6127 , n34985 , n34986 , n6130 , n34988 , n34989 , n6133 , n6134 , n6135 , 
 n6136 , n6137 , n34995 , n6139 , n6140 , n6141 , n34999 , n35000 , n35001 , n35002 , 
 n35003 , n6147 , n6148 , n35006 , n6150 , n6151 , n35009 , n35010 , n6154 , n35012 , 
 n35013 , n6157 , n6158 , n35016 , n35017 , n35018 , n35019 , n6163 , n35021 , n35022 , 
 n35023 , n6167 , n35025 , n6169 , n6170 , n6171 , n35029 , n6173 , n35031 , n35032 , 
 n6176 , n6177 , n35035 , n6179 , n6180 , n35038 , n35039 , n6183 , n35041 , n35042 , 
 n6186 , n35044 , n6188 , n6189 , n35047 , n35048 , n6192 , n6193 , n35051 , n35052 , 
 n6196 , n35054 , n35055 , n6199 , n35057 , n35058 , n35059 , n6203 , n35061 , n35062 , 
 n6206 , n6207 , n35065 , n35066 , n6210 , n35068 , n6212 , n35070 , n35071 , n35072 , 
 n6216 , n6217 , n35075 , n35076 , n35077 , n35078 , n35079 , n6223 , n6224 , n35082 , 
 n6226 , n6227 , n35085 , n35086 , n6230 , n35088 , n35089 , n35090 , n6234 , n6235 , 
 n35093 , n6237 , n6238 , n35096 , n35097 , n6241 , n6242 , n35100 , n35101 , n35102 , 
 n35103 , n35104 , n35105 , n35106 , n35107 , n6257 , n6258 , n35110 , n35111 , n35112 , 
 n6262 , n35114 , n35115 , n6265 , n6266 , n35118 , n6268 , n35120 , n35121 , n6271 , 
 n35123 , n35124 , n6274 , n6275 , n35127 , n6277 , n6278 , n6279 , n35131 , n6281 , 
 n35133 , n35134 , n6284 , n6285 , n6286 , n35138 , n6288 , n6289 , n6290 , n6291 , 
 n6292 , n6293 , n6294 , n6295 , n35147 , n6297 , n6298 , n6299 , n6300 , n6301 , 
 n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , 
 n35163 , n6313 , n6314 , n6315 , n6316 , n35168 , n35169 , n6319 , n6320 , n6321 , 
 n35173 , n35174 , n6324 , n35176 , n6326 , n35178 , n35179 , n6329 , n6330 , n6331 , 
 n6332 , n35184 , n35185 , n6335 , n6336 , n6337 , n35189 , n35190 , n6340 , n35192 , 
 n6342 , n35194 , n6344 , n35196 , n35197 , n6347 , n35199 , n35200 , n6350 , n6351 , 
 n35203 , n6353 , n6354 , n35206 , n35207 , n6357 , n35209 , n35210 , n6360 , n6361 , 
 n35213 , n35214 , n6364 , n6365 , n35217 , n6367 , n35219 , n35220 , n6370 , n35222 , 
 n35223 , n35224 , n6374 , n6375 , n35227 , n6377 , n6378 , n35230 , n35231 , n6381 , 
 n6382 , n35234 , n6384 , n6385 , n6386 , n6387 , n35239 , n6389 , n6390 , n35242 , 
 n35243 , n35244 , n6394 , n6395 , n35247 , n6400 , n35249 , n6402 , n6403 , n35252 , 
 n6408 , n6409 , n35255 , n35256 , n35257 , n35258 , n6414 , n35260 , n35261 , n35262 , 
 n6418 , n6419 , n35265 , n6421 , n6422 , n35268 , n35269 , n6425 , n6426 , n35272 , 
 n35273 , n35274 , n35275 , n6431 , n35277 , n35278 , n6434 , n35280 , n6436 , n35282 , 
 n35283 , n35284 , n6440 , n35286 , n6442 , n35288 , n35289 , n6445 , n35291 , n35292 , 
 n6448 , n6449 , n35295 , n35296 , n6452 , n35298 , n35299 , n6455 , n35301 , n35302 , 
 n35303 , n6459 , n35305 , n6461 , n35307 , n35308 , n35309 , n6465 , n6466 , n35312 , 
 n35313 , n6469 , n6470 , n35316 , n35317 , n6473 , n35319 , n35320 , n35321 , n35322 , 
 n6478 , n35324 , n6480 , n35326 , n35327 , n35328 , n35329 , n6485 , n35331 , n35332 , 
 n35333 , n6489 , n35335 , n6491 , n35337 , n35338 , n6494 , n35340 , n35341 , n6497 , 
 n35343 , n35344 , n6500 , n6501 , n35347 , n6503 , n6504 , n35350 , n35351 , n35352 , 
 n6508 , n6509 , n35355 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , 
 n6518 , n6519 , n6520 , n6521 , n6522 , n35368 , n6524 , n6525 , n6526 , n6527 , 
 n6528 , n35374 , n35375 , n6531 , n35377 , n35378 , n6534 , n6535 , n35381 , n6537 , 
 n35383 , n35384 , n6540 , n6541 , n35387 , n6546 , n35389 , n6548 , n6549 , n35392 , 
 n6554 , n35394 , n35395 , n6557 , n35397 , n6559 , n35399 , n35400 , n6562 , n35402 , 
 n35403 , n6565 , n6566 , n35406 , n6568 , n6569 , n35409 , n6571 , n35411 , n35412 , 
 n6574 , n35414 , n35415 , n35416 , n6578 , n6579 , n35419 , n6581 , n6582 , n35422 , 
 n35423 , n6585 , n6586 , n35426 , n35427 , n6589 , n35429 , n35430 , n6592 , n35432 , 
 n35433 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , 
 n6604 , n6605 , n6606 , n6607 , n6608 , n35448 , n6610 , n6611 , n6612 , n6613 , 
 n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n35461 , n6623 , 
 n6624 , n6625 , n6626 , n6627 , n6628 , n35468 , n6630 , n35470 , n6632 , n6633 , 
 n6634 , n6635 , n6636 , n6637 , n35477 , n35478 , n6640 , n35480 , n35481 , n6643 , 
 n6644 , n6645 , n6646 , n35486 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , 
 n6654 , n6655 , n6656 , n35496 , n35497 , n6659 , n35499 , n6661 , n35501 , n6663 , 
 n35503 , n35504 , n6666 , n6667 , n6668 , n6669 , n6670 , n35510 , n35511 , n6673 , 
 n35513 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n35521 , n35522 , 
 n6684 , n35524 , n35525 , n6690 , n35527 , n6692 , n6693 , n35530 , n6698 , n6699 , 
 n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n35540 , n6708 , n35542 , 
 n6710 , n35544 , n6712 , n35546 , n6714 , n35548 , n6716 , n6717 , n6718 , n6719 , 
 n35553 , n35554 , n6722 , n35556 , n35557 , n6725 , n6726 , n35560 , n6728 , n6729 , 
 n35563 , n6731 , n35565 , n6733 , n35567 , n35568 , n6736 , n6737 , n35571 , n35572 , 
 n6740 , n35574 , n35575 , n35576 , n35577 , n6745 , n35579 , n35580 , n6748 , n35582 , 
 n35583 , n6751 , n35585 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n35592 , 
 n6760 , n6761 , n6762 , n35596 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , 
 n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n35609 , n6777 , n6778 , n6779 , 
 n35613 , n6781 , n6782 , n35616 , n6784 , n35618 , n6786 , n35620 , n35621 , n6789 , 
 n35623 , n6791 , n6792 , n35626 , n6794 , n35628 , n6796 , n6797 , n35631 , n6799 , 
 n35633 , n6801 , n35635 , n35636 , n6804 , n35638 , n6806 , n35640 , n6808 , n35642 , 
 n35643 , n6811 , n6812 , n6813 , n6814 , n35648 , n35649 , n35650 , n6818 , n35652 , 
 n35653 , n6821 , n35655 , n35656 , n6827 , n35658 , n35659 , n6830 , n35661 , n35662 , 
 n6836 , n6837 , n6838 , n6839 , n35667 , n35668 , n6842 , n35670 , n6844 , n6845 , 
 n35673 , n35674 , n6848 , n35676 , n6850 , n35678 , n35679 , n35680 , n35681 , n6855 , 
 n35683 , n35684 , n35685 , n6859 , n35687 , n6861 , n6862 , n6863 , n6864 , n6865 , 
 n35693 , n6867 , n6868 , n6869 , n6870 , n6871 , n35699 , n6873 , n35701 , n35702 , 
 n6876 , n6877 , n6878 , n6879 , n6880 , n35708 , n35709 , n6883 , n6884 , n6885 , 
 n35713 , n35714 , n6888 , n6889 , n6890 , n6891 , n6892 , n35720 , n35721 , n6895 , 
 n35723 , n6897 , n6898 , n6899 , n6900 , n6901 , n35729 , n6903 , n6904 , n6905 , 
 n6906 , n6907 , n6908 , n6909 , n35737 , n6911 , n6912 , n35740 , n35741 , n6915 , 
 n6916 , n6917 , n6918 , n35746 , n35747 , n6921 , n35749 , n6923 , n35751 , n6925 , 
 n35753 , n35754 , n6928 , n35756 , n35757 , n6931 , n6932 , n6933 , n6934 , n6935 , 
 n6936 , n6937 , n6938 , n6939 , n35767 , n6941 , n6942 , n6943 , n6944 , n6945 , 
 n35773 , n35774 , n6948 , n6949 , n35777 , n6954 , n35779 , n6956 , n35781 , n35782 , 
 n6962 , n6963 , n35785 , n35786 , n6966 , n35788 , n35789 , n6969 , n6970 , n6971 , 
 n35793 , n6973 , n6974 , n6975 , n35797 , n6977 , n35799 , n6979 , n6980 , n6981 , 
 n6982 , n6983 , n6984 , n6985 , n35807 , n6987 , n6988 , n6989 , n35811 , n6991 , 
 n35813 , n35814 , n6994 , n6995 , n6996 , n35818 , n35819 , n35820 , n7000 , n35822 , 
 n35823 , n35824 , n7004 , n7005 , n7006 , n7007 , n7008 , n35830 , n7010 , n35832 , 
 n35833 , n35834 , n35835 , n7015 , n35837 , n35838 , n7018 , n35840 , n7020 , n35842 , 
 n7022 , n35844 , n35845 , n35846 , n35847 , n7027 , n35849 , n7029 , n7030 , n7031 , 
 n7032 , n7033 , n35855 , n35856 , n7036 , n35858 , n7038 , n7039 , n35861 , n7041 , 
 n7042 , n7043 , n7044 , n35866 , n7046 , n35868 , n35869 , n7049 , n35871 , n35872 , 
 n7052 , n35874 , n7054 , n35876 , n7056 , n7057 , n35879 , n35880 , n35881 , n7061 , 
 n35883 , n35884 , n35885 , n35886 , n35887 , n35888 , n35889 , n35890 , n7073 , n35892 , 
 n35893 , n7079 , n7080 , n7081 , n7082 , n7083 , n35899 , n35900 , n7086 , n35902 , 
 n35903 , n7089 , n7090 , n7091 , n7092 , n35908 , n35909 , n7095 , n7096 , n35912 , 
 n35913 , n7099 , n35915 , n7101 , n7102 , n7103 , n7104 , n7105 , n35921 , n7107 , 
 n35923 , n7109 , n7110 , n35926 , n35927 , n35928 , n7114 , n35930 , n35931 , n7117 , 
 n35933 , n35934 , n7120 , n35936 , n7122 , n35938 , n7124 , n35940 , n7126 , n7127 , 
 n35943 , n35944 , n35945 , n7131 , n35947 , n35948 , n7134 , n35950 , n35951 , n7137 , 
 n35953 , n7139 , n35955 , n7141 , n7142 , n7143 , n7144 , n35960 , n35961 , n7147 , 
 n7148 , n7149 , n35965 , n35966 , n7152 , n35968 , n7154 , n7155 , n35971 , n7157 , 
 n35973 , n35974 , n7160 , n35976 , n7162 , n35978 , n35979 , n35980 , n35981 , n7167 , 
 n35983 , n35984 , n35985 , n35986 , n35987 , n7173 , n35989 , n35990 , n35991 , n7180 , 
 n7181 , n35994 , n7186 , n35996 , n35997 , n7189 , n35999 , n36000 , n7192 , n36002 , 
 n7194 , n7195 , n7196 , n36006 , n7198 , n7199 , n7200 , n7201 , n36011 , n7203 , 
 n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n36022 , 
 n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , 
 n7224 , n7225 , n7226 , n7227 , n7228 , n36038 , n7230 , n36040 , n7232 , n7233 , 
 n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , 
 n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , 
 n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , 
 n7264 , n7265 , n7266 , n36076 , n36077 , n7269 , n36079 , n36080 , n7275 , n36082 , 
 n36083 , n7278 , n36085 , n7283 , n36087 , n7285 , n36089 , n7287 , n36091 , n7289 , 
 n36093 , n7291 , n36095 , n7293 , n36097 , n7295 , n7296 , n36100 , n36101 , n36102 , 
 n7300 , n36104 , n36105 , n7303 , n36107 , n36108 , n7306 , n36110 , n36111 , n7309 , 
 n36113 , n36114 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n36122 , 
 n36123 , n36124 , n7322 , n36126 , n36127 , n7325 , n36129 , n7327 , n7328 , n7329 , 
 n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n36139 , n7337 , n7338 , n7339 , 
 n7340 , n7341 , n36145 , n36146 , n7344 , n36148 , n36149 , n7347 , n7348 , n7349 , 
 n7350 , n36154 , n36155 , n7353 , n36157 , n7355 , n36159 , n7360 , n36161 , n7362 , 
 n7363 , n36164 , n36165 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , 
 n7376 , n7377 , n7378 , n36176 , n7380 , n7381 , n7382 , n36180 , n36181 , n36182 , 
 n7386 , n36184 , n36185 , n7389 , n36187 , n7391 , n36189 , n7393 , n36191 , n7395 , 
 n36193 , n7397 , n7398 , n36196 , n36197 , n36198 , n7402 , n36200 , n36201 , n7405 , 
 n36203 , n36204 , n7408 , n36206 , n36207 , n7411 , n36209 , n7413 , n7414 , n7415 , 
 n7416 , n7417 , n36215 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n36222 , 
 n7426 , n36224 , n7428 , n36226 , n7433 , n36228 , n7435 , n7436 , n36231 , n7441 , 
 n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , 
 n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n36251 , n7461 , 
 n36253 , n7463 , n36255 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , 
 n36263 , n7473 , n7474 , n7475 , n7476 , n7477 , n36269 , n7479 , n7480 , n7481 , 
 n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , 
 n36283 , n7496 , n36285 , n7498 , n7499 , n36288 , n7504 , n7505 , n36291 , n7507 , 
 n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n36301 , n7517 , 
 n36303 , n36304 , n36305 , n7521 , n36307 , n7523 , n7524 , n36310 , n7526 , n36312 , 
 n7528 , n36314 , n36315 , n7531 , n7532 , n36318 , n36319 , n7535 , n36321 , n36322 , 
 n7538 , n36324 , n7540 , n7541 , n36327 , n36328 , n7547 , n36330 , n7549 , n7550 , 
 n36333 , n7555 , n7556 , n7557 , n36337 , n7559 , n36339 , n36340 , n7562 , n36342 , 
 n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , 
 n7574 , n7575 , n36355 , n7577 , n7578 , n36358 , n7583 , n7584 , n7585 , n7586 , 
 n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n36371 , n36372 , 
 n7597 , n36374 , n7602 , n7603 , n36377 , n7605 , n36379 , n7610 , n36381 , n36382 , 
 n36383 , n36384 , n36385 , n7619 , n36387 , n36388 , n36389 , n7623 , n36391 , n36392 , 
 n7629 , n36394 , n36395 , n7632 , n36397 , n36398 , n36399 , n36400 , n7640 , n7641 , 
 n36403 , n36404 , n36405 , n36406 , n36407 , n36408 , n36409 , n36410 , n36411 , n36412 , 
 n36413 , n36414 , n36415 , n36416 , n36417 , n36418 , n36419 , n36420 , n36421 , n36422 , 
 n36423 , n36424 , n36425 , n36426 , n36427 , n36428 , n36429 , n36430 , n36431 , n36432 , 
 n36433 , n36434 , n36435 , n36436 , n36437 , n36438 , n36439 , n36440 , n36441 , n36442 , 
 n36443 , n36444 , n36445 , n36446 , n36447 , n36448 , n36449 , n36450 , n36451 , n36452 , 
 n36453 , n36454 , n36455 , n36456 , n36457 , n36458 , n36459 , n36460 , n36461 , n36462 , 
 n36463 , n36464 , n36465 , n36466 , n36467 , n36468 , n36469 , n36470 , n36471 , n36472 , 
 n36473 , n36474 , n36475 , n36476 , n36477 , n36478 , n36479 , n36480 , n36481 , n36482 , 
 n36483 , n36484 , n36485 , n36486 , n36487 , n36488 , n36489 , n36490 , n36491 , n36492 , 
 n36493 , n36494 , n36495 , n36496 , n36497 , n36498 , n36499 , n36500 , n36501 , n36502 , 
 n36503 , n36504 , n36505 , n36506 , n36507 , n36508 , n36509 , n36510 , n36511 , n36512 , 
 n36513 , n36514 , n36515 , n36516 , n36517 , n36518 , n36519 , n36520 , n36521 , n36522 , 
 n36523 , n36524 , n36525 , n36526 , n36527 , n36528 , n36529 , n36530 , n36531 , n36532 , 
 n36533 , n36534 , n36535 , n36536 , n36537 , n36538 , n36539 , n36540 , n36541 , n36542 , 
 n36543 , n36544 , n36545 , n36546 , n36547 , n36548 , n36549 , n36550 , n36551 , n36552 , 
 n36553 , n36554 , n36555 , n36556 , n36557 , n36558 , n36559 , n36560 , n36561 , n36562 , 
 n36563 , n36564 , n36565 , n36566 , n36567 , n36568 , n36569 , n36570 , n36571 , n36572 , 
 n36573 , n36574 , n36575 , n36576 , n36577 , n36578 , n36579 , n36580 , n36581 , n36582 , 
 n36583 , n36584 , n36585 , n36586 , n36587 , n36588 , n36589 , n36590 , n36591 , n36592 , 
 n36593 , n36594 , n36595 , n36596 , n36597 , n36598 , n36599 , n36600 , n36601 , n36602 , 
 n36603 , n36604 , n36605 , n36606 , n36607 , n36608 , n36609 , n36610 , n36611 , n36612 , 
 n36613 , n36614 , n36615 , n36616 , n36617 , n36618 , n36619 , n36620 , n36621 , n36622 , 
 n36623 , n36624 , n36625 , n36626 , n36627 , n36628 , n36629 , n36630 , n36631 , n36632 , 
 n36633 , n36634 , n36635 , n36636 , n36637 , n36638 , n36639 , n36640 , n36641 , n36642 , 
 n36643 , n36644 , n36645 , n36646 , n36647 , n36648 , n36649 , n36650 , n36651 , n36652 , 
 n36653 , n36654 , n36655 , n36656 , n36657 , n36658 , n36659 , n36660 , n36661 , n36662 , 
 n36663 , n36664 , n36665 , n36666 , n36667 , n36668 , n36669 , n36670 , n36671 , n36672 , 
 n36673 , n36674 , n36675 , n36676 , n36677 , n36678 , n36679 , n36680 , n36681 , n36682 , 
 n36683 , n36684 , n36685 , n36686 , n36687 , n36688 , n36689 , n36690 , n36691 , n36692 , 
 n36693 , n36694 , n36695 , n36696 , n36697 , n36698 , n36699 , n36700 , n36701 , n36702 , 
 n36703 , n36704 , n36705 , n36706 , n36707 , n36708 , n36709 , n36710 , n36711 , n36712 , 
 n36713 , n36714 , n36715 , n36716 , n36717 , n36718 , n36719 , n36720 , n36721 , n36722 , 
 n36723 , n36724 , n36725 , n36726 , n36727 , n36728 , n36729 , n36730 , n36731 , n36732 , 
 n36733 , n36734 , n36735 , n36736 , n36737 , n36738 , n36739 , n36740 , n36741 , n36742 , 
 n36743 , n36744 , n36745 , n36746 , n36747 , n36748 , n36749 , n36750 , n36751 , n36752 , 
 n36753 , n36754 , n36755 , n36756 , n36757 , n36758 , n36759 , n36760 , n36761 , n36762 , 
 n36763 , n36764 , n36765 , n36766 , n36767 , n36768 , n36769 , n36770 , n36771 , n36772 , 
 n36773 , n36774 , n36775 , n36776 , n36777 , n36778 , n36779 , n36780 , n36781 , n36782 , 
 n36783 , n36784 , n36785 , n36786 , n36787 , n36788 , n36789 , n36790 , n36791 , n36792 , 
 n36793 , n36794 , n36795 , n36796 , n36797 , n36798 , n36799 , n36800 , n36801 , n36802 , 
 n36803 , n36804 , n36805 , n36806 , n36807 , n36808 , n36809 , n36810 , n36811 , n36812 , 
 n36813 , n36814 , n36815 , n36816 , n36817 , n36818 , n36819 , n36820 , n36821 , n36822 , 
 n36823 , n36824 , n36825 , n36826 , n36827 , n36828 , n36829 , n36830 , n36831 , n36832 , 
 n36833 , n36834 , n36835 , n36836 , n36837 , n36838 , n36839 , n36840 , n36841 , n36842 , 
 n36843 , n36844 , n36845 , n36846 , n36847 , n36848 , n36849 , n36850 , n36851 , n36852 , 
 n36853 , n36854 , n36855 , n36856 , n36857 , n36858 , n36859 , n36860 , n36861 , n36862 , 
 n36863 , n36864 , n36865 , n36866 , n36867 , n36868 , n36869 , n36870 , n36871 , n36872 , 
 n36873 , n36874 , n36875 , n36876 , n36877 , n36878 , n36879 , n36880 , n36881 , n36882 , 
 n36883 , n36884 , n36885 , n36886 , n36887 , n36888 , n36889 , n36890 , n36891 , n36892 , 
 n36893 , n36894 , n36895 , n36896 , n36897 , n36898 , n36899 , n36900 , n36901 , n36902 , 
 n36903 , n36904 , n36905 , n36906 , n36907 , n36908 , n36909 , n36910 , n36911 , n36912 , 
 n36913 , n36914 , n36915 , n36916 , n36917 , n36918 , n36919 , n36920 , n36921 , n36922 , 
 n36923 , n36924 , n36925 , n36926 , n36927 , n36928 , n36929 , n36930 , n36931 , n36932 , 
 n36933 , n36934 , n36935 , n36936 , n36937 , n36938 , n36939 , n36940 , n36941 , n36942 , 
 n36943 , n36944 , n36945 , n36946 , n36947 , n36948 , n36949 , n36950 , n36951 , n36952 , 
 n36953 , n36954 , n36955 , n36956 , n36957 , n36958 , n36959 , n36960 , n36961 , n36962 , 
 n36963 , n36964 , n36965 , n36966 , n36967 , n36968 , n36969 , n36970 , n36971 , n36972 , 
 n36973 , n36974 , n36975 , n36976 , n36977 , n36978 , n36979 , n36980 , n36981 , n36982 , 
 n36983 , n36984 , n36985 , n36986 , n36987 , n36988 , n36989 , n36990 , n36991 , n36992 , 
 n36993 , n36994 , n36995 , n36996 , n36997 , n36998 , n36999 , n37000 , n37001 , n37002 , 
 n37003 , n37004 , n37005 , n37006 , n37007 , n37008 , n37009 , n37010 , n37011 , n37012 , 
 n37013 , n37014 , n37015 , n37016 , n37017 , n37018 , n37019 , n37020 , n37021 , n37022 , 
 n37023 , n37024 , n37025 , n37026 , n37027 , n37028 , n37029 , n37030 , n37031 , n37032 , 
 n37033 , n37034 , n37035 , n37036 , n37037 , n37038 , n37039 , n37040 , n37041 , n37042 , 
 n37043 , n37044 , n37045 , n37046 , n37047 , n37048 , n37049 , n37050 , n37051 , n37052 , 
 n37053 , n37054 , n37055 , n37056 , n37057 , n37058 , n37059 , n37060 , n37061 , n37062 , 
 n37063 , n37064 , n37065 , n37066 , n37067 , n37068 , n37069 , n37070 , n37071 , n37072 , 
 n37073 , n37074 , n37075 , n37076 , n37077 , n37078 , n37079 , n37080 , n37081 , n37082 , 
 n37083 , n37084 , n37085 , n37086 , n37087 , n37088 , n37089 , n37090 , n37091 , n37092 , 
 n37093 , n37094 , n37095 , n37096 , n37097 , n37098 , n37099 , n37100 , n37101 , n37102 , 
 n37103 , n37104 , n37105 , n37106 , n37107 , n37108 , n37109 , n37110 , n37111 , n37112 , 
 n37113 , n37114 , n37115 , n37116 , n37117 , n37118 , n37119 , n37120 , n37121 , n37122 , 
 n37123 , n37124 , n37125 , n37126 , n37127 , n37128 , n37129 , n37130 , n37131 , n37132 , 
 n37133 , n37134 , n37135 , n37136 , n37137 , n37138 , n37139 , n37140 , n37141 , n37142 , 
 n37143 , n37144 , n37145 , n37146 , n37147 , n37148 , n37149 , n37150 , n37151 , n37152 , 
 n37153 , n37154 , n37155 , n37156 , n37157 , n37158 , n37159 , n37160 , n37161 , n37162 , 
 n37163 , n37164 , n37165 , n37166 , n37167 , n37168 , n37169 , n37170 , n37171 , n37172 , 
 n37173 , n37174 , n37175 , n37176 , n37177 , n37178 , n37179 , n37180 , n37181 , n37182 , 
 n37183 , n37184 , n37185 , n37186 , n37187 , n37188 , n37189 , n37190 , n37191 , n37192 , 
 n37193 , n37194 , n37195 , n37196 , n37197 , n37198 , n37199 , n37200 , n37201 , n37202 , 
 n37203 , n37204 , n37205 , n37206 , n37207 , n37208 , n37209 , n37210 , n37211 , n37212 , 
 n37213 , n37214 , n37215 , n37216 , n37217 , n37218 , n37219 , n37220 , n37221 , n37222 , 
 n37223 , n37224 , n37225 , n37226 , n37227 , n37228 , n37229 , n37230 , n37231 , n37232 , 
 n37233 , n37234 , n37235 , n37236 , n37237 , n37238 , n37239 , n37240 , n37241 , n37242 , 
 n37243 , n37244 , n37245 , n37246 , n37247 , n37248 , n37249 , n37250 , n37251 , n37252 , 
 n37253 , n37254 , n37255 , n37256 , n37257 , n37258 , n37259 , n37260 , n37261 , n37262 , 
 n37263 , n37264 , n37265 , n37266 , n37267 , n37268 , n37269 , n37270 , n37271 , n37272 , 
 n37273 , n37274 , n37275 , n37276 , n37277 , n37278 , n37279 , n37280 , n37281 , n37282 , 
 n37283 , n37284 , n37285 , n37286 , n37287 , n37288 , n37289 , n37290 , n37291 , n37292 , 
 n37293 , n37294 , n37295 , n37296 , n37297 , n37298 , n37299 , n37300 , n37301 , n37302 , 
 n37303 , n37304 , n37305 , n37306 , n37307 , n37308 , n37309 , n37310 , n37311 , n37312 , 
 n37313 , n37314 , n37315 , n37316 , n37317 , n37318 , n37319 , n37320 , n37321 , n37322 , 
 n37323 , n37324 , n37325 , n37326 , n37327 , n37328 , n37329 , n37330 , n37331 , n37332 , 
 n37333 , n37334 , n37335 , n37336 , n37337 , n37338 , n37339 , n37340 , n37341 , n37342 , 
 n37343 , n37344 , n37345 , n37346 , n37347 , n37348 , n37349 , n37350 , n37351 , n37352 , 
 n37353 , n37354 , n37355 , n37356 , n37357 , n37358 , n37359 , n37360 , n37361 , n37362 , 
 n37363 , n37364 , n37365 , n37366 , n37367 , n37368 , n37369 , n37370 , n37371 , n37372 , 
 n37373 , n37374 , n37375 , n37376 , n37377 , n37378 , n37379 , n37380 , n37381 , n37382 , 
 n37383 , n37384 , n37385 , n37386 , n37387 , n37388 , n37389 , n37390 , n37391 , n37392 , 
 n37393 , n37394 , n37395 , n37396 , n37397 , n37398 , n37399 , n37400 , n37401 , n37402 , 
 n37403 , n37404 , n37405 , n37406 , n37407 , n37408 , n37409 , n37410 , n37411 , n37412 , 
 n37413 , n37414 , n37415 , n37416 , n37417 , n37418 , n37419 , n37420 , n37421 , n37422 , 
 n37423 , n37424 , n37425 , n37426 , n37427 , n37428 , n37429 , n37430 , n37431 , n37432 , 
 n37433 , n37434 , n37435 , n37436 , n37437 , n37438 , n37439 , n37440 , n37441 , n37442 , 
 n37443 , n37444 , n37445 , n37446 , n37447 , n37448 , n37449 , n37450 , n37451 , n37452 , 
 n37453 , n37454 , n37455 , n37456 , n37457 , n37458 , n37459 , n37460 , n37461 , n37462 , 
 n37463 , n37464 , n37465 , n37466 , n37467 , n37468 , n37469 , n37470 , n37471 , n37472 , 
 n37473 , n37474 , n37475 , n37476 , n37477 , n37478 , n37479 , n37480 , n37481 , n37482 , 
 n37483 , n37484 , n37485 , n37486 , n37487 , n37488 , n37489 , n37490 , n37491 , n37492 , 
 n37493 , n37494 , n37495 , n37496 , n37497 , n37498 , n37499 , n37500 , n37501 , n37502 , 
 n37503 , n37504 , n37505 , n37506 , n37507 , n37508 , n37509 , n37510 , n37511 , n37512 , 
 n37513 , n37514 , n37515 , n37516 , n37517 , n37518 , n37519 , n37520 , n37521 , n37522 , 
 n37523 , n37524 , n37525 , n37526 , n37527 , n37528 , n37529 , n37530 , n37531 , n37532 , 
 n37533 , n37534 , n37535 , n37536 , n37537 , n37538 , n37539 , n37540 , n37541 , n37542 , 
 n37543 , n37544 , n37545 , n37546 , n37547 , n37548 , n37549 , n37550 , n37551 , n37552 , 
 n37553 , n37554 , n37555 , n37556 , n37557 , n37558 , n37559 , n37560 , n37561 , n37562 , 
 n37563 , n37564 , n37565 , n37566 , n37567 , n37568 , n37569 , n37570 , n37571 , n37572 , 
 n37573 , n37574 , n37575 , n37576 , n37577 , n37578 , n37579 , n37580 , n37581 , n37582 , 
 n37583 , n37584 , n37585 , n37586 , n37587 , n37588 , n37589 , n37590 , n37591 , n37592 , 
 n37593 , n37594 , n37595 , n37596 , n37597 , n37598 , n37599 , n37600 , n37601 , n37602 , 
 n37603 , n37604 , n37605 , n37606 , n37607 , n37608 , n37609 , n37610 , n37611 , n37612 , 
 n37613 , n37614 , n37615 , n37616 , n37617 , n37618 , n37619 , n37620 , n37621 , n37622 , 
 n37623 , n37624 , n37625 , n37626 , n37627 , n37628 , n37629 , n37630 , n37631 , n37632 , 
 n37633 , n37634 , n37635 , n37636 , n37637 , n37638 , n37639 , n37640 , n37641 , n37642 , 
 n37643 , n37644 , n37645 , n37646 , n37647 , n37648 , n37649 , n37650 , n37651 , n37652 , 
 n37653 , n37654 , n37655 , n37656 , n37657 , n37658 , n37659 , n37660 , n37661 , n37662 , 
 n37663 , n37664 , n37665 , n37666 , n37667 , n37668 , n37669 , n37670 , n37671 , n37672 , 
 n37673 , n37674 , n37675 , n37676 , n37677 , n37678 , n37679 , n37680 , n37681 , n37682 , 
 n37683 , n37684 , n37685 , n37686 , n37687 , n37688 , n37689 , n37690 , n37691 , n37692 , 
 n37693 , n37694 , n37695 , n37696 , n37697 , n37698 , n37699 , n37700 , n37701 , n37702 , 
 n37703 , n37704 , n37705 , n37706 , n37707 , n37708 , n37709 , n37710 , n37711 , n37712 , 
 n37713 , n37714 , n37715 , n37716 , n37717 , n37718 , n37719 , n37720 , n37721 , n37722 , 
 n37723 , n37724 , n37725 , n37726 , n37727 , n37728 , n37729 , n37730 , n37731 , n37732 , 
 n37733 , n37734 , n37735 , n37736 , n37737 , n37738 , n37739 , n37740 , n37741 , n37742 , 
 n37743 , n37744 , n37745 , n37746 , n37747 , n37748 , n37749 , n37750 , n37751 , n37752 , 
 n37753 , n37754 , n37755 , n37756 , n37757 , n37758 , n37759 , n37760 , n37761 , n37762 , 
 n37763 , n37764 , n37765 , n37766 , n37767 , n37768 , n37769 , n37770 , n37771 , n37772 , 
 n37773 , n37774 , n37775 , n37776 , n37777 , n37778 , n37779 , n37780 , n37781 , n37782 , 
 n37783 , n37784 , n37785 , n37786 , n37787 , n37788 , n37789 , n37790 , n37791 , n37792 , 
 n37793 , n37794 , n37795 , n37796 , n37797 , n37798 , n37799 , n37800 , n37801 , n37802 , 
 n37803 , n37804 , n37805 , n37806 , n37807 , n37808 , n37809 , n37810 , n37811 , n37812 , 
 n37813 , n37814 , n37815 , n37816 , n37817 , n37818 , n37819 , n37820 , n37821 , n37822 , 
 n37823 , n37824 , n37825 , n37826 , n37827 , n37828 , n37829 , n37830 , n37831 , n37832 , 
 n37833 , n37834 , n37835 , n37836 , n37837 , n37838 , n37839 , n37840 , n37841 , n37842 , 
 n37843 , n37844 , n37845 , n37846 , n37847 , n37848 , n37849 , n37850 , n37851 , n37852 , 
 n37853 , n37854 , n37855 , n37856 , n37857 , n37858 , n37859 , n37860 , n37861 , n37862 , 
 n37863 , n37864 , n37865 , n37866 , n37867 , n37868 , n37869 , n37870 , n37871 , n37872 , 
 n37873 , n37874 , n37875 , n37876 , n37877 , n37878 , n37879 , n37880 , n37881 , n37882 , 
 n37883 , n37884 , n37885 , n37886 , n37887 , n37888 , n37889 , n37890 , n37891 , n37892 , 
 n37893 , n37894 , n37895 , n37896 , n37897 , n37898 , n37899 , n37900 , n37901 , n37902 , 
 n37903 , n37904 , n37905 , n37906 , n37907 , n37908 , n37909 , n37910 , n37911 , n37912 , 
 n37913 , n37914 , n37915 , n37916 , n37917 , n37918 , n37919 , n37920 , n37921 , n37922 , 
 n37923 , n37924 , n37925 , n37926 , n37927 , n37928 , n37929 , n37930 , n37931 , n37932 , 
 n37933 , n37934 , n37935 , n37936 , n37937 , n37938 , n37939 , n37940 , n37941 , n37942 , 
 n37943 , n37944 , n37945 , n37946 , n37947 , n37948 , n37949 , n37950 , n37951 , n37952 , 
 n37953 , n37954 , n37955 , n37956 , n37957 , n37958 , n37959 , n37960 , n37961 , n37962 , 
 n37963 , n37964 , n37965 , n37966 , n37967 , n37968 , n37969 , n37970 , n37971 , n37972 , 
 n37973 , n37974 , n37975 , n37976 , n37977 , n37978 , n37979 , n37980 , n37981 , n37982 , 
 n37983 , n37984 , n37985 , n37986 , n37987 , n37988 , n37989 , n37990 , n37991 , n37992 , 
 n37993 , n37994 , n37995 , n37996 , n37997 , n37998 , n37999 , n38000 , n38001 , n38002 , 
 n38003 , n38004 , n38005 , n38006 , n38007 , n38008 , n38009 , n38010 , n38011 , n38012 , 
 n38013 , n38014 , n38015 , n38016 , n38017 , n38018 , n38019 , n38020 , n38021 , n38022 , 
 n38023 , n38024 , n38025 , n38026 , n38027 , n38028 , n38029 , n38030 , n38031 , n38032 , 
 n38033 , n38034 , n38035 , n38036 , n38037 , n38038 , n38039 , n38040 , n38041 , n38042 , 
 n38043 , n38044 , n38045 , n38046 , n38047 , n38048 , n38049 , n38050 , n38051 , n38052 , 
 n38053 , n38054 , n38055 , n38056 , n38057 , n38058 , n38059 , n38060 , n38061 , n38062 , 
 n38063 , n38064 , n38065 , n38066 , n38067 , n38068 , n38069 , n38070 , n38071 , n38072 , 
 n38073 , n38074 , n38075 , n38076 , n38077 , n38078 , n38079 , n38080 , n38081 , n38082 , 
 n38083 , n38084 , n38085 , n38086 , n38087 , n38088 , n38089 , n38090 , n38091 , n38092 , 
 n38093 , n38094 , n38095 , n38096 , n38097 , n38098 , n38099 , n38100 , n38101 , n38102 , 
 n38103 , n38104 , n38105 , n38106 , n38107 , n38108 , n38109 , n38110 , n38111 , n38112 , 
 n38113 , n38114 , n38115 , n38116 , n38117 , n38118 , n38119 , n38120 , n38121 , n38122 , 
 n38123 , n38124 , n38125 , n38126 , n38127 , n38128 , n38129 , n38130 , n38131 , n38132 , 
 n38133 , n38134 , n38135 , n38136 , n38137 , n38138 , n38139 , n38140 , n38141 , n38142 , 
 n38143 , n38144 , n38145 , n38146 , n38147 , n38148 , n38149 , n38150 , n38151 , n38152 , 
 n38153 , n38154 , n38155 , n38156 , n38157 , n38158 , n38159 , n38160 , n38161 , n38162 , 
 n38163 , n38164 , n38165 , n38166 , n38167 , n38168 , n38169 , n38170 , n38171 , n38172 , 
 n38173 , n38174 , n38175 , n38176 , n38177 , n38178 , n38179 , n38180 , n38181 , n38182 , 
 n38183 , n38184 , n38185 , n38186 , n38187 , n38188 , n38189 , n38190 , n38191 , n38192 , 
 n38193 , n38194 , n38195 , n38196 , n38197 , n38198 , n38199 , n38200 , n38201 , n38202 , 
 n38203 , n38204 , n38205 , n38206 , n38207 , n38208 , n38209 , n38210 , n38211 , n38212 , 
 n38213 , n38214 , n38215 , n38216 , n38217 , n38218 , n38219 , n38220 , n38221 , n38222 , 
 n38223 , n38224 , n38225 , n38226 , n38227 , n38228 , n38229 , n38230 , n38231 , n38232 , 
 n38233 , n38234 , n38235 , n38236 , n38237 , n38238 , n38239 , n38240 , n38241 , n38242 , 
 n38243 , n38244 , n38245 , n38246 , n38247 , n38248 , n38249 , n38250 , n38251 , n38252 , 
 n38253 , n38254 , n38255 , n38256 , n38257 , n38258 , n38259 , n38260 , n38261 , n38262 , 
 n38263 , n38264 , n38265 , n38266 , n38267 , n38268 , n38269 , n38270 , n38271 , n38272 , 
 n38273 , n38274 , n38275 , n38276 , n38277 , n38278 , n38279 , n38280 , n38281 , n38282 , 
 n38283 , n38284 , n38285 , n38286 , n38287 , n38288 , n38289 , n38290 , n38291 , n38292 , 
 n38293 , n38294 , n38295 , n38296 , n38297 , n38298 , n38299 , n38300 , n38301 , n38302 , 
 n38303 , n38304 , n38305 , n38306 , n38307 , n38308 , n38309 , n38310 , n38311 , n38312 , 
 n38313 , n38314 , n38315 , n38316 , n38317 , n38318 , n38319 , n38320 , n38321 , n38322 , 
 n38323 , n38324 , n38325 , n38326 , n38327 , n38328 , n38329 , n38330 , n38331 , n38332 , 
 n38333 , n38334 , n38335 , n38336 , n38337 , n38338 , n38339 , n38340 , n38341 , n38342 , 
 n38343 , n38344 , n38345 , n38346 , n38347 , n38348 , n38349 , n38350 , n38351 , n38352 , 
 n38353 , n38354 , n38355 , n38356 , n38357 , n38358 , n38359 , n38360 , n38361 , n38362 , 
 n38363 , n38364 , n38365 , n38366 , n38367 , n38368 , n38369 , n38370 , n38371 , n38372 , 
 n38373 , n38374 , n38375 , n38376 , n38377 , n38378 , n38379 , n38380 , n38381 , n38382 , 
 n38383 , n38384 , n38385 , n38386 , n38387 , n38388 , n38389 , n38390 , n38391 , n38392 , 
 n38393 , n38394 , n38395 , n38396 , n38397 , n38398 , n38399 , n38400 , n38401 , n38402 , 
 n38403 , n38404 , n38405 , n38406 , n38407 , n38408 , n38409 , n38410 , n38411 , n38412 , 
 n38413 , n38414 , n38415 , n38416 , n38417 , n38418 , n38419 , n38420 , n38421 , n38422 , 
 n38423 , n38424 , n38425 , n38426 , n38427 , n38428 , n38429 , n38430 , n38431 , n38432 , 
 n38433 , n38434 , n38435 , n38436 , n38437 , n38438 , n38439 , n38440 , n38441 , n38442 , 
 n38443 , n38444 , n38445 , n38446 , n38447 , n38448 , n38449 , n38450 , n38451 , n38452 , 
 n38453 , n38454 , n38455 , n38456 , n38457 , n38458 , n38459 , n38460 , n38461 , n38462 , 
 n38463 , n38464 , n38465 , n38466 , n38467 , n38468 , n38469 , n38470 , n38471 , n38472 , 
 n38473 , n38474 , n38475 , n38476 , n38477 , n38478 , n38479 , n38480 , n38481 , n38482 , 
 n38483 , n38484 , n38485 , n38486 , n38487 , n38488 , n38489 , n38490 , n38491 , n38492 , 
 n38493 , n38494 , n38495 , n38496 , n38497 , n38498 , n38499 , n38500 , n38501 , n38502 , 
 n38503 , n38504 , n38505 , n38506 , n38507 , n38508 , n38509 , n38510 , n38511 , n38512 , 
 n38513 , n38514 , n38515 , n38516 , n38517 , n38518 , n38519 , n38520 , n38521 , n38522 , 
 n38523 , n38524 , n38525 , n38526 , n38527 , n38528 , n38529 , n38530 , n38531 , n38532 , 
 n38533 , n38534 , n38535 , n38536 , n38537 , n38538 , n38539 , n38540 , n38541 , n38542 , 
 n38543 , n38544 , n38545 , n38546 , n38547 , n38548 , n38549 , n38550 , n38551 , n38552 , 
 n38553 , n38554 , n38555 , n38556 , n38557 , n38558 , n38559 , n38560 , n38561 , n38562 , 
 n38563 , n38564 , n38565 , n38566 , n38567 , n38568 , n38569 , n38570 , n38571 , n38572 , 
 n38573 , n38574 , n38575 , n38576 , n38577 , n38578 , n38579 , n38580 , n38581 , n38582 , 
 n38583 , n38584 , n38585 , n38586 , n38587 , n38588 , n38589 , n38590 , n38591 , n38592 , 
 n38593 , n38594 , n38595 , n38596 , n38597 , n38598 , n38599 , n38600 , n38601 , n38602 , 
 n38603 , n38604 , n38605 , n38606 , n38607 , n38608 , n38609 , n38610 , n38611 , n38612 , 
 n38613 , n38614 , n38615 , n38616 , n38617 , n38618 , n38619 , n38620 , n38621 , n38622 , 
 n38623 , n38624 , n38625 , n38626 , n38627 , n38628 , n38629 , n38630 , n38631 , n38632 , 
 n38633 , n38634 , n38635 , n38636 , n38637 , n38638 , n38639 , n38640 , n38641 , n38642 , 
 n38643 , n38644 , n38645 , n38646 , n38647 , n38648 , n38649 , n38650 , n38651 , n38652 , 
 n38653 , n38654 , n38655 , n38656 , n38657 , n38658 , n38659 , n38660 , n38661 , n38662 , 
 n38663 , n38664 , n38665 , n38666 , n38667 , n38668 , n38669 , n38670 , n38671 , n38672 , 
 n38673 , n38674 , n38675 , n38676 , n38677 , n38678 , n38679 , n38680 , n38681 , n38682 , 
 n38683 , n38684 , n38685 , n38686 , n38687 , n38688 , n38689 , n38690 , n38691 , n38692 , 
 n38693 , n38694 , n38695 , n38696 , n38697 , n38698 , n38699 , n38700 , n38701 , n38702 , 
 n38703 , n38704 , n38705 , n38706 , n38707 , n38708 , n38709 , n38710 , n38711 , n38712 , 
 n38713 , n38714 , n38715 , n38716 , n38717 , n38718 , n38719 , n38720 , n38721 , n38722 , 
 n38723 , n38724 , n38725 , n38726 , n38727 , n38728 , n38729 , n38730 , n38731 , n38732 , 
 n38733 , n38734 , n38735 , n38736 , n38737 , n38738 , n38739 , n38740 , n38741 , n38742 , 
 n38743 , n38744 , n38745 , n38746 , n38747 , n38748 , n38749 , n38750 , n38751 , n38752 , 
 n38753 , n38754 , n38755 , n38756 , n38757 , n38758 , n38759 , n38760 , n38761 , n38762 , 
 n38763 , n38764 , n38765 , n38766 , n38767 , n38768 , n38769 , n38770 , n38771 , n38772 , 
 n38773 , n38774 , n38775 , n38776 , n38777 , n38778 , n38779 , n38780 , n38781 , n38782 , 
 n38783 , n38784 , n38785 , n38786 , n38787 , n38788 , n38789 , n38790 , n38791 , n38792 , 
 n38793 , n38794 , n38795 , n38796 , n38797 , n38798 , n38799 , n38800 , n38801 , n38802 , 
 n38803 , n38804 , n38805 , n38806 , n38807 , n38808 , n38809 , n38810 , n38811 , n38812 , 
 n38813 , n38814 , n38815 , n38816 , n38817 , n38818 , n38819 , n38820 , n38821 , n38822 , 
 n38823 , n38824 , n38825 , n38826 , n38827 , n38828 , n38829 , n38830 , n38831 , n38832 , 
 n38833 , n38834 , n38835 , n38836 , n38837 , n38838 , n38839 , n38840 , n38841 , n38842 , 
 n38843 , n38844 , n38845 , n38846 , n38847 , n38848 , n38849 , n38850 , n38851 , n38852 , 
 n38853 , n38854 , n38855 , n38856 , n38857 , n38858 , n38859 , n38860 , n38861 , n38862 , 
 n38863 , n38864 , n38865 , n38866 , n38867 , n38868 , n38869 , n38870 , n38871 , n38872 , 
 n38873 , n38874 , n38875 , n38876 , n38877 , n38878 , n38879 , n38880 , n38881 , n38882 , 
 n38883 , n38884 , n38885 , n38886 , n38887 , n38888 , n38889 , n38890 , n38891 , n38892 , 
 n38893 , n38894 , n38895 , n38896 , n38897 , n38898 , n38899 , n38900 , n38901 , n38902 , 
 n38903 , n38904 , n38905 , n38906 , n38907 , n38908 , n38909 , n38910 , n38911 , n38912 , 
 n38913 , n38914 , n38915 , n38916 , n38917 , n38918 , n38919 , n38920 , n38921 , n38922 , 
 n38923 , n38924 , n38925 , n38926 , n38927 , n38928 , n38929 , n38930 , n38931 , n38932 , 
 n38933 , n38934 , n38935 , n38936 , n38937 , n38938 , n38939 , n38940 , n38941 , n38942 , 
 n38943 , n38944 , n38945 , n38946 , n38947 , n38948 , n38949 , n38950 , n38951 , n38952 , 
 n38953 , n38954 , n38955 , n38956 , n38957 , n38958 , n38959 , n38960 , n38961 , n38962 , 
 n38963 , n38964 , n38965 , n38966 , n38967 , n38968 , n38969 , n38970 , n38971 , n38972 , 
 n38973 , n38974 , n38975 , n38976 , n38977 , n38978 , n38979 , n38980 , n38981 , n38982 , 
 n38983 , n38984 , n38985 , n38986 , n38987 , n38988 , n38989 , n38990 , n38991 , n38992 , 
 n38993 , n38994 , n38995 , n38996 , n38997 , n38998 , n38999 , n39000 , n39001 , n39002 , 
 n39003 , n39004 , n39005 , n39006 , n39007 , n39008 , n39009 , n39010 , n39011 , n39012 , 
 n39013 , n39014 , n39015 , n39016 , n39017 , n39018 , n39019 , n39020 , n39021 , n39022 , 
 n39023 , n39024 , n39025 , n39026 , n39027 , n39028 , n39029 , n39030 , n39031 , n39032 , 
 n39033 , n39034 , n39035 , n39036 , n39037 , n39038 , n39039 , n39040 , n39041 , n39042 , 
 n39043 , n39044 , n39045 , n39046 , n39047 , n39048 , n39049 , n39050 , n39051 , n39052 , 
 n39053 , n39054 , n39055 , n39056 , n39057 , n39058 , n39059 , n39060 , n39061 , n39062 , 
 n39063 , n39064 , n39065 , n39066 , n39067 , n39068 , n39069 , n39070 , n39071 , n39072 , 
 n39073 , n39074 , n39075 , n39076 , n39077 , n39078 , n39079 , n39080 , n39081 , n39082 , 
 n39083 , n39084 , n39085 , n39086 , n39087 , n39088 , n39089 , n39090 , n39091 , n39092 , 
 n39093 , n39094 , n39095 , n39096 , n39097 , n39098 , n39099 , n39100 , n39101 , n39102 , 
 n39103 , n39104 , n39105 , n39106 , n39107 , n39108 , n39109 , n39110 , n39111 , n39112 , 
 n39113 , n39114 , n39115 , n39116 , n39117 , n39118 , n39119 , n39120 , n39121 , n39122 , 
 n39123 , n39124 , n39125 , n39126 , n39127 , n39128 , n39129 , n39130 , n39131 , n39132 , 
 n39133 , n39134 , n39135 , n39136 , n39137 , n39138 , n39139 , n39140 , n39141 , n39142 , 
 n39143 , n39144 , n39145 , n39146 , n39147 , n39148 , n39149 , n39150 , n39151 , n39152 , 
 n39153 , n39154 , n39155 , n39156 , n39157 , n39158 , n39159 , n39160 , n39161 , n39162 , 
 n39163 , n39164 , n39165 , n39166 , n39167 , n39168 , n39169 , n39170 , n39171 , n39172 , 
 n39173 , n39174 , n39175 , n39176 , n39177 , n39178 , n39179 , n39180 , n39181 , n39182 , 
 n39183 , n39184 , n39185 , n39186 , n39187 , n39188 , n39189 , n39190 , n39191 , n39192 , 
 n39193 , n39194 , n39195 , n39196 , n39197 , n39198 , n39199 , n39200 , n39201 , n39202 , 
 n39203 , n39204 , n39205 , n39206 , n39207 , n39208 , n39209 , n39210 , n39211 , n39212 , 
 n39213 , n39214 , n39215 , n39216 , n39217 , n39218 , n39219 , n39220 , n39221 , n39222 , 
 n39223 , n39224 , n39225 , n39226 , n39227 , n39228 , n39229 , n39230 , n39231 , n39232 , 
 n39233 , n39234 , n39235 , n39236 , n39237 , n39238 , n39239 , n39240 , n39241 , n39242 , 
 n39243 , n39244 , n39245 , n39246 , n39247 , n39248 , n39249 , n39250 , n39251 , n39252 , 
 n39253 , n39254 , n39255 , n39256 , n39257 , n39258 , n39259 , n39260 , n39261 , n39262 , 
 n39263 , n39264 , n39265 , n39266 , n39267 , n39268 , n39269 , n39270 , n39271 , n39272 , 
 n39273 , n39274 , n39275 , n39276 , n39277 , n39278 , n39279 , n39280 , n39281 , n39282 , 
 n39283 , n39284 , n39285 , n39286 , n39287 , n39288 , n39289 , n39290 , n39291 , n39292 , 
 n39293 , n39294 , n39295 , n39296 , n39297 , n39298 , n39299 , n39300 , n39301 , n39302 , 
 n39303 , n39304 , n39305 , n39306 , n39307 , n39308 , n39309 , n39310 , n39311 , n39312 , 
 n39313 , n39314 , n39315 , n39316 , n39317 , n39318 , n39319 , n39320 , n39321 , n39322 , 
 n39323 , n39324 , n39325 , n39326 , n39327 , n39328 , n39329 , n39330 , n39331 , n39332 , 
 n39333 , n39334 , n39335 , n39336 , n39337 , n39338 , n39339 , n39340 , n39341 , n39342 , 
 n39343 , n39344 , n39345 , n39346 , n39347 , n39348 , n39349 , n39350 , n39351 , n39352 , 
 n39353 , n39354 , n39355 , n39356 , n39357 , n39358 , n39359 , n39360 , n39361 , n39362 , 
 n39363 , n39364 , n39365 , n39366 , n39367 , n39368 , n39369 , n39370 , n39371 , n39372 , 
 n39373 , n39374 , n39375 , n39376 , n39377 , n39378 , n39379 , n39380 , n39381 , n39382 , 
 n39383 , n39384 , n39385 , n39386 , n39387 , n39388 , n39389 , n39390 , n39391 , n39392 , 
 n39393 , n39394 , n39395 , n39396 , n39397 , n39398 , n39399 , n39400 , n39401 , n39402 , 
 n39403 , n39404 , n39405 , n39406 , n39407 , n39408 , n39409 , n39410 , n39411 , n39412 , 
 n39413 , n39414 , n39415 , n39416 , n39417 , n39418 , n39419 , n39420 , n39421 , n39422 , 
 n39423 , n39424 , n39425 , n39426 , n39427 , n39428 , n39429 , n39430 , n39431 , n39432 , 
 n39433 , n39434 , n39435 , n39436 , n39437 , n39438 , n39439 , n39440 , n39441 , n39442 , 
 n39443 , n39444 , n39445 , n39446 , n39447 , n39448 , n39449 , n39450 , n39451 , n39452 , 
 n39453 , n39454 , n39455 , n39456 , n39457 , n39458 , n39459 , n39460 , n39461 , n39462 , 
 n39463 , n39464 , n39465 , n39466 , n39467 , n39468 , n39469 , n39470 , n39471 , n39472 , 
 n39473 , n39474 , n39475 , n39476 , n39477 , n39478 , n39479 , n39480 , n39481 , n39482 , 
 n39483 , n39484 , n39485 , n39486 , n39487 , n39488 , n39489 , n39490 , n39491 , n39492 , 
 n39493 , n39494 , n39495 , n39496 , n39497 , n39498 , n39499 , n39500 , n39501 , n39502 , 
 n39503 , n39504 , n39505 , n39506 , n39507 , n39508 , n39509 , n39510 , n39511 , n39512 , 
 n39513 , n39514 , n39515 , n39516 , n39517 , n39518 , n39519 , n39520 , n39521 , n39522 , 
 n39523 , n39524 , n39525 , n39526 , n39527 , n39528 , n39529 , n39530 , n39531 , n39532 , 
 n39533 , n39534 , n39535 , n39536 , n39537 , n39538 , n39539 , n39540 , n39541 , n39542 , 
 n39543 , n39544 , n39545 , n39546 , n39547 , n39548 , n39549 , n39550 , n39551 , n39552 , 
 n39553 , n39554 , n39555 , n39556 , n39557 , n39558 , n39559 , n39560 , n39561 , n39562 , 
 n39563 , n39564 , n39565 , n39566 , n39567 , n39568 , n39569 , n39570 , n39571 , n39572 , 
 n39573 , n39574 , n39575 , n39576 , n39577 , n39578 , n39579 , n39580 , n39581 , n39582 , 
 n39583 , n39584 , n39585 , n39586 , n39587 , n39588 , n39589 , n39590 , n39591 , n39592 , 
 n39593 , n39594 , n39595 , n39596 , n39597 , n39598 , n39599 , n39600 , n39601 , n39602 , 
 n39603 , n39604 , n39605 , n39606 , n39607 , n39608 , n39609 , n39610 , n39611 , n39612 , 
 n39613 , n39614 , n39615 , n39616 , n39617 , n39618 , n39619 , n39620 , n39621 , n39622 , 
 n39623 , n39624 , n39625 , n39626 , n39627 , n39628 , n39629 , n39630 , n39631 , n39632 , 
 n39633 , n39634 , n39635 , n39636 , n39637 , n39638 , n39639 , n39640 , n39641 , n39642 , 
 n39643 , n39644 , n39645 , n39646 , n39647 , n39648 , n39649 , n39650 , n39651 , n39652 , 
 n39653 , n39654 , n39655 , n39656 , n39657 , n39658 , n39659 , n39660 , n39661 , n39662 , 
 n39663 , n39664 , n39665 , n39666 , n39667 , n39668 , n39669 , n39670 , n39671 , n39672 , 
 n39673 , n39674 , n39675 , n39676 , n39677 , n39678 , n39679 , n39680 , n39681 , n39682 , 
 n39683 , n39684 , n39685 , n39686 , n39687 , n39688 , n39689 , n39690 , n39691 , n39692 , 
 n39693 , n39694 , n39695 , n39696 , n39697 , n39698 , n39699 , n39700 , n39701 , n39702 , 
 n39703 , n39704 , n39705 , n39706 , n39707 , n39708 , n39709 , n39710 , n39711 , n39712 , 
 n39713 , n39714 , n39715 , n39716 , n39717 , n39718 , n39719 , n39720 , n39721 , n39722 , 
 n39723 , n39724 , n39725 , n39726 , n39727 , n39728 , n39729 , n39730 , n39731 , n39732 , 
 n39733 , n39734 , n39735 , n39736 , n39737 , n39738 , n39739 , n39740 , n39741 , n39742 , 
 n39743 , n39744 , n39745 , n39746 , n39747 , n39748 , n39749 , n39750 , n39751 , n39752 , 
 n39753 , n39754 , n39755 , n39756 , n39757 , n39758 , n39759 , n39760 , n39761 , n39762 , 
 n39763 , n39764 , n39765 , n39766 , n39767 , n39768 , n39769 , n39770 , n39771 , n39772 , 
 n39773 , n39774 , n39775 , n39776 , n39777 , n39778 , n39779 , n39780 , n39781 , n39782 , 
 n39783 , n39784 , n39785 , n39786 , n39787 , n39788 , n39789 , n39790 , n39791 , n39792 , 
 n39793 , n39794 , n39795 , n39796 , n39797 , n39798 , n39799 , n39800 , n39801 , n39802 , 
 n39803 , n39804 , n39805 , n39806 , n39807 , n39808 , n39809 , n39810 , n39811 , n39812 , 
 n39813 , n39814 , n39815 , n39816 , n39817 , n39818 , n39819 , n39820 , n39821 , n39822 , 
 n39823 , n39824 , n39825 , n39826 , n39827 , n39828 , n39829 , n39830 , n39831 , n39832 , 
 n39833 , n39834 , n39835 , n39836 , n39837 , n39838 , n39839 , n39840 , n39841 , n39842 , 
 n39843 , n39844 , n39845 , n39846 , n39847 , n39848 , n39849 , n39850 , n39851 , n39852 , 
 n39853 , n39854 , n39855 , n39856 , n39857 , n39858 , n39859 , n39860 , n39861 , n39862 , 
 n39863 , n39864 , n39865 , n39866 , n39867 , n39868 , n39869 , n39870 , n39871 , n39872 , 
 n39873 , n39874 , n39875 , n39876 , n39877 , n39878 , n39879 , n39880 , n39881 , n39882 , 
 n39883 , n39884 , n39885 , n39886 , n39887 , n39888 , n39889 , n39890 , n39891 , n39892 , 
 n39893 , n39894 , n39895 , n39896 , n39897 , n39898 , n39899 , n39900 , n39901 , n39902 , 
 n39903 , n39904 , n39905 , n39906 , n39907 , n39908 , n39909 , n39910 , n39911 , n39912 , 
 n39913 , n39914 , n39915 , n39916 , n39917 , n39918 , n39919 , n39920 , n39921 , n39922 , 
 n39923 , n39924 , n39925 , n39926 , n39927 , n39928 , n39929 , n39930 , n39931 , n39932 , 
 n39933 , n39934 , n39935 , n39936 , n39937 , n39938 , n39939 , n39940 , n39941 , n39942 , 
 n39943 , n39944 , n39945 , n39946 , n39947 , n39948 , n39949 , n39950 , n39951 , n39952 , 
 n39953 , n39954 , n39955 , n39956 , n39957 , n39958 , n39959 , n39960 , n39961 , n39962 , 
 n39963 , n39964 , n39965 , n39966 , n39967 , n39968 , n39969 , n39970 , n39971 , n39972 , 
 n39973 , n39974 , n39975 , n39976 , n39977 , n39978 , n39979 , n39980 , n39981 , n39982 , 
 n39983 , n39984 , n39985 , n39986 , n39987 , n39988 , n39989 , n39990 , n39991 , n39992 , 
 n39993 , n39994 , n39995 , n39996 , n39997 , n39998 , n39999 , n40000 , n40001 , n40002 , 
 n40003 , n40004 , n40005 , n40006 , n40007 , n40008 , n40009 , n40010 , n40011 , n40012 , 
 n40013 , n40014 , n40015 , n40016 , n40017 , n40018 , n40019 , n40020 , n40021 , n40022 , 
 n40023 , n40024 , n40025 , n40026 , n40027 , n40028 , n40029 , n40030 , n40031 , n40032 , 
 n40033 , n40034 , n40035 , n40036 , n40037 , n40038 , n40039 , n40040 , n40041 , n40042 , 
 n40043 , n40044 , n40045 , n40046 , n40047 , n40048 , n40049 , n40050 , n40051 , n40052 , 
 n40053 , n40054 , n40055 , n40056 , n40057 , n40058 , n40059 , n40060 , n40061 , n40062 , 
 n40063 , n40064 , n40065 , n40066 , n40067 , n40068 , n40069 , n40070 , n40071 , n40072 , 
 n40073 , n40074 , n40075 , n40076 , n40077 , n40078 , n40079 , n40080 , n40081 , n40082 , 
 n40083 , n40084 , n40085 , n40086 , n40087 , n40088 , n40089 , n40090 , n40091 , n40092 , 
 n40093 , n40094 , n40095 , n40096 , n40097 , n40098 , n40099 , n40100 , n40101 , n40102 , 
 n40103 , n40104 , n40105 , n40106 , n40107 , n40108 , n40109 , n40110 , n40111 , n40112 , 
 n40113 , n40114 , n40115 , n40116 , n40117 , n40118 , n40119 , n40120 , n40121 , n40122 , 
 n40123 , n40124 , n40125 , n40126 , n40127 , n40128 , n40129 , n40130 , n40131 , n40132 , 
 n40133 , n40134 , n40135 , n40136 , n40137 , n40138 , n40139 , n40140 , n40141 , n40142 , 
 n40143 , n40144 , n40145 , n40146 , n40147 , n40148 , n40149 , n40150 , n40151 , n40152 , 
 n40153 , n40154 , n40155 , n40156 , n40157 , n40158 , n40159 , n40160 , n40161 , n40162 , 
 n40163 , n40164 , n40165 , n40166 , n40167 , n40168 , n40169 , n40170 , n40171 , n40172 , 
 n40173 , n40174 , n40175 , n40176 , n40177 , n40178 , n40179 , n40180 , n40181 , n40182 , 
 n40183 , n40184 , n40185 , n40186 , n40187 , n40188 , n40189 , n40190 , n40191 , n40192 , 
 n40193 , n40194 , n40195 , n40196 , n40197 , n40198 , n40199 , n40200 , n40201 , n40202 , 
 n40203 , n40204 , n40205 , n40206 , n40207 , n40208 , n40209 , n40210 , n40211 , n40212 , 
 n40213 , n40214 , n40215 , n40216 , n40217 , n40218 , n40219 , n40220 , n40221 , n40222 , 
 n40223 , n40224 , n40225 , n40226 , n40227 , n40228 , n40229 , n40230 , n40231 , n40232 , 
 n40233 , n40234 , n40235 , n40236 , n40237 , n40238 , n40239 , n40240 , n40241 , n40242 , 
 n40243 , n40244 , n40245 , n40246 , n40247 , n40248 , n40249 , n40250 , n40251 , n40252 , 
 n40253 , n40254 , n40255 , n40256 , n40257 , n40258 , n40259 , n40260 , n40261 , n40262 , 
 n40263 , n40264 , n40265 , n40266 , n40267 , n40268 , n40269 , n40270 , n40271 , n40272 , 
 n40273 , n40274 , n40275 , n40276 , n40277 , n40278 , n40279 , n40280 , n40281 , n40282 , 
 n40283 , n40284 , n40285 , n40286 , n40287 , n40288 , n40289 , n40290 , n40291 , n40292 , 
 n40293 , n40294 , n40295 , n40296 , n40297 , n40298 , n40299 , n40300 , n40301 , n40302 , 
 n40303 , n40304 , n40305 , n40306 , n40307 , n40308 , n40309 , n40310 , n40311 , n40312 , 
 n40313 , n40314 , n40315 , n40316 , n40317 , n40318 , n40319 , n40320 , n40321 , n40322 , 
 n40323 , n40324 , n40325 , n40326 , n40327 , n40328 , n40329 , n40330 , n40331 , n40332 , 
 n40333 , n40334 , n40335 , n40336 , n40337 , n40338 , n40339 , n40340 , n40341 , n40342 , 
 n40343 , n40344 , n40345 , n40346 , n40347 , n40348 , n40349 , n40350 , n40351 , n40352 , 
 n40353 , n40354 , n40355 , n40356 , n40357 , n40358 , n40359 , n40360 , n40361 , n40362 , 
 n40363 , n40364 , n40365 , n40366 , n40367 , n40368 , n40369 , n40370 , n40371 , n40372 , 
 n40373 , n40374 , n40375 , n40376 , n40377 , n40378 , n40379 , n40380 , n40381 , n40382 , 
 n40383 , n40384 , n40385 , n40386 , n40387 , n40388 , n40389 , n40390 , n40391 , n40392 , 
 n40393 , n40394 , n40395 , n40396 , n40397 , n40398 , n40399 , n40400 , n40401 , n40402 , 
 n40403 , n40404 , n40405 , n40406 , n40407 , n40408 , n40409 , n40410 , n40411 , n40412 , 
 n40413 , n40414 , n40415 , n40416 , n40417 , n40418 , n40419 , n40420 , n40421 , n40422 , 
 n40423 , n40424 , n40425 , n40426 , n40427 , n40428 , n40429 , n40430 , n40431 , n40432 , 
 n40433 , n40434 , n40435 , n40436 , n40437 , n40438 , n40439 , n40440 , n40441 , n40442 , 
 n40443 , n40444 , n40445 , n40446 , n40447 , n40448 , n40449 , n40450 , n40451 , n40452 , 
 n40453 , n40454 , n40455 , n40456 , n40457 , n40458 , n40459 , n40460 , n40461 , n40462 , 
 n40463 , n40464 , n40465 , n40466 , n40467 , n40468 , n40469 , n40470 , n40471 , n40472 , 
 n40473 , n40474 , n40475 , n40476 , n40477 , n40478 , n40479 , n40480 , n40481 , n40482 , 
 n40483 , n40484 , n40485 , n40486 , n40487 , n40488 , n40489 , n40490 , n40491 , n40492 , 
 n40493 , n40494 , n40495 , n40496 , n40497 , n40498 , n40499 , n40500 , n40501 , n40502 , 
 n40503 , n40504 , n40505 , n40506 , n40507 , n40508 , n40509 , n40510 , n40511 , n40512 , 
 n40513 , n40514 , n40515 , n40516 , n40517 , n40518 , n40519 , n40520 , n40521 , n40522 , 
 n40523 , n40524 , n40525 , n40526 , n40527 , n40528 , n40529 , n40530 , n40531 , n40532 , 
 n40533 , n40534 , n40535 , n40536 , n40537 , n40538 , n40539 , n40540 , n40541 , n40542 , 
 n40543 , n40544 , n40545 , n40546 , n40547 , n40548 , n40549 , n40550 , n40551 , n40552 , 
 n40553 , n40554 , n40555 , n40556 , n40557 , n40558 , n40559 , n40560 , n40561 , n40562 , 
 n40563 , n40564 , n40565 , n40566 , n40567 , n40568 , n40569 , n40570 , n40571 , n40572 , 
 n40573 , n40574 , n40575 , n40576 , n40577 , n40578 , n40579 , n40580 , n40581 , n40582 , 
 n40583 , n40584 , n40585 , n40586 , n40587 , n40588 , n40589 , n40590 , n40591 , n40592 , 
 n40593 , n40594 , n40595 , n40596 , n40597 , n40598 , n40599 , n40600 , n40601 , n40602 , 
 n40603 , n40604 , n40605 , n40606 , n40607 , n40608 , n40609 , n40610 , n40611 , n40612 , 
 n40613 , n40614 , n40615 , n40616 , n40617 , n40618 , n40619 , n40620 , n40621 , n40622 , 
 n40623 , n40624 , n40625 , n40626 , n40627 , n40628 , n40629 , n40630 , n40631 , n40632 , 
 n40633 , n40634 , n40635 , n40636 , n40637 , n40638 , n40639 , n40640 , n40641 , n40642 , 
 n40643 , n40644 , n40645 , n40646 , n40647 , n40648 , n40649 , n40650 , n40651 , n40652 , 
 n40653 , n40654 , n40655 , n40656 , n40657 , n40658 , n40659 , n40660 , n40661 , n40662 , 
 n40663 , n40664 , n40665 , n40666 , n40667 , n40668 , n40669 , n40670 , n40671 , n40672 , 
 n40673 , n40674 , n40675 , n40676 , n40677 , n40678 , n40679 , n40680 , n40681 , n40682 , 
 n40683 , n40684 , n40685 , n40686 , n40687 , n40688 , n40689 , n40690 , n40691 , n40692 , 
 n40693 , n40694 , n40695 , n40696 , n40697 , n40698 , n40699 , n40700 , n40701 , n40702 , 
 n40703 , n40704 , n40705 , n40706 , n40707 , n40708 , n40709 , n40710 , n40711 , n40712 , 
 n40713 , n40714 , n40715 , n40716 , n40717 , n40718 , n40719 , n40720 , n40721 , n40722 , 
 n40723 , n40724 , n40725 , n40726 , n40727 , n40728 , n40729 , n40730 , n40731 , n40732 , 
 n40733 , n40734 , n40735 , n40736 , n40737 , n40738 , n40739 , n40740 , n40741 , n40742 , 
 n40743 , n40744 , n40745 , n40746 , n40747 , n40748 , n40749 , n40750 , n40751 , n40752 , 
 n40753 , n40754 , n40755 , n40756 , n40757 , n40758 , n40759 , n40760 , n40761 , n40762 , 
 n40763 , n40764 , n40765 , n40766 , n40767 , n40768 , n40769 , n40770 , n40771 , n40772 , 
 n40773 , n40774 , n40775 , n40776 , n40777 , n40778 , n40779 , n40780 , n40781 , n40782 , 
 n40783 , n40784 , n40785 , n40786 , n40787 , n40788 , n40789 , n40790 , n40791 , n40792 , 
 n40793 , n40794 , n40795 , n40796 , n40797 , n40798 , n40799 , n40800 , n40801 , n40802 , 
 n40803 , n40804 , n40805 , n40806 , n40807 , n40808 , n40809 , n40810 , n40811 , n40812 , 
 n40813 , n40814 , n40815 , n40816 , n40817 , n40818 , n40819 , n40820 , n40821 , n40822 , 
 n40823 , n40824 , n40825 , n40826 , n40827 , n40828 , n40829 , n40830 , n40831 , n40832 , 
 n40833 , n40834 , n40835 , n40836 , n40837 , n40838 , n40839 , n40840 , n40841 , n40842 , 
 n40843 , n40844 , n40845 , n40846 , n40847 , n40848 , n40849 , n40850 , n40851 , n40852 , 
 n40853 , n40854 , n40855 , n40856 , n40857 , n40858 , n40859 , n40860 , n40861 , n40862 , 
 n40863 , n40864 , n40865 , n40866 , n40867 , n40868 , n40869 , n40870 , n40871 , n40872 , 
 n40873 , n40874 , n40875 , n40876 , n40877 , n40878 , n40879 , n40880 , n40881 , n40882 , 
 n40883 , n40884 , n40885 , n40886 , n40887 , n40888 , n40889 , n40890 , n40891 , n40892 , 
 n40893 , n40894 , n40895 , n40896 , n40897 , n40898 , n40899 , n40900 , n40901 , n40902 , 
 n40903 , n40904 , n40905 , n40906 , n40907 , n40908 , n40909 , n40910 , n40911 , n40912 , 
 n40913 , n40914 , n40915 , n40916 , n40917 , n40918 , n40919 , n40920 , n40921 , n40922 , 
 n40923 , n40924 , n40925 , n40926 , n40927 , n40928 , n40929 , n40930 , n40931 , n40932 , 
 n40933 , n40934 , n40935 , n40936 , n40937 , n40938 , n40939 , n40940 , n40941 , n40942 , 
 n40943 , n40944 , n40945 , n40946 , n40947 , n40948 , n40949 , n40950 , n40951 , n40952 , 
 n40953 , n40954 , n40955 , n40956 , n40957 , n40958 , n40959 , n40960 , n40961 , n40962 , 
 n40963 , n40964 , n40965 , n40966 , n40967 , n40968 , n40969 , n40970 , n40971 , n40972 , 
 n40973 , n40974 , n40975 , n40976 , n40977 , n40978 , n40979 , n40980 , n40981 , n40982 , 
 n40983 , n40984 , n40985 , n40986 , n40987 , n40988 , n40989 , n40990 , n40991 , n40992 , 
 n40993 , n40994 , n40995 , n40996 , n40997 , n40998 , n40999 , n41000 , n41001 , n41002 , 
 n41003 , n41004 , n41005 , n41006 , n41007 , n41008 , n41009 , n41010 , n41011 , n41012 , 
 n41013 , n41014 , n41015 , n41016 , n41017 , n41018 , n41019 , n41020 , n41021 , n41022 , 
 n41023 , n41024 , n41025 , n41026 , n41027 , n41028 , n41029 , n41030 , n41031 , n41032 , 
 n41033 , n41034 , n41035 , n41036 , n41037 , n41038 , n41039 , n41040 , n41041 , n41042 , 
 n41043 , n41044 , n41045 , n41046 , n41047 , n41048 , n41049 , n41050 , n41051 , n41052 , 
 n41053 , n41054 , n41055 , n41056 , n41057 , n41058 , n41059 , n41060 , n41061 , n41062 , 
 n41063 , n41064 , n41065 , n41066 , n41067 , n41068 , n41069 , n41070 , n41071 , n41072 , 
 n41073 , n41074 , n41075 , n41076 , n41077 , n41078 , n41079 , n41080 , n41081 , n41082 , 
 n41083 , n41084 , n41085 , n41086 , n41087 , n41088 , n41089 , n41090 , n41091 , n41092 , 
 n41093 , n41094 , n41095 , n41096 , n41097 , n41098 , n41099 , n41100 , n41101 , n41102 , 
 n41103 , n41104 , n41105 , n41106 , n41107 , n41108 , n41109 , n41110 , n41111 , n41112 , 
 n41113 , n41114 , n41115 , n41116 , n41117 , n41118 , n41119 , n41120 , n41121 , n41122 , 
 n41123 , n41124 , n41125 , n41126 , n41127 , n41128 , n41129 , n41130 , n41131 , n41132 , 
 n41133 , n41134 , n41135 , n41136 , n41137 , n41138 , n41139 , n41140 , n41141 , n41142 , 
 n41143 , n41144 , n41145 , n41146 , n41147 , n41148 , n41149 , n41150 , n41151 , n41152 , 
 n41153 , n41154 , n41155 , n41156 , n41157 , n41158 , n41159 , n41160 , n41161 , n41162 , 
 n41163 , n41164 , n41165 , n41166 , n41167 , n41168 , n41169 , n41170 , n41171 , n41172 , 
 n41173 , n41174 , n41175 , n41176 , n41177 , n41178 , n41179 , n41180 , n41181 , n41182 , 
 n41183 , n41184 , n41185 , n41186 , n41187 , n41188 , n41189 , n41190 , n41191 , n41192 , 
 n41193 , n41194 , n41195 , n41196 , n41197 , n41198 , n41199 , n41200 , n41201 , n41202 , 
 n41203 , n41204 , n41205 , n41206 , n41207 , n41208 , n41209 , n41210 , n41211 , n41212 , 
 n41213 , n41214 , n41215 , n41216 , n41217 , n41218 , n41219 , n41220 , n41221 , n41222 , 
 n41223 , n41224 , n41225 , n41226 , n41227 , n41228 , n41229 , n41230 , n41231 , n41232 , 
 n41233 , n41234 , n41235 , n41236 , n41237 , n41238 , n41239 , n41240 , n41241 , n41242 , 
 n41243 , n41244 , n41245 , n41246 , n41247 , n41248 , n41249 , n41250 , n41251 , n41252 , 
 n41253 , n41254 , n41255 , n41256 , n41257 , n41258 , n41259 , n41260 , n41261 , n41262 , 
 n41263 , n41264 , n41265 , n41266 , n41267 , n41268 , n41269 , n41270 , n41271 , n41272 , 
 n41273 , n41274 , n41275 , n41276 , n41277 , n41278 , n41279 , n41280 , n41281 , n41282 , 
 n41283 , n41284 , n41285 , n41286 , n41287 , n41288 , n41289 , n41290 , n41291 , n41292 , 
 n41293 , n41294 , n41295 , n41296 , n41297 , n41298 , n41299 , n41300 , n41301 , n41302 , 
 n41303 , n41304 , n41305 , n41306 , n41307 , n41308 , n41309 , n41310 , n41311 , n41312 , 
 n41313 , n41314 , n41315 , n41316 , n41317 , n41318 , n41319 , n41320 , n41321 , n41322 , 
 n41323 , n41324 , n41325 , n41326 , n41327 , n41328 , n41329 , n41330 , n41331 , n41332 , 
 n41333 , n41334 , n41335 , n41336 , n41337 , n41338 , n41339 , n41340 , n41341 , n41342 , 
 n41343 , n41344 , n41345 , n41346 , n41347 , n41348 , n41349 , n41350 , n41351 , n41352 , 
 n41353 , n41354 , n41355 , n41356 , n41357 , n41358 , n41359 , n41360 , n41361 , n41362 , 
 n41363 , n41364 , n41365 , n41366 , n41367 , n41368 , n41369 , n41370 , n41371 , n41372 , 
 n41373 , n41374 , n41375 , n41376 , n41377 , n41378 , n41379 , n41380 , n41381 , n41382 , 
 n41383 , n41384 , n41385 , n41386 , n41387 , n41388 , n41389 , n41390 , n41391 , n41392 , 
 n41393 , n41394 , n41395 , n41396 , n41397 , n41398 , n41399 , n41400 , n41401 , n41402 , 
 n41403 , n41404 , n41405 , n41406 , n41407 , n41408 , n41409 , n41410 , n41411 , n41412 , 
 n41413 , n41414 , n41415 , n41416 , n41417 , n41418 , n41419 , n41420 , n41421 , n41422 , 
 n41423 , n41424 , n41425 , n41426 , n41427 , n41428 , n41429 , n41430 , n41431 , n41432 , 
 n41433 , n41434 , n41435 , n41436 , n41437 , n41438 , n41439 , n41440 , n41441 , n41442 , 
 n41443 , n41444 , n41445 , n41446 , n41447 , n41448 , n41449 , n41450 , n41451 , n41452 , 
 n41453 , n41454 , n41455 , n41456 , n41457 , n41458 , n41459 , n41460 , n41461 , n41462 , 
 n41463 , n41464 , n41465 , n41466 , n41467 , n41468 , n41469 , n41470 , n41471 , n41472 , 
 n41473 , n41474 , n41475 , n41476 , n41477 , n41478 , n41479 , n41480 , n41481 , n41482 , 
 n41483 , n41484 , n41485 , n41486 , n41487 , n41488 , n41489 , n41490 , n41491 , n41492 , 
 n41493 , n41494 , n41495 , n41496 , n41497 , n41498 , n41499 , n41500 , n41501 , n41502 , 
 n41503 , n41504 , n41505 , n41506 , n41507 , n41508 , n41509 , n41510 , n41511 , n41512 , 
 n41513 , n41514 , n41515 , n41516 , n41517 , n41518 , n41519 , n41520 , n41521 , n41522 , 
 n41523 , n41524 , n41525 , n41526 , n41527 , n41528 , n41529 , n41530 , n41531 , n41532 , 
 n41533 , n41534 , n41535 , n41536 , n41537 , n41538 , n41539 , n41540 , n41541 , n41542 , 
 n41543 , n41544 , n41545 , n41546 , n41547 , n41548 , n41549 , n41550 , n41551 , n41552 , 
 n41553 , n41554 , n41555 , n41556 , n41557 , n41558 , n41559 , n41560 , n41561 , n41562 , 
 n41563 , n41564 , n41565 , n41566 , n41567 , n41568 , n41569 , n41570 , n41571 , n41572 , 
 n41573 , n41574 , n41575 , n41576 , n41577 , n41578 , n41579 , n41580 , n41581 , n41582 , 
 n41583 , n41584 , n41585 , n41586 , n41587 , n41588 , n41589 , n41590 , n41591 , n41592 , 
 n41593 , n41594 , n41595 , n41596 , n41597 , n41598 , n41599 , n41600 , n41601 , n41602 , 
 n41603 , n41604 , n41605 , n41606 , n41607 , n41608 , n41609 , n41610 , n41611 , n41612 , 
 n41613 , n41614 , n41615 , n41616 , n41617 , n41618 , n41619 , n41620 , n41621 , n41622 , 
 n41623 , n41624 , n41625 , n41626 , n41627 , n41628 , n41629 , n41630 , n41631 , n41632 , 
 n41633 , n41634 , n41635 , n41636 , n41637 , n41638 , n41639 , n41640 , n41641 , n41642 , 
 n41643 , n41644 , n41645 , n41646 , n41647 , n41648 , n41649 , n41650 , n41651 , n41652 , 
 n41653 , n41654 , n41655 , n41656 , n41657 , n41658 , n41659 , n41660 , n41661 , n41662 , 
 n41663 , n41664 , n41665 , n41666 , n41667 , n41668 , n41669 , n41670 , n41671 , n41672 , 
 n41673 , n41674 , n41675 , n41676 , n41677 , n41678 , n41679 , n41680 , n41681 , n41682 , 
 n41683 , n41684 , n41685 , n41686 , n41687 , n41688 , n41689 , n41690 , n41691 , n41692 , 
 n41693 , n41694 , n41695 , n41696 , n41697 , n41698 , n41699 , n41700 , n41701 , n41702 , 
 n41703 , n41704 , n41705 , n41706 , n41707 , n41708 , n41709 , n41710 , n41711 , n41712 , 
 n41713 , n41714 , n41715 , n41716 , n41717 , n41718 , n41719 , n41720 , n41721 , n41722 , 
 n41723 , n41724 , n41725 , n41726 , n41727 , n41728 , n41729 , n41730 , n41731 , n41732 , 
 n41733 , n41734 , n41735 , n41736 , n41737 , n41738 , n41739 , n41740 , n41741 , n41742 , 
 n41743 , n41744 , n41745 , n41746 , n41747 , n41748 , n41749 , n41750 , n41751 , n41752 , 
 n41753 , n41754 , n41755 , n41756 , n41757 , n41758 , n41759 , n41760 , n41761 , n41762 , 
 n41763 , n41764 , n41765 , n41766 , n41767 , n41768 , n41769 , n41770 , n41771 , n41772 , 
 n41773 , n41774 , n41775 , n41776 , n41777 , n41778 , n41779 , n41780 , n41781 , n41782 , 
 n41783 , n41784 , n41785 , n41786 , n41787 , n41788 , n41789 , n41790 , n41791 , n41792 , 
 n41793 , n41794 , n41795 , n41796 , n41797 , n41798 , n41799 , n41800 , n41801 , n41802 , 
 n41803 , n41804 , n41805 , n41806 , n41807 , n41808 , n41809 , n41810 , n41811 , n41812 , 
 n41813 , n41814 , n41815 , n41816 , n41817 , n41818 , n41819 , n41820 , n41821 , n41822 , 
 n41823 , n41824 , n41825 , n41826 , n41827 , n41828 , n41829 , n41830 , n41831 , n41832 , 
 n41833 , n41834 , n41835 , n41836 , n41837 , n41838 , n41839 , n41840 , n41841 , n41842 , 
 n41843 , n41844 , n41845 , n41846 , n41847 , n41848 , n41849 , n41850 , n41851 , n41852 , 
 n41853 , n41854 , n41855 , n41856 , n41857 , n41858 , n41859 , n41860 , n41861 , n41862 , 
 n41863 , n41864 , n41865 , n41866 , n41867 , n41868 , n41869 , n41870 , n41871 , n41872 , 
 n41873 , n41874 , n41875 , n41876 , n41877 , n41878 , n41879 , n41880 , n41881 , n41882 , 
 n41883 , n41884 , n41885 , n41886 , n41887 , n41888 , n41889 , n41890 , n41891 , n41892 , 
 n41893 , n41894 , n41895 , n41896 , n41897 , n41898 , n41899 , n41900 , n41901 , n41902 , 
 n41903 , n41904 , n41905 , n41906 , n41907 , n41908 , n41909 , n41910 , n41911 , n41912 , 
 n41913 , n41914 , n41915 , n41916 , n41917 , n41918 , n41919 , n41920 , n41921 , n41922 , 
 n41923 , n41924 , n41925 , n41926 , n41927 , n41928 , n41929 , n41930 , n41931 , n41932 , 
 n41933 , n41934 , n41935 , n41936 , n41937 , n41938 , n41939 , n41940 , n41941 , n41942 , 
 n41943 , n41944 , n41945 , n41946 , n41947 , n41948 , n41949 , n41950 , n41951 , n41952 , 
 n41953 , n41954 , n41955 , n41956 , n41957 , n41958 , n41959 , n41960 , n41961 , n41962 , 
 n41963 , n41964 , n41965 , n41966 , n41967 , n41968 , n41969 , n41970 , n41971 , n41972 , 
 n41973 , n41974 , n41975 , n41976 , n41977 , n41978 , n41979 , n41980 , n41981 , n41982 , 
 n41983 , n41984 , n41985 , n41986 , n41987 , n41988 , n41989 , n41990 , n41991 , n41992 , 
 n41993 , n41994 , n41995 , n41996 , n41997 , n41998 , n41999 , n42000 , n42001 , n42002 , 
 n42003 , n42004 , n42005 , n42006 , n42007 , n42008 , n42009 , n42010 , n42011 , n42012 , 
 n42013 , n42014 , n42015 , n42016 , n42017 , n42018 , n42019 , n42020 , n42021 , n42022 , 
 n42023 , n42024 , n42025 , n42026 , n42027 , n42028 , n42029 , n42030 , n42031 , n42032 , 
 n42033 , n42034 , n42035 , n42036 , n42037 , n42038 , n42039 , n42040 , n42041 , n42042 , 
 n42043 , n42044 , n42045 , n42046 , n42047 , n42048 , n42049 , n42050 , n42051 , n42052 , 
 n42053 , n42054 , n42055 , n42056 , n42057 , n42058 , n42059 , n42060 , n42061 , n42062 , 
 n42063 , n42064 , n42065 , n42066 , n42067 , n42068 , n42069 , n42070 , n42071 , n42072 , 
 n42073 , n42074 , n42075 , n42076 , n42077 , n42078 , n42079 , n42080 , n42081 , n42082 , 
 n42083 , n42084 , n42085 , n42086 , n42087 , n42088 , n42089 , n42090 , n42091 , n42092 , 
 n42093 , n42094 , n42095 , n42096 , n42097 , n42098 , n42099 , n42100 , n42101 , n42102 , 
 n42103 , n42104 , n42105 , n42106 , n42107 , n42108 , n42109 , n42110 , n42111 , n42112 , 
 n42113 , n42114 , n42115 , n42116 , n42117 , n42118 , n42119 , n42120 , n42121 , n42122 , 
 n42123 , n42124 , n42125 , n42126 , n42127 , n42128 , n42129 , n42130 , n42131 , n42132 , 
 n42133 , n42134 , n42135 , n42136 , n42137 , n42138 , n42139 , n42140 , n42141 , n42142 , 
 n42143 , n42144 , n42145 , n42146 , n42147 , n42148 , n42149 , n42150 , n42151 , n42152 , 
 n42153 , n42154 , n42155 , n42156 , n42157 , n42158 , n42159 , n42160 , n42161 , n42162 , 
 n42163 , n42164 , n42165 , n42166 , n42167 , n42168 , n42169 , n42170 , n42171 , n42172 , 
 n42173 , n42174 , n42175 , n42176 , n42177 , n42178 , n42179 , n42180 , n42181 , n42182 , 
 n42183 , n42184 , n42185 , n42186 , n42187 , n42188 , n42189 , n42190 , n42191 , n42192 , 
 n42193 , n42194 , n42195 , n42196 , n42197 , n42198 , n42199 , n42200 , n42201 , n42202 , 
 n42203 , n42204 , n42205 , n42206 , n42207 , n42208 , n42209 , n42210 , n42211 , n42212 , 
 n42213 , n42214 , n42215 , n42216 , n42217 , n42218 , n42219 , n42220 , n42221 , n42222 , 
 n42223 , n42224 , n42225 , n42226 , n42227 , n42228 , n42229 , n42230 , n42231 , n42232 , 
 n42233 , n42234 , n42235 , n42236 , n42237 , n42238 , n42239 , n42240 , n42241 , n42242 , 
 n42243 , n42244 , n42245 , n42246 , n42247 , n42248 , n42249 , n42250 , n42251 , n42252 , 
 n42253 , n42254 , n42255 , n42256 , n42257 , n42258 , n42259 , n42260 , n42261 , n42262 , 
 n42263 , n42264 , n42265 , n42266 , n42267 , n42268 , n42269 , n42270 , n42271 , n42272 , 
 n42273 , n42274 , n42275 , n42276 , n42277 , n42278 , n42279 , n42280 , n42281 , n42282 , 
 n42283 , n42284 , n42285 , n42286 , n42287 , n42288 , n42289 , n42290 , n42291 , n42292 , 
 n42293 , n42294 , n42295 , n42296 , n42297 , n42298 , n42299 , n42300 , n42301 , n42302 , 
 n42303 , n42304 , n42305 , n42306 , n42307 , n42308 , n42309 , n42310 , n42311 , n42312 , 
 n42313 , n42314 , n42315 , n42316 , n42317 , n42318 , n42319 , n42320 , n42321 , n42322 , 
 n42323 , n42324 , n42325 , n42326 , n42327 , n42328 , n42329 , n42330 , n42331 , n42332 , 
 n42333 , n42334 , n42335 , n42336 , n42337 , n42338 , n42339 , n42340 , n42341 , n42342 , 
 n42343 , n42344 , n42345 , n42346 , n42347 , n42348 , n42349 , n42350 , n42351 , n42352 , 
 n42353 , n42354 , n42355 , n42356 , n42357 , n42358 , n42359 , n42360 , n42361 , n42362 , 
 n42363 , n42364 , n42365 , n42366 , n42367 , n42368 , n42369 , n42370 , n42371 , n42372 , 
 n42373 , n42374 , n42375 , n42376 , n42377 , n42378 , n42379 , n42380 , n42381 , n42382 , 
 n42383 , n42384 , n42385 , n42386 , n42387 , n42388 , n42389 , n42390 , n42391 , n42392 , 
 n42393 , n42394 , n42395 , n42396 , n42397 , n42398 , n42399 , n42400 , n42401 , n42402 , 
 n42403 , n42404 , n42405 , n42406 , n42407 , n42408 , n42409 , n42410 , n42411 , n42412 , 
 n42413 , n42414 , n42415 , n42416 , n42417 , n42418 , n42419 , n42420 , n42421 , n42422 , 
 n42423 , n42424 , n42425 , n42426 , n42427 , n42428 , n42429 , n42430 , n42431 , n42432 , 
 n42433 , n42434 , n42435 , n42436 , n42437 , n42438 , n42439 , n42440 , n42441 , n42442 , 
 n42443 , n42444 , n42445 , n42446 , n42447 , n42448 , n42449 , n42450 , n42451 , n42452 , 
 n42453 , n42454 , n42455 , n42456 , n42457 , n42458 , n42459 , n42460 , n42461 , n42462 , 
 n42463 , n42464 , n42465 , n42466 , n42467 , n42468 , n42469 , n42470 , n42471 , n42472 , 
 n42473 , n42474 , n42475 , n42476 , n42477 , n42478 , n42479 , n42480 , n42481 , n42482 , 
 n42483 , n42484 , n42485 , n42486 , n42487 , n42488 , n42489 , n42490 , n42491 , n42492 , 
 n42493 , n42494 , n42495 , n42496 , n42497 , n42498 , n42499 , n42500 , n42501 , n42502 , 
 n42503 , n42504 , n42505 , n42506 , n42507 , n42508 , n42509 , n42510 , n42511 , n42512 , 
 n42513 , n42514 , n42515 , n42516 , n42517 , n42518 , n42519 , n42520 , n42521 , n42522 , 
 n42523 , n42524 , n42525 , n42526 , n42527 , n42528 , n42529 , n42530 , n42531 , n42532 , 
 n42533 , n42534 , n42535 , n42536 , n42537 , n42538 , n42539 , n42540 , n42541 , n42542 , 
 n42543 , n42544 , n42545 , n42546 , n42547 , n42548 , n42549 , n42550 , n42551 , n42552 , 
 n42553 , n42554 , n42555 , n42556 , n42557 , n42558 , n42559 , n42560 , n42561 , n42562 , 
 n42563 , n42564 , n42565 , n42566 , n42567 , n42568 , n42569 , n42570 , n42571 , n42572 , 
 n42573 , n42574 , n42575 , n42576 , n42577 , n42578 , n42579 , n42580 , n42581 , n42582 , 
 n42583 , n42584 , n42585 , n42586 , n42587 , n42588 , n42589 , n42590 , n42591 , n42592 , 
 n42593 , n42594 , n42595 , n42596 , n42597 , n42598 , n42599 , n42600 , n42601 , n42602 , 
 n42603 , n42604 , n42605 , n42606 , n42607 , n42608 , n42609 , n42610 , n42611 , n42612 , 
 n42613 , n42614 , n42615 , n42616 , n42617 , n42618 , n42619 , n42620 , n42621 , n42622 , 
 n42623 , n42624 , n42625 , n42626 , n42627 , n42628 , n42629 , n42630 , n42631 , n42632 , 
 n42633 , n42634 , n42635 , n42636 , n42637 , n42638 , n42639 , n42640 , n42641 , n42642 , 
 n42643 , n42644 , n42645 , n42646 , n42647 , n42648 , n42649 , n42650 , n42651 , n42652 , 
 n42653 , n42654 , n42655 , n42656 , n42657 , n42658 , n42659 , n42660 , n42661 , n42662 , 
 n42663 , n42664 , n42665 , n42666 , n42667 , n42668 , n42669 , n42670 , n42671 , n42672 , 
 n42673 , n42674 , n42675 , n42676 , n42677 , n42678 , n42679 , n42680 , n42681 , n42682 , 
 n42683 , n42684 , n42685 , n42686 , n42687 , n42688 , n42689 , n42690 , n42691 , n42692 , 
 n42693 , n42694 , n42695 , n42696 , n42697 , n42698 , n42699 , n42700 , n42701 , n42702 , 
 n42703 , n42704 , n42705 , n42706 , n42707 , n42708 , n42709 , n42710 , n42711 , n42712 , 
 n42713 , n42714 , n42715 , n42716 , n42717 , n42718 , n42719 , n42720 , n42721 , n42722 , 
 n42723 , n42724 , n42725 , n42726 , n42727 , n42728 , n42729 , n42730 , n42731 , n42732 , 
 n42733 , n42734 , n42735 , n42736 , n42737 , n42738 , n42739 , n42740 , n42741 , n42742 , 
 n42743 , n42744 , n42745 , n42746 , n42747 , n42748 , n42749 , n42750 , n42751 , n42752 , 
 n42753 , n42754 , n42755 , n42756 , n42757 , n42758 , n42759 , n42760 , n42761 , n42762 , 
 n42763 , n42764 , n42765 , n42766 , n42767 , n42768 , n42769 , n42770 , n42771 , n42772 , 
 n42773 , n42774 , n42775 , n42776 , n42777 , n42778 , n42779 , n42780 , n42781 , n42782 , 
 n42783 , n42784 , n42785 , n42786 , n42787 , n42788 , n42789 , n42790 , n42791 , n42792 , 
 n42793 , n42794 , n42795 , n42796 , n42797 , n42798 , n42799 , n42800 , n42801 , n42802 , 
 n42803 , n42804 , n42805 , n42806 , n42807 , n42808 , n42809 , n42810 , n42811 , n42812 , 
 n42813 , n42814 , n42815 , n42816 , n42817 , n42818 , n42819 , n42820 , n42821 , n42822 , 
 n42823 , n42824 , n42825 , n42826 , n42827 , n42828 , n42829 , n42830 , n42831 , n42832 , 
 n42833 , n42834 , n42835 , n42836 , n42837 , n42838 , n42839 , n42840 , n42841 , n42842 , 
 n42843 , n42844 , n42845 , n42846 , n42847 , n42848 , n42849 , n42850 , n42851 , n42852 , 
 n42853 , n42854 , n42855 , n42856 , n42857 , n42858 , n42859 , n42860 , n42861 , n42862 , 
 n42863 , n42864 , n42865 , n42866 , n42867 , n42868 , n42869 , n42870 , n42871 , n42872 , 
 n42873 , n42874 , n42875 , n42876 , n42877 , n42878 , n42879 , n42880 , n42881 , n42882 , 
 n42883 , n42884 , n42885 , n42886 , n42887 , n42888 , n42889 , n42890 , n42891 , n42892 , 
 n42893 , n42894 , n42895 , n42896 , n42897 , n42898 , n42899 , n42900 , n42901 , n42902 , 
 n42903 , n42904 , n42905 , n42906 , n42907 , n42908 , n42909 , n42910 , n42911 , n42912 , 
 n42913 , n42914 , n42915 , n42916 , n42917 , n42918 , n42919 , n42920 , n42921 , n42922 , 
 n42923 , n42924 , n42925 , n42926 , n42927 , n42928 , n42929 , n42930 , n42931 , n42932 , 
 n42933 , n42934 , n42935 , n42936 , n42937 , n42938 , n42939 , n42940 , n42941 , n42942 , 
 n42943 , n42944 , n42945 , n42946 , n42947 , n42948 , n42949 , n42950 , n42951 , n42952 , 
 n42953 , n42954 , n42955 , n42956 , n42957 , n42958 , n42959 , n42960 , n42961 , n42962 , 
 n42963 , n42964 , n42965 , n42966 , n42967 , n42968 , n42969 , n42970 , n42971 , n42972 , 
 n42973 , n42974 , n42975 , n42976 , n42977 , n42978 , n42979 , n42980 , n42981 , n42982 , 
 n42983 , n42984 , n42985 , n42986 , n42987 , n42988 , n42989 , n42990 , n42991 , n42992 , 
 n42993 , n42994 , n42995 , n42996 , n42997 , n42998 , n42999 , n43000 , n43001 , n43002 , 
 n43003 , n43004 , n43005 , n43006 , n43007 , n43008 , n43009 , n43010 , n43011 , n43012 , 
 n43013 , n43014 , n43015 , n43016 , n43017 , n43018 , n43019 , n43020 , n43021 , n43022 , 
 n43023 , n43024 , n43025 , n43026 , n43027 , n43028 , n43029 , n43030 , n43031 , n43032 , 
 n43033 , n43034 , n43035 , n43036 , n43037 , n43038 , n43039 , n43040 , n43041 , n43042 , 
 n43043 , n43044 , n43045 , n43046 , n43047 , n43048 , n43049 , n43050 , n43051 , n43052 , 
 n43053 , n43054 , n43055 , n43056 , n43057 , n43058 , n43059 , n43060 , n43061 , n43062 , 
 n43063 , n43064 , n43065 , n43066 , n43067 , n43068 , n43069 , n43070 , n43071 , n43072 , 
 n43073 , n43074 , n43075 , n43076 , n43077 , n43078 , n43079 , n43080 , n43081 , n43082 , 
 n43083 , n43084 , n43085 , n43086 , n43087 , n43088 , n43089 , n43090 , n43091 , n43092 , 
 n43093 , n43094 , n43095 , n43096 , n43097 , n43098 , n43099 , n43100 , n43101 , n43102 , 
 n43103 , n43104 , n43105 , n43106 , n43107 , n43108 , n43109 , n43110 , n43111 , n43112 , 
 n43113 , n43114 , n43115 , n43116 , n43117 , n43118 , n43119 , n43120 , n43121 , n43122 , 
 n43123 , n43124 , n43125 , n43126 , n43127 , n43128 , n43129 , n43130 , n43131 , n43132 , 
 n43133 , n43134 , n43135 , n43136 , n43137 , n43138 , n43139 , n43140 , n43141 , n43142 , 
 n43143 , n43144 , n43145 , n43146 , n43147 , n43148 , n43149 , n43150 , n43151 , n43152 , 
 n43153 , n43154 , n43155 , n43156 , n43157 , n43158 , n43159 , n43160 , n43161 , n43162 , 
 n43163 , n43164 , n43165 , n43166 , n43167 , n43168 , n43169 , n43170 , n43171 , n43172 , 
 n43173 , n43174 , n43175 , n43176 , n43177 , n43178 , n43179 , n43180 , n43181 , n43182 , 
 n43183 , n43184 , n43185 , n43186 , n43187 , n43188 , n43189 , n43190 , n43191 , n43192 , 
 n43193 , n43194 , n43195 , n43196 , n43197 , n43198 , n43199 , n43200 , n43201 , n43202 , 
 n43203 , n43204 , n43205 , n43206 , n43207 , n43208 , n43209 , n43210 , n43211 , n43212 , 
 n43213 , n43214 , n43215 , n43216 , n43217 , n43218 , n43219 , n43220 , n43221 , n43222 , 
 n43223 , n43224 , n43225 , n43226 , n43227 , n43228 , n43229 , n43230 , n43231 , n43232 , 
 n43233 , n43234 , n43235 , n43236 , n43237 , n43238 , n43239 , n43240 , n43241 , n43242 , 
 n43243 , n43244 , n43245 , n43246 , n43247 , n43248 , n43249 , n43250 , n43251 , n43252 , 
 n43253 , n43254 , n43255 , n43256 , n43257 , n43258 , n43259 , n43260 , n43261 , n43262 , 
 n43263 , n43264 , n43265 , n43266 , n43267 , n43268 , n43269 , n43270 , n43271 , n43272 , 
 n43273 , n43274 , n43275 , n43276 , n43277 , n43278 , n43279 , n43280 , n43281 , n43282 , 
 n43283 , n43284 , n43285 , n43286 , n43287 , n43288 , n43289 , n43290 , n43291 , n43292 , 
 n43293 , n43294 , n43295 , n43296 , n43297 , n43298 , n43299 , n43300 , n43301 , n43302 , 
 n43303 , n43304 , n43305 , n43306 , n43307 , n43308 , n43309 , n43310 , n43311 , n43312 , 
 n43313 , n43314 , n43315 , n43316 , n43317 , n43318 , n43319 , n43320 , n43321 , n43322 , 
 n43323 , n43324 , n43325 , n43326 , n43327 , n43328 , n43329 , n43330 , n43331 , n43332 , 
 n43333 , n43334 , n43335 , n43336 , n43337 , n43338 , n43339 , n43340 , n43341 , n43342 , 
 n43343 , n43344 , n43345 , n43346 , n43347 , n43348 , n43349 , n43350 , n43351 , n43352 , 
 n43353 , n43354 , n43355 , n43356 , n43357 , n43358 , n43359 , n43360 , n43361 , n43362 , 
 n43363 , n43364 , n43365 , n43366 , n43367 , n43368 , n43369 , n43370 , n43371 , n43372 , 
 n43373 , n43374 , n43375 , n43376 , n43377 , n43378 , n43379 , n43380 , n43381 , n43382 , 
 n43383 , n43384 , n43385 , n43386 , n43387 , n43388 , n43389 , n43390 , n43391 , n43392 , 
 n43393 , n43394 , n43395 , n43396 , n43397 , n43398 , n43399 , n43400 , n43401 , n43402 , 
 n43403 , n43404 , n43405 , n43406 , n43407 , n43408 , n43409 , n43410 , n43411 , n43412 , 
 n43413 , n43414 , n43415 , n43416 , n43417 , n43418 , n43419 , n43420 , n43421 , n43422 , 
 n43423 , n43424 , n43425 , n43426 , n43427 , n43428 , n43429 , n43430 , n43431 , n43432 , 
 n43433 , n43434 , n43435 , n43436 , n43437 , n43438 , n43439 , n43440 , n43441 , n43442 , 
 n43443 , n43444 , n43445 , n43446 , n43447 , n43448 , n43449 , n43450 , n43451 , n43452 , 
 n43453 , n43454 , n43455 , n43456 , n43457 , n43458 , n43459 , n43460 , n43461 , n43462 , 
 n43463 , n43464 , n43465 , n43466 , n43467 , n43468 , n43469 , n43470 , n43471 , n43472 , 
 n43473 , n43474 , n43475 , n43476 , n43477 , n43478 , n43479 , n43480 , n43481 , n43482 , 
 n43483 , n43484 , n43485 , n43486 , n43487 , n43488 , n43489 , n43490 , n43491 , n43492 , 
 n43493 , n43494 , n43495 , n43496 , n43497 , n43498 , n43499 , n43500 , n43501 , n43502 , 
 n43503 , n43504 , n43505 , n43506 , n43507 , n43508 , n43509 , n43510 , n43511 , n43512 , 
 n43513 , n43514 , n43515 , n43516 , n43517 , n43518 , n43519 , n43520 , n43521 , n43522 , 
 n43523 , n43524 , n43525 , n43526 , n43527 , n43528 , n43529 , n43530 , n43531 , n43532 , 
 n43533 , n43534 , n43535 , n43536 , n43537 , n43538 , n43539 , n43540 , n43541 , n43542 , 
 n43543 , n43544 , n43545 , n43546 , n43547 , n43548 , n43549 , n43550 , n43551 , n43552 , 
 n43553 , n43554 , n43555 , n43556 , n43557 , n43558 , n43559 , n43560 , n43561 , n43562 , 
 n43563 , n43564 , n43565 , n43566 , n43567 , n43568 , n43569 , n43570 , n43571 , n43572 , 
 n43573 , n43574 , n43575 , n43576 , n43577 , n43578 , n43579 , n43580 , n43581 , n43582 , 
 n43583 , n43584 , n43585 , n43586 , n43587 , n43588 , n43589 , n43590 , n43591 , n43592 , 
 n43593 , n43594 , n43595 , n43596 , n43597 , n43598 , n43599 , n43600 , n43601 , n43602 , 
 n43603 , n43604 , n43605 , n43606 , n43607 , n43608 , n43609 , n43610 , n43611 , n43612 , 
 n43613 , n43614 , n43615 , n43616 , n43617 , n43618 , n43619 , n43620 , n43621 , n43622 , 
 n43623 , n43624 , n43625 , n43626 , n43627 , n43628 , n43629 , n43630 , n43631 , n43632 , 
 n43633 , n43634 , n43635 , n43636 , n43637 , n43638 , n43639 , n43640 , n43641 , n43642 , 
 n43643 , n43644 , n43645 , n43646 , n43647 , n43648 , n43649 , n43650 , n43651 , n43652 , 
 n43653 , n43654 , n43655 , n43656 , n43657 , n43658 , n43659 , n43660 , n43661 , n43662 , 
 n43663 , n43664 , n43665 , n43666 , n43667 , n43668 , n43669 , n43670 , n43671 , n43672 , 
 n43673 , n43674 , n43675 , n43676 , n43677 , n43678 , n43679 , n43680 , n43681 , n43682 , 
 n43683 , n43684 , n43685 , n43686 , n43687 , n43688 , n43689 , n43690 , n43691 , n43692 , 
 n43693 , n43694 , n43695 , n43696 , n43697 , n43698 , n43699 , n43700 , n43701 , n43702 , 
 n43703 , n43704 , n43705 , n43706 , n43707 , n43708 , n43709 , n43710 , n43711 , n43712 , 
 n43713 , n43714 , n43715 , n43716 , n43717 , n43718 , n43719 , n43720 , n43721 , n43722 , 
 n43723 , n43724 , n43725 , n43726 , n43727 , n43728 , n43729 , n43730 , n43731 , n43732 , 
 n43733 , n43734 , n43735 , n43736 , n43737 , n43738 , n43739 , n43740 , n43741 , n43742 , 
 n43743 , n43744 , n43745 , n43746 , n43747 , n43748 , n43749 , n43750 , n43751 , n43752 , 
 n43753 , n43754 , n43755 , n43756 , n43757 , n43758 , n43759 , n43760 , n43761 , n43762 , 
 n43763 , n43764 , n43765 , n43766 , n43767 , n43768 , n43769 , n43770 , n43771 , n43772 , 
 n43773 , n43774 , n43775 , n43776 , n43777 , n43778 , n43779 , n43780 , n43781 , n43782 , 
 n43783 , n43784 , n43785 , n43786 , n43787 , n43788 , n43789 , n43790 , n43791 , n43792 , 
 n43793 , n43794 , n43795 , n43796 , n43797 , n43798 , n43799 , n43800 , n43801 , n43802 , 
 n43803 , n43804 , n43805 , n43806 , n43807 , n43808 , n43809 , n43810 , n43811 , n43812 , 
 n43813 , n43814 , n43815 , n43816 , n43817 , n43818 , n43819 , n43820 , n43821 , n43822 , 
 n43823 , n43824 , n43825 , n43826 , n43827 , n43828 , n43829 , n43830 , n43831 , n43832 , 
 n43833 , n43834 , n43835 , n43836 , n43837 , n43838 , n43839 , n43840 , n43841 , n43842 , 
 n43843 , n43844 , n43845 , n43846 , n43847 , n43848 , n43849 , n43850 , n43851 , n43852 , 
 n43853 , n43854 , n43855 , n43856 , n43857 , n43858 , n43859 , n43860 , n43861 , n43862 , 
 n43863 , n43864 , n43865 , n43866 , n43867 , n43868 , n43869 , n43870 , n43871 , n43872 , 
 n43873 , n43874 , n43875 , n43876 , n43877 , n43878 , n43879 , n43880 , n43881 , n43882 , 
 n43883 , n43884 , n43885 , n43886 , n43887 , n43888 , n43889 , n43890 , n43891 , n43892 , 
 n43893 , n43894 , n43895 , n43896 , n43897 , n43898 , n43899 , n43900 , n43901 , n43902 , 
 n43903 , n43904 , n43905 , n43906 , n43907 , n43908 , n43909 , n43910 , n43911 , n43912 , 
 n43913 , n43914 , n43915 , n43916 , n43917 , n43918 , n43919 , n43920 , n43921 , n43922 , 
 n43923 , n43924 , n43925 , n43926 , n43927 , n43928 , n43929 , n43930 , n43931 , n43932 , 
 n43933 , n43934 , n43935 , n43936 , n43937 , n43938 , n43939 , n43940 , n43941 , n43942 , 
 n43943 , n43944 , n43945 , n43946 , n43947 , n43948 , n43949 , n43950 , n43951 , n43952 , 
 n43953 , n43954 , n43955 , n43956 , n43957 , n43958 , n43959 , n43960 , n43961 , n43962 , 
 n43963 , n43964 , n43965 , n43966 , n43967 , n43968 , n43969 , n43970 , n43971 , n43972 , 
 n43973 , n43974 , n43975 , n43976 , n43977 , n43978 , n43979 , n43980 , n43981 , n43982 , 
 n43983 , n43984 , n43985 , n43986 , n43987 , n43988 , n43989 , n43990 , n43991 , n43992 , 
 n43993 , n43994 , n43995 , n43996 , n43997 , n43998 , n43999 , n44000 , n44001 , n44002 , 
 n44003 , n44004 , n44005 , n44006 , n44007 , n44008 , n44009 , n44010 , n44011 , n44012 , 
 n44013 , n44014 , n44015 , n44016 , n44017 , n44018 , n44019 , n44020 , n44021 , n44022 , 
 n44023 , n44024 , n44025 , n44026 , n44027 , n44028 , n44029 , n44030 , n44031 , n44032 , 
 n44033 , n44034 , n44035 , n44036 , n44037 , n44038 , n44039 , n44040 , n44041 , n44042 , 
 n44043 , n44044 , n44045 , n44046 , n44047 , n44048 , n44049 , n44050 , n44051 , n44052 , 
 n44053 , n44054 , n44055 , n44056 , n44057 , n44058 , n44059 , n44060 , n44061 , n44062 , 
 n44063 , n44064 , n44065 , n44066 , n44067 , n44068 , n44069 , n44070 , n44071 , n44072 , 
 n44073 , n44074 , n44075 , n44076 , n44077 , n44078 , n44079 , n44080 , n44081 , n44082 , 
 n44083 , n44084 , n44085 , n44086 , n44087 , n44088 , n44089 , n44090 , n44091 , n44092 , 
 n44093 , n44094 , n44095 , n44096 , n44097 , n44098 , n44099 , n44100 , n44101 , n44102 , 
 n44103 , n44104 , n44105 , n44106 , n44107 , n44108 , n44109 , n44110 , n44111 , n44112 , 
 n44113 , n44114 , n44115 , n44116 , n44117 , n44118 , n44119 , n44120 , n44121 , n44122 , 
 n44123 , n44124 , n44125 , n44126 , n44127 , n44128 , n44129 , n44130 , n44131 , n44132 , 
 n44133 , n44134 , n44135 , n44136 , n44137 , n44138 , n44139 , n44140 , n44141 , n44142 , 
 n44143 , n44144 , n44145 , n44146 , n44147 , n44148 , n44149 , n44150 , n44151 , n44152 , 
 n44153 , n44154 , n44155 , n44156 , n44157 , n44158 , n44159 , n44160 , n44161 , n44162 , 
 n44163 , n44164 , n44165 , n44166 , n44167 , n44168 , n44169 , n44170 , n44171 , n44172 , 
 n44173 , n44174 , n44175 , n44176 , n44177 , n44178 , n44179 , n44180 , n44181 , n44182 , 
 n44183 , n44184 , n44185 , n44186 , n44187 , n44188 , n44189 , n44190 , n44191 , n44192 , 
 n44193 , n44194 , n44195 , n44196 , n44197 , n44198 , n44199 , n44200 , n44201 , n44202 , 
 n44203 , n44204 , n44205 , n44206 , n44207 , n44208 , n44209 , n44210 , n44211 , n44212 , 
 n44213 , n44214 , n44215 , n44216 , n44217 , n44218 , n44219 , n44220 , n44221 , n44222 , 
 n44223 , n44224 , n44225 , n44226 , n44227 , n44228 , n44229 , n44230 , n44231 , n44232 , 
 n44233 , n44234 , n44235 , n44236 , n44237 , n44238 , n44239 , n44240 , n44241 , n44242 , 
 n44243 , n44244 , n44245 , n44246 , n44247 , n44248 , n44249 , n44250 , n44251 , n44252 , 
 n44253 , n44254 , n44255 , n44256 , n44257 , n44258 , n44259 , n44260 , n44261 , n44262 , 
 n44263 , n44264 , n44265 , n44266 , n44267 , n44268 , n44269 , n44270 , n44271 , n44272 , 
 n44273 , n44274 , n44275 , n44276 , n44277 , n44278 , n44279 , n44280 , n44281 , n44282 , 
 n44283 , n44284 , n44285 , n44286 , n44287 , n44288 , n44289 , n44290 , n44291 , n44292 , 
 n44293 , n44294 , n44295 , n44296 , n44297 , n44298 , n44299 , n44300 , n44301 , n44302 , 
 n44303 , n44304 , n44305 , n44306 , n44307 , n44308 , n44309 , n44310 , n44311 , n44312 , 
 n44313 , n44314 , n44315 , n44316 , n44317 , n44318 , n44319 , n44320 , n44321 , n44322 , 
 n44323 , n44324 , n44325 , n44326 , n44327 , n44328 , n44329 , n44330 , n44331 , n44332 , 
 n44333 , n44334 , n44335 , n44336 , n44337 , n44338 , n44339 , n44340 , n44341 , n44342 , 
 n44343 , n44344 , n44345 , n44346 , n44347 , n44348 , n44349 , n44350 , n44351 , n44352 , 
 n44353 , n44354 , n44355 , n44356 , n44357 , n44358 , n44359 , n44360 , n44361 , n44362 , 
 n44363 , n44364 , n44365 , n44366 , n44367 , n44368 , n44369 , n44370 , n44371 , n44372 , 
 n44373 , n44374 , n44375 , n44376 , n44377 , n44378 , n44379 , n44380 , n44381 , n44382 , 
 n44383 , n44384 , n44385 , n44386 , n44387 , n44388 , n44389 , n44390 , n44391 , n44392 , 
 n44393 , n44394 , n44395 , n44396 , n44397 , n44398 , n44399 , n44400 , n44401 , n44402 , 
 n44403 , n44404 , n44405 , n44406 , n44407 , n44408 , n44409 , n44410 , n44411 , n44412 , 
 n44413 , n44414 , n44415 , n44416 , n44417 , n44418 , n44419 , n44420 , n44421 , n44422 , 
 n44423 , n44424 , n44425 , n44426 , n44427 , n44428 , n44429 , n44430 , n44431 , n44432 , 
 n44433 , n44434 , n44435 , n44436 , n44437 , n44438 , n44439 , n44440 , n44441 , n44442 , 
 n44443 , n44444 , n44445 , n44446 , n44447 , n44448 , n44449 , n44450 , n44451 , n44452 , 
 n44453 , n44454 , n44455 , n44456 , n44457 , n44458 , n44459 , n44460 , n44461 , n44462 , 
 n44463 , n44464 , n44465 , n44466 , n44467 , n44468 , n44469 , n44470 , n44471 , n44472 , 
 n44473 , n44474 , n44475 , n44476 , n44477 , n44478 , n44479 , n44480 , n44481 , n44482 , 
 n44483 , n44484 , n44485 , n44486 , n44487 , n44488 , n44489 , n44490 , n44491 , n44492 , 
 n44493 , n44494 , n44495 , n44496 , n44497 , n44498 , n44499 , n44500 , n44501 , n44502 , 
 n44503 , n44504 , n44505 , n44506 , n44507 , n44508 , n44509 , n44510 , n44511 , n44512 , 
 n44513 , n44514 , n44515 , n44516 , n44517 , n44518 , n44519 , n44520 , n44521 , n44522 , 
 n44523 , n44524 , n44525 , n44526 , n44527 , n44528 , n44529 , n44530 , n44531 , n44532 , 
 n44533 , n44534 , n44535 , n44536 , n44537 , n44538 , n44539 , n44540 , n44541 , n44542 , 
 n44543 , n44544 , n44545 , n44546 , n44547 , n44548 , n44549 , n44550 , n44551 , n44552 , 
 n44553 , n44554 , n44555 , n44556 , n44557 , n44558 , n44559 , n44560 , n44561 , n44562 , 
 n44563 , n44564 , n44565 , n44566 , n44567 , n44568 , n44569 , n44570 , n44571 , n44572 , 
 n44573 , n44574 , n44575 , n44576 , n44577 , n44578 , n44579 , n44580 , n44581 , n44582 , 
 n44583 , n44584 , n44585 , n44586 , n44587 , n44588 , n44589 , n44590 , n44591 , n44592 , 
 n44593 , n44594 , n44595 , n44596 , n44597 , n44598 , n44599 , n44600 , n44601 , n44602 , 
 n44603 , n44604 , n44605 , n44606 , n44607 , n44608 , n44609 , n44610 , n44611 , n44612 , 
 n44613 , n44614 , n44615 , n44616 , n44617 , n44618 , n44619 , n44620 , n44621 , n44622 , 
 n44623 , n44624 , n44625 , n44626 , n44627 , n44628 , n44629 , n44630 , n44631 , n44632 , 
 n44633 , n44634 , n44635 , n44636 , n44637 , n44638 , n44639 , n44640 , n44641 , n44642 , 
 n44643 , n44644 , n44645 , n44646 , n44647 , n44648 , n44649 , n44650 , n44651 , n44652 , 
 n44653 , n44654 , n44655 , n44656 , n44657 , n44658 , n44659 , n44660 , n44661 , n44662 , 
 n44663 , n44664 , n44665 , n44666 , n44667 , n44668 , n44669 , n44670 , n44671 , n44672 , 
 n44673 , n44674 , n44675 , n44676 , n44677 , n44678 , n44679 , n44680 , n44681 , n44682 , 
 n44683 , n44684 , n44685 , n44686 , n44687 , n44688 , n44689 , n44690 , n44691 , n44692 , 
 n44693 , n44694 , n44695 , n44696 , n44697 , n44698 , n44699 , n44700 , n44701 , n44702 , 
 n44703 , n44704 , n44705 , n44706 , n44707 , n44708 , n44709 , n44710 , n44711 , n44712 , 
 n44713 , n44714 , n44715 , n44716 , n44717 , n44718 , n44719 , n44720 , n44721 , n44722 , 
 n44723 , n44724 , n44725 , n44726 , n44727 , n44728 , n44729 , n44730 , n44731 , n44732 , 
 n44733 , n44734 , n44735 , n44736 , n44737 , n44738 , n44739 , n44740 , n44741 , n44742 , 
 n44743 , n44744 , n44745 , n44746 , n44747 , n44748 , n44749 , n44750 , n44751 , n44752 , 
 n44753 , n44754 , n44755 , n44756 , n44757 , n44758 , n44759 , n44760 , n44761 , n44762 , 
 n44763 , n44764 , n44765 , n44766 , n44767 , n44768 , n44769 , n44770 , n44771 , n44772 , 
 n44773 , n44774 , n44775 , n44776 , n44777 , n44778 , n44779 , n44780 , n44781 , n44782 , 
 n44783 , n44784 , n44785 , n44786 , n44787 , n44788 , n44789 , n44790 , n44791 , n44792 , 
 n44793 , n44794 , n44795 , n44796 , n44797 , n44798 , n44799 , n44800 , n44801 , n44802 , 
 n44803 , n44804 , n44805 , n44806 , n44807 , n44808 , n44809 , n44810 , n44811 , n44812 , 
 n44813 , n44814 , n44815 , n44816 , n44817 , n44818 , n44819 , n44820 , n44821 , n44822 , 
 n44823 , n44824 , n44825 , n44826 , n44827 , n44828 , n44829 , n44830 , n44831 , n44832 , 
 n44833 , n44834 , n44835 , n44836 , n44837 , n44838 , n44839 , n44840 , n44841 , n44842 , 
 n44843 , n44844 , n44845 , n44846 , n44847 , n44848 , n44849 , n44850 , n44851 , n44852 , 
 n44853 , n44854 , n44855 , n44856 , n44857 , n44858 , n44859 , n44860 , n44861 , n44862 , 
 n44863 , n44864 , n44865 , n44866 , n44867 , n44868 , n44869 , n44870 , n44871 , n44872 , 
 n44873 , n44874 , n44875 , n44876 , n44877 , n44878 , n44879 , n44880 , n44881 , n44882 , 
 n44883 , n44884 , n44885 , n44886 , n44887 , n44888 , n44889 , n44890 , n44891 , n44892 , 
 n44893 , n44894 , n44895 , n44896 , n44897 , n44898 , n44899 , n44900 , n44901 , n44902 , 
 n44903 , n44904 , n44905 , n44906 , n44907 , n44908 , n44909 , n44910 , n44911 , n44912 , 
 n44913 , n44914 , n44915 , n44916 , n44917 , n44918 , n44919 , n44920 , n44921 , n44922 , 
 n44923 , n44924 , n44925 , n44926 , n44927 , n44928 , n44929 , n44930 , n44931 , n44932 , 
 n44933 , n44934 , n44935 , n44936 , n44937 , n44938 , n44939 , n44940 , n44941 , n44942 , 
 n44943 , n44944 , n44945 , n44946 , n44947 , n44948 , n44949 , n44950 , n44951 , n44952 , 
 n44953 , n44954 , n44955 , n44956 , n44957 , n44958 , n44959 , n44960 , n44961 , n44962 , 
 n44963 , n44964 , n44965 , n44966 , n44967 , n44968 , n44969 , n44970 , n44971 , n44972 , 
 n44973 , n44974 , n44975 , n44976 , n44977 , n44978 , n44979 , n44980 , n44981 , n44982 , 
 n44983 , n44984 , n44985 , n44986 , n44987 , n44988 , n44989 , n44990 , n44991 , n44992 , 
 n44993 , n44994 , n44995 , n44996 , n44997 , n44998 , n44999 , n45000 , n45001 , n45002 , 
 n45003 , n45004 , n45005 , n45006 , n45007 , n45008 , n45009 , n45010 , n45011 , n45012 , 
 n45013 , n45014 , n45015 , n45016 , n45017 , n45018 , n45019 , n45020 , n45021 , n45022 , 
 n45023 , n45024 , n45025 , n45026 , n45027 , n45028 , n45029 , n45030 , n45031 , n45032 , 
 n45033 , n45034 , n45035 , n45036 , n45037 , n45038 , n45039 , n45040 , n45041 , n45042 , 
 n45043 , n45044 , n45045 , n45046 , n45047 , n45048 , n45049 , n45050 , n45051 , n45052 , 
 n45053 , n45054 , n45055 , n45056 , n45057 , n45058 , n45059 , n45060 , n45061 , n45062 , 
 n45063 , n45064 , n45065 , n45066 , n45067 , n45068 , n45069 , n45070 , n45071 , n45072 , 
 n45073 , n45074 , n45075 , n45076 , n45077 , n45078 , n45079 , n45080 , n45081 , n45082 , 
 n45083 , n45084 , n45085 , n45086 , n45087 , n45088 , n45089 , n45090 , n45091 , n45092 , 
 n45093 , n45094 , n45095 , n45096 , n45097 , n45098 , n45099 , n45100 , n45101 , n45102 , 
 n45103 , n45104 , n45105 , n45106 , n45107 , n45108 , n45109 , n45110 , n45111 , n45112 , 
 n45113 , n45114 , n45115 , n45116 , n45117 , n45118 , n45119 , n45120 , n45121 , n45122 , 
 n45123 , n45124 , n45125 , n45126 , n45127 , n45128 , n45129 , n45130 , n45131 , n45132 , 
 n45133 , n45134 , n45135 , n45136 , n45137 , n45138 , n45139 , n45140 , n45141 , n45142 , 
 n45143 , n45144 , n45145 , n45146 , n45147 , n45148 , n45149 , n45150 , n45151 , n45152 , 
 n45153 , n45154 , n45155 , n45156 , n45157 , n45158 , n45159 , n45160 , n45161 , n45162 , 
 n45163 , n45164 , n45165 , n45166 , n45167 , n45168 , n45169 , n45170 , n45171 , n45172 , 
 n45173 , n45174 , n45175 , n45176 , n45177 , n45178 , n45179 , n45180 , n45181 , n45182 , 
 n45183 , n45184 , n45185 , n45186 , n45187 , n45188 , n45189 , n45190 , n45191 , n45192 , 
 n45193 , n45194 , n45195 , n45196 , n45197 , n45198 , n45199 , n45200 , n45201 , n45202 , 
 n45203 , n45204 , n45205 , n45206 , n45207 , n45208 , n45209 , n45210 , n45211 , n45212 , 
 n45213 , n45214 , n45215 , n45216 , n45217 , n45218 , n45219 , n45220 , n45221 , n45222 , 
 n45223 , n45224 , n45225 , n45226 , n45227 , n45228 , n45229 , n45230 , n45231 , n45232 , 
 n45233 , n45234 , n45235 , n45236 , n45237 , n45238 , n45239 , n45240 , n45241 , n45242 , 
 n45243 , n45244 , n45245 , n45246 , n45247 , n45248 , n45249 , n45250 , n45251 , n45252 , 
 n45253 , n45254 , n45255 , n45256 , n45257 , n45258 , n45259 , n45260 , n45261 , n45262 , 
 n45263 , n45264 , n45265 , n45266 , n45267 , n45268 , n45269 , n45270 , n45271 , n45272 , 
 n45273 , n45274 , n45275 , n45276 , n45277 , n45278 , n45279 , n45280 , n45281 , n45282 , 
 n45283 , n45284 , n45285 , n45286 , n45287 , n45288 , n45289 , n45290 , n45291 , n45292 , 
 n45293 , n45294 , n45295 , n45296 , n45297 , n45298 , n45299 , n45300 , n45301 , n45302 , 
 n45303 , n45304 , n45305 , n45306 , n45307 , n45308 , n45309 , n45310 , n45311 , n45312 , 
 n45313 , n45314 , n45315 , n45316 , n45317 , n45318 , n45319 , n45320 , n45321 , n45322 , 
 n45323 , n45324 , n45325 , n45326 , n45327 , n45328 , n45329 , n45330 , n45331 , n45332 , 
 n45333 , n45334 , n45335 , n45336 , n45337 , n45338 , n45339 , n45340 , n45341 , n45342 , 
 n45343 , n45344 , n45345 , n45346 , n45347 , n45348 , n45349 , n45350 , n45351 , n45352 , 
 n45353 , n45354 , n45355 , n45356 , n45357 , n45358 , n45359 , n45360 , n45361 , n45362 , 
 n45363 , n45364 , n45365 , n45366 , n45367 , n45368 , n45369 , n45370 , n45371 , n45372 , 
 n45373 , n45374 , n45375 , n45376 , n45377 , n45378 , n45379 , n45380 , n45381 , n45382 , 
 n45383 , n45384 , n45385 , n45386 , n45387 , n45388 , n45389 , n45390 , n45391 , n45392 , 
 n45393 , n45394 , n45395 , n45396 , n45397 , n45398 , n45399 , n45400 , n45401 , n45402 , 
 n45403 , n45404 , n45405 , n45406 , n45407 , n45408 , n45409 , n45410 , n45411 , n45412 , 
 n45413 , n45414 , n45415 , n45416 , n45417 , n45418 , n45419 , n45420 , n45421 , n45422 , 
 n45423 , n45424 , n45425 , n45426 , n45427 , n45428 , n45429 , n45430 , n45431 , n45432 , 
 n45433 , n45434 , n45435 , n45436 , n45437 , n45438 , n45439 , n45440 , n45441 , n45442 , 
 n45443 , n45444 , n45445 , n45446 , n45447 , n45448 , n45449 , n45450 , n45451 , n45452 , 
 n45453 , n45454 , n45455 , n45456 , n45457 , n45458 , n45459 , n45460 , n45461 , n45462 , 
 n45463 , n45464 , n45465 , n45466 , n45467 , n45468 , n45469 , n45470 , n45471 , n45472 , 
 n45473 , n45474 , n45475 , n45476 , n45477 , n45478 , n45479 , n45480 , n45481 , n45482 , 
 n45483 , n45484 , n45485 , n45486 , n45487 , n45488 , n45489 , n45490 , n45491 , n45492 , 
 n45493 , n45494 , n45495 , n45496 , n45497 , n45498 , n45499 , n45500 , n45501 , n45502 , 
 n45503 , n45504 , n45505 , n45506 , n45507 , n45508 , n45509 , n45510 , n45511 , n45512 , 
 n45513 , n45514 , n45515 , n45516 , n45517 , n45518 , n45519 , n45520 , n45521 , n45522 , 
 n45523 , n45524 , n45525 , n45526 , n45527 , n45528 , n45529 , n45530 , n45531 , n45532 , 
 n45533 , n45534 , n45535 , n45536 , n45537 , n45538 , n45539 , n45540 , n45541 , n45542 , 
 n45543 , n45544 , n45545 , n45546 , n45547 , n45548 , n45549 , n45550 , n45551 , n45552 , 
 n45553 , n45554 , n45555 , n45556 , n45557 , n45558 , n45559 , n45560 , n45561 , n45562 , 
 n45563 , n45564 , n45565 , n45566 , n45567 , n45568 , n45569 , n45570 , n45571 , n45572 , 
 n45573 , n45574 , n45575 , n45576 , n45577 , n45578 , n45579 , n45580 , n45581 , n45582 , 
 n45583 , n45584 , n45585 , n45586 , n45587 , n45588 , n45589 , n45590 , n45591 , n45592 , 
 n45593 , n45594 , n45595 , n45596 , n45597 , n45598 , n45599 , n45600 , n45601 , n45602 , 
 n45603 , n45604 , n45605 , n45606 , n45607 , n45608 , n45609 , n45610 , n45611 , n45612 , 
 n45613 , n45614 , n45615 , n45616 , n45617 , n45618 , n45619 , n45620 , n45621 , n45622 , 
 n45623 , n45624 , n45625 , n45626 , n45627 , n45628 , n45629 , n45630 , n45631 , n45632 , 
 n45633 , n45634 , n45635 , n45636 , n45637 , n45638 , n45639 , n45640 , n45641 , n45642 , 
 n45643 , n45644 , n45645 , n45646 , n45647 , n45648 , n45649 , n45650 , n45651 , n45652 , 
 n45653 , n45654 , n45655 , n45656 , n45657 , n45658 , n45659 , n45660 , n45661 , n45662 , 
 n45663 , n45664 , n45665 , n45666 , n45667 , n45668 , n45669 , n45670 , n45671 , n45672 , 
 n45673 , n45674 , n45675 , n45676 , n45677 , n45678 , n45679 , n45680 , n45681 , n45682 , 
 n45683 , n45684 , n45685 , n45686 , n45687 , n45688 , n45689 , n45690 , n45691 , n45692 , 
 n45693 , n45694 , n45695 , n45696 , n45697 , n45698 , n45699 , n45700 , n45701 , n45702 , 
 n45703 , n45704 , n45705 , n45706 , n45707 , n45708 , n45709 , n45710 , n45711 , n45712 , 
 n45713 , n45714 , n45715 , n45716 , n45717 , n45718 , n45719 , n45720 , n45721 , n45722 , 
 n45723 , n45724 , n45725 , n45726 , n45727 , n45728 , n45729 , n45730 , n45731 , n45732 , 
 n45733 , n45734 , n45735 , n45736 , n45737 , n45738 , n45739 , n45740 , n45741 , n45742 , 
 n45743 , n45744 , n45745 , n45746 , n45747 , n45748 , n45749 , n45750 , n45751 , n45752 , 
 n45753 , n45754 , n45755 , n45756 , n45757 , n45758 , n45759 , n45760 , n45761 , n45762 , 
 n45763 , n45764 , n45765 , n45766 , n45767 , n45768 , n45769 , n45770 , n45771 , n45772 , 
 C0n , C0 , C1n , C1 ;
buf ( n454 , n0 );
buf ( n455 , n1 );
buf ( n456 , n2 );
buf ( n457 , n3 );
buf ( n458 , n4 );
buf ( n459 , n5 );
buf ( n460 , n6 );
buf ( n461 , n7 );
buf ( n462 , n8 );
buf ( n463 , n9 );
buf ( n464 , n10 );
buf ( n465 , n11 );
buf ( n466 , n12 );
buf ( n467 , n13 );
buf ( n468 , n14 );
buf ( n469 , n15 );
buf ( n470 , n16 );
buf ( n471 , n17 );
buf ( n472 , n18 );
buf ( n473 , n19 );
buf ( n474 , n20 );
buf ( n475 , n21 );
buf ( n476 , n22 );
buf ( n477 , n23 );
buf ( n478 , n24 );
buf ( n479 , n25 );
buf ( n480 , n26 );
buf ( n481 , n27 );
buf ( n482 , n28 );
buf ( n483 , n29 );
buf ( n484 , n30 );
buf ( n485 , n31 );
buf ( n486 , n32 );
buf ( n487 , n33 );
buf ( n488 , n34 );
buf ( n489 , n35 );
buf ( n490 , n36 );
buf ( n491 , n37 );
buf ( n492 , n38 );
buf ( n493 , n39 );
buf ( n494 , n40 );
buf ( n495 , n41 );
buf ( n496 , n42 );
buf ( n497 , n43 );
buf ( n498 , n44 );
buf ( n499 , n45 );
buf ( n500 , n46 );
buf ( n501 , n47 );
buf ( n502 , n48 );
buf ( n503 , n49 );
buf ( n504 , n50 );
buf ( n505 , n51 );
buf ( n506 , n52 );
buf ( n507 , n53 );
buf ( n508 , n54 );
buf ( n509 , n55 );
buf ( n510 , n56 );
buf ( n511 , n57 );
buf ( n512 , n58 );
buf ( n513 , n59 );
buf ( n514 , n60 );
buf ( n515 , n61 );
buf ( n516 , n62 );
buf ( n517 , n63 );
buf ( n518 , n64 );
buf ( n519 , n65 );
buf ( n520 , n66 );
buf ( n521 , n67 );
buf ( n522 , n68 );
buf ( n523 , n69 );
buf ( n524 , n70 );
buf ( n525 , n71 );
buf ( n526 , n72 );
buf ( n527 , n73 );
buf ( n528 , n74 );
buf ( n529 , n75 );
buf ( n530 , n76 );
buf ( n531 , n77 );
buf ( n532 , n78 );
buf ( n533 , n79 );
buf ( n534 , n80 );
buf ( n535 , n81 );
buf ( n536 , n82 );
buf ( n537 , n83 );
buf ( n538 , n84 );
buf ( n539 , n85 );
buf ( n540 , n86 );
buf ( n541 , n87 );
buf ( n542 , n88 );
buf ( n543 , n89 );
buf ( n544 , n90 );
buf ( n545 , n91 );
buf ( n546 , n92 );
buf ( n547 , n93 );
buf ( n548 , n94 );
buf ( n549 , n95 );
buf ( n550 , n96 );
buf ( n551 , n97 );
buf ( n552 , n98 );
buf ( n99 , n553 );
buf ( n100 , n554 );
buf ( n101 , n555 );
buf ( n102 , n556 );
buf ( n103 , n557 );
buf ( n104 , n558 );
buf ( n105 , n559 );
buf ( n106 , n560 );
buf ( n107 , n561 );
buf ( n108 , n562 );
buf ( n109 , n563 );
buf ( n110 , n564 );
buf ( n111 , n565 );
buf ( n112 , n566 );
buf ( n113 , n567 );
buf ( n114 , n568 );
buf ( n115 , n569 );
buf ( n116 , n570 );
buf ( n117 , n571 );
buf ( n118 , n572 );
buf ( n119 , n573 );
buf ( n120 , n574 );
buf ( n121 , n575 );
buf ( n122 , n576 );
buf ( n123 , n577 );
buf ( n124 , n578 );
buf ( n125 , n579 );
buf ( n126 , n580 );
buf ( n127 , n581 );
buf ( n128 , n582 );
buf ( n129 , n583 );
buf ( n130 , n584 );
buf ( n131 , n585 );
buf ( n132 , n586 );
buf ( n133 , n587 );
buf ( n134 , n588 );
buf ( n135 , n589 );
buf ( n136 , n590 );
buf ( n137 , n591 );
buf ( n138 , n592 );
buf ( n139 , n593 );
buf ( n140 , n594 );
buf ( n141 , n595 );
buf ( n142 , n596 );
buf ( n143 , n597 );
buf ( n144 , n598 );
buf ( n145 , n599 );
buf ( n146 , n600 );
buf ( n147 , n601 );
buf ( n148 , n602 );
buf ( n149 , n603 );
buf ( n150 , n604 );
buf ( n151 , n605 );
buf ( n152 , n606 );
buf ( n153 , n607 );
buf ( n154 , n608 );
buf ( n155 , n609 );
buf ( n156 , n610 );
buf ( n157 , n611 );
buf ( n158 , n612 );
buf ( n159 , n613 );
buf ( n160 , n614 );
buf ( n161 , n615 );
buf ( n162 , n616 );
buf ( n163 , n617 );
buf ( n164 , n618 );
buf ( n165 , n619 );
buf ( n166 , n620 );
buf ( n167 , n621 );
buf ( n168 , n622 );
buf ( n169 , n623 );
buf ( n170 , n624 );
buf ( n171 , n625 );
buf ( n172 , n626 );
buf ( n173 , n627 );
buf ( n174 , n628 );
buf ( n175 , n629 );
buf ( n176 , n630 );
buf ( n177 , n631 );
buf ( n178 , n632 );
buf ( n179 , n633 );
buf ( n180 , n634 );
buf ( n181 , n635 );
buf ( n182 , n636 );
buf ( n183 , n637 );
buf ( n184 , n638 );
buf ( n185 , n639 );
buf ( n186 , n640 );
buf ( n187 , n641 );
buf ( n188 , n642 );
buf ( n189 , n643 );
buf ( n190 , n644 );
buf ( n191 , n645 );
buf ( n192 , n646 );
buf ( n193 , n647 );
buf ( n194 , n648 );
buf ( n195 , n649 );
buf ( n196 , n650 );
buf ( n197 , n651 );
buf ( n198 , n652 );
buf ( n199 , n653 );
buf ( n200 , n654 );
buf ( n201 , n655 );
buf ( n202 , n656 );
buf ( n203 , n657 );
buf ( n204 , n658 );
buf ( n205 , n659 );
buf ( n206 , n660 );
buf ( n207 , n661 );
buf ( n208 , n662 );
buf ( n209 , n663 );
buf ( n210 , n664 );
buf ( n211 , n665 );
buf ( n212 , n666 );
buf ( n213 , n667 );
buf ( n214 , n668 );
buf ( n215 , n669 );
buf ( n216 , n670 );
buf ( n217 , n671 );
buf ( n218 , n672 );
buf ( n219 , n673 );
buf ( n220 , n674 );
buf ( n221 , n675 );
buf ( n222 , n676 );
buf ( n223 , n677 );
buf ( n224 , n678 );
buf ( n225 , n679 );
buf ( n226 , n680 );
buf ( n553 , C0 );
buf ( n554 , C0 );
buf ( n555 , C0 );
buf ( n556 , C0 );
buf ( n557 , C0 );
buf ( n558 , C0 );
buf ( n559 , C0 );
buf ( n560 , C0 );
buf ( n561 , C0 );
buf ( n562 , C0 );
buf ( n563 , C0 );
buf ( n564 , C0 );
buf ( n565 , C0 );
buf ( n566 , C0 );
buf ( n567 , C0 );
buf ( n568 , C0 );
buf ( n569 , C0 );
buf ( n570 , C0 );
buf ( n571 , C0 );
buf ( n572 , C0 );
buf ( n573 , C0 );
buf ( n574 , C0 );
buf ( n575 , C0 );
buf ( n576 , C0 );
buf ( n577 , C0 );
buf ( n578 , C0 );
buf ( n579 , C0 );
buf ( n580 , C0 );
buf ( n581 , C0 );
buf ( n582 , C0 );
buf ( n583 , C0 );
buf ( n584 , n45646 );
buf ( n585 , n45525 );
buf ( n586 , n45633 );
buf ( n587 , n45442 );
buf ( n588 , n45648 );
buf ( n589 , n45277 );
buf ( n590 , n45370 );
buf ( n591 , n45394 );
buf ( n592 , n45473 );
buf ( n593 , n45564 );
buf ( n594 , n45332 );
buf ( n595 , n45532 );
buf ( n596 , n45636 );
buf ( n597 , n45631 );
buf ( n598 , n42086 );
buf ( n599 , n41028 );
buf ( n600 , n40945 );
buf ( n601 , n40879 );
buf ( n602 , n42140 );
buf ( n603 , n42142 );
buf ( n604 , n40917 );
buf ( n605 , n40931 );
buf ( n606 , n40895 );
buf ( n607 , n40906 );
buf ( n608 , n3832 );
buf ( n609 , n3898 );
buf ( n610 , n3888 );
buf ( n611 , n3877 );
buf ( n612 , n45743 );
buf ( n613 , n44992 );
buf ( n614 , n44998 );
buf ( n615 , n45680 );
buf ( n616 , n45132 );
buf ( n617 , C0 );
buf ( n618 , C0 );
buf ( n619 , C0 );
buf ( n620 , C0 );
buf ( n621 , C0 );
buf ( n622 , C0 );
buf ( n623 , C0 );
buf ( n624 , C0 );
buf ( n625 , C0 );
buf ( n626 , C0 );
buf ( n627 , C0 );
buf ( n628 , C0 );
buf ( n629 , C0 );
buf ( n630 , C0 );
buf ( n631 , C0 );
buf ( n632 , C0 );
buf ( n633 , C0 );
buf ( n634 , C0 );
buf ( n635 , C0 );
buf ( n636 , C0 );
buf ( n637 , C0 );
buf ( n638 , C0 );
buf ( n639 , C0 );
buf ( n640 , C0 );
buf ( n641 , C0 );
buf ( n642 , C0 );
buf ( n643 , C0 );
buf ( n644 , C0 );
buf ( n645 , C0 );
buf ( n646 , C0 );
buf ( n647 , C0 );
buf ( n648 , C0 );
buf ( n649 , C0 );
buf ( n650 , C0 );
buf ( n651 , n42904 );
buf ( n652 , n45757 );
buf ( n653 , n45752 );
buf ( n654 , n45528 );
buf ( n655 , n45772 );
buf ( n656 , n45766 );
buf ( n657 , n45722 );
buf ( n658 , n45669 );
buf ( n659 , n45749 );
buf ( n660 , n45598 );
buf ( n661 , n45630 );
buf ( n662 , n45579 );
buf ( n663 , n45547 );
buf ( n664 , n42058 );
buf ( n665 , n45708 );
buf ( n666 , n42138 );
buf ( n667 , n42110 );
buf ( n668 , n45695 );
buf ( n669 , n45732 );
buf ( n670 , n42084 );
buf ( n671 , n42157 );
buf ( n672 , n42917 );
buf ( n673 , n45736 );
buf ( n674 , n42170 );
buf ( n675 , n42183 );
buf ( n676 , n42933 );
buf ( n677 , n3996 );
buf ( n678 , n45700 );
buf ( n679 , n42926 );
buf ( n680 , n42910 );
and ( n29489 , n456 , n468 );
not ( n29490 , n456 );
and ( n29491 , n29490 , n484 );
nor ( n29492 , n29489 , n29491 );
not ( n29493 , n29492 );
buf ( n29494 , n29493 );
and ( n29495 , n456 , n458 );
not ( n29496 , n456 );
and ( n29497 , n29496 , n474 );
nor ( n29498 , n29495 , n29497 );
not ( n29499 , n29498 );
buf ( n29500 , n29499 );
not ( n29501 , n456 );
nand ( n29502 , n29501 , n479 );
nand ( n29503 , n456 , n463 );
nand ( n29504 , n29502 , n29503 );
buf ( n29505 , n29504 );
buf ( n29506 , n29505 );
and ( n29507 , n456 , n461 );
not ( n29508 , n456 );
and ( n29509 , n29508 , n477 );
nor ( n29510 , n29507 , n29509 );
not ( n29511 , n29510 );
buf ( n29512 , n29511 );
xnor ( n29513 , n454 , n456 );
and ( n29514 , n29513 , n455 );
not ( n29515 , n29513 );
not ( n29516 , n455 );
and ( n29517 , n29515 , n29516 );
or ( n29518 , n29514 , n29517 );
not ( n29519 , n29518 );
not ( n29520 , n29519 );
not ( n29521 , n29520 );
xor ( n29522 , n494 , n495 );
not ( n29523 , n29522 );
buf ( n29524 , n493 );
not ( n29525 , n29524 );
and ( n29526 , n456 , n471 );
not ( n29527 , n456 );
and ( n29528 , n29527 , n487 );
nor ( n29529 , n29526 , n29528 );
buf ( n29530 , n29529 );
not ( n29531 , n29530 );
or ( n29532 , n29525 , n29531 );
buf ( n29533 , n29529 );
not ( n29534 , n29533 );
buf ( n29535 , n29534 );
buf ( n29536 , n29535 );
not ( n29537 , n493 );
buf ( n29538 , n29537 );
nand ( n29539 , n29536 , n29538 );
buf ( n29540 , n29539 );
buf ( n29541 , n29540 );
nand ( n29542 , n29532 , n29541 );
buf ( n29543 , n29542 );
not ( n29544 , n29543 );
or ( n29545 , n29523 , n29544 );
buf ( n29546 , n493 );
not ( n29547 , n29546 );
and ( n29548 , n456 , n472 );
not ( n29549 , n456 );
and ( n29550 , n29549 , n488 );
nor ( n29551 , n29548 , n29550 );
buf ( n29552 , n29551 );
not ( n29553 , n29552 );
or ( n29554 , n29547 , n29553 );
buf ( n29555 , n29551 );
not ( n29556 , n29555 );
buf ( n29557 , n29556 );
buf ( n29558 , n29557 );
buf ( n29559 , n29537 );
nand ( n29560 , n29558 , n29559 );
buf ( n29561 , n29560 );
buf ( n29562 , n29561 );
nand ( n29563 , n29554 , n29562 );
buf ( n29564 , n29563 );
buf ( n29565 , n29564 );
not ( n29566 , n493 );
not ( n29567 , n495 );
not ( n29568 , n494 );
nand ( n29569 , n29567 , n29568 );
not ( n29570 , n29569 );
or ( n29571 , n29566 , n29570 );
not ( n29572 , n493 );
nand ( n29573 , n494 , n495 );
nand ( n29574 , n29572 , n29573 );
nand ( n29575 , n29571 , n29574 );
not ( n29576 , n29575 );
buf ( n29577 , n29576 );
nand ( n29578 , n29565 , n29577 );
buf ( n29579 , n29578 );
nand ( n29580 , n29545 , n29579 );
xor ( n29581 , n501 , n500 );
not ( n29582 , n29581 );
not ( n29583 , n29582 );
buf ( n29584 , n29583 );
not ( n29585 , n29584 );
buf ( n29586 , n499 );
not ( n29587 , n29586 );
and ( n29588 , n456 , n465 );
not ( n29589 , n456 );
and ( n29590 , n29589 , n481 );
nor ( n29591 , n29588 , n29590 );
buf ( n29592 , n29591 );
not ( n29593 , n29592 );
or ( n29594 , n29587 , n29593 );
or ( n29595 , n456 , n481 );
not ( n29596 , n499 );
not ( n29597 , n465 );
nand ( n29598 , n29597 , n456 );
nand ( n29599 , n29595 , n29596 , n29598 );
buf ( n29600 , n29599 );
nand ( n29601 , n29594 , n29600 );
buf ( n29602 , n29601 );
buf ( n29603 , n29602 );
not ( n29604 , n29603 );
or ( n29605 , n29585 , n29604 );
not ( n29606 , n499 );
and ( n29607 , n456 , n466 );
not ( n29608 , n456 );
and ( n29609 , n29608 , n482 );
nor ( n29610 , n29607 , n29609 );
not ( n29611 , n29610 );
or ( n29612 , n29606 , n29611 );
not ( n29613 , n29610 );
buf ( n29614 , n29613 );
buf ( n29615 , n29596 );
nand ( n29616 , n29614 , n29615 );
buf ( n29617 , n29616 );
nand ( n29618 , n29612 , n29617 );
buf ( n29619 , n499 );
buf ( n29620 , n500 );
xnor ( n29621 , n29619 , n29620 );
buf ( n29622 , n29621 );
nor ( n29623 , n29581 , n29622 );
buf ( n29624 , n29623 );
nand ( n29625 , n29618 , n29624 );
buf ( n29626 , n29625 );
nand ( n29627 , n29605 , n29626 );
buf ( n29628 , n29627 );
xor ( n29629 , n29580 , n29628 );
not ( n29630 , n501 );
not ( n29631 , n29505 );
not ( n29632 , n29631 );
or ( n29633 , n29630 , n29632 );
buf ( n29634 , n29505 );
not ( n29635 , n501 );
buf ( n29636 , n29635 );
nand ( n29637 , n29634 , n29636 );
buf ( n29638 , n29637 );
nand ( n29639 , n29633 , n29638 );
not ( n29640 , n29639 );
not ( n29641 , n502 );
not ( n29642 , n503 );
not ( n29643 , n29642 );
or ( n29644 , n29641 , n29643 );
not ( n29645 , n502 );
nand ( n29646 , n29645 , n503 );
nand ( n29647 , n29644 , n29646 );
not ( n29648 , n29647 );
or ( n29649 , n29640 , n29648 );
not ( n29650 , n501 );
and ( n29651 , n456 , n464 );
not ( n29652 , n456 );
and ( n29653 , n29652 , n480 );
nor ( n29654 , n29651 , n29653 );
not ( n29655 , n29654 );
or ( n29656 , n29650 , n29655 );
buf ( n29657 , n29635 );
not ( n29658 , n29654 );
buf ( n29659 , n29658 );
nand ( n29660 , n29657 , n29659 );
buf ( n29661 , n29660 );
nand ( n29662 , n29656 , n29661 );
xor ( n29663 , n501 , n502 );
buf ( n29664 , n29663 );
and ( n29665 , n502 , n503 );
not ( n29666 , n502 );
and ( n29667 , n29666 , n29642 );
nor ( n29668 , n29665 , n29667 );
not ( n29669 , n29668 );
nand ( n29670 , n29664 , n29669 );
not ( n29671 , n29670 );
nand ( n29672 , n29662 , n29671 );
nand ( n29673 , n29649 , n29672 );
and ( n29674 , n456 , n472 );
not ( n29675 , n456 );
and ( n29676 , n29675 , n488 );
nor ( n29677 , n29674 , n29676 );
not ( n29678 , n29677 );
buf ( n29679 , n29678 );
buf ( n29680 , n29679 );
buf ( n29681 , n29680 );
buf ( n29682 , n29681 );
buf ( n29683 , n494 );
and ( n29684 , n29682 , n29683 );
buf ( n29685 , n29537 );
nor ( n29686 , n29684 , n29685 );
buf ( n29687 , n29686 );
buf ( n29688 , n29687 );
buf ( n29689 , n29678 );
not ( n29690 , n29689 );
buf ( n29691 , n29690 );
buf ( n29692 , n29691 );
not ( n29693 , n29692 );
buf ( n29694 , n29693 );
buf ( n29695 , n29694 );
buf ( n29696 , n494 );
or ( n29697 , n29695 , n29696 );
buf ( n29698 , n495 );
nand ( n29699 , n29697 , n29698 );
buf ( n29700 , n29699 );
buf ( n29701 , n29700 );
nand ( n29702 , n29688 , n29701 );
buf ( n29703 , n29702 );
xnor ( n29704 , n29673 , n29703 );
xor ( n29705 , n29629 , n29704 );
not ( n29706 , n497 );
not ( n29707 , n496 );
nand ( n29708 , n29707 , n29551 );
not ( n29709 , n29708 );
or ( n29710 , n29706 , n29709 );
buf ( n29711 , n29681 );
buf ( n29712 , n496 );
and ( n29713 , n29711 , n29712 );
buf ( n29714 , n495 );
not ( n29715 , n29714 );
buf ( n29716 , n29715 );
buf ( n29717 , n29716 );
nor ( n29718 , n29713 , n29717 );
buf ( n29719 , n29718 );
nand ( n29720 , n29710 , n29719 );
not ( n29721 , n29720 );
buf ( n29722 , n29721 );
buf ( n29723 , n29671 );
not ( n29724 , n29723 );
not ( n29725 , n29635 );
not ( n29726 , n29613 );
or ( n29727 , n29725 , n29726 );
and ( n29728 , n456 , n466 );
not ( n29729 , n456 );
and ( n29730 , n29729 , n482 );
nor ( n29731 , n29728 , n29730 );
nand ( n29732 , n29731 , n501 );
nand ( n29733 , n29727 , n29732 );
buf ( n29734 , n29733 );
not ( n29735 , n29734 );
or ( n29736 , n29724 , n29735 );
xor ( n29737 , n502 , n503 );
not ( n29738 , n501 );
and ( n29739 , n456 , n465 );
not ( n29740 , n456 );
and ( n29741 , n29740 , n481 );
nor ( n29742 , n29739 , n29741 );
not ( n29743 , n29742 );
or ( n29744 , n29738 , n29743 );
and ( n29745 , n456 , n465 );
not ( n29746 , n456 );
and ( n29747 , n29746 , n481 );
nor ( n29748 , n29745 , n29747 );
not ( n29749 , n29748 );
buf ( n29750 , n29749 );
buf ( n29751 , n29635 );
nand ( n29752 , n29750 , n29751 );
buf ( n29753 , n29752 );
nand ( n29754 , n29744 , n29753 );
nand ( n29755 , n29737 , n29754 );
buf ( n29756 , n29755 );
nand ( n29757 , n29736 , n29756 );
buf ( n29758 , n29757 );
buf ( n29759 , n29758 );
and ( n29760 , n29722 , n29759 );
buf ( n29761 , n29760 );
buf ( n29762 , n29691 );
not ( n29763 , n29762 );
buf ( n29764 , n29763 );
and ( n29765 , n29764 , n29522 );
not ( n684 , n29668 );
not ( n29767 , n29662 );
or ( n686 , n684 , n29767 );
nand ( n687 , n29642 , n502 );
not ( n29770 , n687 );
not ( n689 , n503 );
not ( n690 , n29645 );
or ( n691 , n689 , n690 );
nand ( n692 , n691 , n29663 );
nor ( n693 , n29770 , n692 );
nand ( n29776 , n29754 , n693 );
nand ( n695 , n686 , n29776 );
xor ( n696 , n29765 , n695 );
xor ( n697 , n498 , n499 );
not ( n698 , n697 );
not ( n699 , n497 );
or ( n700 , n699 , n498 );
not ( n701 , n498 );
or ( n29784 , n701 , n497 );
nand ( n703 , n700 , n29784 );
and ( n29786 , n698 , n703 );
not ( n705 , n29786 );
not ( n706 , n497 );
not ( n707 , n706 );
and ( n708 , n456 , n469 );
not ( n709 , n456 );
and ( n29792 , n709 , n485 );
nor ( n711 , n708 , n29792 );
not ( n712 , n711 );
buf ( n29795 , n712 );
not ( n714 , n29795 );
buf ( n29797 , n714 );
not ( n716 , n29797 );
not ( n717 , n716 );
or ( n718 , n707 , n717 );
buf ( n29801 , n712 );
not ( n720 , n29801 );
buf ( n29803 , n720 );
nand ( n722 , n29803 , n497 );
nand ( n723 , n718 , n722 );
not ( n724 , n723 );
or ( n725 , n705 , n724 );
buf ( n29808 , n497 );
not ( n727 , n29808 );
buf ( n29810 , n29492 );
not ( n729 , n29810 );
or ( n730 , n727 , n729 );
and ( n731 , n456 , n468 );
not ( n732 , n456 );
and ( n733 , n732 , n484 );
nor ( n734 , n731 , n733 );
buf ( n29817 , n734 );
not ( n736 , n29817 );
buf ( n29819 , n736 );
buf ( n29820 , n29819 );
buf ( n29821 , n706 );
nand ( n743 , n29820 , n29821 );
buf ( n29823 , n743 );
buf ( n29824 , n29823 );
nand ( n29825 , n730 , n29824 );
buf ( n29826 , n29825 );
buf ( n29827 , n697 );
buf ( n29828 , n29827 );
buf ( n29829 , n29828 );
nand ( n751 , n29826 , n29829 );
nand ( n752 , n725 , n751 );
xor ( n753 , n696 , n752 );
xor ( n754 , n29761 , n753 );
not ( n758 , n495 );
nand ( n29835 , n758 , n496 );
not ( n760 , n29835 );
not ( n761 , n496 );
nand ( n762 , n761 , n495 );
not ( n763 , n762 );
or ( n764 , n760 , n763 );
xor ( n765 , n496 , n497 );
not ( n766 , n765 );
nand ( n770 , n764 , n766 );
not ( n29844 , n770 );
buf ( n29845 , n29844 );
not ( n29846 , n29845 );
and ( n774 , n456 , n472 );
not ( n775 , n456 );
and ( n776 , n775 , n488 );
or ( n777 , n774 , n776 );
and ( n778 , n495 , n777 );
not ( n782 , n495 );
buf ( n29853 , n29678 );
not ( n784 , n29853 );
buf ( n29855 , n784 );
and ( n786 , n782 , n29855 );
nor ( n787 , n778 , n786 );
buf ( n29858 , n787 );
not ( n789 , n29858 );
or ( n790 , n29846 , n789 );
and ( n791 , n456 , n471 );
not ( n792 , n456 );
and ( n793 , n792 , n487 );
nor ( n794 , n791 , n793 );
not ( n795 , n794 );
nand ( n796 , n795 , n29716 );
not ( n797 , n796 );
nand ( n798 , n794 , n495 );
not ( n799 , n798 );
or ( n800 , n797 , n799 );
buf ( n29871 , n765 );
buf ( n802 , n29871 );
buf ( n29873 , n802 );
nand ( n804 , n800 , n29873 );
buf ( n29875 , n804 );
nand ( n806 , n790 , n29875 );
buf ( n29877 , n806 );
buf ( n29878 , n29877 );
not ( n809 , n29829 );
not ( n29880 , n723 );
or ( n814 , n809 , n29880 );
buf ( n29882 , n497 );
not ( n29883 , n29882 );
and ( n817 , n456 , n470 );
not ( n818 , n456 );
and ( n819 , n818 , n486 );
nor ( n820 , n817 , n819 );
buf ( n29888 , n820 );
not ( n822 , n29888 );
or ( n823 , n29883 , n822 );
and ( n824 , n456 , n470 );
not ( n825 , n456 );
and ( n29893 , n825 , n486 );
nor ( n827 , n824 , n29893 );
not ( n828 , n827 );
nand ( n829 , n828 , n706 );
buf ( n29897 , n829 );
nand ( n831 , n823 , n29897 );
buf ( n29899 , n831 );
buf ( n29900 , n29899 );
nand ( n834 , n698 , n703 );
not ( n835 , n834 );
buf ( n29903 , n835 );
nand ( n29904 , n29900 , n29903 );
buf ( n29905 , n29904 );
nand ( n842 , n814 , n29905 );
buf ( n29907 , n842 );
xor ( n844 , n29878 , n29907 );
not ( n845 , n504 );
nand ( n846 , n845 , n503 );
not ( n847 , n846 );
buf ( n29912 , n847 );
not ( n849 , n29912 );
buf ( n29914 , n503 );
not ( n851 , n29914 );
and ( n852 , n456 , n464 );
not ( n29917 , n456 );
and ( n854 , n29917 , n480 );
nor ( n855 , n852 , n854 );
buf ( n29920 , n855 );
not ( n857 , n29920 );
or ( n858 , n851 , n857 );
buf ( n29923 , n855 );
not ( n860 , n29923 );
buf ( n29925 , n860 );
buf ( n29926 , n29925 );
not ( n863 , n503 );
buf ( n29928 , n863 );
nand ( n868 , n29926 , n29928 );
buf ( n29930 , n868 );
buf ( n29931 , n29930 );
nand ( n871 , n858 , n29931 );
buf ( n29933 , n871 );
buf ( n29934 , n29933 );
not ( n29935 , n29934 );
or ( n875 , n849 , n29935 );
xor ( n876 , n863 , n29505 );
buf ( n29938 , n876 );
not ( n878 , n29938 );
buf ( n29940 , n504 );
nand ( n29941 , n878 , n29940 );
buf ( n29942 , n29941 );
buf ( n29943 , n29942 );
nand ( n883 , n875 , n29943 );
buf ( n29945 , n883 );
buf ( n29946 , n29945 );
and ( n886 , n844 , n29946 );
and ( n887 , n29878 , n29907 );
or ( n888 , n886 , n887 );
buf ( n29950 , n888 );
and ( n890 , n754 , n29950 );
and ( n891 , n29761 , n753 );
or ( n892 , n890 , n891 );
xor ( n893 , n29705 , n892 );
xor ( n894 , n29765 , n695 );
and ( n895 , n894 , n752 );
and ( n896 , n29765 , n695 );
or ( n897 , n895 , n896 );
buf ( n29959 , n29873 );
not ( n899 , n29959 );
not ( n900 , n29716 );
not ( n901 , n820 );
not ( n902 , n901 );
or ( n903 , n900 , n902 );
nand ( n904 , n820 , n495 );
nand ( n29966 , n903 , n904 );
buf ( n29967 , n29966 );
not ( n907 , n29967 );
or ( n908 , n899 , n907 );
not ( n909 , n798 );
not ( n910 , n796 );
or ( n914 , n909 , n910 );
nand ( n29973 , n914 , n29844 );
buf ( n29974 , n29973 );
nand ( n917 , n908 , n29974 );
buf ( n29976 , n917 );
not ( n919 , n29976 );
buf ( n29978 , n503 );
not ( n29979 , n29978 );
and ( n922 , n456 , n462 );
not ( n923 , n456 );
and ( n924 , n923 , n478 );
nor ( n925 , n922 , n924 );
buf ( n29984 , n925 );
not ( n927 , n29984 );
or ( n928 , n29979 , n927 );
not ( n929 , n456 );
not ( n930 , n478 );
nand ( n931 , n929 , n930 );
not ( n932 , n462 );
nand ( n933 , n932 , n456 );
nand ( n934 , n863 , n931 , n933 );
buf ( n29993 , n934 );
nand ( n936 , n928 , n29993 );
buf ( n29995 , n936 );
buf ( n29996 , n29995 );
not ( n939 , n29996 );
buf ( n29998 , n939 );
not ( n941 , n29998 );
not ( n942 , n504 );
not ( n943 , n942 );
and ( n944 , n941 , n943 );
nand ( n945 , n942 , n503 );
nor ( n30004 , n876 , n945 );
nor ( n950 , n944 , n30004 );
buf ( n30006 , n950 );
not ( n952 , n30006 );
buf ( n30008 , n952 );
not ( n954 , n30008 );
or ( n955 , n919 , n954 );
not ( n956 , n950 );
not ( n957 , n29976 );
not ( n30013 , n957 );
or ( n959 , n956 , n30013 );
buf ( n30015 , n29583 );
not ( n961 , n30015 );
buf ( n30017 , n29618 );
not ( n963 , n30017 );
or ( n964 , n961 , n963 );
buf ( n30020 , n29624 );
buf ( n30021 , n499 );
not ( n967 , n30021 );
and ( n30023 , n456 , n467 );
not ( n969 , n456 );
and ( n970 , n969 , n483 );
nor ( n971 , n30023 , n970 );
buf ( n30027 , n971 );
not ( n973 , n30027 );
or ( n974 , n967 , n973 );
buf ( n30030 , n971 );
not ( n976 , n30030 );
buf ( n30032 , n976 );
buf ( n30033 , n30032 );
buf ( n30034 , n29596 );
nand ( n980 , n30033 , n30034 );
buf ( n30036 , n980 );
buf ( n30037 , n30036 );
nand ( n30038 , n974 , n30037 );
buf ( n30039 , n30038 );
buf ( n30040 , n30039 );
nand ( n986 , n30020 , n30040 );
buf ( n30042 , n986 );
buf ( n30043 , n30042 );
nand ( n989 , n964 , n30043 );
buf ( n30045 , n989 );
nand ( n994 , n959 , n30045 );
nand ( n30047 , n955 , n994 );
xor ( n996 , n897 , n30047 );
buf ( n30049 , n504 );
not ( n998 , n30049 );
and ( n999 , n456 , n461 );
not ( n1000 , n456 );
and ( n1001 , n1000 , n477 );
or ( n1002 , n999 , n1001 );
and ( n1003 , n1002 , n863 );
not ( n1004 , n1002 );
and ( n30057 , n1004 , n503 );
or ( n1006 , n1003 , n30057 );
buf ( n30059 , n1006 );
not ( n1008 , n30059 );
or ( n1009 , n998 , n1008 );
buf ( n30062 , n29995 );
buf ( n30063 , n847 );
nand ( n1012 , n30062 , n30063 );
buf ( n30065 , n1012 );
buf ( n30066 , n30065 );
nand ( n1015 , n1009 , n30066 );
buf ( n30068 , n1015 );
buf ( n30069 , n30068 );
buf ( n30070 , n770 );
not ( n1019 , n30070 );
buf ( n30072 , n1019 );
not ( n1024 , n30072 );
not ( n1025 , n29966 );
or ( n30075 , n1024 , n1025 );
not ( n1027 , n29716 );
not ( n1028 , n712 );
or ( n1029 , n1027 , n1028 );
and ( n1030 , n456 , n469 );
not ( n1031 , n456 );
and ( n30081 , n1031 , n485 );
nor ( n1033 , n1030 , n30081 );
nand ( n1034 , n1033 , n495 );
nand ( n1035 , n1029 , n1034 );
nand ( n1036 , n1035 , n29873 );
nand ( n1037 , n30075 , n1036 );
buf ( n30087 , n1037 );
xor ( n1039 , n30069 , n30087 );
buf ( n30089 , n29829 );
not ( n1041 , n30089 );
buf ( n30091 , n497 );
not ( n1043 , n30091 );
buf ( n30093 , n971 );
not ( n1045 , n30093 );
or ( n1046 , n1043 , n1045 );
buf ( n30096 , n30032 );
buf ( n30097 , n706 );
nand ( n1049 , n30096 , n30097 );
buf ( n30099 , n1049 );
buf ( n30100 , n30099 );
nand ( n1052 , n1046 , n30100 );
buf ( n30102 , n1052 );
buf ( n30103 , n30102 );
not ( n1055 , n30103 );
or ( n1056 , n1041 , n1055 );
buf ( n30106 , n29826 );
buf ( n30107 , n835 );
nand ( n1059 , n30106 , n30107 );
buf ( n30109 , n1059 );
buf ( n30110 , n30109 );
nand ( n1062 , n1056 , n30110 );
buf ( n30112 , n1062 );
buf ( n30113 , n30112 );
xor ( n1065 , n1039 , n30113 );
buf ( n30115 , n1065 );
xor ( n1067 , n996 , n30115 );
xor ( n1068 , n893 , n1067 );
not ( n1069 , n1068 );
buf ( n30119 , n30008 );
buf ( n30120 , n29976 );
xor ( n1072 , n30119 , n30120 );
buf ( n30122 , n1072 );
buf ( n30123 , n30122 );
buf ( n30124 , n30045 );
xor ( n1076 , n30123 , n30124 );
buf ( n30126 , n1076 );
buf ( n30127 , n30126 );
buf ( n30128 , n29624 );
not ( n1080 , n30128 );
buf ( n30130 , n499 );
not ( n1085 , n30130 );
buf ( n30132 , n734 );
not ( n1087 , n30132 );
or ( n1088 , n1085 , n1087 );
buf ( n30135 , n29493 );
buf ( n30136 , n29596 );
nand ( n1091 , n30135 , n30136 );
buf ( n30138 , n1091 );
buf ( n30139 , n30138 );
nand ( n1094 , n1088 , n30139 );
buf ( n30141 , n1094 );
buf ( n30142 , n30141 );
not ( n1097 , n30142 );
or ( n1098 , n1080 , n1097 );
buf ( n30145 , n30039 );
buf ( n30146 , n29583 );
nand ( n1101 , n30145 , n30146 );
buf ( n30148 , n1101 );
buf ( n30149 , n30148 );
nand ( n1104 , n1098 , n30149 );
buf ( n30151 , n1104 );
buf ( n30152 , n30151 );
xor ( n1107 , n29722 , n29759 );
buf ( n30154 , n1107 );
buf ( n30155 , n30154 );
xor ( n1110 , n30152 , n30155 );
buf ( n30157 , n29557 );
buf ( n30158 , n765 );
and ( n1113 , n30157 , n30158 );
buf ( n30160 , n1113 );
buf ( n30161 , n30160 );
not ( n1116 , n29786 );
buf ( n30163 , n497 );
not ( n1118 , n30163 );
buf ( n30165 , n29529 );
not ( n1120 , n30165 );
or ( n1121 , n1118 , n1120 );
buf ( n30168 , n29535 );
buf ( n30169 , n706 );
nand ( n1127 , n30168 , n30169 );
buf ( n30171 , n1127 );
buf ( n30172 , n30171 );
nand ( n1130 , n1121 , n30172 );
buf ( n30174 , n1130 );
not ( n1132 , n30174 );
or ( n1133 , n1116 , n1132 );
buf ( n30177 , n29899 );
buf ( n30178 , n29829 );
nand ( n30179 , n30177 , n30178 );
buf ( n30180 , n30179 );
nand ( n1138 , n1133 , n30180 );
buf ( n30182 , n1138 );
xor ( n1140 , n30161 , n30182 );
buf ( n30184 , n504 );
not ( n1142 , n30184 );
buf ( n30186 , n29933 );
not ( n1144 , n30186 );
or ( n1145 , n1142 , n1144 );
not ( n30189 , n863 );
not ( n1147 , n29749 );
buf ( n30191 , n1147 );
not ( n1149 , n30191 );
buf ( n30193 , n1149 );
not ( n1151 , n30193 );
or ( n1152 , n30189 , n1151 );
not ( n1153 , n456 );
nand ( n1154 , n1153 , n481 );
nand ( n1155 , n456 , n465 );
nand ( n1156 , n1154 , n1155 , n503 );
nand ( n1157 , n1152 , n1156 );
nand ( n1158 , n1157 , n847 );
buf ( n30202 , n1158 );
nand ( n1160 , n1145 , n30202 );
buf ( n30204 , n1160 );
buf ( n30205 , n30204 );
and ( n1163 , n1140 , n30205 );
and ( n1164 , n30161 , n30182 );
or ( n1165 , n1163 , n1164 );
buf ( n30209 , n1165 );
buf ( n30210 , n30209 );
and ( n1168 , n1110 , n30210 );
and ( n30212 , n30152 , n30155 );
or ( n1170 , n1168 , n30212 );
buf ( n30214 , n1170 );
buf ( n30215 , n30214 );
xor ( n1173 , n30127 , n30215 );
xor ( n1174 , n29761 , n753 );
xor ( n1175 , n1174 , n29950 );
buf ( n30219 , n1175 );
and ( n1177 , n1173 , n30219 );
and ( n1178 , n30127 , n30215 );
or ( n1179 , n1177 , n1178 );
buf ( n30223 , n1179 );
not ( n1181 , n30223 );
nand ( n1182 , n1069 , n1181 );
nand ( n1183 , n1068 , n30223 );
nand ( n1187 , n1182 , n1183 );
not ( n30228 , n1187 );
not ( n1189 , n30228 );
xor ( n1190 , n30127 , n30215 );
xor ( n1191 , n1190 , n30219 );
buf ( n30232 , n1191 );
buf ( n30233 , n29671 );
not ( n1194 , n30233 );
buf ( n30235 , n501 );
not ( n1196 , n30235 );
buf ( n30237 , n971 );
not ( n1198 , n30237 );
or ( n1199 , n1196 , n1198 );
and ( n1200 , n456 , n467 );
not ( n1201 , n456 );
and ( n1202 , n1201 , n483 );
nor ( n1203 , n1200 , n1202 );
not ( n1204 , n1203 );
buf ( n30245 , n1204 );
buf ( n30246 , n29635 );
nand ( n1207 , n30245 , n30246 );
buf ( n30248 , n1207 );
buf ( n30249 , n30248 );
nand ( n1210 , n1199 , n30249 );
buf ( n30251 , n1210 );
buf ( n30252 , n30251 );
not ( n1213 , n30252 );
or ( n1214 , n1194 , n1213 );
buf ( n30255 , n29733 );
buf ( n30256 , n29647 );
nand ( n30257 , n30255 , n30256 );
buf ( n30258 , n30257 );
buf ( n30259 , n30258 );
nand ( n1223 , n1214 , n30259 );
buf ( n30261 , n1223 );
buf ( n30262 , n30261 );
buf ( n30263 , n29583 );
not ( n30264 , n30263 );
buf ( n30265 , n30141 );
not ( n1229 , n30265 );
or ( n1230 , n30264 , n1229 );
buf ( n30268 , n499 );
not ( n1232 , n30268 );
buf ( n30270 , n29803 );
not ( n1234 , n30270 );
or ( n1235 , n1232 , n1234 );
buf ( n30273 , n1033 );
not ( n30274 , n30273 );
buf ( n30275 , n29596 );
nand ( n1239 , n30274 , n30275 );
buf ( n30277 , n1239 );
buf ( n30278 , n30277 );
nand ( n1242 , n1235 , n30278 );
buf ( n30280 , n1242 );
buf ( n30281 , n30280 );
buf ( n30282 , n29624 );
nand ( n1246 , n30281 , n30282 );
buf ( n30284 , n1246 );
buf ( n30285 , n30284 );
nand ( n1249 , n1230 , n30285 );
buf ( n30287 , n1249 );
buf ( n30288 , n30287 );
xor ( n1252 , n30262 , n30288 );
not ( n1253 , n504 );
not ( n1254 , n1157 );
or ( n1255 , n1253 , n1254 );
not ( n1256 , n863 );
and ( n1257 , n456 , n466 );
not ( n1258 , n456 );
and ( n1259 , n1258 , n482 );
nor ( n1260 , n1257 , n1259 );
not ( n1261 , n1260 );
not ( n1262 , n1261 );
or ( n1263 , n1256 , n1262 );
nand ( n1264 , n29610 , n503 );
nand ( n1265 , n1263 , n1264 );
nand ( n1266 , n1265 , n847 );
nand ( n1267 , n1255 , n1266 );
buf ( n30305 , n1267 );
nor ( n1269 , n29694 , n498 );
not ( n1270 , n1269 );
not ( n1271 , n29596 );
and ( n1272 , n1270 , n1271 );
buf ( n30310 , n498 );
not ( n1274 , n30310 );
buf ( n30312 , n29681 );
not ( n1276 , n30312 );
or ( n1277 , n1274 , n1276 );
buf ( n30315 , n497 );
nand ( n1279 , n1277 , n30315 );
buf ( n30317 , n1279 );
nor ( n1281 , n1272 , n30317 );
buf ( n30319 , n1281 );
and ( n1283 , n30305 , n30319 );
buf ( n30321 , n1283 );
buf ( n30322 , n30321 );
and ( n1286 , n1252 , n30322 );
and ( n1287 , n30262 , n30288 );
or ( n1288 , n1286 , n1287 );
buf ( n30326 , n1288 );
buf ( n30327 , n30326 );
xor ( n1291 , n29878 , n29907 );
xor ( n30329 , n1291 , n29946 );
buf ( n30330 , n30329 );
buf ( n30331 , n30330 );
xor ( n1295 , n30327 , n30331 );
xor ( n1296 , n30152 , n30155 );
xor ( n1297 , n1296 , n30210 );
buf ( n30335 , n1297 );
buf ( n30336 , n30335 );
and ( n1300 , n1295 , n30336 );
and ( n1301 , n30327 , n30331 );
or ( n1302 , n1300 , n1301 );
buf ( n30340 , n1302 );
or ( n1304 , n30232 , n30340 );
not ( n1305 , n1304 );
xor ( n1309 , n30327 , n30331 );
xor ( n30344 , n1309 , n30336 );
buf ( n30345 , n30344 );
xor ( n1312 , n30161 , n30182 );
xor ( n1313 , n1312 , n30205 );
buf ( n30348 , n1313 );
buf ( n30349 , n30348 );
and ( n1316 , n497 , n29691 );
not ( n1317 , n497 );
and ( n1318 , n1317 , n29764 );
or ( n1319 , n1316 , n1318 );
not ( n1320 , n1319 );
not ( n1321 , n835 );
or ( n1322 , n1320 , n1321 );
nand ( n1323 , n30174 , n29829 );
nand ( n1324 , n1322 , n1323 );
buf ( n30359 , n1324 );
buf ( n30360 , n29624 );
not ( n1327 , n30360 );
not ( n1328 , n499 );
and ( n1329 , n456 , n470 );
not ( n1330 , n456 );
and ( n1331 , n1330 , n486 );
nor ( n1332 , n1329 , n1331 );
not ( n1333 , n1332 );
or ( n1334 , n1328 , n1333 );
buf ( n30369 , n901 );
buf ( n30370 , n29596 );
nand ( n1337 , n30369 , n30370 );
buf ( n30372 , n1337 );
nand ( n1342 , n1334 , n30372 );
buf ( n30374 , n1342 );
not ( n1344 , n30374 );
or ( n1345 , n1327 , n1344 );
buf ( n30377 , n30280 );
buf ( n30378 , n29583 );
nand ( n30379 , n30377 , n30378 );
buf ( n30380 , n30379 );
buf ( n30381 , n30380 );
nand ( n1351 , n1345 , n30381 );
buf ( n30383 , n1351 );
buf ( n30384 , n30383 );
xor ( n1354 , n30359 , n30384 );
and ( n1355 , n29664 , n29669 );
buf ( n30387 , n1355 );
not ( n1357 , n30387 );
not ( n1358 , n29635 );
not ( n1359 , n29819 );
or ( n1360 , n1358 , n1359 );
and ( n1361 , n456 , n468 );
not ( n1362 , n456 );
and ( n1363 , n1362 , n484 );
nor ( n1364 , n1361 , n1363 );
nand ( n1365 , n1364 , n501 );
nand ( n1366 , n1360 , n1365 );
buf ( n30398 , n1366 );
not ( n1368 , n30398 );
or ( n1369 , n1357 , n1368 );
buf ( n30401 , n30251 );
buf ( n30402 , n29737 );
nand ( n1372 , n30401 , n30402 );
buf ( n30404 , n1372 );
buf ( n30405 , n30404 );
nand ( n1375 , n1369 , n30405 );
buf ( n30407 , n1375 );
buf ( n30408 , n30407 );
and ( n1378 , n1354 , n30408 );
and ( n30410 , n30359 , n30384 );
or ( n1380 , n1378 , n30410 );
buf ( n30412 , n1380 );
buf ( n30413 , n30412 );
xor ( n1383 , n30349 , n30413 );
xor ( n1384 , n30262 , n30288 );
xor ( n1385 , n1384 , n30322 );
buf ( n30417 , n1385 );
buf ( n30418 , n30417 );
and ( n1388 , n1383 , n30418 );
and ( n1389 , n30349 , n30413 );
or ( n1390 , n1388 , n1389 );
buf ( n30422 , n1390 );
nand ( n1392 , n30345 , n30422 );
xor ( n1393 , n30349 , n30413 );
xor ( n1394 , n1393 , n30418 );
buf ( n30426 , n1394 );
buf ( n30427 , n1267 );
buf ( n30428 , n1281 );
xor ( n1398 , n30427 , n30428 );
buf ( n30430 , n1398 );
buf ( n30431 , n30430 );
and ( n1401 , n456 , n469 );
not ( n1402 , n456 );
and ( n1403 , n1402 , n485 );
nor ( n1404 , n1401 , n1403 );
not ( n1405 , n1404 );
and ( n1409 , n1405 , n29635 );
not ( n30438 , n1405 );
and ( n1411 , n30438 , n501 );
or ( n1412 , n1409 , n1411 );
not ( n1413 , n1412 );
not ( n1414 , n1355 );
or ( n1415 , n1413 , n1414 );
buf ( n30444 , n1366 );
buf ( n30445 , n29737 );
nand ( n1418 , n30444 , n30445 );
buf ( n30447 , n1418 );
nand ( n1420 , n1415 , n30447 );
not ( n1421 , n1420 );
not ( n1422 , n504 );
not ( n1423 , n1265 );
or ( n1424 , n1422 , n1423 );
buf ( n30453 , n503 );
not ( n1426 , n30453 );
buf ( n30455 , n971 );
not ( n1428 , n30455 );
or ( n1429 , n1426 , n1428 );
buf ( n30458 , n30032 );
buf ( n30459 , n863 );
nand ( n1432 , n30458 , n30459 );
buf ( n30461 , n1432 );
buf ( n30462 , n30461 );
nand ( n1435 , n1429 , n30462 );
buf ( n30464 , n1435 );
buf ( n30465 , n30464 );
buf ( n30466 , n847 );
nand ( n1439 , n30465 , n30466 );
buf ( n30468 , n1439 );
nand ( n1441 , n1424 , n30468 );
not ( n1442 , n1441 );
nand ( n1443 , n29694 , n29829 );
nand ( n1444 , n1442 , n1443 );
not ( n1445 , n1444 );
or ( n1446 , n1421 , n1445 );
not ( n1447 , n1443 );
nand ( n1448 , n1447 , n1441 );
nand ( n1449 , n1446 , n1448 );
buf ( n30478 , n1449 );
xor ( n1451 , n30431 , n30478 );
xor ( n1452 , n30359 , n30384 );
xor ( n1453 , n1452 , n30408 );
buf ( n30482 , n1453 );
buf ( n30483 , n30482 );
and ( n1459 , n1451 , n30483 );
and ( n1460 , n30431 , n30478 );
or ( n1461 , n1459 , n1460 );
buf ( n30487 , n1461 );
nand ( n1463 , n30426 , n30487 );
nand ( n1464 , n1392 , n1463 );
not ( n1465 , n30345 );
not ( n1466 , n30422 );
nand ( n1467 , n1465 , n1466 );
and ( n30493 , n1464 , n1467 );
not ( n1469 , n30493 );
not ( n1470 , n30426 );
not ( n1471 , n30487 );
nand ( n1472 , n1470 , n1471 );
and ( n1473 , n1467 , n1472 );
buf ( n30499 , n29583 );
not ( n1475 , n30499 );
buf ( n30501 , n1342 );
not ( n1477 , n30501 );
or ( n1478 , n1475 , n1477 );
buf ( n30504 , n499 );
not ( n1480 , n30504 );
and ( n1481 , n456 , n471 );
not ( n1482 , n456 );
and ( n1483 , n1482 , n487 );
nor ( n1484 , n1481 , n1483 );
buf ( n30510 , n1484 );
not ( n1486 , n30510 );
or ( n1487 , n1480 , n1486 );
not ( n1488 , n1484 );
buf ( n30514 , n1488 );
buf ( n30515 , n29596 );
nand ( n1491 , n30514 , n30515 );
buf ( n30517 , n1491 );
buf ( n30518 , n30517 );
nand ( n1494 , n1487 , n30518 );
buf ( n30520 , n1494 );
buf ( n30521 , n30520 );
buf ( n30522 , n29624 );
nand ( n1498 , n30521 , n30522 );
buf ( n30524 , n1498 );
buf ( n30525 , n30524 );
nand ( n1501 , n1478 , n30525 );
buf ( n30527 , n1501 );
buf ( n30528 , n847 );
not ( n1504 , n30528 );
buf ( n30530 , n503 );
not ( n1506 , n30530 );
buf ( n30532 , n29492 );
not ( n1508 , n30532 );
or ( n1509 , n1506 , n1508 );
buf ( n30535 , n29819 );
buf ( n30536 , n863 );
nand ( n1512 , n30535 , n30536 );
buf ( n30538 , n1512 );
buf ( n30539 , n30538 );
nand ( n1515 , n1509 , n30539 );
buf ( n30541 , n1515 );
buf ( n30542 , n30541 );
not ( n1518 , n30542 );
or ( n1519 , n1504 , n1518 );
buf ( n30545 , n30464 );
buf ( n30546 , n504 );
nand ( n1522 , n30545 , n30546 );
buf ( n30548 , n1522 );
buf ( n30549 , n30548 );
nand ( n30550 , n1519 , n30549 );
buf ( n30551 , n30550 );
buf ( n30552 , n30551 );
buf ( n30553 , n29694 );
buf ( n30554 , n500 );
and ( n1530 , n30553 , n30554 );
buf ( n30556 , n29596 );
nor ( n1532 , n1530 , n30556 );
buf ( n30558 , n1532 );
buf ( n30559 , n30558 );
buf ( n30560 , n29764 );
buf ( n30561 , n500 );
or ( n1537 , n30560 , n30561 );
buf ( n30563 , n501 );
nand ( n1539 , n1537 , n30563 );
buf ( n30565 , n1539 );
buf ( n30566 , n30565 );
and ( n1542 , n30559 , n30566 );
buf ( n30568 , n1542 );
buf ( n30569 , n30568 );
and ( n1545 , n30552 , n30569 );
buf ( n30571 , n1545 );
xor ( n1547 , n30527 , n30571 );
xor ( n1548 , n1443 , n1441 );
xnor ( n1549 , n1548 , n1420 );
xor ( n1550 , n1547 , n1549 );
buf ( n30576 , n29583 );
not ( n1552 , n30576 );
buf ( n30578 , n30520 );
not ( n1554 , n30578 );
or ( n1555 , n1552 , n1554 );
buf ( n30581 , n29694 );
buf ( n30582 , n29596 );
nand ( n1558 , n30581 , n30582 );
buf ( n30584 , n1558 );
buf ( n30585 , n30584 );
not ( n1561 , n30585 );
buf ( n30587 , n29551 );
buf ( n30588 , n499 );
nand ( n1564 , n30587 , n30588 );
buf ( n30590 , n1564 );
buf ( n30591 , n30590 );
not ( n1567 , n30591 );
or ( n1568 , n1561 , n1567 );
buf ( n30594 , n29624 );
nand ( n1573 , n1568 , n30594 );
buf ( n30596 , n1573 );
buf ( n30597 , n30596 );
nand ( n1576 , n1555 , n30597 );
buf ( n30599 , n1576 );
buf ( n30600 , n30599 );
buf ( n30601 , n29737 );
not ( n1580 , n30601 );
buf ( n30603 , n1412 );
not ( n1582 , n30603 );
or ( n1583 , n1580 , n1582 );
buf ( n30606 , n501 );
not ( n1585 , n30606 );
buf ( n30608 , n1332 );
not ( n1587 , n30608 );
or ( n1588 , n1585 , n1587 );
buf ( n30611 , n901 );
buf ( n30612 , n29635 );
nand ( n1591 , n30611 , n30612 );
buf ( n30614 , n1591 );
buf ( n30615 , n30614 );
nand ( n1594 , n1588 , n30615 );
buf ( n30617 , n1594 );
buf ( n30618 , n30617 );
buf ( n30619 , n1355 );
nand ( n1598 , n30618 , n30619 );
buf ( n30621 , n1598 );
buf ( n30622 , n30621 );
nand ( n1604 , n1583 , n30622 );
buf ( n30624 , n1604 );
buf ( n30625 , n30624 );
xor ( n1607 , n30600 , n30625 );
xor ( n1608 , n30552 , n30569 );
buf ( n30628 , n1608 );
buf ( n30629 , n30628 );
and ( n1611 , n1607 , n30629 );
and ( n1612 , n30600 , n30625 );
or ( n1613 , n1611 , n1612 );
buf ( n30633 , n1613 );
nor ( n1615 , n1550 , n30633 );
xor ( n1616 , n30431 , n30478 );
xor ( n1617 , n1616 , n30483 );
buf ( n30637 , n1617 );
xor ( n1619 , n30527 , n30571 );
and ( n1620 , n1619 , n1549 );
and ( n1621 , n30527 , n30571 );
or ( n1622 , n1620 , n1621 );
nor ( n1623 , n30637 , n1622 );
nor ( n1624 , n1615 , n1623 );
not ( n1625 , n1624 );
buf ( n30645 , n29694 );
not ( n1627 , n29582 );
buf ( n30647 , n1627 );
and ( n30648 , n30645 , n30647 );
buf ( n30649 , n30648 );
buf ( n30650 , n30649 );
buf ( n30651 , n29737 );
not ( n1633 , n30651 );
buf ( n30653 , n30617 );
not ( n1635 , n30653 );
or ( n1636 , n1633 , n1635 );
buf ( n30656 , n501 );
not ( n1638 , n30656 );
buf ( n30658 , n1484 );
not ( n1640 , n30658 );
or ( n1641 , n1638 , n1640 );
buf ( n30661 , n1488 );
buf ( n30662 , n29635 );
nand ( n1644 , n30661 , n30662 );
buf ( n30664 , n1644 );
buf ( n30665 , n30664 );
nand ( n1647 , n1641 , n30665 );
buf ( n30667 , n1647 );
nand ( n1649 , n30667 , n1355 );
buf ( n30669 , n1649 );
nand ( n1651 , n1636 , n30669 );
buf ( n30671 , n1651 );
buf ( n30672 , n30671 );
xor ( n30673 , n30650 , n30672 );
buf ( n30674 , n504 );
not ( n1656 , n30674 );
buf ( n30676 , n30541 );
not ( n1658 , n30676 );
or ( n1659 , n1656 , n1658 );
buf ( n30679 , n503 );
not ( n1661 , n30679 );
buf ( n30681 , n29803 );
not ( n1663 , n30681 );
or ( n1664 , n1661 , n1663 );
buf ( n30684 , n1405 );
buf ( n30685 , n863 );
nand ( n1667 , n30684 , n30685 );
buf ( n30687 , n1667 );
buf ( n30688 , n30687 );
nand ( n1670 , n1664 , n30688 );
buf ( n30690 , n1670 );
buf ( n30691 , n30690 );
buf ( n30692 , n847 );
nand ( n1677 , n30691 , n30692 );
buf ( n30694 , n1677 );
buf ( n30695 , n30694 );
nand ( n1680 , n1659 , n30695 );
buf ( n30697 , n1680 );
buf ( n30698 , n30697 );
xor ( n1683 , n30673 , n30698 );
buf ( n30700 , n1683 );
not ( n1685 , n30700 );
buf ( n30702 , n29681 );
buf ( n30703 , n502 );
and ( n1688 , n30702 , n30703 );
buf ( n30705 , n29635 );
nor ( n1690 , n1688 , n30705 );
buf ( n30707 , n1690 );
buf ( n30708 , n30707 );
buf ( n30709 , n29694 );
buf ( n30710 , n502 );
or ( n1695 , n30709 , n30710 );
buf ( n30712 , n503 );
nand ( n1697 , n1695 , n30712 );
buf ( n30714 , n1697 );
buf ( n30715 , n30714 );
and ( n1700 , n30708 , n30715 );
buf ( n30717 , n1700 );
buf ( n30718 , n30717 );
buf ( n30719 , n504 );
not ( n1704 , n30719 );
buf ( n30721 , n30690 );
not ( n1706 , n30721 );
or ( n1707 , n1704 , n1706 );
buf ( n30724 , n503 );
not ( n1709 , n30724 );
buf ( n30726 , n1332 );
not ( n1711 , n30726 );
or ( n1712 , n1709 , n1711 );
buf ( n30729 , n901 );
buf ( n30730 , n863 );
nand ( n1715 , n30729 , n30730 );
buf ( n30732 , n1715 );
buf ( n30733 , n30732 );
nand ( n1718 , n1712 , n30733 );
buf ( n30735 , n1718 );
buf ( n30736 , n30735 );
buf ( n30737 , n847 );
nand ( n1722 , n30736 , n30737 );
buf ( n30739 , n1722 );
buf ( n30740 , n30739 );
nand ( n1725 , n1707 , n30740 );
buf ( n30742 , n1725 );
buf ( n30743 , n30742 );
and ( n1728 , n30718 , n30743 );
buf ( n30745 , n1728 );
not ( n1730 , n30745 );
nand ( n1731 , n1685 , n1730 );
not ( n1732 , n1731 );
xor ( n1733 , n30718 , n30743 );
buf ( n30750 , n1733 );
buf ( n30751 , n501 );
not ( n30752 , n30751 );
buf ( n30753 , n29551 );
not ( n1741 , n30753 );
or ( n1742 , n30752 , n1741 );
buf ( n30756 , n29681 );
buf ( n30757 , n29635 );
nand ( n1745 , n30756 , n30757 );
buf ( n30759 , n1745 );
buf ( n30760 , n30759 );
nand ( n1748 , n1742 , n30760 );
buf ( n30762 , n1748 );
not ( n1750 , n30762 );
not ( n1751 , n1355 );
or ( n30765 , n1750 , n1751 );
buf ( n30766 , n30667 );
buf ( n30767 , n29737 );
nand ( n1755 , n30766 , n30767 );
buf ( n30769 , n1755 );
nand ( n1757 , n30765 , n30769 );
nand ( n1758 , n30750 , n1757 );
or ( n1759 , n30750 , n1757 );
buf ( n30773 , n504 );
not ( n1761 , n30773 );
buf ( n30775 , n30735 );
not ( n1763 , n30775 );
or ( n1764 , n1761 , n1763 );
buf ( n30778 , n794 );
buf ( n30779 , n847 );
nand ( n1767 , n30778 , n30779 );
buf ( n30781 , n1767 );
buf ( n30782 , n30781 );
nand ( n1770 , n1764 , n30782 );
buf ( n30784 , n1770 );
not ( n1772 , n30784 );
not ( n1773 , n794 );
nor ( n1774 , n1773 , n29681 , n863 );
buf ( n30788 , n29737 );
not ( n1776 , n30788 );
buf ( n30790 , n29551 );
nor ( n1778 , n1776 , n30790 );
buf ( n30792 , n1778 );
nor ( n1780 , n1774 , n30792 );
nor ( n1781 , n1772 , n1780 );
nand ( n1782 , n1759 , n1781 );
nand ( n1783 , n1758 , n1782 );
not ( n1784 , n1783 );
or ( n1785 , n1732 , n1784 );
buf ( n1786 , n30700 );
nand ( n1787 , n1786 , n30745 );
nand ( n1788 , n1785 , n1787 );
xor ( n1789 , n30600 , n30625 );
xor ( n1790 , n1789 , n30629 );
buf ( n30804 , n1790 );
not ( n1792 , n30804 );
xor ( n1793 , n30650 , n30672 );
and ( n1794 , n1793 , n30698 );
and ( n1795 , n30650 , n30672 );
or ( n1796 , n1794 , n1795 );
buf ( n30810 , n1796 );
not ( n1798 , n30810 );
nand ( n1799 , n1792 , n1798 );
nand ( n1800 , n1788 , n1799 );
nand ( n1801 , n1550 , n30633 );
nand ( n1802 , n30804 , n30810 );
nand ( n1803 , n1800 , n1801 , n1802 );
not ( n1804 , n1803 );
or ( n1805 , n1625 , n1804 );
buf ( n1806 , n30637 );
nand ( n1807 , n1806 , n1622 );
nand ( n1808 , n1805 , n1807 );
nand ( n1809 , n1473 , n1808 );
nand ( n1810 , n1469 , n1809 );
not ( n1811 , n1810 );
or ( n1812 , n1305 , n1811 );
nand ( n1813 , n30232 , n30340 );
buf ( n1814 , n1813 );
nand ( n1815 , n1812 , n1814 );
not ( n1816 , n1815 );
or ( n30830 , n1189 , n1816 );
not ( n1818 , n1469 );
not ( n1819 , n1809 );
or ( n1820 , n1818 , n1819 );
nand ( n1821 , n1820 , n1304 );
and ( n1822 , n1187 , n1814 );
and ( n1823 , n1821 , n1822 );
nor ( n1824 , n1823 , n29516 );
nand ( n1825 , n30830 , n1824 );
not ( n30839 , n1825 );
buf ( n30840 , n520 );
buf ( n30841 , n502 );
or ( n1829 , n30840 , n30841 );
buf ( n30843 , n503 );
nand ( n1831 , n1829 , n30843 );
buf ( n30845 , n1831 );
buf ( n30846 , n30845 );
buf ( n30847 , n520 );
buf ( n30848 , n502 );
nand ( n1836 , n30847 , n30848 );
buf ( n30850 , n1836 );
buf ( n30851 , n30850 );
buf ( n30852 , n501 );
and ( n1840 , n30846 , n30851 , n30852 );
buf ( n30854 , n1840 );
buf ( n30855 , n30854 );
xor ( n1843 , n503 , n518 );
buf ( n30857 , n1843 );
not ( n1845 , n30857 );
not ( n1846 , n503 );
nor ( n1847 , n1846 , n504 );
buf ( n30861 , n1847 );
not ( n1849 , n30861 );
or ( n1850 , n1845 , n1849 );
buf ( n30864 , n517 );
buf ( n30865 , n503 );
xor ( n1853 , n30864 , n30865 );
buf ( n30867 , n1853 );
buf ( n30868 , n30867 );
buf ( n30869 , n504 );
nand ( n1857 , n30868 , n30869 );
buf ( n30871 , n1857 );
buf ( n30872 , n30871 );
nand ( n1860 , n1850 , n30872 );
buf ( n30874 , n1860 );
buf ( n30875 , n30874 );
and ( n1863 , n30855 , n30875 );
buf ( n30877 , n1863 );
xor ( n1865 , n500 , n501 );
buf ( n30879 , n1865 );
not ( n1870 , n30879 );
buf ( n30881 , n1870 );
buf ( n30882 , n30881 );
not ( n1873 , n30882 );
buf ( n30884 , n1873 );
buf ( n30885 , n30884 );
buf ( n30886 , n520 );
and ( n1877 , n30885 , n30886 );
buf ( n30888 , n1877 );
buf ( n30889 , n30867 );
not ( n1880 , n30889 );
and ( n1881 , n942 , n503 );
buf ( n30892 , n1881 );
not ( n1883 , n30892 );
or ( n1884 , n1880 , n1883 );
xor ( n1885 , n503 , n516 );
buf ( n30896 , n1885 );
buf ( n30897 , n504 );
nand ( n1888 , n30896 , n30897 );
buf ( n30899 , n1888 );
buf ( n30900 , n30899 );
nand ( n1891 , n1884 , n30900 );
buf ( n30902 , n1891 );
xor ( n1893 , n30888 , n30902 );
buf ( n30904 , n501 );
buf ( n30905 , n519 );
xor ( n1896 , n30904 , n30905 );
buf ( n30907 , n1896 );
not ( n1898 , n30907 );
buf ( n30909 , n501 );
buf ( n30910 , n502 );
xnor ( n30911 , n30909 , n30910 );
buf ( n30912 , n30911 );
not ( n1906 , n30912 );
xor ( n1907 , n502 , n503 );
not ( n1908 , n1907 );
nand ( n1909 , n1906 , n1908 );
buf ( n30917 , n1909 );
not ( n1911 , n30917 );
buf ( n30919 , n1911 );
not ( n1913 , n30919 );
or ( n1914 , n1898 , n1913 );
buf ( n1915 , n1907 );
buf ( n30923 , n1915 );
xor ( n1917 , n501 , n518 );
buf ( n30925 , n1917 );
nand ( n1919 , n30923 , n30925 );
buf ( n30927 , n1919 );
nand ( n1921 , n1914 , n30927 );
xor ( n1922 , n1893 , n1921 );
xor ( n1923 , n30877 , n1922 );
xor ( n1924 , n30855 , n30875 );
buf ( n30932 , n1924 );
buf ( n30933 , n501 );
buf ( n30934 , n520 );
xor ( n1928 , n30933 , n30934 );
buf ( n30936 , n1928 );
buf ( n30937 , n30936 );
not ( n1931 , n30937 );
buf ( n30939 , n30919 );
not ( n1933 , n30939 );
or ( n1934 , n1931 , n1933 );
buf ( n1935 , n1915 );
buf ( n30943 , n1935 );
buf ( n30944 , n30907 );
nand ( n1938 , n30943 , n30944 );
buf ( n30946 , n1938 );
buf ( n30947 , n30946 );
nand ( n1941 , n1934 , n30947 );
buf ( n30949 , n1941 );
or ( n1943 , n30932 , n30949 );
not ( n1944 , n519 );
buf ( n30952 , n1944 );
not ( n1946 , n30952 );
buf ( n30954 , n1847 );
not ( n1948 , n30954 );
or ( n1949 , n1946 , n1948 );
buf ( n30957 , n1843 );
buf ( n30958 , n504 );
nand ( n1952 , n30957 , n30958 );
buf ( n30960 , n1952 );
buf ( n30961 , n30960 );
nand ( n1955 , n1949 , n30961 );
buf ( n30963 , n1955 );
not ( n1957 , n30963 );
and ( n1958 , n520 , n1935 );
not ( n1959 , n520 );
not ( n1960 , n1881 );
nand ( n1961 , n1960 , n519 );
and ( n1962 , n1961 , n503 );
and ( n1963 , n1959 , n1962 );
nor ( n1964 , n1958 , n1963 );
nor ( n1965 , n1957 , n1964 );
nand ( n1966 , n1943 , n1965 );
nand ( n1967 , n30932 , n30949 );
nand ( n1968 , n1966 , n1967 );
and ( n1969 , n1923 , n1968 );
and ( n1970 , n30877 , n1922 );
or ( n1971 , n1969 , n1970 );
not ( n1972 , n1917 );
not ( n1973 , n30919 );
or ( n1974 , n1972 , n1973 );
buf ( n30982 , n1935 );
buf ( n30983 , n517 );
buf ( n30984 , n501 );
xor ( n30985 , n30983 , n30984 );
buf ( n30986 , n30985 );
buf ( n30987 , n30986 );
nand ( n1981 , n30982 , n30987 );
buf ( n30989 , n1981 );
nand ( n1983 , n1974 , n30989 );
buf ( n30991 , n499 );
buf ( n30992 , n520 );
xor ( n1986 , n30991 , n30992 );
buf ( n30994 , n1986 );
buf ( n30995 , n30994 );
not ( n30996 , n30995 );
not ( n1993 , n499 );
nor ( n1994 , n500 , n501 );
not ( n1995 , n1994 );
or ( n1996 , n1993 , n1995 );
not ( n1997 , n499 );
nand ( n1998 , n1997 , n500 , n501 );
nand ( n1999 , n1996 , n1998 );
not ( n2000 , n1999 );
not ( n2001 , n2000 );
buf ( n31006 , n2001 );
not ( n2003 , n31006 );
or ( n2004 , n30996 , n2003 );
buf ( n31009 , n30881 );
not ( n2006 , n31009 );
buf ( n31011 , n2006 );
buf ( n31012 , n31011 );
buf ( n31013 , n519 );
buf ( n31014 , n499 );
xor ( n2011 , n31013 , n31014 );
buf ( n31016 , n2011 );
buf ( n31017 , n31016 );
nand ( n2014 , n31012 , n31017 );
buf ( n31019 , n2014 );
buf ( n31020 , n31019 );
nand ( n2017 , n2004 , n31020 );
buf ( n31022 , n2017 );
xor ( n2019 , n1983 , n31022 );
xor ( n2020 , n503 , n515 );
not ( n2021 , n2020 );
not ( n2022 , n504 );
or ( n2023 , n2021 , n2022 );
nand ( n2024 , n1885 , n942 , n503 );
nand ( n2025 , n2023 , n2024 );
and ( n2026 , n520 , n500 );
nor ( n2027 , n2026 , n29596 );
or ( n2028 , n520 , n500 );
nand ( n2029 , n2028 , n501 );
and ( n2030 , n2027 , n2029 );
xor ( n2031 , n2025 , n2030 );
xor ( n2032 , n2019 , n2031 );
not ( n2033 , n2032 );
xor ( n2034 , n30888 , n30902 );
and ( n2035 , n2034 , n1921 );
and ( n2036 , n30888 , n30902 );
or ( n2037 , n2035 , n2036 );
not ( n2038 , n2037 );
nand ( n2039 , n2033 , n2038 );
nand ( n2040 , n1971 , n2039 );
xor ( n2041 , n1983 , n31022 );
and ( n2042 , n2041 , n2031 );
and ( n2043 , n1983 , n31022 );
or ( n2044 , n2042 , n2043 );
buf ( n31049 , n31016 );
not ( n2046 , n31049 );
buf ( n31051 , n2001 );
not ( n2048 , n31051 );
or ( n2049 , n2046 , n2048 );
buf ( n31054 , n31011 );
xor ( n2051 , n499 , n518 );
buf ( n31056 , n2051 );
nand ( n2053 , n31054 , n31056 );
buf ( n31058 , n2053 );
buf ( n31059 , n31058 );
nand ( n2056 , n2049 , n31059 );
buf ( n31061 , n2056 );
and ( n2058 , n2025 , n2030 );
not ( n31063 , n2058 );
xor ( n2063 , n31061 , n31063 );
buf ( n31065 , n30986 );
not ( n2065 , n31065 );
buf ( n31067 , n30919 );
not ( n2067 , n31067 );
or ( n2068 , n2065 , n2067 );
buf ( n31070 , n1935 );
buf ( n31071 , n516 );
buf ( n31072 , n501 );
xor ( n2072 , n31071 , n31072 );
buf ( n31074 , n2072 );
buf ( n31075 , n31074 );
nand ( n2075 , n31070 , n31075 );
buf ( n31077 , n2075 );
buf ( n31078 , n31077 );
nand ( n2078 , n2068 , n31078 );
buf ( n31080 , n2078 );
xor ( n2080 , n498 , n499 );
buf ( n2081 , n2080 );
buf ( n31083 , n2081 );
buf ( n31084 , n520 );
and ( n2084 , n31083 , n31084 );
buf ( n31086 , n2084 );
not ( n2086 , n31086 );
buf ( n31088 , n2020 );
not ( n2088 , n31088 );
buf ( n31090 , n1881 );
not ( n2090 , n31090 );
or ( n2091 , n2088 , n2090 );
xor ( n2092 , n503 , n514 );
buf ( n31094 , n2092 );
buf ( n31095 , n504 );
nand ( n2095 , n31094 , n31095 );
buf ( n31097 , n2095 );
buf ( n31098 , n31097 );
nand ( n2098 , n2091 , n31098 );
buf ( n31100 , n2098 );
not ( n2100 , n31100 );
and ( n2101 , n2086 , n2100 );
not ( n2102 , n2086 );
and ( n2103 , n2102 , n31100 );
nor ( n2104 , n2101 , n2103 );
xor ( n2105 , n31080 , n2104 );
xnor ( n2106 , n2063 , n2105 );
nand ( n2107 , n2044 , n2106 );
nand ( n2108 , n2032 , n2037 );
nand ( n2109 , n2040 , n2107 , n2108 );
not ( n2110 , n2109 );
buf ( n31112 , n520 );
buf ( n31113 , n498 );
or ( n2113 , n31112 , n31113 );
buf ( n31115 , n499 );
nand ( n2115 , n2113 , n31115 );
buf ( n31117 , n2115 );
buf ( n31118 , n31117 );
buf ( n31119 , n520 );
buf ( n31120 , n498 );
nand ( n2120 , n31119 , n31120 );
buf ( n31122 , n2120 );
buf ( n31123 , n31122 );
buf ( n31124 , n497 );
and ( n2124 , n31118 , n31123 , n31124 );
buf ( n31126 , n2124 );
not ( n2126 , n31126 );
not ( n2127 , n2126 );
not ( n2128 , n2092 );
not ( n2129 , n1881 );
or ( n2130 , n2128 , n2129 );
buf ( n31132 , n513 );
buf ( n31133 , n503 );
xor ( n2133 , n31132 , n31133 );
buf ( n31135 , n2133 );
buf ( n31136 , n31135 );
buf ( n31137 , n504 );
nand ( n2137 , n31136 , n31137 );
buf ( n31139 , n2137 );
nand ( n2139 , n2130 , n31139 );
not ( n2140 , n2139 );
or ( n2141 , n2127 , n2140 );
or ( n2142 , n2126 , n2139 );
nand ( n2143 , n2141 , n2142 );
buf ( n2144 , n2143 );
not ( n2145 , n2144 );
nand ( n2146 , n2100 , n2086 );
not ( n2147 , n2146 );
not ( n2148 , n31080 );
or ( n2149 , n2147 , n2148 );
nand ( n31151 , n31100 , n31086 );
nand ( n2151 , n2149 , n31151 );
not ( n2152 , n2151 );
not ( n2153 , n2152 );
or ( n2154 , n2145 , n2153 );
not ( n2155 , n2143 );
nand ( n2156 , n2155 , n2151 );
nand ( n2157 , n2154 , n2156 );
buf ( n31159 , n31074 );
not ( n2159 , n31159 );
nor ( n2160 , n30912 , n1907 );
buf ( n31162 , n2160 );
buf ( n2162 , n31162 );
buf ( n31164 , n2162 );
buf ( n31165 , n31164 );
not ( n2165 , n31165 );
or ( n2166 , n2159 , n2165 );
buf ( n31168 , n1915 );
buf ( n31169 , n515 );
buf ( n31170 , n501 );
xor ( n2170 , n31169 , n31170 );
buf ( n31172 , n2170 );
buf ( n31173 , n31172 );
nand ( n2173 , n31168 , n31173 );
buf ( n31175 , n2173 );
buf ( n31176 , n31175 );
nand ( n2176 , n2166 , n31176 );
buf ( n31178 , n2176 );
buf ( n31179 , n31178 );
buf ( n31180 , n2051 );
not ( n2180 , n31180 );
buf ( n31182 , n2001 );
not ( n2182 , n31182 );
or ( n31184 , n2180 , n2182 );
buf ( n31185 , n31011 );
buf ( n31186 , n517 );
buf ( n31187 , n499 );
xor ( n2187 , n31186 , n31187 );
buf ( n31189 , n2187 );
buf ( n31190 , n31189 );
nand ( n2190 , n31185 , n31190 );
buf ( n31192 , n2190 );
buf ( n31193 , n31192 );
nand ( n2193 , n31184 , n31193 );
buf ( n31195 , n2193 );
buf ( n31196 , n31195 );
xor ( n2196 , n31179 , n31196 );
buf ( n31198 , n520 );
buf ( n31199 , n497 );
xor ( n2199 , n31198 , n31199 );
buf ( n31201 , n2199 );
buf ( n31202 , n31201 );
not ( n2202 , n31202 );
not ( n2206 , n497 );
nor ( n31205 , n498 , n499 );
not ( n2208 , n31205 );
or ( n2209 , n2206 , n2208 );
not ( n2210 , n497 );
nand ( n2211 , n2210 , n498 , n499 );
nand ( n2212 , n2209 , n2211 );
buf ( n2213 , n2212 );
buf ( n31212 , n2213 );
not ( n2215 , n31212 );
or ( n2216 , n2202 , n2215 );
buf ( n31215 , n519 );
buf ( n31216 , n497 );
xnor ( n2219 , n31215 , n31216 );
buf ( n31218 , n2219 );
buf ( n31219 , n31218 );
not ( n2222 , n31219 );
buf ( n31221 , n2081 );
nand ( n2224 , n2222 , n31221 );
buf ( n31223 , n2224 );
buf ( n31224 , n31223 );
nand ( n2227 , n2216 , n31224 );
buf ( n31226 , n2227 );
buf ( n31227 , n31226 );
xor ( n2230 , n2196 , n31227 );
buf ( n31229 , n2230 );
and ( n2232 , n2157 , n31229 );
not ( n2233 , n2157 );
not ( n2234 , n31229 );
and ( n2235 , n2233 , n2234 );
nor ( n2236 , n2232 , n2235 );
not ( n2237 , n31061 );
nand ( n2238 , n2237 , n31063 );
not ( n2239 , n2238 );
not ( n2240 , n2105 );
or ( n2241 , n2239 , n2240 );
nand ( n2242 , n31061 , n2058 );
nand ( n31241 , n2241 , n2242 );
nor ( n2247 , n2236 , n31241 );
nor ( n2248 , n2106 , n2044 );
nor ( n2249 , n2247 , n2248 );
not ( n2250 , n2249 );
or ( n2251 , n2110 , n2250 );
nand ( n2252 , n2236 , n31241 );
nand ( n2253 , n2251 , n2252 );
not ( n2254 , n2253 );
or ( n2255 , n2151 , n2144 );
not ( n2256 , n2255 );
not ( n2257 , n31229 );
or ( n2258 , n2256 , n2257 );
nand ( n2259 , n2144 , n2151 );
nand ( n2260 , n2258 , n2259 );
not ( n2261 , n2260 );
not ( n2262 , n2261 );
buf ( n31258 , n512 );
buf ( n31259 , n503 );
xor ( n2265 , n31258 , n31259 );
buf ( n31261 , n2265 );
not ( n2267 , n31261 );
not ( n2268 , n504 );
or ( n2269 , n2267 , n2268 );
nand ( n2270 , n31135 , n1881 );
nand ( n2271 , n2269 , n2270 );
buf ( n31267 , n2271 );
buf ( n31268 , n496 );
buf ( n31269 , n497 );
xor ( n2275 , n31268 , n31269 );
buf ( n31271 , n2275 );
buf ( n31272 , n31271 );
buf ( n31273 , n520 );
and ( n2279 , n31272 , n31273 );
buf ( n31275 , n2279 );
buf ( n31276 , n31275 );
xor ( n2282 , n31267 , n31276 );
buf ( n31278 , n2213 );
not ( n2284 , n31278 );
buf ( n31280 , n2284 );
buf ( n31281 , n31280 );
buf ( n31282 , n31218 );
or ( n2288 , n31281 , n31282 );
buf ( n31284 , n2081 );
not ( n2290 , n31284 );
buf ( n31286 , n2290 );
buf ( n31287 , n31286 );
buf ( n31288 , n518 );
buf ( n31289 , n497 );
xor ( n2295 , n31288 , n31289 );
buf ( n31291 , n2295 );
buf ( n31292 , n31291 );
not ( n2298 , n31292 );
buf ( n31294 , n2298 );
buf ( n31295 , n31294 );
or ( n2301 , n31287 , n31295 );
nand ( n2302 , n2288 , n2301 );
buf ( n31298 , n2302 );
buf ( n31299 , n31298 );
xor ( n2305 , n2282 , n31299 );
buf ( n31301 , n2305 );
buf ( n31302 , n31301 );
xor ( n2308 , n31179 , n31196 );
and ( n2309 , n2308 , n31227 );
and ( n2310 , n31179 , n31196 );
or ( n2311 , n2309 , n2310 );
buf ( n31307 , n2311 );
buf ( n31308 , n31307 );
xor ( n2314 , n31302 , n31308 );
buf ( n31310 , n31189 );
not ( n2316 , n31310 );
buf ( n31312 , n2001 );
not ( n2318 , n31312 );
or ( n2319 , n2316 , n2318 );
buf ( n31315 , n30884 );
buf ( n31316 , n516 );
buf ( n31317 , n499 );
xor ( n2323 , n31316 , n31317 );
buf ( n31319 , n2323 );
buf ( n31320 , n31319 );
nand ( n2326 , n31315 , n31320 );
buf ( n31322 , n2326 );
buf ( n31323 , n31322 );
nand ( n2329 , n2319 , n31323 );
buf ( n31325 , n2329 );
not ( n2331 , n31325 );
nand ( n2332 , n2139 , n31126 );
not ( n2333 , n2332 );
and ( n2334 , n2331 , n2333 );
not ( n2335 , n2331 );
and ( n2336 , n2335 , n2332 );
nor ( n2337 , n2334 , n2336 );
buf ( n31333 , n31172 );
not ( n2339 , n31333 );
buf ( n31335 , n30919 );
not ( n2341 , n31335 );
or ( n2342 , n2339 , n2341 );
buf ( n31338 , n1935 );
buf ( n31339 , n514 );
buf ( n31340 , n501 );
xor ( n2346 , n31339 , n31340 );
buf ( n31342 , n2346 );
buf ( n31343 , n31342 );
nand ( n2349 , n31338 , n31343 );
buf ( n31345 , n2349 );
buf ( n31346 , n31345 );
nand ( n2352 , n2342 , n31346 );
buf ( n31348 , n2352 );
not ( n2354 , n31348 );
and ( n2355 , n2337 , n2354 );
not ( n2356 , n2337 );
and ( n2357 , n2356 , n31348 );
nor ( n2358 , n2355 , n2357 );
buf ( n31354 , n2358 );
xor ( n2360 , n2314 , n31354 );
buf ( n31356 , n2360 );
not ( n2362 , n31356 );
not ( n2363 , n2362 );
or ( n2364 , n2262 , n2363 );
xor ( n2365 , n31302 , n31308 );
and ( n2366 , n2365 , n31354 );
and ( n2367 , n31302 , n31308 );
or ( n2368 , n2366 , n2367 );
buf ( n31364 , n2368 );
not ( n2370 , n31364 );
nand ( n2371 , n2332 , n2331 );
not ( n2372 , n2371 );
not ( n2373 , n31348 );
or ( n2374 , n2372 , n2373 );
nand ( n2375 , n2333 , n31325 );
nand ( n2376 , n2374 , n2375 );
buf ( n31372 , n31261 );
not ( n2378 , n31372 );
buf ( n31374 , n1847 );
not ( n2380 , n31374 );
or ( n2381 , n2378 , n2380 );
buf ( n31377 , n511 );
buf ( n31378 , n503 );
xor ( n2384 , n31377 , n31378 );
buf ( n31380 , n2384 );
buf ( n31381 , n31380 );
buf ( n31382 , n504 );
nand ( n2388 , n31381 , n31382 );
buf ( n31384 , n2388 );
buf ( n31385 , n31384 );
nand ( n2391 , n2381 , n31385 );
buf ( n31387 , n2391 );
buf ( n31388 , n31387 );
buf ( n31389 , n520 );
buf ( n31390 , n495 );
xor ( n2396 , n31389 , n31390 );
buf ( n31392 , n2396 );
buf ( n31393 , n31392 );
not ( n2399 , n31393 );
nand ( n2400 , n758 , n496 );
not ( n2401 , n2400 );
not ( n2402 , n496 );
nand ( n2403 , n2402 , n495 );
not ( n2404 , n2403 );
or ( n31400 , n2401 , n2404 );
xnor ( n2409 , n496 , n497 );
nand ( n2410 , n31400 , n2409 );
buf ( n2411 , n2410 );
not ( n2412 , n2411 );
buf ( n31405 , n2412 );
not ( n2414 , n31405 );
or ( n2415 , n2399 , n2414 );
buf ( n31408 , n31271 );
buf ( n31409 , n519 );
buf ( n31410 , n495 );
xor ( n2419 , n31409 , n31410 );
buf ( n31412 , n2419 );
buf ( n31413 , n31412 );
nand ( n2422 , n31408 , n31413 );
buf ( n31415 , n2422 );
buf ( n31416 , n31415 );
nand ( n2425 , n2415 , n31416 );
buf ( n31418 , n2425 );
buf ( n31419 , n31418 );
xor ( n2428 , n31388 , n31419 );
buf ( n31421 , n31291 );
not ( n2430 , n31421 );
buf ( n31423 , n2213 );
not ( n2432 , n31423 );
or ( n2433 , n2430 , n2432 );
buf ( n31426 , n2081 );
buf ( n31427 , n517 );
buf ( n31428 , n497 );
xor ( n2437 , n31427 , n31428 );
buf ( n31430 , n2437 );
buf ( n31431 , n31430 );
nand ( n2440 , n31426 , n31431 );
buf ( n31433 , n2440 );
buf ( n31434 , n31433 );
nand ( n2443 , n2433 , n31434 );
buf ( n31436 , n2443 );
buf ( n31437 , n31436 );
xor ( n2446 , n2428 , n31437 );
buf ( n31439 , n2446 );
not ( n2448 , n31439 );
and ( n2449 , n2376 , n2448 );
not ( n2450 , n2376 );
and ( n2451 , n2450 , n31439 );
nor ( n2452 , n2449 , n2451 );
not ( n2453 , n2452 );
buf ( n31446 , n31319 );
not ( n2455 , n31446 );
buf ( n31448 , n2001 );
not ( n2457 , n31448 );
or ( n2458 , n2455 , n2457 );
buf ( n31451 , n30884 );
buf ( n31452 , n515 );
buf ( n31453 , n499 );
xor ( n2462 , n31452 , n31453 );
buf ( n31455 , n2462 );
buf ( n31456 , n31455 );
nand ( n2465 , n31451 , n31456 );
buf ( n31458 , n2465 );
buf ( n31459 , n31458 );
nand ( n2468 , n2458 , n31459 );
buf ( n31461 , n2468 );
buf ( n31462 , n31461 );
buf ( n31463 , n520 );
buf ( n31464 , n496 );
or ( n2473 , n31463 , n31464 );
buf ( n31466 , n497 );
nand ( n2475 , n2473 , n31466 );
buf ( n31468 , n2475 );
buf ( n31469 , n520 );
buf ( n31470 , n496 );
nand ( n2479 , n31469 , n31470 );
buf ( n31472 , n2479 );
and ( n2481 , n31468 , n31472 , n495 );
not ( n2482 , n31342 );
not ( n2483 , n30919 );
or ( n2484 , n2482 , n2483 );
buf ( n31477 , n1915 );
buf ( n31478 , n513 );
buf ( n31479 , n501 );
xor ( n31480 , n31478 , n31479 );
buf ( n31481 , n31480 );
buf ( n31482 , n31481 );
nand ( n2491 , n31477 , n31482 );
buf ( n31484 , n2491 );
nand ( n2493 , n2484 , n31484 );
xor ( n2494 , n2481 , n2493 );
buf ( n31487 , n2494 );
xor ( n2496 , n31462 , n31487 );
xor ( n2497 , n31267 , n31276 );
and ( n2498 , n2497 , n31299 );
and ( n2499 , n31267 , n31276 );
or ( n2500 , n2498 , n2499 );
buf ( n31493 , n2500 );
buf ( n31494 , n31493 );
xor ( n2503 , n2496 , n31494 );
buf ( n31496 , n2503 );
not ( n2505 , n31496 );
nand ( n2506 , n2453 , n2505 );
nand ( n2507 , n2452 , n31496 );
nand ( n2508 , n2370 , n2506 , n2507 );
nand ( n2509 , n2364 , n2508 );
not ( n2510 , n2509 );
not ( n2511 , n2510 );
or ( n2512 , n2254 , n2511 );
nand ( n2513 , n31356 , n2260 );
not ( n2514 , n2513 );
not ( n2515 , n2505 );
not ( n2516 , n2453 );
or ( n2517 , n2515 , n2516 );
nand ( n2518 , n2517 , n2507 );
nand ( n2519 , n31364 , n2518 );
not ( n2520 , n2519 );
or ( n2521 , n2514 , n2520 );
not ( n2522 , n2518 );
not ( n2523 , n31364 );
nand ( n2524 , n2522 , n2523 );
nand ( n2525 , n2521 , n2524 );
nand ( n2526 , n2512 , n2525 );
buf ( n31519 , n31380 );
not ( n2528 , n31519 );
buf ( n31521 , n1847 );
not ( n2530 , n31521 );
or ( n2531 , n2528 , n2530 );
buf ( n31524 , n510 );
buf ( n31525 , n503 );
xor ( n2534 , n31524 , n31525 );
buf ( n31527 , n2534 );
buf ( n31528 , n31527 );
buf ( n31529 , n504 );
nand ( n2538 , n31528 , n31529 );
buf ( n31531 , n2538 );
buf ( n31532 , n31531 );
nand ( n2541 , n2531 , n31532 );
buf ( n31534 , n2541 );
buf ( n31535 , n31534 );
buf ( n31536 , n31455 );
not ( n2545 , n31536 );
buf ( n31538 , n2001 );
not ( n2547 , n31538 );
or ( n2548 , n2545 , n2547 );
buf ( n31541 , n31011 );
buf ( n31542 , n514 );
buf ( n31543 , n499 );
xor ( n2552 , n31542 , n31543 );
buf ( n31545 , n2552 );
buf ( n31546 , n31545 );
nand ( n2555 , n31541 , n31546 );
buf ( n31548 , n2555 );
buf ( n31549 , n31548 );
nand ( n2558 , n2548 , n31549 );
buf ( n31551 , n2558 );
buf ( n31552 , n31551 );
xor ( n2561 , n31535 , n31552 );
not ( n2562 , n31271 );
xor ( n2563 , n495 , n518 );
not ( n2564 , n2563 );
or ( n2565 , n2562 , n2564 );
buf ( n31558 , n31412 );
not ( n2567 , n31558 );
buf ( n31560 , n2567 );
or ( n31561 , n31560 , n2411 );
nand ( n2573 , n2565 , n31561 );
buf ( n31563 , n2573 );
xor ( n2575 , n2561 , n31563 );
buf ( n31565 , n2575 );
not ( n2577 , n31565 );
not ( n2578 , n2577 );
xor ( n2579 , n31462 , n31487 );
and ( n2580 , n2579 , n31494 );
and ( n2581 , n31462 , n31487 );
or ( n2582 , n2580 , n2581 );
buf ( n31572 , n2582 );
not ( n2584 , n31572 );
not ( n2585 , n2584 );
or ( n2586 , n2578 , n2585 );
nand ( n2587 , n31572 , n31565 );
nand ( n2588 , n2586 , n2587 );
and ( n2589 , n2481 , n2493 );
xor ( n2590 , n494 , n495 );
buf ( n2591 , n2590 );
buf ( n31581 , n2591 );
buf ( n31582 , n520 );
and ( n2594 , n31581 , n31582 );
buf ( n31584 , n2594 );
buf ( n31585 , n31430 );
not ( n2597 , n31585 );
buf ( n31587 , n2213 );
not ( n2599 , n31587 );
or ( n2600 , n2597 , n2599 );
buf ( n31590 , n2081 );
buf ( n31591 , n516 );
buf ( n31592 , n497 );
xor ( n2604 , n31591 , n31592 );
buf ( n31594 , n2604 );
buf ( n31595 , n31594 );
nand ( n2607 , n31590 , n31595 );
buf ( n31597 , n2607 );
buf ( n31598 , n31597 );
nand ( n2610 , n2600 , n31598 );
buf ( n31600 , n2610 );
xor ( n2612 , n31584 , n31600 );
buf ( n31602 , n31481 );
not ( n2614 , n31602 );
buf ( n31604 , n31164 );
not ( n2616 , n31604 );
or ( n2617 , n2614 , n2616 );
buf ( n31607 , n1915 );
buf ( n31608 , n512 );
buf ( n31609 , n501 );
xor ( n2621 , n31608 , n31609 );
buf ( n31611 , n2621 );
buf ( n31612 , n31611 );
nand ( n2624 , n31607 , n31612 );
buf ( n31614 , n2624 );
buf ( n31615 , n31614 );
nand ( n2627 , n2617 , n31615 );
buf ( n31617 , n2627 );
xor ( n2629 , n2612 , n31617 );
xor ( n2630 , n2589 , n2629 );
xor ( n2631 , n31388 , n31419 );
and ( n2632 , n2631 , n31437 );
and ( n2633 , n31388 , n31419 );
or ( n2634 , n2632 , n2633 );
buf ( n31624 , n2634 );
xor ( n2636 , n2630 , n31624 );
not ( n2637 , n2636 );
and ( n2638 , n2588 , n2637 );
not ( n2639 , n2588 );
and ( n2640 , n2639 , n2636 );
nor ( n2641 , n2638 , n2640 );
not ( n2642 , n2641 );
buf ( n2643 , n2448 );
not ( n2644 , n2643 );
not ( n2645 , n2505 );
or ( n2646 , n2644 , n2645 );
nand ( n2647 , n2646 , n2376 );
not ( n2648 , n2643 );
nand ( n2649 , n2648 , n31496 );
nand ( n2650 , n2647 , n2649 );
not ( n31640 , n2650 );
nand ( n2652 , n2642 , n31640 );
nand ( n2653 , n2526 , n2652 );
nand ( n2654 , n2650 , n2641 );
and ( n2655 , n2653 , n2654 );
buf ( n31645 , n520 );
buf ( n31646 , n493 );
xor ( n2658 , n31645 , n31646 );
buf ( n31648 , n2658 );
buf ( n31649 , n31648 );
not ( n2661 , n31649 );
not ( n2662 , n2590 );
and ( n2663 , n493 , n494 );
not ( n2664 , n493 );
and ( n2665 , n2664 , n29568 );
nor ( n2666 , n2663 , n2665 );
nand ( n2667 , n2662 , n2666 );
not ( n2668 , n2667 );
buf ( n31658 , n2668 );
buf ( n2670 , n31658 );
buf ( n31660 , n2670 );
buf ( n31661 , n31660 );
not ( n2673 , n31661 );
or ( n2674 , n2661 , n2673 );
buf ( n31664 , n2591 );
xor ( n2676 , n493 , n519 );
buf ( n31666 , n2676 );
nand ( n2678 , n31664 , n31666 );
buf ( n31668 , n2678 );
buf ( n31669 , n31668 );
nand ( n2681 , n2674 , n31669 );
buf ( n31671 , n2681 );
buf ( n31672 , n31671 );
buf ( n31673 , n31545 );
not ( n2685 , n31673 );
buf ( n31675 , n2001 );
not ( n2687 , n31675 );
or ( n2688 , n2685 , n2687 );
buf ( n31678 , n31011 );
buf ( n31679 , n499 );
buf ( n31680 , n513 );
xor ( n2692 , n31679 , n31680 );
buf ( n31682 , n2692 );
buf ( n31683 , n31682 );
nand ( n2695 , n31678 , n31683 );
buf ( n31685 , n2695 );
buf ( n31686 , n31685 );
nand ( n2698 , n2688 , n31686 );
buf ( n31688 , n2698 );
buf ( n31689 , n31688 );
xor ( n2701 , n31672 , n31689 );
buf ( n31691 , n520 );
buf ( n31692 , n494 );
or ( n2704 , n31691 , n31692 );
buf ( n31694 , n495 );
nand ( n2706 , n2704 , n31694 );
buf ( n31696 , n2706 );
buf ( n31697 , n31696 );
buf ( n31698 , n520 );
buf ( n31699 , n494 );
nand ( n2711 , n31698 , n31699 );
buf ( n31701 , n2711 );
buf ( n31702 , n31701 );
buf ( n31703 , n493 );
and ( n2715 , n31697 , n31702 , n31703 );
buf ( n31705 , n2715 );
buf ( n31706 , n31705 );
buf ( n31707 , n31611 );
not ( n2719 , n31707 );
buf ( n31709 , n31164 );
not ( n2721 , n31709 );
or ( n2722 , n2719 , n2721 );
buf ( n31712 , n1915 );
xor ( n2724 , n501 , n511 );
buf ( n31714 , n2724 );
nand ( n2726 , n31712 , n31714 );
buf ( n31716 , n2726 );
buf ( n31717 , n31716 );
nand ( n2729 , n2722 , n31717 );
buf ( n31719 , n2729 );
buf ( n31720 , n31719 );
xor ( n2732 , n31706 , n31720 );
buf ( n31722 , n2732 );
buf ( n31723 , n31722 );
xor ( n2738 , n2701 , n31723 );
buf ( n31725 , n2738 );
xor ( n2740 , n2589 , n2629 );
and ( n2741 , n2740 , n31624 );
and ( n2742 , n2589 , n2629 );
or ( n2743 , n2741 , n2742 );
xor ( n2744 , n31725 , n2743 );
xor ( n2745 , n31584 , n31600 );
and ( n2746 , n2745 , n31617 );
and ( n2747 , n31584 , n31600 );
or ( n2748 , n2746 , n2747 );
xor ( n2749 , n31535 , n31552 );
and ( n2750 , n2749 , n31563 );
and ( n2751 , n31535 , n31552 );
or ( n2752 , n2750 , n2751 );
buf ( n31739 , n2752 );
xor ( n2754 , n2748 , n31739 );
buf ( n31741 , n31527 );
not ( n2756 , n31741 );
buf ( n31743 , n1847 );
not ( n2758 , n31743 );
or ( n2759 , n2756 , n2758 );
xor ( n2760 , n503 , n509 );
buf ( n31747 , n2760 );
buf ( n31748 , n504 );
nand ( n2763 , n31747 , n31748 );
buf ( n31750 , n2763 );
buf ( n31751 , n31750 );
nand ( n2766 , n2759 , n31751 );
buf ( n31753 , n2766 );
buf ( n31754 , n31594 );
not ( n2769 , n31754 );
buf ( n31756 , n2213 );
not ( n2771 , n31756 );
or ( n2772 , n2769 , n2771 );
buf ( n31759 , n2081 );
xor ( n2774 , n497 , n515 );
buf ( n31761 , n2774 );
nand ( n2776 , n31759 , n31761 );
buf ( n31763 , n2776 );
buf ( n31764 , n31763 );
nand ( n2779 , n2772 , n31764 );
buf ( n31766 , n2779 );
not ( n2781 , n31766 );
xor ( n2782 , n31753 , n2781 );
buf ( n31769 , n2563 );
not ( n2784 , n31769 );
buf ( n31771 , n2412 );
not ( n2786 , n31771 );
or ( n2787 , n2784 , n2786 );
buf ( n31774 , n31271 );
buf ( n31775 , n517 );
buf ( n31776 , n495 );
xor ( n2791 , n31775 , n31776 );
buf ( n31778 , n2791 );
buf ( n31779 , n31778 );
nand ( n2794 , n31774 , n31779 );
buf ( n31781 , n2794 );
buf ( n31782 , n31781 );
nand ( n2797 , n2787 , n31782 );
buf ( n31784 , n2797 );
xnor ( n2799 , n2782 , n31784 );
xor ( n2800 , n2754 , n2799 );
xor ( n2801 , n2744 , n2800 );
not ( n2802 , n31565 );
not ( n2803 , n31572 );
or ( n2804 , n2802 , n2803 );
not ( n2805 , n2577 );
not ( n2806 , n2584 );
or ( n2807 , n2805 , n2806 );
nand ( n2808 , n2807 , n2636 );
nand ( n2809 , n2804 , n2808 );
nand ( n2810 , n2801 , n2809 );
not ( n2811 , n2801 );
not ( n31798 , n2809 );
nand ( n2813 , n2811 , n31798 );
nand ( n2814 , n2810 , n2813 );
not ( n2815 , n455 );
nand ( n2816 , n2814 , n2815 );
nor ( n2817 , n2655 , n2816 );
nand ( n2818 , n2815 , n2654 );
nor ( n2819 , n2814 , n2818 );
and ( n2820 , n2653 , n2819 );
nor ( n2821 , n2817 , n2820 );
not ( n2822 , n2821 );
or ( n2823 , n30839 , n2822 );
nand ( n2824 , n2823 , n454 );
buf ( n31811 , n467 );
buf ( n31812 , n536 );
buf ( n31813 , n548 );
or ( n2828 , n31812 , n31813 );
buf ( n31815 , n549 );
nand ( n2830 , n2828 , n31815 );
buf ( n31817 , n2830 );
buf ( n31818 , n31817 );
buf ( n31819 , n536 );
buf ( n31820 , n548 );
nand ( n2835 , n31819 , n31820 );
buf ( n31822 , n2835 );
buf ( n31823 , n31822 );
buf ( n31824 , n547 );
and ( n2839 , n31818 , n31823 , n31824 );
buf ( n31826 , n2839 );
buf ( n31827 , n31826 );
and ( n2842 , n31811 , n31827 );
buf ( n31829 , n2842 );
buf ( n31830 , n31829 );
not ( n2845 , n552 );
nand ( n2846 , n2845 , n551 );
buf ( n31833 , n2846 );
not ( n2848 , n551 );
buf ( n31835 , n2848 );
buf ( n31836 , n531 );
and ( n2851 , n31835 , n31836 );
buf ( n31838 , n531 );
not ( n2853 , n31838 );
buf ( n31840 , n2853 );
buf ( n31841 , n31840 );
buf ( n31842 , n551 );
and ( n2857 , n31841 , n31842 );
nor ( n2858 , n2851 , n2857 );
buf ( n31845 , n2858 );
buf ( n31846 , n31845 );
or ( n2861 , n31833 , n31846 );
buf ( n31848 , n2848 );
buf ( n31849 , n530 );
and ( n2864 , n31848 , n31849 );
buf ( n31851 , n530 );
not ( n2866 , n31851 );
buf ( n31853 , n2866 );
buf ( n31854 , n31853 );
buf ( n31855 , n551 );
and ( n2870 , n31854 , n31855 );
nor ( n2871 , n2864 , n2870 );
buf ( n31858 , n2871 );
buf ( n31859 , n31858 );
buf ( n31860 , n2845 );
or ( n2875 , n31859 , n31860 );
nand ( n2876 , n2861 , n2875 );
buf ( n31863 , n2876 );
buf ( n31864 , n31863 );
xor ( n2879 , n31830 , n31864 );
buf ( n31866 , n549 );
not ( n2881 , n31866 );
buf ( n31868 , n2881 );
buf ( n31869 , n31868 );
buf ( n31870 , n533 );
and ( n2885 , n31869 , n31870 );
buf ( n31872 , n533 );
not ( n2887 , n31872 );
buf ( n31874 , n2887 );
buf ( n31875 , n31874 );
buf ( n31876 , n549 );
and ( n2894 , n31875 , n31876 );
nor ( n2895 , n2885 , n2894 );
buf ( n31879 , n2895 );
buf ( n31880 , n31879 );
not ( n2898 , n31880 );
buf ( n31882 , n2898 );
buf ( n31883 , n31882 );
not ( n2901 , n31883 );
xor ( n2902 , n549 , n550 );
not ( n2903 , n2848 );
buf ( n31887 , n550 );
not ( n2905 , n31887 );
buf ( n31889 , n2905 );
not ( n2907 , n31889 );
or ( n2908 , n2903 , n2907 );
nand ( n2909 , n550 , n551 );
nand ( n2910 , n2908 , n2909 );
nand ( n2911 , n2902 , n2910 );
buf ( n31895 , n2911 );
not ( n2913 , n31895 );
buf ( n31897 , n2913 );
buf ( n31898 , n31897 );
not ( n2916 , n31898 );
or ( n2917 , n2901 , n2916 );
xnor ( n2918 , n550 , n551 );
buf ( n31902 , n2918 );
buf ( n31903 , n31868 );
buf ( n31904 , n532 );
and ( n2922 , n31903 , n31904 );
buf ( n31906 , n532 );
not ( n2924 , n31906 );
buf ( n31908 , n2924 );
buf ( n31909 , n31908 );
buf ( n31910 , n549 );
and ( n2928 , n31909 , n31910 );
nor ( n2929 , n2922 , n2928 );
buf ( n31913 , n2929 );
buf ( n31914 , n31913 );
or ( n2932 , n31902 , n31914 );
nand ( n2933 , n2917 , n2932 );
buf ( n31917 , n2933 );
buf ( n31918 , n31917 );
and ( n2936 , n2879 , n31918 );
and ( n2937 , n31830 , n31864 );
or ( n2938 , n2936 , n2937 );
buf ( n31922 , n2938 );
buf ( n31923 , n31922 );
buf ( n31924 , n465 );
buf ( n31925 , n536 );
buf ( n31926 , n546 );
or ( n2944 , n31925 , n31926 );
buf ( n31928 , n547 );
nand ( n2946 , n2944 , n31928 );
buf ( n31930 , n2946 );
buf ( n31931 , n31930 );
buf ( n31932 , n536 );
buf ( n31933 , n546 );
nand ( n2951 , n31932 , n31933 );
buf ( n31935 , n2951 );
buf ( n31936 , n31935 );
buf ( n31937 , n545 );
and ( n2955 , n31931 , n31936 , n31937 );
buf ( n31939 , n2955 );
buf ( n31940 , n31939 );
xor ( n2958 , n31924 , n31940 );
buf ( n31942 , n2958 );
buf ( n31943 , n31942 );
not ( n2961 , n2846 );
not ( n2962 , n2961 );
buf ( n31946 , n2962 );
buf ( n31947 , n31858 );
or ( n31948 , n31946 , n31947 );
buf ( n31949 , n2848 );
buf ( n31950 , n529 );
and ( n2968 , n31949 , n31950 );
not ( n2969 , n529 );
buf ( n31953 , n2969 );
buf ( n31954 , n551 );
and ( n2972 , n31953 , n31954 );
nor ( n2973 , n2968 , n2972 );
buf ( n31957 , n2973 );
buf ( n31958 , n31957 );
buf ( n31959 , n2845 );
or ( n2977 , n31958 , n31959 );
nand ( n2978 , n31948 , n2977 );
buf ( n31962 , n2978 );
buf ( n31963 , n31962 );
xor ( n2981 , n31943 , n31963 );
buf ( n31965 , n547 );
buf ( n31966 , n533 );
and ( n2984 , n31965 , n31966 );
not ( n2985 , n31965 );
buf ( n31969 , n31874 );
and ( n2987 , n2985 , n31969 );
nor ( n2988 , n2984 , n2987 );
buf ( n31972 , n2988 );
buf ( n31973 , n31972 );
not ( n2991 , n31973 );
buf ( n31975 , n548 );
buf ( n31976 , n549 );
xnor ( n2994 , n31975 , n31976 );
buf ( n31978 , n2994 );
buf ( n31979 , n31978 );
not ( n2997 , n31979 );
buf ( n31981 , n2997 );
buf ( n31982 , n31981 );
not ( n3000 , n31982 );
or ( n3001 , n2991 , n3000 );
buf ( n31985 , n548 );
buf ( n31986 , n549 );
xnor ( n3004 , n31985 , n31986 );
buf ( n31988 , n3004 );
buf ( n31989 , n31988 );
buf ( n31990 , n547 );
not ( n3008 , n31990 );
buf ( n31992 , n548 );
not ( n3010 , n31992 );
and ( n3011 , n3008 , n3010 );
buf ( n31995 , n547 );
buf ( n31996 , n548 );
and ( n3014 , n31995 , n31996 );
nor ( n3015 , n3011 , n3014 );
buf ( n31999 , n3015 );
buf ( n32000 , n31999 );
nand ( n3018 , n31989 , n32000 );
buf ( n32002 , n3018 );
buf ( n3020 , n32002 );
buf ( n32004 , n3020 );
buf ( n32005 , n547 );
buf ( n32006 , n534 );
not ( n3024 , n32006 );
buf ( n32008 , n3024 );
buf ( n32009 , n32008 );
and ( n3027 , n32005 , n32009 );
not ( n3028 , n32005 );
buf ( n32012 , n534 );
and ( n3030 , n3028 , n32012 );
nor ( n3031 , n3027 , n3030 );
buf ( n32015 , n3031 );
buf ( n32016 , n32015 );
or ( n3034 , n32004 , n32016 );
nand ( n3035 , n3001 , n3034 );
buf ( n32019 , n3035 );
buf ( n32020 , n32019 );
xor ( n3041 , n2981 , n32020 );
buf ( n32022 , n3041 );
buf ( n32023 , n32022 );
xor ( n3044 , n31923 , n32023 );
buf ( n3045 , n2911 );
buf ( n32026 , n3045 );
buf ( n32027 , n31913 );
or ( n3048 , n32026 , n32027 );
buf ( n32029 , n2918 );
buf ( n32030 , n31868 );
buf ( n32031 , n531 );
and ( n3052 , n32030 , n32031 );
buf ( n32033 , n31840 );
buf ( n32034 , n549 );
and ( n3055 , n32033 , n32034 );
nor ( n3056 , n3052 , n3055 );
buf ( n32037 , n3056 );
buf ( n32038 , n32037 );
or ( n3059 , n32029 , n32038 );
nand ( n3060 , n3048 , n3059 );
buf ( n32041 , n3060 );
buf ( n32042 , n32041 );
xor ( n3063 , n546 , n547 );
not ( n3064 , n3063 );
buf ( n32045 , n545 );
buf ( n32046 , n546 );
xor ( n3067 , n32045 , n32046 );
buf ( n32048 , n3067 );
nand ( n3069 , n3064 , n32048 );
buf ( n32050 , n3069 );
buf ( n32051 , n545 );
not ( n3072 , n32051 );
buf ( n32053 , n3072 );
buf ( n32054 , n32053 );
buf ( n32055 , n536 );
and ( n3076 , n32054 , n32055 );
buf ( n32057 , n536 );
not ( n3078 , n32057 );
buf ( n32059 , n3078 );
buf ( n32060 , n32059 );
buf ( n32061 , n545 );
and ( n3082 , n32060 , n32061 );
nor ( n3083 , n3076 , n3082 );
buf ( n32064 , n3083 );
buf ( n32065 , n32064 );
or ( n3086 , n32050 , n32065 );
not ( n3087 , n3063 );
buf ( n32068 , n3087 );
buf ( n32069 , n32053 );
buf ( n32070 , n535 );
and ( n3091 , n32069 , n32070 );
buf ( n32072 , n535 );
not ( n3093 , n32072 );
buf ( n32074 , n3093 );
buf ( n32075 , n32074 );
buf ( n32076 , n545 );
and ( n3097 , n32075 , n32076 );
nor ( n3098 , n3091 , n3097 );
buf ( n32079 , n3098 );
buf ( n32080 , n32079 );
or ( n3101 , n32068 , n32080 );
nand ( n3102 , n3086 , n3101 );
buf ( n32083 , n3102 );
buf ( n32084 , n32083 );
xor ( n32085 , n32042 , n32084 );
buf ( n32086 , n3087 );
buf ( n32087 , n32059 );
nor ( n3108 , n32086 , n32087 );
buf ( n32089 , n3108 );
xor ( n3110 , n32089 , n466 );
buf ( n32091 , n3020 );
buf ( n32092 , n547 );
buf ( n32093 , n32074 );
and ( n3114 , n32092 , n32093 );
not ( n3115 , n32092 );
buf ( n32096 , n535 );
and ( n3117 , n3115 , n32096 );
nor ( n3118 , n3114 , n3117 );
buf ( n32099 , n3118 );
buf ( n32100 , n32099 );
or ( n3121 , n32091 , n32100 );
buf ( n32102 , n31978 );
buf ( n32103 , n32015 );
or ( n3124 , n32102 , n32103 );
nand ( n3125 , n3121 , n3124 );
buf ( n32106 , n3125 );
and ( n3127 , n3110 , n32106 );
and ( n3128 , n32089 , n466 );
or ( n3129 , n3127 , n3128 );
buf ( n32110 , n3129 );
xor ( n3131 , n32085 , n32110 );
buf ( n32112 , n3131 );
buf ( n32113 , n32112 );
and ( n3134 , n3044 , n32113 );
and ( n3135 , n31923 , n32023 );
or ( n3136 , n3134 , n3135 );
buf ( n32117 , n3136 );
not ( n3138 , n454 );
nand ( n3139 , n32117 , n3138 );
not ( n3140 , n3139 );
and ( n3141 , n454 , n544 );
not ( n3142 , n454 );
or ( n3143 , n32079 , n3069 );
buf ( n32124 , n32053 );
buf ( n32125 , n534 );
and ( n3146 , n32124 , n32125 );
buf ( n32127 , n32008 );
buf ( n32128 , n545 );
and ( n3149 , n32127 , n32128 );
nor ( n3150 , n3146 , n3149 );
buf ( n32131 , n3150 );
or ( n3152 , n32131 , n3087 );
nand ( n3153 , n3143 , n3152 );
and ( n3154 , n31924 , n31940 );
buf ( n32135 , n3154 );
xor ( n3156 , n3153 , n32135 );
buf ( n32137 , n3020 );
buf ( n32138 , n31972 );
not ( n3159 , n32138 );
buf ( n32140 , n3159 );
buf ( n32141 , n32140 );
or ( n3162 , n32137 , n32141 );
buf ( n32143 , n31978 );
buf ( n32144 , n547 );
buf ( n32145 , n31908 );
and ( n3166 , n32144 , n32145 );
not ( n3167 , n32144 );
buf ( n32148 , n532 );
and ( n3169 , n3167 , n32148 );
nor ( n3170 , n3166 , n3169 );
buf ( n32151 , n3170 );
buf ( n32152 , n32151 );
or ( n3176 , n32143 , n32152 );
nand ( n3177 , n3162 , n3176 );
buf ( n32155 , n3177 );
xor ( n3179 , n3156 , n32155 );
xor ( n3180 , n32042 , n32084 );
and ( n3181 , n3180 , n32110 );
and ( n3182 , n32042 , n32084 );
or ( n3183 , n3181 , n3182 );
buf ( n32161 , n3183 );
xnor ( n3185 , n544 , n545 );
buf ( n32163 , n3185 );
not ( n3187 , n32163 );
buf ( n32165 , n3187 );
buf ( n32166 , n32165 );
buf ( n32167 , n536 );
and ( n3191 , n32166 , n32167 );
buf ( n32169 , n3191 );
xor ( n3193 , n32169 , n464 );
buf ( n32171 , n31957 );
not ( n3195 , n32171 );
buf ( n32173 , n3195 );
buf ( n32174 , n32173 );
not ( n3198 , n32174 );
not ( n3199 , n2846 );
buf ( n32177 , n3199 );
not ( n3201 , n32177 );
or ( n3202 , n3198 , n3201 );
buf ( n32180 , n551 );
buf ( n32181 , n528 );
not ( n3205 , n32181 );
buf ( n32183 , n3205 );
buf ( n32184 , n32183 );
and ( n3208 , n32180 , n32184 );
not ( n3209 , n32180 );
buf ( n32187 , n528 );
and ( n3211 , n3209 , n32187 );
nor ( n3212 , n3208 , n3211 );
buf ( n32190 , n3212 );
buf ( n32191 , n32190 );
buf ( n32192 , n2845 );
or ( n3216 , n32191 , n32192 );
nand ( n3217 , n3202 , n3216 );
buf ( n32195 , n3217 );
xor ( n3219 , n3193 , n32195 );
buf ( n32197 , n3045 );
buf ( n32198 , n32037 );
or ( n3222 , n32197 , n32198 );
buf ( n32200 , n2918 );
buf ( n32201 , n31868 );
buf ( n32202 , n530 );
and ( n3226 , n32201 , n32202 );
buf ( n32204 , n31853 );
buf ( n32205 , n549 );
and ( n3229 , n32204 , n32205 );
nor ( n3230 , n3226 , n3229 );
buf ( n32208 , n3230 );
buf ( n32209 , n32208 );
or ( n3233 , n32200 , n32209 );
nand ( n3234 , n3222 , n3233 );
buf ( n32212 , n3234 );
xor ( n3236 , n31943 , n31963 );
and ( n32214 , n3236 , n32020 );
and ( n3238 , n31943 , n31963 );
or ( n3239 , n32214 , n3238 );
buf ( n32217 , n3239 );
xor ( n3241 , n32212 , n32217 );
xor ( n3242 , n3219 , n3241 );
xor ( n3243 , n32161 , n3242 );
xor ( n3244 , n3179 , n3243 );
and ( n3245 , n3142 , n3244 );
or ( n3246 , n3141 , n3245 );
nor ( n3247 , n3140 , n3246 );
and ( n3248 , n2824 , n3247 );
not ( n3249 , n3248 );
nand ( n3250 , n2824 , n3139 );
nand ( n3251 , n3246 , n3250 );
nand ( n3252 , n3249 , n3251 );
not ( n3253 , n3252 );
nand ( n3254 , n2362 , n2261 );
nand ( n3255 , n3254 , n2513 );
buf ( n3256 , n2253 );
not ( n3257 , n3256 );
xor ( n3258 , n3255 , n3257 );
nand ( n3259 , n3258 , n2815 );
not ( n3260 , n3259 );
buf ( n3261 , n1472 );
nand ( n3262 , n3261 , n1463 );
not ( n3263 , n3262 );
xor ( n3264 , n1808 , n3263 );
nand ( n3265 , n3264 , n455 );
not ( n3266 , n3265 );
or ( n3267 , n3260 , n3266 );
nand ( n3268 , n3267 , n454 );
buf ( n32246 , n3045 );
buf ( n32247 , n31868 );
buf ( n32248 , n535 );
and ( n3272 , n32247 , n32248 );
buf ( n32250 , n32074 );
buf ( n32251 , n549 );
and ( n3275 , n32250 , n32251 );
nor ( n3276 , n3272 , n3275 );
buf ( n32254 , n3276 );
buf ( n32255 , n32254 );
or ( n3279 , n32246 , n32255 );
buf ( n32257 , n2918 );
buf ( n32258 , n31868 );
buf ( n32259 , n534 );
and ( n3283 , n32258 , n32259 );
buf ( n32261 , n32008 );
buf ( n32262 , n549 );
and ( n3286 , n32261 , n32262 );
nor ( n3287 , n3283 , n3286 );
buf ( n32265 , n3287 );
buf ( n32266 , n32265 );
or ( n3290 , n32257 , n32266 );
nand ( n3291 , n3279 , n3290 );
buf ( n32269 , n3291 );
buf ( n32270 , n32269 );
buf ( n32271 , n2962 );
buf ( n32272 , n2848 );
buf ( n32273 , n533 );
and ( n3297 , n32272 , n32273 );
buf ( n32275 , n31874 );
buf ( n32276 , n551 );
and ( n3303 , n32275 , n32276 );
nor ( n3304 , n3297 , n3303 );
buf ( n32279 , n3304 );
buf ( n32280 , n32279 );
or ( n3307 , n32271 , n32280 );
buf ( n32282 , n2848 );
buf ( n32283 , n532 );
and ( n3310 , n32282 , n32283 );
buf ( n32285 , n31908 );
buf ( n32286 , n551 );
and ( n3313 , n32285 , n32286 );
nor ( n3314 , n3310 , n3313 );
buf ( n32289 , n3314 );
buf ( n32290 , n32289 );
buf ( n32291 , n2845 );
or ( n3318 , n32290 , n32291 );
nand ( n3319 , n3307 , n3318 );
buf ( n32294 , n3319 );
buf ( n32295 , n32294 );
xor ( n3322 , n32270 , n32295 );
buf ( n32297 , n31978 );
buf ( n32298 , n32059 );
nor ( n3325 , n32297 , n32298 );
buf ( n32300 , n3325 );
buf ( n32301 , n32300 );
buf ( n32302 , n468 );
xor ( n3329 , n32301 , n32302 );
buf ( n32304 , n469 );
buf ( n32305 , n536 );
buf ( n32306 , n550 );
and ( n3333 , n32305 , n32306 );
buf ( n32308 , n32059 );
buf ( n32309 , n31889 );
and ( n3336 , n32308 , n32309 );
buf ( n32311 , n2848 );
nor ( n3338 , n3336 , n32311 );
buf ( n32313 , n3338 );
buf ( n32314 , n32313 );
buf ( n32315 , n31868 );
nor ( n3342 , n3333 , n32314 , n32315 );
buf ( n32317 , n3342 );
buf ( n32318 , n32317 );
and ( n3345 , n32304 , n32318 );
buf ( n32320 , n3345 );
buf ( n32321 , n32320 );
xor ( n3348 , n3329 , n32321 );
buf ( n32323 , n3348 );
buf ( n32324 , n32323 );
and ( n3351 , n3322 , n32324 );
and ( n3352 , n32270 , n32295 );
or ( n3353 , n3351 , n3352 );
buf ( n32328 , n3353 );
buf ( n32329 , n32328 );
buf ( n32330 , n3138 );
nand ( n32331 , n32329 , n32330 );
buf ( n32332 , n32331 );
not ( n3359 , n32332 );
not ( n3360 , n454 );
not ( n3361 , n3360 );
buf ( n32336 , n3045 );
buf ( n32337 , n32265 );
or ( n3364 , n32336 , n32337 );
buf ( n32339 , n2918 );
buf ( n32340 , n31879 );
or ( n3367 , n32339 , n32340 );
nand ( n3368 , n3364 , n3367 );
buf ( n32343 , n3368 );
xor ( n3370 , n31811 , n31827 );
buf ( n32345 , n3370 );
buf ( n32346 , n32289 );
buf ( n32347 , n2846 );
or ( n3374 , n32346 , n32347 );
buf ( n32349 , n31845 );
buf ( n32350 , n552 );
not ( n3377 , n32350 );
buf ( n32352 , n3377 );
buf ( n32353 , n32352 );
or ( n3380 , n32349 , n32353 );
nand ( n3381 , n3374 , n3380 );
buf ( n32356 , n3381 );
and ( n3383 , n32345 , n32356 );
not ( n3384 , n32345 );
not ( n3385 , n32356 );
and ( n3386 , n3384 , n3385 );
or ( n3387 , n3383 , n3386 );
buf ( n32362 , n3020 );
buf ( n32363 , n547 );
buf ( n32364 , n32059 );
and ( n3391 , n32363 , n32364 );
not ( n3392 , n32363 );
buf ( n32367 , n536 );
and ( n3394 , n3392 , n32367 );
nor ( n3395 , n3391 , n3394 );
buf ( n32370 , n3395 );
buf ( n32371 , n32370 );
or ( n3398 , n32362 , n32371 );
buf ( n32373 , n31978 );
buf ( n32374 , n32099 );
or ( n3401 , n32373 , n32374 );
nand ( n3402 , n3398 , n3401 );
buf ( n32377 , n3402 );
xnor ( n3404 , n3387 , n32377 );
xor ( n3405 , n32343 , n3404 );
xor ( n3406 , n32301 , n32302 );
and ( n3407 , n3406 , n32321 );
and ( n3408 , n32301 , n32302 );
or ( n3409 , n3407 , n3408 );
buf ( n32384 , n3409 );
xor ( n3411 , n3405 , n32384 );
not ( n32386 , n3411 );
or ( n3416 , n3361 , n32386 );
nand ( n3417 , n547 , n454 );
nand ( n3418 , n3416 , n3417 );
nor ( n3419 , n3359 , n3418 );
nand ( n3420 , n3268 , n3419 );
not ( n3421 , n3420 );
xor ( n3422 , n32304 , n32318 );
buf ( n32394 , n3422 );
buf ( n32395 , n32394 );
buf ( n32396 , n2962 );
buf ( n32397 , n2848 );
buf ( n32398 , n534 );
and ( n3428 , n32397 , n32398 );
buf ( n32400 , n32008 );
buf ( n32401 , n551 );
and ( n3431 , n32400 , n32401 );
nor ( n3432 , n3428 , n3431 );
buf ( n32404 , n3432 );
buf ( n32405 , n32404 );
or ( n3435 , n32396 , n32405 );
buf ( n32407 , n32279 );
buf ( n32408 , n32352 );
or ( n3438 , n32407 , n32408 );
nand ( n3439 , n3435 , n3438 );
buf ( n32411 , n3439 );
buf ( n32412 , n32411 );
xor ( n3442 , n32395 , n32412 );
buf ( n32414 , n31868 );
buf ( n32415 , n536 );
and ( n3445 , n32414 , n32415 );
buf ( n32417 , n32059 );
buf ( n32418 , n549 );
and ( n3448 , n32417 , n32418 );
nor ( n3449 , n3445 , n3448 );
buf ( n32421 , n3449 );
or ( n3451 , n32421 , n3045 );
or ( n3452 , n2918 , n32254 );
nand ( n3453 , n3451 , n3452 );
buf ( n32425 , n3453 );
and ( n3455 , n3442 , n32425 );
and ( n3456 , n32395 , n32412 );
or ( n3457 , n3455 , n3456 );
buf ( n32429 , n3457 );
nand ( n3459 , n32429 , n3138 );
not ( n3460 , n3459 );
not ( n3461 , n2815 );
not ( n3462 , n2248 );
not ( n3463 , n3462 );
nand ( n3464 , n2040 , n2108 );
not ( n3465 , n3464 );
or ( n3466 , n3463 , n3465 );
nand ( n32438 , n3466 , n2107 );
not ( n3468 , n2252 );
nor ( n3469 , n3468 , n2247 );
xor ( n3470 , n32438 , n3469 );
not ( n3471 , n3470 );
or ( n3472 , n3461 , n3471 );
not ( n3473 , n1615 );
not ( n3474 , n3473 );
nand ( n3475 , n1800 , n1802 );
not ( n3476 , n3475 );
or ( n3477 , n3474 , n3476 );
nand ( n3478 , n3477 , n1801 );
not ( n3479 , n3478 );
not ( n3480 , n1623 );
nand ( n3481 , n3480 , n1807 );
nand ( n3482 , n3479 , n3481 );
not ( n3483 , n3481 );
nand ( n3484 , n3483 , n3478 );
nand ( n3485 , n3482 , n3484 , n455 );
nand ( n3486 , n3472 , n3485 );
nand ( n3487 , n3486 , n454 );
not ( n3488 , n3487 );
or ( n3489 , n3460 , n3488 );
and ( n3490 , n454 , n548 );
not ( n3491 , n454 );
xor ( n3492 , n32270 , n32295 );
xor ( n3493 , n3492 , n32324 );
buf ( n32465 , n3493 );
and ( n3495 , n3491 , n32465 );
or ( n3496 , n3490 , n3495 );
nand ( n3497 , n3489 , n3496 );
or ( n3498 , n3421 , n3497 );
not ( n3499 , n32332 );
not ( n3500 , n3268 );
or ( n3501 , n3499 , n3500 );
nand ( n3502 , n3501 , n3418 );
nand ( n3503 , n3498 , n3502 );
not ( n3504 , n3261 );
not ( n3505 , n1808 );
or ( n3506 , n3504 , n3505 );
nand ( n3507 , n3506 , n1463 );
and ( n3508 , n1467 , n1392 );
and ( n3509 , n3507 , n3508 );
not ( n3510 , n3507 );
not ( n3511 , n3508 );
and ( n3512 , n3510 , n3511 );
nor ( n3513 , n3509 , n3512 );
and ( n3514 , n454 , n455 );
and ( n3515 , n3513 , n3514 );
xor ( n3516 , n32343 , n3404 );
and ( n3517 , n3516 , n32384 );
and ( n32489 , n32343 , n3404 );
or ( n3522 , n3517 , n32489 );
and ( n3523 , n3522 , n3138 );
nor ( n3524 , n3515 , n3523 );
not ( n3525 , n3524 );
nand ( n3526 , n2524 , n2519 );
not ( n3527 , n3526 );
not ( n3528 , n3527 );
not ( n3529 , n3256 );
and ( n3530 , n3529 , n2513 );
not ( n3531 , n3254 );
nand ( n3532 , n3531 , n2513 );
not ( n3533 , n3532 );
nor ( n3534 , n3530 , n3533 );
not ( n3535 , n3534 );
or ( n3536 , n3528 , n3535 );
and ( n3537 , n2513 , n3526 );
and ( n3538 , n3537 , n3529 );
or ( n3539 , n3527 , n3532 );
nand ( n3540 , n3539 , n2815 );
nor ( n3541 , n3538 , n3540 );
nand ( n3542 , n3536 , n3541 );
not ( n3543 , n454 );
nor ( n3544 , n3542 , n3543 );
nor ( n3545 , n3525 , n3544 );
buf ( n32514 , n454 );
buf ( n32515 , n546 );
and ( n3548 , n32514 , n32515 );
not ( n3549 , n32514 );
xor ( n3550 , n32089 , n466 );
xor ( n3551 , n3550 , n32106 );
not ( n3552 , n32345 );
nand ( n3553 , n3552 , n3385 );
not ( n3554 , n3553 );
not ( n3555 , n32377 );
or ( n3556 , n3554 , n3555 );
nand ( n3557 , n32356 , n32345 );
nand ( n3558 , n3556 , n3557 );
xor ( n3559 , n31830 , n31864 );
xor ( n3560 , n3559 , n31918 );
buf ( n32529 , n3560 );
xor ( n3562 , n3558 , n32529 );
xor ( n3563 , n3551 , n3562 );
buf ( n32532 , n3563 );
and ( n3565 , n3549 , n32532 );
or ( n3566 , n3548 , n3565 );
buf ( n32535 , n3566 );
not ( n3568 , n32535 );
nand ( n3569 , n3545 , n3568 );
not ( n3570 , n455 );
nand ( n3571 , n1304 , n1814 );
not ( n3572 , n3571 );
and ( n3573 , n1810 , n3572 );
not ( n3574 , n1810 );
and ( n3575 , n3574 , n3571 );
nor ( n3576 , n3573 , n3575 );
not ( n3577 , n3576 );
or ( n3578 , n3570 , n3577 );
nand ( n3579 , n2652 , n2654 );
not ( n3580 , n3579 );
and ( n3581 , n2526 , n3580 );
not ( n3582 , n2526 );
and ( n3583 , n3582 , n3579 );
nor ( n3584 , n3581 , n3583 );
nand ( n3585 , n3584 , n2815 );
nand ( n3586 , n3578 , n3585 );
and ( n3587 , n3586 , n454 );
xor ( n3588 , n31923 , n32023 );
xor ( n3589 , n3588 , n32113 );
buf ( n32558 , n3589 );
buf ( n32559 , n32558 );
buf ( n32560 , n3360 );
nand ( n3593 , n32559 , n32560 );
buf ( n32562 , n3593 );
nand ( n3595 , n545 , n454 );
and ( n3596 , n32562 , n3595 );
xor ( n3597 , n32089 , n466 );
xor ( n3598 , n3597 , n32106 );
and ( n3599 , n3558 , n3598 );
xor ( n3600 , n32089 , n466 );
xor ( n3601 , n3600 , n32106 );
and ( n3602 , n32529 , n3601 );
and ( n3603 , n3558 , n32529 );
or ( n3604 , n3599 , n3602 , n3603 );
nand ( n3605 , n3604 , n3138 );
and ( n3606 , n3596 , n3605 );
not ( n3607 , n3606 );
nor ( n3608 , n3587 , n3607 );
not ( n3609 , n3608 );
nand ( n3610 , n3503 , n3569 , n3609 );
not ( n3611 , n3419 );
not ( n32580 , n3268 );
or ( n3616 , n3611 , n32580 );
nand ( n3617 , n3487 , n3459 );
or ( n3618 , n3496 , n3617 );
nand ( n3619 , n3616 , n3618 );
xor ( n3620 , n30877 , n1922 );
xor ( n3621 , n3620 , n1968 );
nand ( n3622 , n3621 , n2815 , n454 );
buf ( n32588 , n2848 );
buf ( n32589 , n535 );
and ( n3625 , n32588 , n32589 );
buf ( n32591 , n32074 );
buf ( n32592 , n551 );
and ( n3628 , n32591 , n32592 );
nor ( n3629 , n3625 , n3628 );
buf ( n32595 , n3629 );
buf ( n32596 , n32595 );
buf ( n32597 , n32352 );
or ( n3633 , n32596 , n32597 );
buf ( n32599 , n2962 );
buf ( n32600 , n536 );
or ( n3636 , n32599 , n32600 );
nand ( n3637 , n3633 , n3636 );
buf ( n32603 , n3637 );
nand ( n3639 , n32603 , n3138 );
and ( n3640 , n3622 , n3639 );
nand ( n3641 , n1731 , n1787 );
buf ( n3642 , n1783 );
not ( n3643 , n3642 );
and ( n3644 , n3641 , n3643 );
not ( n3645 , n3641 );
and ( n3646 , n3645 , n3642 );
nor ( n3647 , n3644 , n3646 );
and ( n3648 , n455 , n454 );
nand ( n3649 , n3647 , n3648 );
nand ( n3650 , n3640 , n3649 );
not ( n3651 , n3650 );
and ( n3652 , n454 , n551 );
not ( n3653 , n454 );
buf ( n32619 , n471 );
buf ( n32620 , n2848 );
buf ( n32621 , n536 );
buf ( n32622 , n552 );
and ( n3658 , n32621 , n32622 );
buf ( n32624 , n3658 );
buf ( n32625 , n32624 );
nor ( n3661 , n32620 , n32625 );
buf ( n32627 , n3661 );
buf ( n32628 , n32627 );
xor ( n3664 , n32619 , n32628 );
buf ( n32630 , n3664 );
and ( n3666 , n3653 , n32630 );
or ( n3667 , n3652 , n3666 );
not ( n3668 , n3667 );
nand ( n3669 , n3651 , n3668 );
not ( n3670 , n3669 );
or ( n3671 , n30949 , n30932 );
nand ( n3672 , n3671 , n1967 );
xnor ( n3673 , n3672 , n1965 );
nand ( n3674 , n2815 , n3673 );
not ( n3675 , n3674 );
not ( n3676 , n1781 );
or ( n3677 , n1757 , n30750 );
nand ( n3678 , n3677 , n1758 );
not ( n3679 , n3678 );
or ( n3680 , n3676 , n3679 );
or ( n3681 , n3678 , n1781 );
nand ( n3682 , n3680 , n3681 );
nand ( n3683 , n3682 , n455 );
not ( n3684 , n3683 );
or ( n3685 , n3675 , n3684 );
nand ( n3686 , n3685 , n454 );
buf ( n32652 , n3686 );
buf ( n32653 , n3138 );
buf ( n32654 , n472 );
nand ( n3690 , n32653 , n32654 );
buf ( n32656 , n3690 );
buf ( n32657 , n32656 );
nand ( n3693 , n32652 , n32657 );
buf ( n32659 , n3693 );
buf ( n32660 , n454 );
buf ( n32661 , n552 );
and ( n3697 , n32660 , n32661 );
not ( n32663 , n32660 );
buf ( n32664 , n32624 );
and ( n3703 , n32663 , n32664 );
or ( n3704 , n3697 , n3703 );
buf ( n32667 , n3704 );
and ( n3706 , n32659 , n32667 );
not ( n3707 , n3706 );
or ( n3708 , n3670 , n3707 );
nand ( n3709 , n3667 , n3650 );
nand ( n3710 , n3708 , n3709 );
not ( n3711 , n454 );
not ( n3712 , n1798 );
not ( n3713 , n1792 );
or ( n3714 , n3712 , n3713 );
nand ( n3715 , n3714 , n1802 );
and ( n3716 , n3715 , n1788 );
not ( n3717 , n3715 );
not ( n3718 , n1788 );
and ( n3719 , n3717 , n3718 );
nor ( n3720 , n3716 , n3719 );
and ( n3721 , n455 , n3720 );
not ( n3722 , n455 );
nand ( n3723 , n2039 , n2108 );
xor ( n3724 , n1971 , n3723 );
and ( n3725 , n3722 , n3724 );
nor ( n3726 , n3721 , n3725 );
not ( n3727 , n3726 );
or ( n3728 , n3711 , n3727 );
or ( n3729 , n32404 , n2845 );
or ( n3730 , n32595 , n2962 );
nand ( n3731 , n3729 , n3730 );
nand ( n3732 , n3731 , n3138 );
nand ( n3733 , n3728 , n3732 );
buf ( n32696 , n454 );
buf ( n32697 , n550 );
and ( n3736 , n32696 , n32697 );
not ( n32699 , n32696 );
buf ( n32700 , n2918 );
buf ( n32701 , n32059 );
nor ( n3740 , n32700 , n32701 );
buf ( n32703 , n3740 );
buf ( n32704 , n32703 );
buf ( n32705 , n470 );
xor ( n3744 , n32704 , n32705 );
and ( n3745 , n32619 , n32628 );
buf ( n32708 , n3745 );
buf ( n32709 , n32708 );
xor ( n3748 , n3744 , n32709 );
buf ( n32711 , n3748 );
buf ( n32712 , n32711 );
and ( n3751 , n32699 , n32712 );
or ( n3752 , n3736 , n3751 );
buf ( n32715 , n3752 );
nand ( n3754 , n3733 , n32715 );
not ( n3755 , n3754 );
or ( n3756 , n3710 , n3755 );
not ( n3757 , n3733 );
not ( n3758 , n32715 );
nand ( n3759 , n3757 , n3758 );
nand ( n3760 , n3756 , n3759 );
not ( n3761 , n3760 );
not ( n3762 , n2815 );
nand ( n3763 , n3462 , n2107 );
not ( n3764 , n3763 );
not ( n3765 , n3464 );
or ( n3766 , n3764 , n3765 );
or ( n3767 , n3464 , n3763 );
nand ( n3768 , n3766 , n3767 );
not ( n3769 , n3768 );
or ( n3770 , n3762 , n3769 );
buf ( n3771 , n1801 );
nand ( n32734 , n3771 , n3473 );
not ( n3776 , n32734 );
and ( n3777 , n3475 , n3776 );
not ( n3778 , n3475 );
and ( n3779 , n3778 , n32734 );
nor ( n3780 , n3777 , n3779 );
nand ( n3781 , n3780 , n455 );
nand ( n3782 , n3770 , n3781 );
and ( n3783 , n3782 , n454 );
xor ( n3784 , n32704 , n32705 );
and ( n3785 , n3784 , n32709 );
and ( n3786 , n32704 , n32705 );
or ( n3787 , n3785 , n3786 );
buf ( n32747 , n3787 );
and ( n3789 , n32747 , n3138 );
nor ( n3790 , n3783 , n3789 );
not ( n3791 , n3790 );
not ( n3792 , n549 );
not ( n3793 , n454 );
or ( n3794 , n3792 , n3793 );
xor ( n3795 , n32395 , n32412 );
xor ( n3796 , n3795 , n32425 );
buf ( n32756 , n3796 );
buf ( n32757 , n32756 );
buf ( n32758 , n3360 );
nand ( n3800 , n32757 , n32758 );
buf ( n32760 , n3800 );
nand ( n3802 , n3794 , n32760 );
nand ( n3803 , n3791 , n3802 );
not ( n3804 , n3803 );
or ( n3805 , n3761 , n3804 );
not ( n3806 , n3802 );
nand ( n32766 , n3806 , n3790 );
nand ( n3808 , n3805 , n32766 );
nor ( n3809 , n3619 , n3808 );
not ( n3810 , n454 );
not ( n3811 , n3586 );
or ( n3812 , n3810 , n3811 );
nand ( n3813 , n3812 , n3606 );
nand ( n3814 , n3809 , n3569 , n3813 );
not ( n3815 , n3524 );
not ( n3816 , n3544 );
not ( n3817 , n3816 );
or ( n3818 , n3815 , n3817 );
nand ( n3819 , n3818 , n32535 );
not ( n3820 , n3819 );
and ( n3821 , n3813 , n3820 );
nand ( n3822 , n3586 , n454 );
and ( n3823 , n3822 , n3605 );
nor ( n3824 , n3823 , n3596 );
nor ( n3825 , n3821 , n3824 );
nand ( n3826 , n3610 , n3814 , n3825 );
buf ( n3827 , n3826 );
not ( n3828 , n3827 );
or ( n3829 , n3253 , n3828 );
not ( n3830 , n3826 );
nand ( n3831 , n3830 , n3251 , n3249 );
nand ( n3832 , n3829 , n3831 );
or ( n3833 , n3832 , n469 );
nand ( n3834 , n3832 , n469 );
nand ( n3835 , n3833 , n3834 );
not ( n3836 , n3835 );
buf ( n3837 , n3503 );
not ( n32797 , n3837 );
buf ( n3842 , n3569 );
not ( n3843 , n3842 );
or ( n3844 , n32797 , n3843 );
not ( n3845 , n3820 );
nand ( n3846 , n3844 , n3845 );
not ( n3847 , n3846 );
nor ( n3848 , n3619 , n3808 );
buf ( n3849 , n3848 );
nand ( n3850 , n3842 , n3849 );
and ( n3851 , n3822 , n3605 );
nor ( n3852 , n3851 , n3596 );
or ( n3853 , n3852 , n3608 );
not ( n3854 , n3853 );
nand ( n3855 , n3847 , n3850 , n3854 );
not ( n3856 , n3850 );
or ( n3857 , n3856 , n3846 );
nand ( n3858 , n3857 , n3853 );
not ( n3859 , n470 );
nand ( n3860 , n3855 , n3858 , n3859 );
buf ( n3861 , n3860 );
not ( n3862 , n3861 );
not ( n3863 , n3459 );
nor ( n3864 , n3863 , n3496 );
nand ( n3865 , n3487 , n3864 );
not ( n3866 , n3865 );
not ( n32823 , n3808 );
not ( n3868 , n32823 );
or ( n3869 , n3866 , n3868 );
nand ( n3870 , n3869 , n3497 );
not ( n3871 , n3421 );
nand ( n3872 , n3871 , n3502 );
not ( n3873 , n3872 );
and ( n3874 , n3870 , n3873 );
not ( n3875 , n3870 );
and ( n3876 , n3875 , n3872 );
nor ( n3877 , n3874 , n3876 );
nand ( n3878 , n3877 , n472 );
not ( n3879 , n3878 );
xor ( n3880 , n471 , n3879 );
nand ( n3881 , n3842 , n3845 );
not ( n3882 , n3881 );
nor ( n3883 , n3849 , n3837 );
not ( n3884 , n3883 );
not ( n3885 , n3884 );
or ( n3886 , n3882 , n3885 );
or ( n3887 , n3881 , n3884 );
nand ( n3888 , n3886 , n3887 );
and ( n3889 , n3880 , n3888 );
and ( n3890 , n471 , n3879 );
or ( n3891 , n3889 , n3890 );
buf ( n32848 , n3891 );
not ( n3896 , n32848 );
or ( n3897 , n3862 , n3896 );
nand ( n3898 , n3855 , n3858 );
and ( n3899 , n3898 , n470 );
not ( n3900 , n3899 );
nand ( n3901 , n3897 , n3900 );
not ( n3902 , n3901 );
or ( n3903 , n3836 , n3902 );
or ( n3904 , n3835 , n3901 );
nand ( n3905 , n3903 , n3904 );
not ( n3906 , n3905 );
or ( n3907 , n29521 , n3906 );
xnor ( n3908 , n1405 , n29494 );
not ( n3909 , n29494 );
and ( n3910 , n456 , n467 );
not ( n3911 , n456 );
and ( n3912 , n3911 , n483 );
nor ( n3913 , n3910 , n3912 );
not ( n3914 , n3913 );
or ( n3915 , n3909 , n3914 );
not ( n3916 , n3913 );
not ( n32870 , n29494 );
nand ( n3918 , n3916 , n32870 );
nand ( n3919 , n3915 , n3918 );
nand ( n3920 , n3908 , n3919 );
not ( n3921 , n3916 );
and ( n3922 , n504 , n3921 );
not ( n3923 , n504 );
and ( n3924 , n3923 , n3916 );
nor ( n3925 , n3922 , n3924 );
or ( n3926 , n3920 , n3925 );
xnor ( n3927 , n503 , n3916 );
or ( n3928 , n3927 , n3908 );
nand ( n3929 , n3926 , n3928 );
not ( n3930 , n32870 );
buf ( n3931 , n1404 );
not ( n3932 , n3931 );
or ( n3933 , n3930 , n3932 );
nand ( n3934 , n3933 , n504 );
and ( n3935 , n456 , n469 );
not ( n3936 , n456 );
and ( n3937 , n3936 , n485 );
or ( n32891 , n3935 , n3937 );
nand ( n3942 , n32891 , n29494 );
and ( n3943 , n3934 , n3942 , n3916 );
buf ( n3944 , n901 );
not ( n3945 , n3944 );
and ( n3946 , n3945 , n32891 );
not ( n3947 , n3946 );
not ( n3948 , n502 );
not ( n3949 , n3931 );
or ( n3950 , n3948 , n3949 );
not ( n3951 , n502 );
nand ( n3952 , n32891 , n3951 );
nand ( n3953 , n3950 , n3952 );
not ( n3954 , n3953 );
or ( n3955 , n3947 , n3954 );
not ( n3956 , n501 );
not ( n32907 , n3931 );
or ( n3958 , n3956 , n32907 );
not ( n3959 , n501 );
nand ( n3960 , n32891 , n3959 );
nand ( n3961 , n3958 , n3960 );
nand ( n3962 , n3961 , n3944 );
nand ( n3963 , n3955 , n3962 );
xor ( n3964 , n3943 , n3963 );
xor ( n3965 , n3929 , n3964 );
not ( n3966 , n3944 );
not ( n3967 , n3953 );
or ( n3968 , n3966 , n3967 );
not ( n3969 , n503 );
not ( n3970 , n3931 );
or ( n3971 , n3969 , n3970 );
not ( n32922 , n503 );
nand ( n3976 , n32891 , n32922 );
nand ( n32924 , n3971 , n3976 );
nand ( n3978 , n32924 , n3946 );
nand ( n32926 , n3968 , n3978 );
not ( n3980 , n3908 );
and ( n3981 , n3980 , n504 );
nor ( n3982 , n32926 , n3981 );
not ( n32930 , n3946 );
not ( n32931 , n942 );
or ( n3985 , n32930 , n32931 );
nand ( n32933 , n32924 , n3944 );
nand ( n3987 , n3985 , n32933 );
nand ( n32935 , n3944 , n504 );
and ( n3989 , n32935 , n32891 );
nand ( n3990 , n3987 , n3989 );
or ( n3991 , n3982 , n3990 );
nand ( n3992 , n32926 , n3981 );
nand ( n32940 , n3991 , n3992 );
xor ( n3994 , n3965 , n32940 );
nand ( n3995 , n3994 , n29519 );
nand ( n3996 , n3907 , n3995 );
not ( n3997 , n29520 );
not ( n3998 , n454 );
buf ( n32946 , n3045 );
buf ( n32947 , n31868 );
buf ( n32948 , n529 );
and ( n32949 , n32947 , n32948 );
buf ( n32950 , n2969 );
buf ( n32951 , n549 );
and ( n4005 , n32950 , n32951 );
nor ( n4006 , n32949 , n4005 );
buf ( n32954 , n4006 );
buf ( n32955 , n32954 );
or ( n4009 , n32946 , n32955 );
buf ( n32957 , n2918 );
buf ( n32958 , n31868 );
buf ( n32959 , n528 );
and ( n4013 , n32958 , n32959 );
buf ( n32961 , n32183 );
buf ( n32962 , n549 );
and ( n4016 , n32961 , n32962 );
nor ( n4017 , n4013 , n4016 );
buf ( n32965 , n4017 );
buf ( n32966 , n32965 );
or ( n4020 , n32957 , n32966 );
nand ( n4021 , n4009 , n4020 );
buf ( n32969 , n4021 );
buf ( n32970 , n32969 );
buf ( n32971 , n543 );
buf ( n32972 , n544 );
nor ( n4026 , n32971 , n32972 );
buf ( n32974 , n4026 );
not ( n4028 , n32974 );
nand ( n4029 , n543 , n544 );
nand ( n4030 , n4028 , n3185 , n4029 );
buf ( n32978 , n4030 );
buf ( n32979 , n543 );
not ( n4033 , n32979 );
buf ( n32981 , n4033 );
and ( n4035 , n535 , n32981 );
and ( n32983 , n32074 , n543 );
nor ( n4037 , n4035 , n32983 );
buf ( n32985 , n4037 );
or ( n4039 , n32978 , n32985 );
buf ( n4040 , n3185 );
buf ( n32988 , n4040 );
buf ( n32989 , n543 );
buf ( n32990 , n32008 );
and ( n4044 , n32989 , n32990 );
not ( n4045 , n32989 );
buf ( n32993 , n534 );
and ( n4047 , n4045 , n32993 );
nor ( n4048 , n4044 , n4047 );
buf ( n32996 , n4048 );
buf ( n32997 , n32996 );
or ( n4051 , n32988 , n32997 );
nand ( n32999 , n4039 , n4051 );
buf ( n33000 , n32999 );
buf ( n33001 , n33000 );
xor ( n4055 , n32970 , n33001 );
buf ( n33003 , n2846 );
buf ( n33004 , n32190 );
or ( n4058 , n33003 , n33004 );
buf ( n33006 , n551 );
buf ( n33007 , n527 );
not ( n4061 , n33007 );
buf ( n33009 , n4061 );
buf ( n33010 , n33009 );
and ( n4064 , n33006 , n33010 );
not ( n4065 , n33006 );
buf ( n33013 , n527 );
and ( n4067 , n4065 , n33013 );
nor ( n4068 , n4064 , n4067 );
buf ( n33016 , n4068 );
buf ( n33017 , n33016 );
buf ( n33018 , n32352 );
or ( n4072 , n33017 , n33018 );
nand ( n4073 , n4058 , n4072 );
buf ( n33021 , n4073 );
buf ( n33022 , n463 );
buf ( n33023 , n536 );
buf ( n33024 , n544 );
or ( n4078 , n33023 , n33024 );
buf ( n33026 , n545 );
nand ( n4080 , n4078 , n33026 );
buf ( n33028 , n4080 );
buf ( n33029 , n33028 );
buf ( n33030 , n536 );
buf ( n33031 , n544 );
nand ( n4085 , n33030 , n33031 );
buf ( n33033 , n4085 );
buf ( n33034 , n33033 );
buf ( n33035 , n543 );
and ( n4089 , n33029 , n33034 , n33035 );
buf ( n33037 , n4089 );
buf ( n33038 , n33037 );
xor ( n4092 , n33022 , n33038 );
buf ( n33040 , n4092 );
xor ( n4094 , n33021 , n33040 );
buf ( n33042 , n3020 );
buf ( n33043 , n32151 );
or ( n4097 , n33042 , n33043 );
buf ( n33045 , n31978 );
buf ( n33046 , n547 );
buf ( n33047 , n31840 );
and ( n4101 , n33046 , n33047 );
not ( n4102 , n33046 );
buf ( n33050 , n531 );
and ( n4104 , n4102 , n33050 );
nor ( n4105 , n4101 , n4104 );
buf ( n33053 , n4105 );
buf ( n33054 , n33053 );
or ( n4108 , n33045 , n33054 );
nand ( n4109 , n4097 , n4108 );
buf ( n33057 , n4109 );
and ( n4111 , n4094 , n33057 );
and ( n4112 , n33021 , n33040 );
or ( n4113 , n4111 , n4112 );
buf ( n33061 , n4113 );
xor ( n4115 , n4055 , n33061 );
buf ( n33063 , n4115 );
buf ( n33064 , n33063 );
buf ( n33065 , n3020 );
buf ( n33066 , n33053 );
or ( n4120 , n33065 , n33066 );
buf ( n33068 , n31978 );
buf ( n33069 , n547 );
buf ( n33070 , n31853 );
and ( n4124 , n33069 , n33070 );
not ( n4125 , n33069 );
buf ( n33073 , n530 );
and ( n4127 , n4125 , n33073 );
nor ( n4128 , n4124 , n4127 );
buf ( n33076 , n4128 );
buf ( n33077 , n33076 );
or ( n4131 , n33068 , n33077 );
nand ( n4132 , n4120 , n4131 );
buf ( n33080 , n4132 );
buf ( n33081 , n33080 );
and ( n33082 , n33022 , n33038 );
buf ( n33083 , n33082 );
buf ( n33084 , n33083 );
xor ( n33085 , n33081 , n33084 );
buf ( n33086 , n3069 );
buf ( n33087 , n32053 );
buf ( n33088 , n533 );
and ( n33089 , n33087 , n33088 );
buf ( n33090 , n31874 );
buf ( n33091 , n545 );
and ( n33092 , n33090 , n33091 );
nor ( n4146 , n33089 , n33092 );
buf ( n33094 , n4146 );
buf ( n33095 , n33094 );
or ( n4149 , n33086 , n33095 );
buf ( n33097 , n3087 );
buf ( n33098 , n545 );
buf ( n33099 , n31908 );
and ( n4153 , n33098 , n33099 );
not ( n4154 , n33098 );
buf ( n33102 , n532 );
and ( n4156 , n4154 , n33102 );
nor ( n4157 , n4153 , n4156 );
buf ( n33105 , n4157 );
buf ( n33106 , n33105 );
or ( n4160 , n33097 , n33106 );
nand ( n4161 , n4149 , n4160 );
buf ( n33109 , n4161 );
buf ( n33110 , n33109 );
xor ( n4164 , n33085 , n33110 );
buf ( n33112 , n4164 );
buf ( n33113 , n33112 );
and ( n4170 , n542 , n543 );
not ( n33115 , n542 );
and ( n33116 , n33115 , n32981 );
nor ( n4173 , n4170 , n33116 );
not ( n33118 , n4173 );
buf ( n33119 , n33118 );
buf ( n33120 , n32059 );
nor ( n4180 , n33119 , n33120 );
buf ( n33122 , n4180 );
buf ( n33123 , n33122 );
buf ( n33124 , n462 );
xor ( n4184 , n33123 , n33124 );
buf ( n33126 , n551 );
buf ( n33127 , n526 );
xor ( n33128 , n33126 , n33127 );
buf ( n33129 , n33128 );
buf ( n33130 , n33129 );
not ( n4190 , n33130 );
buf ( n33132 , n552 );
not ( n4192 , n33132 );
or ( n4193 , n4190 , n4192 );
buf ( n33135 , n2846 );
buf ( n33136 , n33016 );
or ( n4196 , n33135 , n33136 );
nand ( n4197 , n4193 , n4196 );
buf ( n33139 , n4197 );
buf ( n33140 , n33139 );
xor ( n4200 , n4184 , n33140 );
buf ( n33142 , n4200 );
buf ( n33143 , n33142 );
xor ( n4203 , n33113 , n33143 );
buf ( n33145 , n2911 );
buf ( n33146 , n32208 );
or ( n4206 , n33145 , n33146 );
buf ( n33148 , n2918 );
buf ( n33149 , n32954 );
or ( n33150 , n33148 , n33149 );
nand ( n4210 , n4206 , n33150 );
buf ( n33152 , n4210 );
buf ( n33153 , n33152 );
not ( n4213 , n32974 );
nand ( n4214 , n4213 , n3185 , n4029 );
and ( n33156 , n32059 , n543 );
and ( n4216 , n32981 , n536 );
nor ( n4217 , n33156 , n4216 );
or ( n4218 , n4214 , n4217 );
or ( n4219 , n4037 , n3185 );
nand ( n4220 , n4218 , n4219 );
buf ( n33162 , n4220 );
xor ( n4222 , n33153 , n33162 );
or ( n4223 , n32131 , n3069 );
or ( n4224 , n33094 , n3087 );
nand ( n4225 , n4223 , n4224 );
buf ( n33167 , n4225 );
and ( n4227 , n4222 , n33167 );
and ( n4228 , n33153 , n33162 );
or ( n4229 , n4227 , n4228 );
buf ( n33171 , n4229 );
buf ( n33172 , n33171 );
xor ( n4232 , n4203 , n33172 );
buf ( n33174 , n4232 );
buf ( n33175 , n33174 );
xor ( n4235 , n33064 , n33175 );
xor ( n33177 , n32169 , n464 );
and ( n33178 , n33177 , n32195 );
and ( n33179 , n32169 , n464 );
or ( n4239 , n33178 , n33179 );
xor ( n4240 , n33021 , n33040 );
xor ( n4241 , n4240 , n33057 );
and ( n4242 , n4239 , n4241 );
xor ( n4243 , n3153 , n32135 );
and ( n4244 , n4243 , n32155 );
and ( n33186 , n3153 , n32135 );
or ( n4249 , n4244 , n33186 );
xor ( n33188 , n33021 , n33040 );
xor ( n33189 , n33188 , n33057 );
and ( n4252 , n4249 , n33189 );
and ( n4253 , n4239 , n4249 );
or ( n4254 , n4242 , n4252 , n4253 );
buf ( n33193 , n4254 );
and ( n4259 , n4235 , n33193 );
and ( n4260 , n33064 , n33175 );
or ( n33196 , n4259 , n4260 );
buf ( n33197 , n33196 );
buf ( n33198 , n33197 );
buf ( n33199 , n3138 );
nand ( n4265 , n33198 , n33199 );
buf ( n33201 , n4265 );
nand ( n4267 , n3998 , n33201 );
not ( n4268 , n4267 );
or ( n4269 , n520 , n492 );
nand ( n4270 , n4269 , n493 );
nand ( n4271 , n520 , n492 );
and ( n4272 , n4270 , n4271 , n491 );
xor ( n33208 , n503 , n508 );
nand ( n4274 , n33208 , n942 , n503 );
and ( n4275 , n503 , n507 );
not ( n4276 , n503 );
buf ( n33212 , n507 );
not ( n4278 , n33212 );
buf ( n33214 , n4278 );
and ( n4280 , n4276 , n33214 );
nor ( n4281 , n4275 , n4280 );
nand ( n4282 , n4281 , n504 );
nand ( n4283 , n4274 , n4282 );
xor ( n4284 , n4272 , n4283 );
buf ( n33220 , n4284 );
xor ( n4286 , n492 , n493 );
buf ( n33222 , n4286 );
buf ( n33223 , n520 );
and ( n4289 , n33222 , n33223 );
buf ( n33225 , n4289 );
buf ( n33226 , n33225 );
xor ( n4292 , n501 , n510 );
not ( n4293 , n4292 );
not ( n4294 , n1915 );
or ( n4295 , n4293 , n4294 );
nand ( n4296 , n2160 , n2724 );
nand ( n4297 , n4295 , n4296 );
buf ( n33233 , n4297 );
xor ( n4299 , n33226 , n33233 );
xor ( n4300 , n497 , n514 );
buf ( n33236 , n4300 );
not ( n4302 , n33236 );
buf ( n33238 , n2081 );
not ( n4304 , n33238 );
or ( n4305 , n4302 , n4304 );
buf ( n33241 , n2213 );
buf ( n33242 , n2774 );
nand ( n4308 , n33241 , n33242 );
buf ( n33244 , n4308 );
buf ( n33245 , n33244 );
nand ( n4311 , n4305 , n33245 );
buf ( n33247 , n4311 );
buf ( n33248 , n33247 );
and ( n4314 , n4299 , n33248 );
and ( n4315 , n33226 , n33233 );
or ( n4316 , n4314 , n4315 );
buf ( n33252 , n4316 );
buf ( n33253 , n33252 );
xor ( n4319 , n33220 , n33253 );
buf ( n33255 , n2760 );
not ( n4321 , n33255 );
buf ( n33257 , n1847 );
not ( n4323 , n33257 );
or ( n4324 , n4321 , n4323 );
buf ( n33260 , n33208 );
buf ( n33261 , n504 );
nand ( n4327 , n33260 , n33261 );
buf ( n33263 , n4327 );
buf ( n33264 , n33263 );
nand ( n33265 , n4324 , n33264 );
buf ( n33266 , n33265 );
buf ( n33267 , n33266 );
xor ( n4333 , n495 , n516 );
buf ( n33269 , n4333 );
not ( n4335 , n33269 );
buf ( n33271 , n31271 );
not ( n33272 , n33271 );
or ( n4341 , n4335 , n33272 );
buf ( n33274 , n2411 );
buf ( n33275 , n31778 );
not ( n4344 , n33275 );
buf ( n33277 , n4344 );
buf ( n33278 , n33277 );
or ( n4347 , n33274 , n33278 );
nand ( n4348 , n4341 , n4347 );
buf ( n33281 , n4348 );
buf ( n33282 , n33281 );
xor ( n4354 , n33267 , n33282 );
buf ( n33284 , n2676 );
not ( n4356 , n33284 );
buf ( n33286 , n2668 );
not ( n4358 , n33286 );
or ( n4359 , n4356 , n4358 );
buf ( n33289 , n2591 );
buf ( n33290 , n518 );
buf ( n33291 , n493 );
xor ( n4363 , n33290 , n33291 );
buf ( n33293 , n4363 );
buf ( n33294 , n33293 );
nand ( n4366 , n33289 , n33294 );
buf ( n33296 , n4366 );
buf ( n33297 , n33296 );
nand ( n4369 , n4359 , n33297 );
buf ( n33299 , n4369 );
buf ( n33300 , n33299 );
and ( n4372 , n4354 , n33300 );
and ( n4373 , n33267 , n33282 );
or ( n4374 , n4372 , n4373 );
buf ( n33304 , n4374 );
buf ( n33305 , n33304 );
xor ( n4377 , n4319 , n33305 );
buf ( n33307 , n4377 );
buf ( n33308 , n33307 );
xor ( n4380 , n33267 , n33282 );
xor ( n33310 , n4380 , n33300 );
buf ( n33311 , n33310 );
buf ( n33312 , n33311 );
xor ( n4384 , n33226 , n33233 );
xor ( n4385 , n4384 , n33248 );
buf ( n33315 , n4385 );
buf ( n33316 , n33315 );
xor ( n4388 , n33312 , n33316 );
xor ( n4389 , n31672 , n31689 );
and ( n4390 , n4389 , n31723 );
and ( n4391 , n31672 , n31689 );
or ( n4392 , n4390 , n4391 );
buf ( n33322 , n4392 );
buf ( n33323 , n33322 );
and ( n4395 , n4388 , n33323 );
and ( n4396 , n33312 , n33316 );
or ( n4397 , n4395 , n4396 );
buf ( n33327 , n4397 );
buf ( n33328 , n33327 );
xor ( n4400 , n33308 , n33328 );
buf ( n33330 , n4300 );
not ( n4402 , n33330 );
buf ( n33332 , n2213 );
not ( n4404 , n33332 );
or ( n4405 , n4402 , n4404 );
buf ( n33335 , n2081 );
buf ( n33336 , n513 );
buf ( n33337 , n497 );
xor ( n4409 , n33336 , n33337 );
buf ( n33339 , n4409 );
buf ( n33340 , n33339 );
nand ( n33341 , n33335 , n33340 );
buf ( n33342 , n33341 );
buf ( n33343 , n33342 );
nand ( n4415 , n4405 , n33343 );
buf ( n33345 , n4415 );
not ( n33346 , n33345 );
buf ( n33347 , n4292 );
not ( n4419 , n33347 );
buf ( n33349 , n31164 );
not ( n4421 , n33349 );
or ( n33351 , n4419 , n4421 );
buf ( n33352 , n1915 );
buf ( n33353 , n509 );
buf ( n33354 , n501 );
xor ( n4426 , n33353 , n33354 );
buf ( n33356 , n4426 );
buf ( n33357 , n33356 );
nand ( n4429 , n33352 , n33357 );
buf ( n33359 , n4429 );
buf ( n33360 , n33359 );
nand ( n33361 , n33351 , n33360 );
buf ( n33362 , n33361 );
not ( n33363 , n33362 );
not ( n4435 , n33363 );
or ( n4436 , n33346 , n4435 );
not ( n4437 , n33345 );
nand ( n4438 , n4437 , n33362 );
nand ( n4439 , n4436 , n4438 );
buf ( n33369 , n4333 );
not ( n33370 , n33369 );
buf ( n33371 , n2410 );
not ( n33372 , n33371 );
buf ( n33373 , n33372 );
buf ( n33374 , n33373 );
not ( n4449 , n33374 );
or ( n4450 , n33370 , n4449 );
buf ( n33377 , n31271 );
xor ( n4452 , n495 , n515 );
buf ( n33379 , n4452 );
nand ( n33380 , n33377 , n33379 );
buf ( n33381 , n33380 );
buf ( n33382 , n33381 );
nand ( n33383 , n4450 , n33382 );
buf ( n33384 , n33383 );
and ( n4462 , n4439 , n33384 );
not ( n4463 , n4439 );
not ( n4464 , n33384 );
and ( n4465 , n4463 , n4464 );
nor ( n4466 , n4462 , n4465 );
buf ( n33390 , n33293 );
not ( n4468 , n33390 );
buf ( n33392 , n2668 );
not ( n33393 , n33392 );
or ( n4471 , n4468 , n33393 );
buf ( n33395 , n2591 );
buf ( n33396 , n517 );
buf ( n33397 , n493 );
xor ( n4475 , n33396 , n33397 );
buf ( n33399 , n4475 );
buf ( n33400 , n33399 );
nand ( n4478 , n33395 , n33400 );
buf ( n33402 , n4478 );
buf ( n33403 , n33402 );
nand ( n33404 , n4471 , n33403 );
buf ( n33405 , n33404 );
buf ( n33406 , n33405 );
xor ( n4484 , n499 , n512 );
not ( n4485 , n4484 );
not ( n4486 , n2001 );
or ( n4487 , n4485 , n4486 );
buf ( n33411 , n30884 );
buf ( n33412 , n511 );
buf ( n33413 , n499 );
xor ( n4491 , n33412 , n33413 );
buf ( n33415 , n4491 );
buf ( n33416 , n33415 );
nand ( n4494 , n33411 , n33416 );
buf ( n33418 , n4494 );
nand ( n4496 , n4487 , n33418 );
buf ( n33420 , n4496 );
xor ( n4498 , n33406 , n33420 );
buf ( n33422 , n491 );
buf ( n33423 , n520 );
xor ( n4501 , n33422 , n33423 );
buf ( n33425 , n4501 );
buf ( n33426 , n33425 );
not ( n4504 , n33426 );
not ( n4505 , n4286 );
and ( n4506 , n491 , n492 );
not ( n4507 , n491 );
not ( n4508 , n492 );
and ( n4509 , n4507 , n4508 );
nor ( n4510 , n4506 , n4509 );
nand ( n4511 , n4505 , n4510 );
not ( n4512 , n4511 );
buf ( n33436 , n4512 );
buf ( n4514 , n33436 );
buf ( n33438 , n4514 );
buf ( n33439 , n33438 );
not ( n4517 , n33439 );
or ( n4518 , n4504 , n4517 );
xor ( n4519 , n492 , n493 );
buf ( n33443 , n4519 );
buf ( n33444 , n519 );
buf ( n33445 , n491 );
xor ( n4523 , n33444 , n33445 );
buf ( n33447 , n4523 );
buf ( n33448 , n33447 );
nand ( n4526 , n33443 , n33448 );
buf ( n33450 , n4526 );
buf ( n33451 , n33450 );
nand ( n4529 , n4518 , n33451 );
buf ( n33453 , n4529 );
buf ( n33454 , n33453 );
xor ( n4532 , n4498 , n33454 );
buf ( n33456 , n4532 );
xor ( n4534 , n4466 , n33456 );
not ( n4535 , n31753 );
nand ( n4536 , n4535 , n2781 );
not ( n4537 , n4536 );
not ( n4538 , n31784 );
or ( n4539 , n4537 , n4538 );
not ( n4540 , n2781 );
nand ( n4541 , n4540 , n31753 );
nand ( n4542 , n4539 , n4541 );
not ( n4543 , n4542 );
and ( n4544 , n31706 , n31720 );
buf ( n33468 , n4544 );
not ( n33469 , n33468 );
and ( n33470 , n31011 , n4484 );
and ( n33471 , n2001 , n31682 );
nor ( n4549 , n33470 , n33471 );
nand ( n4550 , n33469 , n4549 );
not ( n4551 , n4550 );
or ( n4552 , n4543 , n4551 );
not ( n4553 , n4549 );
nand ( n4554 , n33468 , n4553 );
nand ( n33478 , n4552 , n4554 );
xor ( n4559 , n4534 , n33478 );
buf ( n33480 , n4559 );
xor ( n4561 , n4400 , n33480 );
buf ( n33482 , n4561 );
xor ( n4563 , n2748 , n31739 );
and ( n4564 , n4563 , n2799 );
and ( n4565 , n2748 , n31739 );
or ( n33486 , n4564 , n4565 );
buf ( n33487 , n33486 );
nand ( n4571 , n33469 , n4553 );
nor ( n4572 , n4542 , n4571 );
not ( n4573 , n4572 );
not ( n4574 , n4554 );
nand ( n4575 , n4574 , n4542 );
not ( n33493 , n4550 );
nand ( n4577 , n33493 , n4542 );
not ( n4578 , n4542 );
and ( n4579 , n4549 , n33468 );
nand ( n4580 , n4578 , n4579 );
nand ( n4581 , n4573 , n4575 , n4577 , n4580 );
buf ( n33499 , n4581 );
xor ( n4583 , n33487 , n33499 );
xor ( n4584 , n33312 , n33316 );
xor ( n4585 , n4584 , n33323 );
buf ( n33503 , n4585 );
buf ( n33504 , n33503 );
and ( n4588 , n4583 , n33504 );
and ( n4589 , n33487 , n33499 );
or ( n4590 , n4588 , n4589 );
buf ( n33508 , n4590 );
nor ( n4592 , n33482 , n33508 );
xor ( n4593 , n33487 , n33499 );
xor ( n4594 , n4593 , n33504 );
buf ( n33512 , n4594 );
xor ( n4596 , n31725 , n2743 );
and ( n4597 , n4596 , n2800 );
and ( n4598 , n31725 , n2743 );
or ( n4599 , n4597 , n4598 );
nor ( n4600 , n33512 , n4599 );
nor ( n4601 , n4592 , n4600 );
not ( n4602 , n4601 );
not ( n4603 , n2253 );
not ( n4604 , n2510 );
or ( n4605 , n4603 , n4604 );
nand ( n4606 , n4605 , n2525 );
not ( n33524 , n2801 );
not ( n4608 , n2809 );
and ( n4609 , n33524 , n4608 );
nor ( n4610 , n2641 , n2650 );
nor ( n4611 , n4609 , n4610 );
nand ( n4612 , n4606 , n4611 );
not ( n4613 , n2810 );
not ( n4614 , n2654 );
or ( n4615 , n4613 , n4614 );
nand ( n4616 , n4615 , n2813 );
nand ( n4617 , n4612 , n4616 );
not ( n4618 , n4617 );
or ( n4619 , n4602 , n4618 );
nand ( n4620 , n33512 , n4599 );
or ( n4621 , n4592 , n4620 );
nand ( n4622 , n33482 , n33508 );
nand ( n4623 , n4621 , n4622 );
not ( n4624 , n4623 );
nand ( n4625 , n4619 , n4624 );
xor ( n4626 , n490 , n491 );
buf ( n33544 , n4626 );
buf ( n33545 , n520 );
and ( n4629 , n33544 , n33545 );
buf ( n33547 , n4629 );
not ( n4631 , n504 );
buf ( n33549 , n506 );
buf ( n33550 , n503 );
xor ( n4634 , n33549 , n33550 );
buf ( n33552 , n4634 );
not ( n4636 , n33552 );
or ( n4637 , n4631 , n4636 );
not ( n4638 , n503 );
nor ( n4639 , n4638 , n504 );
nand ( n4640 , n4281 , n4639 );
nand ( n4641 , n4637 , n4640 );
xor ( n4642 , n33547 , n4641 );
buf ( n33560 , n33356 );
not ( n33561 , n33560 );
buf ( n33562 , n501 );
buf ( n33563 , n502 );
xnor ( n4647 , n33562 , n33563 );
buf ( n33565 , n4647 );
buf ( n33566 , n33565 );
buf ( n33567 , n1907 );
nor ( n4651 , n33566 , n33567 );
buf ( n33569 , n4651 );
buf ( n33570 , n33569 );
not ( n33571 , n33570 );
or ( n4655 , n33561 , n33571 );
buf ( n33573 , n1915 );
xor ( n4657 , n501 , n508 );
buf ( n33575 , n4657 );
nand ( n4659 , n33573 , n33575 );
buf ( n33577 , n4659 );
buf ( n33578 , n33577 );
nand ( n4662 , n4655 , n33578 );
buf ( n33580 , n4662 );
xor ( n4664 , n4642 , n33580 );
buf ( n33582 , n4664 );
buf ( n33583 , n33362 );
not ( n4667 , n33583 );
buf ( n33585 , n33384 );
not ( n33586 , n33585 );
or ( n33587 , n4667 , n33586 );
buf ( n33588 , n33384 );
buf ( n33589 , n33362 );
or ( n4673 , n33588 , n33589 );
buf ( n33591 , n33345 );
nand ( n4675 , n4673 , n33591 );
buf ( n33593 , n4675 );
buf ( n33594 , n33593 );
nand ( n4681 , n33587 , n33594 );
buf ( n33596 , n4681 );
buf ( n33597 , n33596 );
xor ( n4684 , n33582 , n33597 );
xor ( n33599 , n33406 , n33420 );
and ( n4689 , n33599 , n33454 );
and ( n4690 , n33406 , n33420 );
or ( n4691 , n4689 , n4690 );
buf ( n33603 , n4691 );
buf ( n33604 , n33603 );
xor ( n4694 , n4684 , n33604 );
buf ( n33606 , n4694 );
buf ( n33607 , n33606 );
buf ( n33608 , n33399 );
not ( n4698 , n33608 );
buf ( n33610 , n2668 );
not ( n4700 , n33610 );
or ( n4701 , n4698 , n4700 );
buf ( n33613 , n2591 );
xor ( n4703 , n493 , n516 );
buf ( n33615 , n4703 );
nand ( n4705 , n33613 , n33615 );
buf ( n33617 , n4705 );
buf ( n33618 , n33617 );
nand ( n4708 , n4701 , n33618 );
buf ( n33620 , n4708 );
buf ( n33621 , n33620 );
buf ( n33622 , n518 );
buf ( n33623 , n491 );
xor ( n4713 , n33622 , n33623 );
buf ( n33625 , n4713 );
not ( n4715 , n33625 );
not ( n4716 , n4519 );
or ( n4717 , n4715 , n4716 );
nand ( n4718 , n4512 , n33447 );
nand ( n4719 , n4717 , n4718 );
buf ( n33631 , n4719 );
xor ( n4721 , n33621 , n33631 );
and ( n33633 , n4272 , n4283 );
buf ( n33634 , n33633 );
xor ( n4724 , n4721 , n33634 );
buf ( n33636 , n4724 );
buf ( n33637 , n33636 );
buf ( n33638 , n33339 );
not ( n4728 , n33638 );
buf ( n33640 , n2213 );
not ( n4730 , n33640 );
or ( n4731 , n4728 , n4730 );
buf ( n33643 , n2081 );
buf ( n33644 , n512 );
buf ( n33645 , n497 );
xor ( n4735 , n33644 , n33645 );
buf ( n33647 , n4735 );
buf ( n33648 , n33647 );
nand ( n4738 , n33643 , n33648 );
buf ( n33650 , n4738 );
buf ( n33651 , n33650 );
nand ( n4741 , n4731 , n33651 );
buf ( n33653 , n4741 );
buf ( n33654 , n33653 );
not ( n4744 , n2001 );
not ( n4745 , n33415 );
or ( n4746 , n4744 , n4745 );
buf ( n33658 , n31011 );
and ( n4748 , n499 , n510 );
not ( n4749 , n499 );
not ( n4750 , n510 );
and ( n4751 , n4749 , n4750 );
nor ( n4752 , n4748 , n4751 );
buf ( n33664 , n4752 );
nand ( n4754 , n33658 , n33664 );
buf ( n33666 , n4754 );
nand ( n4756 , n4746 , n33666 );
buf ( n33668 , n4756 );
xor ( n4758 , n33654 , n33668 );
xnor ( n4759 , n514 , n495 );
buf ( n33671 , n4759 );
not ( n4761 , n33671 );
buf ( n33673 , n31271 );
nand ( n4763 , n4761 , n33673 );
buf ( n33675 , n4763 );
nand ( n4765 , n2412 , n4452 );
nand ( n4766 , n33675 , n4765 );
buf ( n33678 , n4766 );
xor ( n4768 , n4758 , n33678 );
buf ( n33680 , n4768 );
buf ( n33681 , n33680 );
xor ( n4771 , n33637 , n33681 );
xor ( n4772 , n33220 , n33253 );
and ( n4773 , n4772 , n33305 );
and ( n4774 , n33220 , n33253 );
or ( n33686 , n4773 , n4774 );
buf ( n33687 , n33686 );
buf ( n33688 , n33687 );
xor ( n4778 , n4771 , n33688 );
buf ( n33690 , n4778 );
buf ( n33691 , n33690 );
xor ( n4781 , n33607 , n33691 );
xor ( n4782 , n4466 , n33456 );
and ( n4783 , n4782 , n33478 );
and ( n4784 , n4466 , n33456 );
or ( n4785 , n4783 , n4784 );
buf ( n33697 , n4785 );
xor ( n4787 , n4781 , n33697 );
buf ( n33699 , n4787 );
not ( n4789 , n33699 );
xor ( n4790 , n33308 , n33328 );
and ( n4791 , n4790 , n33480 );
and ( n4792 , n33308 , n33328 );
or ( n4793 , n4791 , n4792 );
buf ( n33705 , n4793 );
not ( n4795 , n33705 );
nor ( n4796 , n4789 , n4795 );
not ( n33708 , n4796 );
not ( n33709 , n33699 );
nand ( n33710 , n33709 , n4795 );
nand ( n4800 , n33708 , n33710 );
not ( n4801 , n4800 );
and ( n4802 , n4625 , n4801 );
not ( n4803 , n4625 );
and ( n4804 , n4803 , n4800 );
nor ( n4805 , n4802 , n4804 );
and ( n33717 , n4805 , n29516 );
not ( n4810 , n33201 );
nor ( n33719 , n33717 , n4810 );
buf ( n33720 , n29681 );
not ( n4813 , n493 );
nand ( n33722 , n4813 , n492 );
not ( n4818 , n492 );
nand ( n4819 , n4818 , n493 );
nand ( n33725 , n33722 , n4819 );
buf ( n4821 , n33725 );
buf ( n33727 , n4821 );
and ( n4823 , n33720 , n33727 );
buf ( n33729 , n4823 );
buf ( n33730 , n33729 );
not ( n33731 , n29671 );
not ( n4827 , n29639 );
or ( n4828 , n33731 , n4827 );
not ( n4829 , n501 );
not ( n4830 , n925 );
or ( n4831 , n4829 , n4830 );
and ( n4832 , n456 , n462 );
not ( n4833 , n456 );
and ( n4834 , n4833 , n478 );
nor ( n4835 , n4832 , n4834 );
not ( n4836 , n4835 );
nand ( n4837 , n4836 , n29635 );
nand ( n4838 , n4831 , n4837 );
nand ( n4839 , n4838 , n29737 );
nand ( n4840 , n4828 , n4839 );
buf ( n33746 , n4840 );
xor ( n4842 , n33730 , n33746 );
buf ( n33748 , n835 );
not ( n4844 , n33748 );
buf ( n33750 , n30102 );
not ( n4846 , n33750 );
or ( n4847 , n4844 , n4846 );
not ( n4848 , n497 );
not ( n4849 , n29610 );
or ( n4850 , n4848 , n4849 );
nand ( n4851 , n706 , n1261 );
nand ( n4852 , n4850 , n4851 );
buf ( n33758 , n4852 );
buf ( n33759 , n29829 );
nand ( n4855 , n33758 , n33759 );
buf ( n33761 , n4855 );
buf ( n33762 , n33761 );
nand ( n4858 , n4847 , n33762 );
buf ( n33764 , n4858 );
buf ( n33765 , n33764 );
xor ( n4861 , n4842 , n33765 );
buf ( n33767 , n4861 );
not ( n4863 , n29580 );
not ( n4864 , n29628 );
or ( n33770 , n4863 , n4864 );
not ( n4866 , n29580 );
not ( n4867 , n4866 );
not ( n4868 , n29628 );
not ( n4869 , n4868 );
or ( n4870 , n4867 , n4869 );
nand ( n4871 , n4870 , n29704 );
nand ( n4872 , n33770 , n4871 );
xor ( n4873 , n33767 , n4872 );
not ( n4874 , n29844 );
not ( n4875 , n1035 );
or ( n4876 , n4874 , n4875 );
buf ( n33782 , n495 );
not ( n4878 , n33782 );
buf ( n33784 , n29493 );
not ( n33785 , n33784 );
buf ( n33786 , n33785 );
buf ( n33787 , n33786 );
not ( n4883 , n33787 );
or ( n4884 , n4878 , n4883 );
buf ( n33790 , n29493 );
buf ( n33791 , n29716 );
nand ( n4887 , n33790 , n33791 );
buf ( n33793 , n4887 );
buf ( n33794 , n33793 );
nand ( n33795 , n4884 , n33794 );
buf ( n33796 , n33795 );
buf ( n33797 , n33796 );
buf ( n33798 , n29873 );
nand ( n4894 , n33797 , n33798 );
buf ( n33800 , n4894 );
nand ( n4896 , n4876 , n33800 );
not ( n4897 , n4896 );
not ( n4898 , n504 );
or ( n4899 , n456 , n476 );
not ( n4900 , n460 );
nand ( n4901 , n4900 , n456 );
nand ( n4902 , n4899 , n863 , n4901 );
and ( n4903 , n456 , n460 );
not ( n4904 , n456 );
and ( n4905 , n4904 , n476 );
nor ( n4906 , n4903 , n4905 );
nand ( n4907 , n4906 , n503 );
nand ( n4908 , n4902 , n4907 );
not ( n4909 , n4908 );
or ( n4910 , n4898 , n4909 );
not ( n4911 , n945 );
nand ( n4912 , n1006 , n4911 );
nand ( n4913 , n4910 , n4912 );
not ( n4914 , n4913 );
not ( n4915 , n4914 );
or ( n4916 , n4897 , n4915 );
or ( n4917 , n4914 , n4896 );
nand ( n4918 , n4916 , n4917 );
buf ( n33824 , n29576 );
not ( n4920 , n33824 );
buf ( n33826 , n29543 );
not ( n4922 , n33826 );
or ( n4923 , n4920 , n4922 );
buf ( n33829 , n493 );
not ( n4925 , n33829 );
buf ( n33831 , n820 );
not ( n4927 , n33831 );
or ( n4928 , n4925 , n4927 );
or ( n4929 , n456 , n486 );
nand ( n4930 , n3859 , n456 );
nand ( n4931 , n4929 , n29537 , n4930 );
buf ( n33837 , n4931 );
nand ( n4933 , n4928 , n33837 );
buf ( n33839 , n4933 );
buf ( n33840 , n33839 );
buf ( n33841 , n29522 );
nand ( n33842 , n33840 , n33841 );
buf ( n33843 , n33842 );
buf ( n33844 , n33843 );
nand ( n4940 , n4923 , n33844 );
buf ( n33846 , n4940 );
and ( n4942 , n4918 , n33846 );
not ( n4943 , n4918 );
not ( n4944 , n33846 );
and ( n33850 , n4943 , n4944 );
nor ( n4949 , n4942 , n33850 );
xor ( n33852 , n4873 , n4949 );
not ( n4951 , n33852 );
not ( n4952 , n4951 );
buf ( n33855 , n29624 );
not ( n4957 , n33855 );
buf ( n33857 , n29602 );
not ( n4959 , n33857 );
or ( n4960 , n4957 , n4959 );
buf ( n33860 , n499 );
not ( n4962 , n33860 );
and ( n4963 , n456 , n464 );
not ( n4964 , n456 );
and ( n4965 , n4964 , n480 );
nor ( n4966 , n4963 , n4965 );
buf ( n33866 , n4966 );
not ( n4968 , n33866 );
or ( n4969 , n4962 , n4968 );
buf ( n33869 , n29925 );
buf ( n33870 , n29596 );
nand ( n4972 , n33869 , n33870 );
buf ( n33872 , n4972 );
buf ( n33873 , n33872 );
nand ( n4975 , n4969 , n33873 );
buf ( n33875 , n4975 );
buf ( n33876 , n33875 );
buf ( n33877 , n29583 );
nand ( n4979 , n33876 , n33877 );
buf ( n33879 , n4979 );
buf ( n33880 , n33879 );
nand ( n4982 , n4960 , n33880 );
buf ( n33882 , n4982 );
buf ( n33883 , n33882 );
buf ( n33884 , n29673 );
not ( n4986 , n33884 );
buf ( n33886 , n29703 );
nor ( n4988 , n4986 , n33886 );
buf ( n33888 , n4988 );
buf ( n33889 , n33888 );
xor ( n4991 , n33883 , n33889 );
xor ( n4992 , n30069 , n30087 );
and ( n4993 , n4992 , n30113 );
and ( n4994 , n30069 , n30087 );
or ( n4995 , n4993 , n4994 );
buf ( n33895 , n4995 );
buf ( n33896 , n33895 );
xor ( n4998 , n4991 , n33896 );
buf ( n33898 , n4998 );
not ( n33899 , n33898 );
xor ( n5001 , n897 , n30047 );
and ( n5002 , n5001 , n30115 );
and ( n5003 , n897 , n30047 );
or ( n5004 , n5002 , n5003 );
not ( n5005 , n5004 );
not ( n5006 , n5005 );
or ( n5007 , n33899 , n5006 );
not ( n5008 , n33898 );
nand ( n5009 , n5008 , n5004 );
nand ( n5010 , n5007 , n5009 );
not ( n5011 , n5010 );
nand ( n5012 , n4952 , n5011 );
nand ( n5013 , n5010 , n4951 );
xor ( n5014 , n29705 , n892 );
and ( n33914 , n5014 , n1067 );
and ( n5016 , n29705 , n892 );
or ( n5017 , n33914 , n5016 );
not ( n5018 , n5017 );
and ( n5019 , n5012 , n5013 , n5018 );
buf ( n33919 , n4508 );
not ( n33920 , n33919 );
buf ( n33921 , n29691 );
not ( n5023 , n33921 );
or ( n5024 , n33920 , n5023 );
buf ( n33924 , n493 );
nand ( n5026 , n5024 , n33924 );
buf ( n33926 , n5026 );
buf ( n33927 , n33926 );
buf ( n33928 , n29855 );
not ( n5030 , n33928 );
buf ( n33930 , n5030 );
buf ( n33931 , n33930 );
buf ( n33932 , n492 );
and ( n5034 , n33931 , n33932 );
buf ( n33934 , n491 );
not ( n5036 , n33934 );
buf ( n33936 , n5036 );
buf ( n33937 , n33936 );
nor ( n5039 , n5034 , n33937 );
buf ( n33939 , n5039 );
buf ( n33940 , n33939 );
nand ( n5042 , n33927 , n33940 );
buf ( n33942 , n5042 );
buf ( n33943 , n33942 );
not ( n5045 , n33943 );
buf ( n33945 , n847 );
not ( n5047 , n33945 );
buf ( n33947 , n4908 );
not ( n5049 , n33947 );
or ( n5050 , n5047 , n5049 );
and ( n5051 , n456 , n459 );
not ( n5052 , n456 );
and ( n5053 , n5052 , n475 );
nor ( n5054 , n5051 , n5053 );
nand ( n5055 , n5054 , n503 );
not ( n5056 , n5055 );
not ( n5057 , n459 );
and ( n5058 , n456 , n5057 );
not ( n5059 , n456 );
not ( n5060 , n475 );
and ( n5061 , n5059 , n5060 );
nor ( n5062 , n5058 , n5061 );
buf ( n33962 , n5062 );
buf ( n33963 , n863 );
nand ( n5065 , n33962 , n33963 );
buf ( n33965 , n5065 );
not ( n5067 , n33965 );
or ( n5068 , n5056 , n5067 );
nand ( n5069 , n5068 , n504 );
buf ( n33969 , n5069 );
nand ( n5071 , n5050 , n33969 );
buf ( n33971 , n5071 );
buf ( n33972 , n33971 );
not ( n5074 , n33972 );
or ( n5075 , n5045 , n5074 );
buf ( n33975 , n33971 );
buf ( n33976 , n33942 );
or ( n5078 , n33975 , n33976 );
nand ( n5079 , n5075 , n5078 );
buf ( n33979 , n5079 );
buf ( n33980 , n33979 );
nor ( n5082 , n4896 , n4913 );
or ( n5083 , n4944 , n5082 );
nand ( n5084 , n4896 , n4913 );
nand ( n33984 , n5083 , n5084 );
buf ( n33985 , n33984 );
xor ( n33986 , n33980 , n33985 );
xor ( n5088 , n33730 , n33746 );
and ( n5089 , n5088 , n33765 );
and ( n5090 , n33730 , n33746 );
or ( n5091 , n5089 , n5090 );
buf ( n33991 , n5091 );
buf ( n33992 , n33991 );
xor ( n33993 , n33986 , n33992 );
buf ( n33994 , n33993 );
xor ( n33995 , n33767 , n4872 );
and ( n5100 , n33995 , n4949 );
and ( n5101 , n33767 , n4872 );
or ( n33998 , n5100 , n5101 );
xor ( n5106 , n33994 , n33998 );
buf ( n34000 , n29522 );
not ( n5108 , n34000 );
buf ( n34002 , n493 );
not ( n5110 , n34002 );
buf ( n34004 , n1033 );
not ( n34005 , n34004 );
or ( n5113 , n5110 , n34005 );
buf ( n34007 , n712 );
buf ( n34008 , n29537 );
nand ( n5116 , n34007 , n34008 );
buf ( n34010 , n5116 );
buf ( n34011 , n34010 );
nand ( n5119 , n5113 , n34011 );
buf ( n34013 , n5119 );
buf ( n34014 , n34013 );
not ( n34015 , n34014 );
or ( n5123 , n5108 , n34015 );
nand ( n5124 , n33839 , n29576 );
buf ( n34018 , n5124 );
nand ( n5126 , n5123 , n34018 );
buf ( n34020 , n5126 );
buf ( n34021 , n34020 );
and ( n5129 , n491 , n492 );
not ( n5130 , n491 );
not ( n5131 , n492 );
and ( n5132 , n5130 , n5131 );
nor ( n5133 , n5129 , n5132 );
not ( n5134 , n5133 );
nor ( n5135 , n33725 , n5134 );
buf ( n34029 , n5135 );
buf ( n5137 , n34029 );
buf ( n34031 , n5137 );
buf ( n34032 , n34031 );
not ( n5140 , n34032 );
buf ( n34034 , n33936 );
buf ( n34035 , n29551 );
and ( n5143 , n34034 , n34035 );
not ( n5144 , n34034 );
buf ( n34038 , n29764 );
and ( n5146 , n5144 , n34038 );
nor ( n5147 , n5143 , n5146 );
buf ( n34041 , n5147 );
buf ( n34042 , n34041 );
not ( n5150 , n34042 );
or ( n5151 , n5140 , n5150 );
buf ( n34045 , n491 );
not ( n5153 , n34045 );
buf ( n34047 , n1484 );
not ( n5155 , n34047 );
or ( n5156 , n5153 , n5155 );
buf ( n34050 , n29535 );
buf ( n34051 , n33936 );
nand ( n5159 , n34050 , n34051 );
buf ( n34053 , n5159 );
buf ( n34054 , n34053 );
nand ( n5162 , n5156 , n34054 );
buf ( n34056 , n5162 );
buf ( n34057 , n34056 );
buf ( n34058 , n4821 );
nand ( n5166 , n34057 , n34058 );
buf ( n34060 , n5166 );
buf ( n34061 , n34060 );
nand ( n5169 , n5151 , n34061 );
buf ( n34063 , n5169 );
buf ( n34064 , n34063 );
xor ( n5172 , n34021 , n34064 );
buf ( n34066 , n29624 );
not ( n5174 , n34066 );
buf ( n34068 , n33875 );
not ( n5176 , n34068 );
or ( n5177 , n5174 , n5176 );
buf ( n34071 , n29505 );
not ( n5179 , n34071 );
buf ( n34073 , n5179 );
nand ( n5181 , n34073 , n499 );
not ( n5182 , n5181 );
not ( n5183 , n29631 );
nand ( n5184 , n5183 , n29596 );
not ( n5185 , n5184 );
or ( n5186 , n5182 , n5185 );
nand ( n5187 , n5186 , n1627 );
buf ( n34081 , n5187 );
nand ( n5189 , n5177 , n34081 );
buf ( n34083 , n5189 );
buf ( n34084 , n34083 );
xor ( n5192 , n5172 , n34084 );
buf ( n34086 , n5192 );
buf ( n34087 , n34086 );
not ( n5195 , n29873 );
buf ( n34089 , n495 );
not ( n5197 , n34089 );
buf ( n34091 , n971 );
not ( n5199 , n34091 );
or ( n5200 , n5197 , n5199 );
buf ( n34094 , n1204 );
buf ( n34095 , n29716 );
nand ( n5203 , n34094 , n34095 );
buf ( n34097 , n5203 );
buf ( n34098 , n34097 );
nand ( n5206 , n5200 , n34098 );
buf ( n34100 , n5206 );
not ( n5208 , n34100 );
or ( n5209 , n5195 , n5208 );
buf ( n34103 , n495 );
not ( n5211 , n34103 );
buf ( n34105 , n33786 );
not ( n5213 , n34105 );
or ( n5214 , n5211 , n5213 );
buf ( n34108 , n33793 );
nand ( n5216 , n5214 , n34108 );
buf ( n34110 , n5216 );
nand ( n5218 , n34110 , n29844 );
nand ( n34112 , n5209 , n5218 );
not ( n5220 , n29647 );
buf ( n34114 , n501 );
not ( n5222 , n34114 );
and ( n5223 , n456 , n461 );
not ( n34117 , n456 );
and ( n5225 , n34117 , n477 );
nor ( n5226 , n5223 , n5225 );
buf ( n34120 , n5226 );
not ( n5228 , n34120 );
or ( n34122 , n5222 , n5228 );
buf ( n34123 , n29511 );
buf ( n34124 , n29635 );
nand ( n5232 , n34123 , n34124 );
buf ( n34126 , n5232 );
buf ( n34127 , n34126 );
nand ( n5235 , n34122 , n34127 );
buf ( n34129 , n5235 );
not ( n5237 , n34129 );
or ( n5238 , n5220 , n5237 );
nand ( n5239 , n4838 , n29671 );
nand ( n5240 , n5238 , n5239 );
xor ( n5241 , n34112 , n5240 );
not ( n5242 , n835 );
not ( n5243 , n4852 );
or ( n34137 , n5242 , n5243 );
buf ( n34138 , n497 );
not ( n34139 , n34138 );
buf ( n34140 , n1147 );
not ( n5248 , n34140 );
or ( n5249 , n34139 , n5248 );
buf ( n34143 , n29749 );
buf ( n34144 , n706 );
nand ( n5252 , n34143 , n34144 );
buf ( n34146 , n5252 );
buf ( n34147 , n34146 );
nand ( n34148 , n5249 , n34147 );
buf ( n34149 , n34148 );
buf ( n34150 , n34149 );
buf ( n34151 , n29829 );
nand ( n5265 , n34150 , n34151 );
buf ( n34153 , n5265 );
nand ( n5267 , n34137 , n34153 );
xor ( n5268 , n5241 , n5267 );
buf ( n34156 , n5268 );
xor ( n5270 , n34087 , n34156 );
xor ( n34158 , n33883 , n33889 );
and ( n5272 , n34158 , n33896 );
and ( n5273 , n33883 , n33889 );
or ( n5274 , n5272 , n5273 );
buf ( n34162 , n5274 );
buf ( n34163 , n34162 );
xor ( n5277 , n5270 , n34163 );
buf ( n34165 , n5277 );
xor ( n5279 , n5106 , n34165 );
nand ( n5280 , n5005 , n5008 );
not ( n5281 , n5280 );
not ( n5282 , n33852 );
or ( n5283 , n5281 , n5282 );
nand ( n5284 , n5004 , n33898 );
nand ( n5285 , n5283 , n5284 );
nor ( n5286 , n5279 , n5285 );
nor ( n5287 , n5019 , n5286 );
not ( n5288 , n5287 );
not ( n5289 , n30232 );
not ( n5290 , n30340 );
nand ( n5291 , n5289 , n5290 );
nand ( n5292 , n1069 , n1181 );
nand ( n5293 , n5291 , n5292 , n1808 , n1473 );
nand ( n5294 , n30493 , n5292 , n5291 );
not ( n5295 , n1813 );
not ( n5296 , n1183 );
or ( n5297 , n5295 , n5296 );
nand ( n5298 , n5297 , n1182 );
nand ( n5299 , n5293 , n5294 , n5298 );
not ( n5300 , n5299 );
or ( n5301 , n5288 , n5300 );
nand ( n34189 , n5279 , n5285 );
not ( n5303 , n34189 );
nand ( n5304 , n5011 , n4951 );
nand ( n5305 , n5010 , n33852 );
nand ( n5306 , n5304 , n5305 , n5017 );
not ( n5307 , n5306 );
or ( n5308 , n5303 , n5307 );
not ( n5309 , n5286 );
nand ( n5310 , n5308 , n5309 );
buf ( n5311 , n5310 );
nand ( n5312 , n5301 , n5311 );
buf ( n34200 , n5240 );
not ( n5314 , n34200 );
buf ( n34202 , n5314 );
not ( n5316 , n34202 );
buf ( n34204 , n34112 );
not ( n34205 , n34204 );
buf ( n34206 , n34205 );
not ( n5320 , n34206 );
and ( n5321 , n5316 , n5320 );
nand ( n5322 , n34206 , n34202 );
and ( n5323 , n5322 , n5267 );
nor ( n5324 , n5321 , n5323 );
buf ( n34212 , n5324 );
not ( n5326 , n34212 );
buf ( n34214 , n29678 );
xor ( n5328 , n490 , n491 );
buf ( n34216 , n5328 );
and ( n5330 , n34214 , n34216 );
buf ( n34218 , n5330 );
not ( n5332 , n4911 );
nand ( n5333 , n33965 , n5055 );
not ( n5334 , n5333 );
or ( n5335 , n5332 , n5334 );
not ( n5336 , n503 );
not ( n5337 , n29498 );
or ( n5338 , n5336 , n5337 );
buf ( n34226 , n29499 );
buf ( n34227 , n863 );
nand ( n5341 , n34226 , n34227 );
buf ( n34229 , n5341 );
nand ( n5343 , n5338 , n34229 );
nand ( n5344 , n504 , n5343 );
nand ( n5345 , n5335 , n5344 );
xor ( n34233 , n34218 , n5345 );
buf ( n34234 , n29671 );
not ( n5348 , n34234 );
buf ( n34236 , n34129 );
not ( n5350 , n34236 );
or ( n5351 , n5348 , n5350 );
nand ( n5352 , n4906 , n501 );
not ( n5353 , n5352 );
not ( n5354 , n501 );
not ( n5355 , n460 );
and ( n5356 , n5355 , n456 );
nor ( n5357 , n456 , n476 );
nor ( n5358 , n5356 , n5357 );
nand ( n5359 , n5354 , n5358 );
not ( n5360 , n5359 );
or ( n5361 , n5353 , n5360 );
nand ( n34249 , n5361 , n29647 );
buf ( n34250 , n34249 );
nand ( n5364 , n5351 , n34250 );
buf ( n34252 , n5364 );
xnor ( n34253 , n34233 , n34252 );
buf ( n34254 , n34253 );
not ( n5368 , n34254 );
buf ( n34256 , n5368 );
buf ( n34257 , n34256 );
not ( n5371 , n34257 );
or ( n5372 , n5326 , n5371 );
buf ( n34260 , n5324 );
buf ( n34261 , n34256 );
or ( n5375 , n34260 , n34261 );
nand ( n5376 , n5372 , n5375 );
buf ( n34264 , n5376 );
buf ( n34265 , n34264 );
xor ( n5379 , n34021 , n34064 );
and ( n5380 , n5379 , n34084 );
and ( n5381 , n34021 , n34064 );
or ( n5382 , n5380 , n5381 );
buf ( n34270 , n5382 );
buf ( n34271 , n34270 );
and ( n5385 , n34265 , n34271 );
not ( n5386 , n34265 );
buf ( n34274 , n34270 );
not ( n5388 , n34274 );
buf ( n34276 , n5388 );
buf ( n34277 , n34276 );
and ( n5391 , n5386 , n34277 );
nor ( n5392 , n5385 , n5391 );
buf ( n34280 , n5392 );
xor ( n5394 , n34087 , n34156 );
and ( n5395 , n5394 , n34163 );
and ( n5396 , n34087 , n34156 );
or ( n5397 , n5395 , n5396 );
buf ( n34285 , n5397 );
xor ( n5399 , n34280 , n34285 );
buf ( n34287 , n4821 );
not ( n5401 , n34287 );
buf ( n34289 , n491 );
not ( n5403 , n34289 );
buf ( n34291 , n820 );
not ( n5405 , n34291 );
or ( n5406 , n5403 , n5405 );
buf ( n34294 , n901 );
buf ( n34295 , n33936 );
nand ( n5409 , n34294 , n34295 );
buf ( n34297 , n5409 );
buf ( n34298 , n34297 );
nand ( n5412 , n5406 , n34298 );
buf ( n34300 , n5412 );
buf ( n34301 , n34300 );
not ( n34302 , n34301 );
or ( n5416 , n5401 , n34302 );
buf ( n34304 , n34056 );
buf ( n34305 , n34031 );
nand ( n5419 , n34304 , n34305 );
buf ( n34307 , n5419 );
buf ( n34308 , n34307 );
nand ( n34309 , n5416 , n34308 );
buf ( n34310 , n34309 );
buf ( n34311 , n34310 );
not ( n5428 , n29576 );
not ( n5429 , n34013 );
or ( n34314 , n5428 , n5429 );
not ( n5434 , n493 );
not ( n5435 , n1364 );
or ( n5436 , n5434 , n5435 );
not ( n5437 , n468 );
nand ( n5438 , n5437 , n456 );
not ( n5439 , n484 );
not ( n5440 , n456 );
nand ( n5441 , n5439 , n5440 );
nand ( n5442 , n5438 , n5441 , n29537 );
nand ( n5443 , n5436 , n5442 );
buf ( n34325 , n5443 );
buf ( n34326 , n29522 );
nand ( n5446 , n34325 , n34326 );
buf ( n34328 , n5446 );
nand ( n5448 , n34314 , n34328 );
buf ( n34330 , n5448 );
xor ( n5450 , n34311 , n34330 );
not ( n5451 , n847 );
not ( n5452 , n4908 );
or ( n5453 , n5451 , n5452 );
nand ( n5454 , n5453 , n5069 );
not ( n5455 , n5454 );
nor ( n5456 , n5455 , n33942 );
buf ( n34338 , n5456 );
xor ( n5458 , n5450 , n34338 );
buf ( n34340 , n5458 );
buf ( n34341 , n34340 );
buf ( n34342 , n29829 );
not ( n5462 , n34342 );
buf ( n34344 , n497 );
not ( n5464 , n34344 );
buf ( n34346 , n4966 );
not ( n5466 , n34346 );
or ( n5467 , n5464 , n5466 );
buf ( n34349 , n29658 );
buf ( n34350 , n706 );
nand ( n5470 , n34349 , n34350 );
buf ( n34352 , n5470 );
buf ( n34353 , n34352 );
nand ( n5473 , n5467 , n34353 );
buf ( n34355 , n5473 );
buf ( n34356 , n34355 );
not ( n5476 , n34356 );
or ( n5477 , n5462 , n5476 );
and ( n5478 , n29749 , n706 );
not ( n5479 , n29749 );
and ( n5480 , n5479 , n497 );
or ( n5481 , n5478 , n5480 );
nand ( n5482 , n5481 , n29786 );
buf ( n34364 , n5482 );
nand ( n5484 , n5477 , n34364 );
buf ( n34366 , n5484 );
buf ( n34367 , n29844 );
not ( n5487 , n34367 );
buf ( n34369 , n34100 );
not ( n5489 , n34369 );
or ( n5490 , n5487 , n5489 );
buf ( n34372 , n495 );
not ( n5492 , n34372 );
buf ( n34374 , n29731 );
not ( n5494 , n34374 );
or ( n5495 , n5492 , n5494 );
buf ( n34377 , n29613 );
buf ( n34378 , n29716 );
nand ( n5498 , n34377 , n34378 );
buf ( n34380 , n5498 );
buf ( n34381 , n34380 );
nand ( n34382 , n5495 , n34381 );
buf ( n34383 , n34382 );
buf ( n34384 , n34383 );
buf ( n34385 , n29873 );
nand ( n5505 , n34384 , n34385 );
buf ( n34387 , n5505 );
buf ( n34388 , n34387 );
nand ( n5508 , n5490 , n34388 );
buf ( n34390 , n5508 );
xor ( n5510 , n34366 , n34390 );
buf ( n34392 , n5510 );
nand ( n5512 , n5181 , n5184 );
and ( n5513 , n29624 , n5512 );
not ( n5514 , n499 );
not ( n5515 , n925 );
or ( n5516 , n5514 , n5515 );
and ( n5517 , n5440 , n930 );
and ( n5518 , n932 , n456 );
nor ( n5519 , n5517 , n5518 );
nand ( n5520 , n5519 , n29596 );
nand ( n5521 , n5516 , n5520 );
and ( n5522 , n5521 , n1627 );
nor ( n5523 , n5513 , n5522 );
buf ( n34405 , n5523 );
xnor ( n5525 , n34392 , n34405 );
buf ( n34407 , n5525 );
buf ( n34408 , n34407 );
xor ( n5528 , n34341 , n34408 );
xor ( n5529 , n33980 , n33985 );
and ( n5530 , n5529 , n33992 );
and ( n5531 , n33980 , n33985 );
or ( n5532 , n5530 , n5531 );
buf ( n34414 , n5532 );
buf ( n34415 , n34414 );
xor ( n5535 , n5528 , n34415 );
buf ( n34417 , n5535 );
xor ( n5537 , n5399 , n34417 );
not ( n5538 , n5537 );
xor ( n5539 , n33994 , n33998 );
and ( n5540 , n5539 , n34165 );
and ( n5541 , n33994 , n33998 );
or ( n5542 , n5540 , n5541 );
not ( n5543 , n5542 );
nor ( n5544 , n5538 , n5543 );
not ( n5545 , n5544 );
not ( n5546 , n5537 );
nand ( n5547 , n5546 , n5543 );
nand ( n5548 , n5545 , n5547 );
not ( n5549 , n5548 );
and ( n5550 , n5312 , n5549 );
not ( n5551 , n5312 );
and ( n5552 , n5551 , n5548 );
nor ( n5553 , n5550 , n5552 );
nand ( n5554 , n5553 , n455 );
nand ( n5555 , n33719 , n5554 );
not ( n5556 , n5555 );
or ( n5557 , n4268 , n5556 );
not ( n5558 , n541 );
not ( n5559 , n454 );
or ( n5560 , n5558 , n5559 );
xor ( n5561 , n33113 , n33143 );
and ( n5562 , n5561 , n33172 );
and ( n5563 , n33113 , n33143 );
or ( n5564 , n5562 , n5563 );
buf ( n34446 , n5564 );
buf ( n34447 , n34446 );
xor ( n5567 , n33123 , n33124 );
and ( n5568 , n5567 , n33140 );
and ( n5569 , n33123 , n33124 );
or ( n5570 , n5568 , n5569 );
buf ( n34452 , n5570 );
buf ( n34453 , n34452 );
nand ( n5573 , n32981 , n542 );
not ( n5574 , n542 );
nand ( n5575 , n5574 , n543 );
and ( n5576 , n542 , n541 );
not ( n5577 , n542 );
not ( n5578 , n541 );
and ( n5579 , n5577 , n5578 );
nor ( n5580 , n5576 , n5579 );
nand ( n5581 , n5573 , n5575 , n5580 );
buf ( n5582 , n5581 );
buf ( n34464 , n5582 );
buf ( n34465 , n541 );
buf ( n34466 , n32059 );
and ( n5586 , n34465 , n34466 );
not ( n5587 , n34465 );
buf ( n34469 , n536 );
and ( n5589 , n5587 , n34469 );
nor ( n34471 , n5586 , n5589 );
buf ( n34472 , n34471 );
buf ( n34473 , n34472 );
or ( n5596 , n34464 , n34473 );
buf ( n34475 , n33118 );
buf ( n34476 , n541 );
buf ( n34477 , n32074 );
and ( n5603 , n34476 , n34477 );
not ( n5604 , n34476 );
buf ( n34480 , n535 );
and ( n5606 , n5604 , n34480 );
nor ( n5607 , n5603 , n5606 );
buf ( n34483 , n5607 );
buf ( n34484 , n34483 );
or ( n5610 , n34475 , n34484 );
nand ( n5611 , n5596 , n5610 );
buf ( n34487 , n5611 );
buf ( n34488 , n34487 );
xor ( n5614 , n34453 , n34488 );
xor ( n5615 , n33081 , n33084 );
and ( n5616 , n5615 , n33110 );
and ( n5617 , n33081 , n33084 );
or ( n5618 , n5616 , n5617 );
buf ( n34494 , n5618 );
buf ( n34495 , n34494 );
xor ( n5621 , n5614 , n34495 );
buf ( n34497 , n5621 );
buf ( n34498 , n34497 );
xor ( n5624 , n34447 , n34498 );
or ( n5625 , n3069 , n33105 );
buf ( n34501 , n545 );
buf ( n34502 , n31840 );
and ( n34503 , n34501 , n34502 );
not ( n5629 , n34501 );
buf ( n34505 , n531 );
and ( n5631 , n5629 , n34505 );
nor ( n5632 , n34503 , n5631 );
buf ( n34508 , n5632 );
or ( n5634 , n34508 , n3087 );
nand ( n5635 , n5625 , n5634 );
buf ( n5636 , n4214 );
buf ( n34512 , n5636 );
buf ( n34513 , n32996 );
or ( n5639 , n34512 , n34513 );
buf ( n34515 , n4040 );
buf ( n34516 , n543 );
buf ( n34517 , n31874 );
and ( n5643 , n34516 , n34517 );
not ( n5644 , n34516 );
buf ( n34520 , n533 );
and ( n5646 , n5644 , n34520 );
nor ( n5647 , n5643 , n5646 );
buf ( n34523 , n5647 );
buf ( n34524 , n34523 );
or ( n5650 , n34515 , n34524 );
nand ( n5651 , n5639 , n5650 );
buf ( n34527 , n5651 );
xor ( n34528 , n5635 , n34527 );
buf ( n34529 , n3045 );
buf ( n34530 , n32965 );
or ( n5656 , n34529 , n34530 );
buf ( n34532 , n2918 );
buf ( n34533 , n31868 );
buf ( n34534 , n527 );
and ( n5660 , n34533 , n34534 );
buf ( n34536 , n33009 );
buf ( n34537 , n549 );
and ( n5663 , n34536 , n34537 );
nor ( n5664 , n5660 , n5663 );
buf ( n34540 , n5664 );
buf ( n34541 , n34540 );
or ( n5667 , n34532 , n34541 );
nand ( n5668 , n5656 , n5667 );
buf ( n34544 , n5668 );
xor ( n5670 , n34528 , n34544 );
buf ( n34546 , n33129 );
not ( n5672 , n34546 );
buf ( n34548 , n3199 );
not ( n5674 , n34548 );
or ( n5675 , n5672 , n5674 );
buf ( n34551 , n551 );
buf ( n34552 , n525 );
and ( n5678 , n34551 , n34552 );
not ( n5679 , n34551 );
buf ( n34555 , n525 );
not ( n5681 , n34555 );
buf ( n34557 , n5681 );
buf ( n34558 , n34557 );
and ( n5684 , n5679 , n34558 );
nor ( n5685 , n5678 , n5684 );
buf ( n34561 , n5685 );
buf ( n34562 , n34561 );
buf ( n34563 , n552 );
nand ( n5689 , n34562 , n34563 );
buf ( n34565 , n5689 );
buf ( n34566 , n34565 );
nand ( n5692 , n5675 , n34566 );
buf ( n34568 , n5692 );
buf ( n34569 , n34568 );
buf ( n34570 , n461 );
buf ( n34571 , n536 );
buf ( n34572 , n542 );
or ( n5698 , n34571 , n34572 );
buf ( n34574 , n543 );
nand ( n5700 , n5698 , n34574 );
buf ( n34576 , n5700 );
buf ( n34577 , n34576 );
buf ( n34578 , n536 );
buf ( n34579 , n542 );
nand ( n5705 , n34578 , n34579 );
buf ( n34581 , n5705 );
buf ( n34582 , n34581 );
buf ( n34583 , n541 );
and ( n5709 , n34577 , n34582 , n34583 );
buf ( n34585 , n5709 );
buf ( n34586 , n34585 );
xor ( n5712 , n34570 , n34586 );
buf ( n34588 , n5712 );
buf ( n34589 , n34588 );
xor ( n5715 , n34569 , n34589 );
or ( n5716 , n33076 , n3020 );
not ( n5717 , n31988 );
and ( n5718 , n547 , n529 );
not ( n5719 , n547 );
and ( n5720 , n5719 , n2969 );
nor ( n5721 , n5718 , n5720 );
nand ( n5722 , n5717 , n5721 );
nand ( n5723 , n5716 , n5722 );
buf ( n34599 , n5723 );
xor ( n5725 , n5715 , n34599 );
buf ( n34601 , n5725 );
xor ( n5727 , n32970 , n33001 );
and ( n5728 , n5727 , n33061 );
and ( n5729 , n32970 , n33001 );
or ( n5730 , n5728 , n5729 );
buf ( n34606 , n5730 );
xor ( n5732 , n34601 , n34606 );
xor ( n5733 , n5670 , n5732 );
buf ( n34609 , n5733 );
xor ( n5735 , n5624 , n34609 );
buf ( n34611 , n5735 );
buf ( n34612 , n34611 );
buf ( n34613 , n3360 );
nand ( n5739 , n34612 , n34613 );
buf ( n34615 , n5739 );
nand ( n5741 , n5560 , n34615 );
not ( n5742 , n5741 );
nand ( n5743 , n5557 , n5742 );
not ( n5744 , n542 );
not ( n34620 , n454 );
or ( n34621 , n5744 , n34620 );
xor ( n5747 , n33064 , n33175 );
xor ( n5748 , n5747 , n33193 );
buf ( n34624 , n5748 );
buf ( n34625 , n34624 );
buf ( n34626 , n3360 );
nand ( n5755 , n34625 , n34626 );
buf ( n34628 , n5755 );
nand ( n34629 , n34621 , n34628 );
not ( n5761 , n34629 );
or ( n5762 , n33512 , n4599 );
not ( n5763 , n5762 );
not ( n5764 , n4617 );
or ( n5765 , n5763 , n5764 );
nand ( n5766 , n5765 , n4620 );
not ( n34636 , n4592 );
nand ( n5768 , n34636 , n4622 );
not ( n5769 , n5768 );
and ( n5770 , n5766 , n5769 );
not ( n5771 , n5766 );
and ( n5772 , n5771 , n5768 );
nor ( n34642 , n5770 , n5772 );
and ( n5774 , n2815 , n454 );
and ( n5775 , n34642 , n5774 );
xor ( n5776 , n32169 , n464 );
xor ( n5777 , n5776 , n32195 );
and ( n5778 , n32212 , n5777 );
xor ( n5779 , n32169 , n464 );
xor ( n5780 , n5779 , n32195 );
and ( n5781 , n32217 , n5780 );
and ( n5782 , n32212 , n32217 );
or ( n5783 , n5778 , n5781 , n5782 );
buf ( n34653 , n5783 );
xor ( n5785 , n33153 , n33162 );
xor ( n5786 , n5785 , n33167 );
buf ( n34656 , n5786 );
buf ( n34657 , n34656 );
xor ( n5789 , n34653 , n34657 );
xor ( n5790 , n33021 , n33040 );
xor ( n5791 , n5790 , n33057 );
xor ( n5792 , n4239 , n4249 );
xor ( n5793 , n5791 , n5792 );
buf ( n34663 , n5793 );
and ( n5795 , n5789 , n34663 );
and ( n5796 , n34653 , n34657 );
or ( n5797 , n5795 , n5796 );
buf ( n34667 , n5797 );
and ( n5799 , n34667 , n3138 );
nor ( n5800 , n5775 , n5799 );
not ( n5801 , n5019 );
not ( n5802 , n5801 );
nand ( n5803 , n5293 , n5294 , n5298 );
not ( n5804 , n5803 );
or ( n5805 , n5802 , n5804 );
buf ( n5806 , n5306 );
nand ( n5807 , n5805 , n5806 );
nand ( n5808 , n5309 , n34189 );
not ( n5809 , n5808 );
and ( n5810 , n5807 , n5809 );
not ( n5811 , n5807 );
and ( n5812 , n5811 , n5808 );
nor ( n5813 , n5810 , n5812 );
nand ( n5814 , n5813 , n455 , n454 );
nand ( n5815 , n5761 , n5800 , n5814 );
not ( n5816 , n454 );
not ( n5817 , n2815 );
nand ( n5818 , n5762 , n4620 );
not ( n5819 , n5818 );
and ( n5820 , n4617 , n5819 );
not ( n5821 , n4617 );
and ( n5822 , n5821 , n5818 );
nor ( n5823 , n5820 , n5822 );
not ( n5824 , n5823 );
or ( n5825 , n5817 , n5824 );
not ( n5826 , n5803 );
nand ( n5827 , n5806 , n5801 );
and ( n5828 , n5826 , n5827 );
not ( n5829 , n5826 );
not ( n5830 , n5827 );
and ( n5831 , n5829 , n5830 );
nor ( n5832 , n5828 , n5831 );
nand ( n5833 , n455 , n5832 );
nand ( n5834 , n5825 , n5833 );
not ( n5835 , n5834 );
or ( n5836 , n5816 , n5835 );
xor ( n5837 , n3153 , n32135 );
xor ( n34707 , n5837 , n32155 );
and ( n5839 , n32161 , n34707 );
xor ( n5840 , n3153 , n32135 );
xor ( n5841 , n5840 , n32155 );
and ( n5842 , n3242 , n5841 );
and ( n5843 , n32161 , n3242 );
or ( n5844 , n5839 , n5842 , n5843 );
nand ( n5845 , n5844 , n3138 );
not ( n5846 , n5845 );
not ( n5847 , n454 );
not ( n5848 , n5847 );
xor ( n5849 , n34653 , n34657 );
xor ( n5850 , n5849 , n34663 );
buf ( n34720 , n5850 );
not ( n5852 , n34720 );
or ( n5853 , n5848 , n5852 );
nand ( n5854 , n454 , n543 );
nand ( n5855 , n5853 , n5854 );
nor ( n5856 , n5846 , n5855 );
nand ( n5857 , n5836 , n5856 );
not ( n5858 , n5857 );
nor ( n5859 , n5858 , n3248 );
and ( n5860 , n5743 , n5815 , n5859 );
not ( n5861 , n5860 );
not ( n5862 , n3827 );
or ( n5863 , n5861 , n5862 );
not ( n5864 , n4267 );
not ( n5865 , n5555 );
or ( n5866 , n5864 , n5865 );
nand ( n5867 , n5866 , n5742 );
not ( n5868 , n454 );
not ( n5869 , n5834 );
or ( n5870 , n5868 , n5869 );
nand ( n5871 , n5870 , n5856 );
buf ( n5872 , n3246 );
nand ( n5873 , n5871 , n3250 , n5872 );
not ( n5874 , n5845 );
nand ( n5875 , n5834 , n454 );
not ( n5876 , n5875 );
or ( n5877 , n5874 , n5876 );
nand ( n5878 , n5877 , n5855 );
nand ( n5879 , n5873 , n5878 );
nand ( n5880 , n5867 , n5879 , n5815 );
not ( n5881 , n5800 );
not ( n5882 , n5814 );
or ( n5883 , n5881 , n5882 );
nand ( n5884 , n5883 , n34629 );
not ( n5885 , n5884 );
nand ( n5886 , n5867 , n5885 );
buf ( n5887 , n5555 );
and ( n5888 , n5741 , n4267 );
nand ( n5889 , n5887 , n5888 );
nand ( n5890 , n5880 , n5886 , n5889 );
not ( n5891 , n5890 );
nand ( n5892 , n5863 , n5891 );
buf ( n34762 , n2911 );
buf ( n34763 , n31868 );
buf ( n34764 , n525 );
and ( n5896 , n34763 , n34764 );
buf ( n34766 , n34557 );
buf ( n34767 , n549 );
and ( n5899 , n34766 , n34767 );
nor ( n5900 , n5896 , n5899 );
buf ( n34770 , n5900 );
buf ( n34771 , n34770 );
or ( n5903 , n34762 , n34771 );
buf ( n34773 , n2918 );
buf ( n34774 , n31868 );
buf ( n34775 , n524 );
and ( n5907 , n34774 , n34775 );
buf ( n34777 , n524 );
not ( n5909 , n34777 );
buf ( n34779 , n5909 );
buf ( n34780 , n34779 );
buf ( n34781 , n549 );
and ( n5913 , n34780 , n34781 );
nor ( n5914 , n5907 , n5913 );
buf ( n34784 , n5914 );
buf ( n34785 , n34784 );
or ( n34786 , n34773 , n34785 );
nand ( n34787 , n5903 , n34786 );
buf ( n34788 , n34787 );
buf ( n34789 , n459 );
buf ( n34790 , n536 );
buf ( n34791 , n540 );
or ( n34792 , n34790 , n34791 );
buf ( n34793 , n541 );
nand ( n5928 , n34792 , n34793 );
buf ( n34795 , n5928 );
buf ( n34796 , n34795 );
buf ( n34797 , n536 );
buf ( n34798 , n540 );
nand ( n5936 , n34797 , n34798 );
buf ( n34800 , n5936 );
buf ( n34801 , n34800 );
buf ( n34802 , n539 );
and ( n5940 , n34796 , n34801 , n34802 );
buf ( n34804 , n5940 );
buf ( n34805 , n34804 );
and ( n5943 , n34789 , n34805 );
buf ( n34807 , n5943 );
xor ( n5945 , n34788 , n34807 );
buf ( n34809 , n5636 );
buf ( n34810 , n32981 );
buf ( n34811 , n531 );
and ( n5949 , n34810 , n34811 );
buf ( n34813 , n31840 );
buf ( n34814 , n543 );
and ( n5952 , n34813 , n34814 );
nor ( n5953 , n5949 , n5952 );
buf ( n34817 , n5953 );
buf ( n34818 , n34817 );
or ( n5956 , n34809 , n34818 );
buf ( n34820 , n4040 );
buf ( n34821 , n543 );
buf ( n34822 , n31853 );
and ( n5960 , n34821 , n34822 );
not ( n5961 , n34821 );
buf ( n34825 , n530 );
and ( n5963 , n5961 , n34825 );
nor ( n5964 , n5960 , n5963 );
buf ( n34828 , n5964 );
buf ( n34829 , n34828 );
or ( n5967 , n34820 , n34829 );
nand ( n5968 , n5956 , n5967 );
buf ( n34832 , n5968 );
xor ( n5970 , n5945 , n34832 );
xor ( n5971 , n34789 , n34805 );
buf ( n34835 , n5971 );
buf ( n34836 , n34835 );
buf ( n34837 , n551 );
buf ( n34838 , n524 );
and ( n5976 , n34837 , n34838 );
not ( n5977 , n34837 );
buf ( n34841 , n34779 );
and ( n5979 , n5977 , n34841 );
nor ( n5980 , n5976 , n5979 );
buf ( n34844 , n5980 );
buf ( n34845 , n34844 );
not ( n5983 , n34845 );
buf ( n34847 , n5983 );
buf ( n34848 , n34847 );
buf ( n34849 , n2846 );
or ( n5987 , n34848 , n34849 );
or ( n5988 , n523 , n551 );
nand ( n5989 , n523 , n551 );
nand ( n5990 , n5988 , n5989 );
buf ( n34854 , n5990 );
buf ( n34855 , n32352 );
or ( n5993 , n34854 , n34855 );
nand ( n5994 , n5987 , n5993 );
buf ( n34858 , n5994 );
buf ( n34859 , n34858 );
xor ( n5997 , n34836 , n34859 );
buf ( n34861 , n32059 );
buf ( n34862 , n539 );
or ( n6000 , n34861 , n34862 );
not ( n6001 , n539 );
buf ( n34865 , n6001 );
buf ( n34866 , n536 );
or ( n6004 , n34865 , n34866 );
nand ( n6005 , n6000 , n6004 );
buf ( n34869 , n6005 );
buf ( n34870 , n34869 );
not ( n6008 , n34870 );
xor ( n6009 , n540 , n541 );
not ( n6010 , n6009 );
buf ( n34874 , n539 );
buf ( n34875 , n540 );
xor ( n6013 , n34874 , n34875 );
buf ( n34877 , n6013 );
nand ( n6015 , n6010 , n34877 );
not ( n6016 , n6015 );
buf ( n34880 , n6016 );
not ( n6018 , n34880 );
or ( n6019 , n6008 , n6018 );
buf ( n34883 , n6010 );
buf ( n34884 , n6001 );
buf ( n34885 , n535 );
and ( n6023 , n34884 , n34885 );
buf ( n34887 , n32074 );
buf ( n34888 , n539 );
and ( n6026 , n34887 , n34888 );
nor ( n6027 , n6023 , n6026 );
buf ( n34891 , n6027 );
buf ( n34892 , n34891 );
or ( n6030 , n34883 , n34892 );
nand ( n6031 , n6019 , n6030 );
buf ( n34895 , n6031 );
buf ( n34896 , n34895 );
and ( n6034 , n5997 , n34896 );
and ( n6035 , n34836 , n34859 );
or ( n6036 , n6034 , n6035 );
buf ( n34900 , n6036 );
buf ( n34901 , n3020 );
buf ( n34902 , n547 );
buf ( n34903 , n33009 );
and ( n6041 , n34902 , n34903 );
not ( n6042 , n34902 );
buf ( n34906 , n527 );
and ( n6044 , n6042 , n34906 );
nor ( n6045 , n6041 , n6044 );
buf ( n34909 , n6045 );
buf ( n34910 , n34909 );
or ( n6048 , n34901 , n34910 );
buf ( n34912 , n31978 );
buf ( n34913 , n547 );
buf ( n34914 , n526 );
xnor ( n6052 , n34913 , n34914 );
buf ( n34916 , n6052 );
buf ( n34917 , n34916 );
or ( n6055 , n34912 , n34917 );
nand ( n6056 , n6048 , n6055 );
buf ( n34920 , n6056 );
buf ( n34921 , n34920 );
buf ( n34922 , n6015 );
buf ( n34923 , n34891 );
or ( n6061 , n34922 , n34923 );
buf ( n34925 , n6010 );
and ( n6063 , n539 , n32008 );
not ( n6064 , n539 );
and ( n6065 , n6064 , n534 );
nor ( n6066 , n6063 , n6065 );
buf ( n34930 , n6066 );
or ( n6068 , n34925 , n34930 );
nand ( n6069 , n6061 , n6068 );
buf ( n34933 , n6069 );
buf ( n34934 , n34933 );
xor ( n6072 , n34921 , n34934 );
buf ( n34936 , n3069 );
buf ( n34937 , n32053 );
buf ( n34938 , n529 );
and ( n6076 , n34937 , n34938 );
buf ( n34940 , n2969 );
buf ( n34941 , n545 );
and ( n6079 , n34940 , n34941 );
nor ( n6080 , n6076 , n6079 );
buf ( n34944 , n6080 );
buf ( n34945 , n34944 );
or ( n34946 , n34936 , n34945 );
buf ( n34947 , n3087 );
or ( n6088 , n32053 , n528 );
or ( n34949 , n545 , n32183 );
nand ( n6093 , n6088 , n34949 );
not ( n6094 , n6093 );
buf ( n34952 , n6094 );
or ( n6096 , n34947 , n34952 );
nand ( n6097 , n34946 , n6096 );
buf ( n34955 , n6097 );
buf ( n34956 , n34955 );
xor ( n6100 , n6072 , n34956 );
buf ( n34958 , n6100 );
xor ( n6102 , n34900 , n34958 );
xor ( n6103 , n5970 , n6102 );
xor ( n6104 , n34569 , n34589 );
and ( n6105 , n6104 , n34599 );
and ( n6106 , n34569 , n34589 );
or ( n6107 , n6105 , n6106 );
buf ( n34965 , n6107 );
buf ( n34966 , n34965 );
buf ( n34967 , n6009 );
buf ( n34968 , n536 );
and ( n6112 , n34967 , n34968 );
buf ( n34970 , n6112 );
buf ( n34971 , n34970 );
buf ( n34972 , n460 );
xor ( n6116 , n34971 , n34972 );
buf ( n34974 , n34561 );
not ( n6118 , n34974 );
buf ( n34976 , n3199 );
not ( n6120 , n34976 );
or ( n6121 , n6118 , n6120 );
buf ( n34979 , n34844 );
buf ( n34980 , n552 );
nand ( n6124 , n34979 , n34980 );
buf ( n34982 , n6124 );
buf ( n34983 , n34982 );
nand ( n6127 , n6121 , n34983 );
buf ( n34985 , n6127 );
buf ( n34986 , n34985 );
xor ( n6130 , n6116 , n34986 );
buf ( n34988 , n6130 );
buf ( n34989 , n34988 );
xor ( n6133 , n34966 , n34989 );
xor ( n6134 , n5635 , n34527 );
and ( n6135 , n6134 , n34544 );
and ( n6136 , n5635 , n34527 );
or ( n6137 , n6135 , n6136 );
buf ( n34995 , n6137 );
and ( n6139 , n6133 , n34995 );
and ( n6140 , n34966 , n34989 );
or ( n6141 , n6139 , n6140 );
buf ( n34999 , n6141 );
buf ( n35000 , n34999 );
buf ( n35001 , n3020 );
buf ( n35002 , n547 );
buf ( n35003 , n32183 );
and ( n6147 , n35002 , n35003 );
not ( n6148 , n35002 );
buf ( n35006 , n528 );
and ( n6150 , n6148 , n35006 );
nor ( n6151 , n6147 , n6150 );
buf ( n35009 , n6151 );
buf ( n35010 , n35009 );
or ( n6154 , n35001 , n35010 );
buf ( n35012 , n31978 );
buf ( n35013 , n34909 );
or ( n6157 , n35012 , n35013 );
nand ( n6158 , n6154 , n6157 );
buf ( n35016 , n6158 );
buf ( n35017 , n35016 );
buf ( n35018 , n32053 );
buf ( n35019 , n530 );
and ( n6163 , n35018 , n35019 );
buf ( n35021 , n31853 );
buf ( n35022 , n545 );
and ( n35023 , n35021 , n35022 );
nor ( n6167 , n6163 , n35023 );
buf ( n35025 , n6167 );
or ( n6169 , n35025 , n3069 );
or ( n6170 , n34944 , n3087 );
nand ( n6171 , n6169 , n6170 );
buf ( n35029 , n6171 );
xor ( n6173 , n35017 , n35029 );
buf ( n35031 , n526 );
buf ( n35032 , n31868 );
and ( n6176 , n35031 , n35032 );
not ( n6177 , n35031 );
buf ( n35035 , n549 );
and ( n6179 , n6177 , n35035 );
nor ( n6180 , n6176 , n6179 );
buf ( n35038 , n6180 );
buf ( n35039 , n35038 );
not ( n6183 , n35039 );
buf ( n35041 , n6183 );
buf ( n35042 , n35041 );
not ( n6186 , n35042 );
buf ( n35044 , n31897 );
not ( n6188 , n35044 );
or ( n6189 , n6186 , n6188 );
buf ( n35047 , n2918 );
buf ( n35048 , n34770 );
or ( n6192 , n35047 , n35048 );
nand ( n6193 , n6189 , n6192 );
buf ( n35051 , n6193 );
buf ( n35052 , n35051 );
xor ( n6196 , n6173 , n35052 );
buf ( n35054 , n6196 );
buf ( n35055 , n35054 );
xor ( n6199 , n35000 , n35055 );
buf ( n35057 , n4030 );
buf ( n35058 , n32981 );
buf ( n35059 , n532 );
and ( n6203 , n35058 , n35059 );
buf ( n35061 , n31908 );
buf ( n35062 , n543 );
and ( n6206 , n35061 , n35062 );
nor ( n6207 , n6203 , n6206 );
buf ( n35065 , n6207 );
buf ( n35066 , n35065 );
or ( n6210 , n35057 , n35066 );
buf ( n35068 , n32165 );
not ( n6212 , n35068 );
buf ( n35070 , n6212 );
buf ( n35071 , n35070 );
buf ( n35072 , n34817 );
or ( n6216 , n35071 , n35072 );
nand ( n6217 , n6210 , n6216 );
buf ( n35075 , n6217 );
buf ( n35076 , n35075 );
buf ( n35077 , n5582 );
buf ( n35078 , n541 );
buf ( n35079 , n32008 );
and ( n6223 , n35078 , n35079 );
not ( n6224 , n35078 );
buf ( n35082 , n534 );
and ( n6226 , n6224 , n35082 );
nor ( n6227 , n6223 , n6226 );
buf ( n35085 , n6227 );
buf ( n35086 , n35085 );
or ( n6230 , n35077 , n35086 );
buf ( n35088 , n33118 );
buf ( n35089 , n541 );
buf ( n35090 , n31874 );
and ( n6234 , n35089 , n35090 );
not ( n6235 , n35089 );
buf ( n35093 , n533 );
and ( n6237 , n6235 , n35093 );
nor ( n6238 , n6234 , n6237 );
buf ( n35096 , n6238 );
buf ( n35097 , n35096 );
or ( n6241 , n35088 , n35097 );
nand ( n6242 , n6230 , n6241 );
buf ( n35100 , n6242 );
buf ( n35101 , n35100 );
xor ( n35102 , n35076 , n35101 );
buf ( n35103 , n2911 );
buf ( n35104 , n34540 );
or ( n35105 , n35103 , n35104 );
buf ( n35106 , n2918 );
buf ( n35107 , n35038 );
or ( n6257 , n35106 , n35107 );
nand ( n6258 , n35105 , n6257 );
buf ( n35110 , n6258 );
buf ( n35111 , n5582 );
buf ( n35112 , n34483 );
or ( n6262 , n35111 , n35112 );
buf ( n35114 , n33118 );
buf ( n35115 , n35085 );
or ( n6265 , n35114 , n35115 );
nand ( n6266 , n6262 , n6265 );
buf ( n35118 , n6266 );
xor ( n6268 , n35110 , n35118 );
buf ( n35120 , n4030 );
buf ( n35121 , n34523 );
or ( n6271 , n35120 , n35121 );
buf ( n35123 , n4040 );
buf ( n35124 , n35065 );
or ( n6274 , n35123 , n35124 );
nand ( n6275 , n6271 , n6274 );
buf ( n35127 , n6275 );
and ( n6277 , n6268 , n35127 );
and ( n6278 , n35110 , n35118 );
or ( n6279 , n6277 , n6278 );
buf ( n35131 , n6279 );
xor ( n6281 , n35102 , n35131 );
buf ( n35133 , n6281 );
buf ( n35134 , n35133 );
and ( n6284 , n6199 , n35134 );
and ( n6285 , n35000 , n35055 );
or ( n6286 , n6284 , n6285 );
buf ( n35138 , n6286 );
xor ( n6288 , n6103 , n35138 );
buf ( n6289 , n31988 );
or ( n6290 , n35009 , n6289 );
not ( n6291 , n32002 );
nand ( n6292 , n6291 , n5721 );
nand ( n6293 , n6290 , n6292 );
not ( n6294 , n6293 );
and ( n6295 , n34570 , n34586 );
buf ( n35147 , n6295 );
not ( n6297 , n35147 );
nand ( n6298 , n6294 , n6297 );
not ( n6299 , n6298 );
not ( n6300 , n3063 );
not ( n6301 , n35025 );
not ( n6302 , n6301 );
or ( n6303 , n6300 , n6302 );
not ( n6304 , n34508 );
not ( n6305 , n3069 );
nand ( n6306 , n6304 , n6305 );
nand ( n6307 , n6303 , n6306 );
not ( n6308 , n6307 );
or ( n6309 , n6299 , n6308 );
nand ( n6310 , n35147 , n6293 );
nand ( n6311 , n6309 , n6310 );
buf ( n35163 , n6311 );
xor ( n6313 , n34971 , n34972 );
and ( n6314 , n6313 , n34986 );
and ( n6315 , n34971 , n34972 );
or ( n6316 , n6314 , n6315 );
buf ( n35168 , n6316 );
buf ( n35169 , n35168 );
xor ( n6319 , n35163 , n35169 );
xor ( n6320 , n34836 , n34859 );
xor ( n6321 , n6320 , n34896 );
buf ( n35173 , n6321 );
buf ( n35174 , n35173 );
and ( n6324 , n6319 , n35174 );
and ( n35176 , n35163 , n35169 );
or ( n6326 , n6324 , n35176 );
buf ( n35178 , n6326 );
buf ( n35179 , n35178 );
xor ( n6329 , n35076 , n35101 );
and ( n6330 , n6329 , n35131 );
and ( n6331 , n35076 , n35101 );
or ( n6332 , n6330 , n6331 );
buf ( n35184 , n6332 );
buf ( n35185 , n35184 );
xor ( n6335 , n35179 , n35185 );
xor ( n6336 , n539 , n538 );
not ( n6337 , n6336 );
buf ( n35189 , n6337 );
buf ( n35190 , n32059 );
nor ( n6340 , n35189 , n35190 );
buf ( n35192 , n6340 );
xor ( n6342 , n35192 , n458 );
buf ( n35194 , n552 );
not ( n6344 , n35194 );
buf ( n35196 , n551 );
buf ( n35197 , n522 );
not ( n6347 , n35197 );
buf ( n35199 , n6347 );
buf ( n35200 , n35199 );
and ( n6350 , n35196 , n35200 );
not ( n6351 , n35196 );
buf ( n35203 , n522 );
and ( n6353 , n6351 , n35203 );
nor ( n6354 , n6350 , n6353 );
buf ( n35206 , n6354 );
buf ( n35207 , n35206 );
not ( n6357 , n35207 );
buf ( n35209 , n6357 );
buf ( n35210 , n35209 );
not ( n6360 , n35210 );
or ( n6361 , n6344 , n6360 );
buf ( n35213 , n2962 );
buf ( n35214 , n5990 );
or ( n6364 , n35213 , n35214 );
nand ( n6365 , n6361 , n6364 );
buf ( n35217 , n6365 );
xor ( n6367 , n6342 , n35217 );
buf ( n35219 , n5582 );
buf ( n35220 , n35096 );
or ( n6370 , n35219 , n35220 );
buf ( n35222 , n33118 );
buf ( n35223 , n541 );
buf ( n35224 , n31908 );
and ( n6374 , n35223 , n35224 );
not ( n6375 , n35223 );
buf ( n35227 , n532 );
and ( n6377 , n6375 , n35227 );
nor ( n6378 , n6374 , n6377 );
buf ( n35230 , n6378 );
buf ( n35231 , n35230 );
or ( n6381 , n35222 , n35231 );
nand ( n6382 , n6370 , n6381 );
buf ( n35234 , n6382 );
xor ( n6384 , n35017 , n35029 );
and ( n6385 , n6384 , n35052 );
and ( n6386 , n35017 , n35029 );
or ( n6387 , n6385 , n6386 );
buf ( n35239 , n6387 );
xor ( n6389 , n35234 , n35239 );
xor ( n6390 , n6367 , n6389 );
buf ( n35242 , n6390 );
xor ( n35243 , n6335 , n35242 );
buf ( n35244 , n35243 );
and ( n6394 , n6288 , n35244 );
and ( n6395 , n6103 , n35138 );
or ( n35247 , n6394 , n6395 );
nand ( n6400 , n35247 , n3138 );
not ( n35249 , n6400 );
not ( n6402 , n5847 );
xor ( n6403 , n35179 , n35185 );
and ( n35252 , n6403 , n35242 );
and ( n6408 , n35179 , n35185 );
or ( n6409 , n35252 , n6408 );
buf ( n35255 , n6409 );
buf ( n35256 , n35255 );
buf ( n35257 , n5636 );
buf ( n35258 , n34828 );
or ( n6414 , n35257 , n35258 );
buf ( n35260 , n4040 );
buf ( n35261 , n543 );
buf ( n35262 , n2969 );
and ( n6418 , n35261 , n35262 );
not ( n6419 , n35261 );
buf ( n35265 , n529 );
and ( n6421 , n6419 , n35265 );
nor ( n6422 , n6418 , n6421 );
buf ( n35268 , n6422 );
buf ( n35269 , n35268 );
or ( n6425 , n35260 , n35269 );
nand ( n6426 , n6414 , n6425 );
buf ( n35272 , n6426 );
buf ( n35273 , n35272 );
buf ( n35274 , n5582 );
buf ( n35275 , n35230 );
or ( n6431 , n35274 , n35275 );
buf ( n35277 , n33118 );
buf ( n35278 , n541 );
not ( n6434 , n35278 );
buf ( n35280 , n531 );
nor ( n6436 , n6434 , n35280 );
buf ( n35282 , n6436 );
buf ( n35283 , n35282 );
buf ( n35284 , n531 );
not ( n6440 , n35284 );
buf ( n35286 , n541 );
nor ( n6442 , n6440 , n35286 );
buf ( n35288 , n6442 );
buf ( n35289 , n35288 );
nor ( n6445 , n35283 , n35289 );
buf ( n35291 , n6445 );
buf ( n35292 , n35291 );
or ( n6448 , n35277 , n35292 );
nand ( n6449 , n6431 , n6448 );
buf ( n35295 , n6449 );
buf ( n35296 , n35295 );
xor ( n6452 , n35273 , n35296 );
buf ( n35298 , n3045 );
buf ( n35299 , n34784 );
or ( n6455 , n35298 , n35299 );
buf ( n35301 , n2918 );
buf ( n35302 , n31868 );
buf ( n35303 , n523 );
and ( n6459 , n35302 , n35303 );
buf ( n35305 , n523 );
not ( n6461 , n35305 );
buf ( n35307 , n6461 );
buf ( n35308 , n35307 );
buf ( n35309 , n549 );
and ( n6465 , n35308 , n35309 );
nor ( n6466 , n6459 , n6465 );
buf ( n35312 , n6466 );
buf ( n35313 , n35312 );
or ( n6469 , n35301 , n35313 );
nand ( n6470 , n6455 , n6469 );
buf ( n35316 , n6470 );
buf ( n35317 , n35316 );
xor ( n6473 , n6452 , n35317 );
buf ( n35319 , n6473 );
buf ( n35320 , n35319 );
buf ( n35321 , n536 );
buf ( n35322 , n538 );
or ( n6478 , n35321 , n35322 );
buf ( n35324 , n539 );
nand ( n6480 , n6478 , n35324 );
buf ( n35326 , n6480 );
buf ( n35327 , n35326 );
buf ( n35328 , n536 );
buf ( n35329 , n538 );
nand ( n6485 , n35328 , n35329 );
buf ( n35331 , n6485 );
buf ( n35332 , n35331 );
buf ( n35333 , n537 );
and ( n6489 , n35327 , n35332 , n35333 );
buf ( n35335 , n6489 );
xor ( n6491 , n457 , n35335 );
buf ( n35337 , n2846 );
buf ( n35338 , n35206 );
or ( n6494 , n35337 , n35338 );
buf ( n35340 , n551 );
buf ( n35341 , n521 );
not ( n6497 , n35341 );
buf ( n35343 , n6497 );
buf ( n35344 , n35343 );
and ( n6500 , n35340 , n35344 );
not ( n6501 , n35340 );
buf ( n35347 , n521 );
and ( n6503 , n6501 , n35347 );
nor ( n6504 , n6500 , n6503 );
buf ( n35350 , n6504 );
buf ( n35351 , n35350 );
buf ( n35352 , n32352 );
or ( n6508 , n35351 , n35352 );
nand ( n6509 , n6494 , n6508 );
buf ( n35355 , n6509 );
and ( n6511 , n6491 , n35355 );
not ( n6512 , n6491 );
not ( n6513 , n35355 );
and ( n6514 , n6512 , n6513 );
nor ( n6515 , n6511 , n6514 );
or ( n6516 , n6094 , n3069 );
and ( n6517 , n33009 , n545 );
and ( n6518 , n32053 , n527 );
nor ( n6519 , n6517 , n6518 );
or ( n6520 , n6519 , n3064 );
nand ( n6521 , n6516 , n6520 );
xor ( n6522 , n6515 , n6521 );
buf ( n35368 , n6522 );
xor ( n6524 , n35320 , n35368 );
not ( n6525 , n6066 );
not ( n6526 , n6525 );
not ( n6527 , n6016 );
or ( n6528 , n6526 , n6527 );
buf ( n35374 , n6001 );
buf ( n35375 , n533 );
and ( n6531 , n35374 , n35375 );
buf ( n35377 , n31874 );
buf ( n35378 , n539 );
and ( n6534 , n35377 , n35378 );
nor ( n6535 , n6531 , n6534 );
buf ( n35381 , n6535 );
or ( n6537 , n6010 , n35381 );
nand ( n35383 , n6528 , n6537 );
buf ( n35384 , n35383 );
not ( n6540 , n535 );
not ( n6541 , n537 );
not ( n35387 , n6541 );
or ( n6546 , n6540 , n35387 );
nand ( n35389 , n537 , n32074 );
nand ( n6548 , n6546 , n35389 );
not ( n6549 , n6548 );
not ( n35392 , n6336 );
or ( n6554 , n6549 , n35392 );
buf ( n35394 , n538 );
buf ( n35395 , n537 );
xor ( n6557 , n35394 , n35395 );
buf ( n35397 , n6557 );
nand ( n6559 , n35397 , n6337 );
buf ( n35399 , n6541 );
buf ( n35400 , n536 );
and ( n6562 , n35399 , n35400 );
buf ( n35402 , n32059 );
buf ( n35403 , n537 );
and ( n6565 , n35402 , n35403 );
nor ( n6566 , n6562 , n6565 );
buf ( n35406 , n6566 );
or ( n6568 , n6559 , n35406 );
nand ( n6569 , n6554 , n6568 );
buf ( n35409 , n6569 );
xor ( n6571 , n35384 , n35409 );
buf ( n35411 , n3020 );
buf ( n35412 , n34916 );
or ( n6574 , n35411 , n35412 );
buf ( n35414 , n31978 );
buf ( n35415 , n547 );
buf ( n35416 , n34557 );
and ( n6578 , n35415 , n35416 );
not ( n6579 , n35415 );
buf ( n35419 , n525 );
and ( n6581 , n6579 , n35419 );
nor ( n6582 , n6578 , n6581 );
buf ( n35422 , n6582 );
buf ( n35423 , n35422 );
or ( n6585 , n35414 , n35423 );
nand ( n6586 , n6574 , n6585 );
buf ( n35426 , n6586 );
buf ( n35427 , n35426 );
xor ( n6589 , n6571 , n35427 );
buf ( n35429 , n6589 );
buf ( n35430 , n35429 );
xor ( n6592 , n6524 , n35430 );
buf ( n35432 , n6592 );
buf ( n35433 , n35432 );
xor ( n6595 , n35256 , n35433 );
xor ( n6596 , n34788 , n34807 );
and ( n6597 , n6596 , n34832 );
and ( n6598 , n34788 , n34807 );
or ( n6599 , n6597 , n6598 );
xor ( n6600 , n35192 , n458 );
and ( n6601 , n6600 , n35217 );
and ( n6602 , n35192 , n458 );
or ( n6603 , n6601 , n6602 );
xor ( n6604 , n6599 , n6603 );
xor ( n6605 , n34921 , n34934 );
and ( n6606 , n6605 , n34956 );
and ( n6607 , n34921 , n34934 );
or ( n6608 , n6606 , n6607 );
buf ( n35448 , n6608 );
xor ( n6610 , n6604 , n35448 );
xor ( n6611 , n35192 , n458 );
xor ( n6612 , n6611 , n35217 );
and ( n6613 , n35234 , n6612 );
xor ( n6614 , n35192 , n458 );
xor ( n6615 , n6614 , n35217 );
and ( n6616 , n35239 , n6615 );
and ( n6617 , n35234 , n35239 );
or ( n6618 , n6613 , n6616 , n6617 );
xor ( n6619 , n34788 , n34807 );
xor ( n6620 , n6619 , n34832 );
and ( n6621 , n34900 , n6620 );
xor ( n35461 , n34788 , n34807 );
xor ( n6623 , n35461 , n34832 );
and ( n6624 , n34958 , n6623 );
and ( n6625 , n34900 , n34958 );
or ( n6626 , n6621 , n6624 , n6625 );
xor ( n6627 , n6618 , n6626 );
xor ( n6628 , n6610 , n6627 );
buf ( n35468 , n6628 );
xor ( n6630 , n6595 , n35468 );
buf ( n35470 , n6630 );
not ( n6632 , n35470 );
or ( n6633 , n6402 , n6632 );
nand ( n6634 , n454 , n537 );
nand ( n6635 , n6633 , n6634 );
nor ( n6636 , n35249 , n6635 );
not ( n6637 , n6636 );
buf ( n35477 , n520 );
buf ( n35478 , n489 );
and ( n6640 , n35477 , n35478 );
buf ( n35480 , n6640 );
buf ( n35481 , n35480 );
not ( n6643 , n503 );
not ( n6644 , n505 );
nor ( n6645 , n6644 , n504 );
nor ( n6646 , n6643 , n6645 );
buf ( n35486 , n6646 );
xor ( n6648 , n35481 , n35486 );
and ( n6649 , n501 , n507 );
not ( n6650 , n501 );
and ( n6651 , n6650 , n33214 );
nor ( n6652 , n6649 , n6651 );
not ( n6653 , n6652 );
not ( n6654 , n33569 );
or ( n6655 , n6653 , n6654 );
xor ( n6656 , n501 , n506 );
buf ( n35496 , n6656 );
buf ( n35497 , n1907 );
nand ( n6659 , n35496 , n35497 );
buf ( n35499 , n6659 );
nand ( n6661 , n6655 , n35499 );
buf ( n35501 , n6661 );
xor ( n6663 , n6648 , n35501 );
buf ( n35503 , n6663 );
buf ( n35504 , n35503 );
not ( n6666 , n497 );
not ( n6667 , n31205 );
or ( n6668 , n6666 , n6667 );
nand ( n6669 , n6668 , n2211 );
not ( n6670 , n6669 );
buf ( n35510 , n511 );
buf ( n35511 , n497 );
xor ( n6673 , n35510 , n35511 );
buf ( n35513 , n6673 );
not ( n6675 , n35513 );
or ( n6676 , n6670 , n6675 );
and ( n6677 , n510 , n497 );
not ( n6678 , n510 );
and ( n6679 , n6678 , n699 );
nor ( n6680 , n6677 , n6679 );
nand ( n6681 , n6680 , n2081 );
nand ( n35521 , n6676 , n6681 );
buf ( n35522 , n35521 );
not ( n6684 , n35522 );
buf ( n35524 , n6684 );
not ( n35525 , n35524 );
not ( n6690 , n489 );
not ( n35527 , n1944 );
or ( n6692 , n6690 , n35527 );
not ( n6693 , n489 );
nand ( n35530 , n6693 , n519 );
nand ( n6698 , n6692 , n35530 );
not ( n6699 , n6698 );
nor ( n6700 , n489 , n490 );
not ( n6701 , n6700 );
nand ( n6702 , n489 , n490 );
nand ( n6703 , n6701 , n6702 );
nor ( n6704 , n6703 , n4626 );
not ( n6705 , n6704 );
or ( n6706 , n6699 , n6705 );
buf ( n35540 , n4626 );
xor ( n6708 , n489 , n518 );
buf ( n35542 , n6708 );
nand ( n6710 , n35540 , n35542 );
buf ( n35544 , n6710 );
nand ( n6712 , n6706 , n35544 );
buf ( n35546 , n6712 );
not ( n6714 , n35546 );
buf ( n35548 , n6714 );
not ( n6716 , n35548 );
or ( n6717 , n35525 , n6716 );
nand ( n6718 , n35521 , n6712 );
nand ( n6719 , n6717 , n6718 );
buf ( n35553 , n513 );
buf ( n35554 , n495 );
xor ( n6722 , n35553 , n35554 );
buf ( n35556 , n6722 );
buf ( n35557 , n35556 );
not ( n6725 , n35557 );
nand ( n6726 , n699 , n496 );
buf ( n35560 , n6726 );
not ( n6728 , n496 );
nand ( n6729 , n6728 , n497 );
buf ( n35563 , n6729 );
nand ( n6731 , n2403 , n2400 );
buf ( n35565 , n6731 );
and ( n6733 , n35560 , n35563 , n35565 );
buf ( n35567 , n6733 );
buf ( n35568 , n35567 );
not ( n6736 , n35568 );
or ( n6737 , n6725 , n6736 );
buf ( n35571 , n496 );
buf ( n35572 , n497 );
xor ( n6740 , n35571 , n35572 );
buf ( n35574 , n6740 );
buf ( n35575 , n35574 );
buf ( n35576 , n512 );
buf ( n35577 , n495 );
xor ( n6745 , n35576 , n35577 );
buf ( n35579 , n6745 );
buf ( n35580 , n35579 );
nand ( n6748 , n35575 , n35580 );
buf ( n35582 , n6748 );
buf ( n35583 , n35582 );
nand ( n6751 , n6737 , n35583 );
buf ( n35585 , n6751 );
buf ( n6753 , n35585 );
not ( n6754 , n6753 );
and ( n6755 , n6719 , n6754 );
not ( n6756 , n6719 );
and ( n6757 , n6756 , n6753 );
nor ( n6758 , n6755 , n6757 );
buf ( n35592 , n6758 );
xor ( n6760 , n35504 , n35592 );
xor ( n6761 , n493 , n515 );
not ( n6762 , n6761 );
and ( n35596 , n494 , n493 );
not ( n6764 , n494 );
not ( n6765 , n493 );
and ( n6766 , n6764 , n6765 );
nor ( n6767 , n35596 , n6766 );
not ( n6768 , n6767 );
nor ( n6769 , n6768 , n2590 );
not ( n6770 , n6769 );
or ( n6771 , n6762 , n6770 );
xor ( n6772 , n493 , n514 );
nand ( n6773 , n6772 , n2591 );
nand ( n6774 , n6771 , n6773 );
xor ( n6775 , n491 , n517 );
buf ( n35609 , n6775 );
not ( n6777 , n35609 );
not ( n6778 , n4510 );
nor ( n6779 , n6778 , n4286 );
buf ( n35613 , n6779 );
not ( n6781 , n35613 );
or ( n6782 , n6777 , n6781 );
buf ( n35616 , n4286 );
xor ( n6784 , n491 , n516 );
buf ( n35618 , n6784 );
nand ( n6786 , n35616 , n35618 );
buf ( n35620 , n6786 );
buf ( n35621 , n35620 );
nand ( n6789 , n6782 , n35621 );
buf ( n35623 , n6789 );
xor ( n6791 , n6774 , n35623 );
xor ( n6792 , n499 , n509 );
buf ( n35626 , n6792 );
not ( n6794 , n35626 );
buf ( n35628 , n1999 );
not ( n6796 , n35628 );
or ( n6797 , n6794 , n6796 );
buf ( n35631 , n30884 );
xor ( n6799 , n499 , n508 );
buf ( n35633 , n6799 );
nand ( n6801 , n35631 , n35633 );
buf ( n35635 , n6801 );
buf ( n35636 , n35635 );
nand ( n6804 , n6797 , n35636 );
buf ( n35638 , n6804 );
xor ( n6806 , n6791 , n35638 );
buf ( n35640 , n6806 );
xor ( n6808 , n6760 , n35640 );
buf ( n35642 , n6808 );
buf ( n35643 , n35642 );
xor ( n6811 , n33621 , n33631 );
and ( n6812 , n6811 , n33634 );
and ( n6813 , n33621 , n33631 );
or ( n6814 , n6812 , n6813 );
buf ( n35648 , n6814 );
buf ( n35649 , n35648 );
buf ( n35650 , n33625 );
not ( n6818 , n35650 );
buf ( n35652 , n4512 );
not ( n35653 , n35652 );
or ( n6821 , n6818 , n35653 );
buf ( n35655 , n4519 );
buf ( n35656 , n6775 );
nand ( n6827 , n35655 , n35656 );
buf ( n35658 , n6827 );
buf ( n35659 , n35658 );
nand ( n6830 , n6821 , n35659 );
buf ( n35661 , n6830 );
buf ( n35662 , n35661 );
not ( n6836 , n1881 );
not ( n6837 , n33552 );
or ( n6838 , n6836 , n6837 );
xor ( n6839 , n503 , n505 );
buf ( n35667 , n6839 );
buf ( n35668 , n504 );
nand ( n6842 , n35667 , n35668 );
buf ( n35670 , n6842 );
nand ( n6844 , n6838 , n35670 );
not ( n6845 , n6844 );
buf ( n35673 , n520 );
buf ( n35674 , n490 );
or ( n6848 , n35673 , n35674 );
buf ( n35676 , n491 );
nand ( n6850 , n6848 , n35676 );
buf ( n35678 , n6850 );
buf ( n35679 , n35678 );
buf ( n35680 , n520 );
buf ( n35681 , n490 );
nand ( n6855 , n35680 , n35681 );
buf ( n35683 , n6855 );
buf ( n35684 , n35683 );
buf ( n35685 , n489 );
and ( n6859 , n35679 , n35684 , n35685 );
buf ( n35687 , n6859 );
not ( n6861 , n35687 );
not ( n6862 , n6861 );
or ( n6863 , n6845 , n6862 );
or ( n6864 , n6861 , n6844 );
nand ( n6865 , n6863 , n6864 );
buf ( n35693 , n6865 );
xor ( n6867 , n35662 , n35693 );
xor ( n6868 , n33547 , n4641 );
and ( n6869 , n6868 , n33580 );
and ( n6870 , n33547 , n4641 );
or ( n6871 , n6869 , n6870 );
buf ( n35699 , n6871 );
xor ( n6873 , n6867 , n35699 );
buf ( n35701 , n6873 );
buf ( n35702 , n35701 );
xor ( n6876 , n35649 , n35702 );
xor ( n6877 , n33582 , n33597 );
and ( n6878 , n6877 , n33604 );
and ( n6879 , n33582 , n33597 );
or ( n6880 , n6878 , n6879 );
buf ( n35708 , n6880 );
buf ( n35709 , n35708 );
and ( n6883 , n6876 , n35709 );
and ( n6884 , n35649 , n35702 );
or ( n6885 , n6883 , n6884 );
buf ( n35713 , n6885 );
buf ( n35714 , n35713 );
xor ( n6888 , n35643 , n35714 );
xor ( n6889 , n35662 , n35693 );
and ( n6890 , n6889 , n35699 );
and ( n6891 , n35662 , n35693 );
or ( n6892 , n6890 , n6891 );
buf ( n35720 , n6892 );
buf ( n35721 , n35720 );
and ( n6895 , n6844 , n35687 );
buf ( n35723 , n6895 );
not ( n6897 , n4657 );
not ( n6898 , n33569 );
or ( n6899 , n6897 , n6898 );
nand ( n6900 , n6652 , n1907 );
nand ( n6901 , n6899 , n6900 );
buf ( n35729 , n6901 );
not ( n6903 , n35729 );
xor ( n6904 , n489 , n520 );
not ( n6905 , n6904 );
not ( n6906 , n6704 );
or ( n6907 , n6905 , n6906 );
nand ( n6908 , n4626 , n6698 );
nand ( n6909 , n6907 , n6908 );
buf ( n35737 , n6909 );
not ( n6911 , n35737 );
or ( n6912 , n6903 , n6911 );
buf ( n35740 , n6909 );
buf ( n35741 , n6901 );
or ( n6915 , n35740 , n35741 );
not ( n6916 , n33647 );
not ( n6917 , n2213 );
or ( n6918 , n6916 , n6917 );
buf ( n35746 , n2081 );
buf ( n35747 , n35513 );
nand ( n6921 , n35746 , n35747 );
buf ( n35749 , n6921 );
nand ( n6923 , n6918 , n35749 );
buf ( n35751 , n6923 );
nand ( n6925 , n6915 , n35751 );
buf ( n35753 , n6925 );
buf ( n35754 , n35753 );
nand ( n6928 , n6912 , n35754 );
buf ( n35756 , n6928 );
buf ( n35757 , n35756 );
xor ( n6931 , n35723 , n35757 );
xor ( n6932 , n499 , n500 );
not ( n6933 , n6932 );
not ( n6934 , n4752 );
nor ( n6935 , n6934 , n1865 );
not ( n6936 , n6935 );
or ( n6937 , n6933 , n6936 );
nand ( n6938 , n6792 , n1865 );
nand ( n6939 , n6937 , n6938 );
buf ( n35767 , n6939 );
not ( n6941 , n4703 );
not ( n6942 , n6769 );
or ( n6943 , n6941 , n6942 );
nand ( n6944 , n2591 , n6761 );
nand ( n6945 , n6943 , n6944 );
buf ( n35773 , n6945 );
xor ( n35774 , n35767 , n35773 );
not ( n6948 , n31271 );
not ( n6949 , n35556 );
or ( n35777 , n6948 , n6949 );
not ( n6954 , n4759 );
nand ( n35779 , n6954 , n6731 , n2409 );
nand ( n6956 , n35777 , n35779 );
buf ( n35781 , n6956 );
and ( n35782 , n35774 , n35781 );
and ( n6962 , n35767 , n35773 );
or ( n6963 , n35782 , n6962 );
buf ( n35785 , n6963 );
buf ( n35786 , n35785 );
xor ( n6966 , n6931 , n35786 );
buf ( n35788 , n6966 );
buf ( n35789 , n35788 );
xor ( n6969 , n35721 , n35789 );
xor ( n6970 , n35767 , n35773 );
xor ( n6971 , n6970 , n35781 );
buf ( n35793 , n6971 );
xor ( n6973 , n6901 , n6909 );
and ( n6974 , n6973 , n6923 );
not ( n6975 , n6973 );
buf ( n35797 , n6923 );
not ( n6977 , n35797 );
buf ( n35799 , n6977 );
and ( n6979 , n6975 , n35799 );
nor ( n6980 , n6974 , n6979 );
xor ( n6981 , n35793 , n6980 );
xor ( n6982 , n33654 , n33668 );
and ( n6983 , n6982 , n33678 );
and ( n6984 , n33654 , n33668 );
or ( n6985 , n6983 , n6984 );
buf ( n35807 , n6985 );
and ( n6987 , n6981 , n35807 );
and ( n6988 , n35793 , n6980 );
or ( n6989 , n6987 , n6988 );
buf ( n35811 , n6989 );
xor ( n6991 , n6969 , n35811 );
buf ( n35813 , n6991 );
buf ( n35814 , n35813 );
and ( n6994 , n6888 , n35814 );
and ( n6995 , n35643 , n35714 );
or ( n6996 , n6994 , n6995 );
buf ( n35818 , n6996 );
buf ( n35819 , n519 );
buf ( n35820 , n489 );
and ( n7000 , n35819 , n35820 );
buf ( n35822 , n7000 );
buf ( n35823 , n35822 );
buf ( n35824 , n32922 );
xor ( n7004 , n35823 , n35824 );
not ( n7005 , n6704 );
not ( n7006 , n6708 );
or ( n7007 , n7005 , n7006 );
xnor ( n7008 , n490 , n491 );
buf ( n35830 , n7008 );
not ( n7010 , n35830 );
buf ( n35832 , n7010 );
buf ( n35833 , n35832 );
buf ( n35834 , n517 );
buf ( n35835 , n489 );
xor ( n7015 , n35834 , n35835 );
buf ( n35837 , n7015 );
buf ( n35838 , n35837 );
nand ( n7018 , n35833 , n35838 );
buf ( n35840 , n7018 );
nand ( n7020 , n7007 , n35840 );
buf ( n35842 , n7020 );
xor ( n7022 , n7004 , n35842 );
buf ( n35844 , n7022 );
buf ( n35845 , n35844 );
buf ( n35846 , n505 );
buf ( n35847 , n501 );
xor ( n7027 , n35846 , n35847 );
buf ( n35849 , n7027 );
not ( n7029 , n35849 );
not ( n7030 , n1915 );
or ( n7031 , n7029 , n7030 );
nand ( n7032 , n33569 , n6656 );
nand ( n7033 , n7031 , n7032 );
buf ( n35855 , n7033 );
buf ( n35856 , n35579 );
not ( n7036 , n35856 );
buf ( n35858 , n35567 );
not ( n7038 , n35858 );
or ( n7039 , n7036 , n7038 );
buf ( n35861 , n35574 );
and ( n7041 , n511 , n495 );
not ( n7042 , n511 );
and ( n7043 , n7042 , n758 );
nor ( n7044 , n7041 , n7043 );
buf ( n35866 , n7044 );
nand ( n7046 , n35861 , n35866 );
buf ( n35868 , n7046 );
buf ( n35869 , n35868 );
nand ( n7049 , n7039 , n35869 );
buf ( n35871 , n7049 );
buf ( n35872 , n35871 );
xor ( n7052 , n35855 , n35872 );
buf ( n35874 , n6799 );
not ( n7054 , n35874 );
buf ( n35876 , n2001 );
not ( n7056 , n35876 );
or ( n7057 , n7054 , n7056 );
buf ( n35879 , n31011 );
buf ( n35880 , n507 );
buf ( n35881 , n499 );
xor ( n7061 , n35880 , n35881 );
buf ( n35883 , n7061 );
buf ( n35884 , n35883 );
nand ( n35885 , n35879 , n35884 );
buf ( n35886 , n35885 );
buf ( n35887 , n35886 );
nand ( n35888 , n7057 , n35887 );
buf ( n35889 , n35888 );
buf ( n35890 , n35889 );
xor ( n7073 , n7052 , n35890 );
buf ( n35892 , n7073 );
buf ( n35893 , n35892 );
xor ( n7079 , n35845 , n35893 );
xor ( n7080 , n35723 , n35757 );
and ( n7081 , n7080 , n35786 );
and ( n7082 , n35723 , n35757 );
or ( n7083 , n7081 , n7082 );
buf ( n35899 , n7083 );
buf ( n35900 , n35899 );
xor ( n7086 , n7079 , n35900 );
buf ( n35902 , n7086 );
buf ( n35903 , n35902 );
xor ( n7089 , n35721 , n35789 );
and ( n7090 , n7089 , n35811 );
and ( n7091 , n35721 , n35789 );
or ( n7092 , n7090 , n7091 );
buf ( n35908 , n7092 );
buf ( n35909 , n35908 );
xor ( n7095 , n35903 , n35909 );
not ( n7096 , n2081 );
buf ( n35912 , n509 );
buf ( n35913 , n497 );
xor ( n7099 , n35912 , n35913 );
buf ( n35915 , n7099 );
not ( n7101 , n35915 );
or ( n7102 , n7096 , n7101 );
nand ( n7103 , n6680 , n6669 );
nand ( n7104 , n7102 , n7103 );
not ( n7105 , n7104 );
buf ( n35921 , n6784 );
not ( n7107 , n35921 );
buf ( n35923 , n33438 );
not ( n7109 , n35923 );
or ( n7110 , n7107 , n7109 );
buf ( n35926 , n4519 );
buf ( n35927 , n515 );
buf ( n35928 , n491 );
xor ( n7114 , n35927 , n35928 );
buf ( n35930 , n7114 );
buf ( n35931 , n35930 );
nand ( n7117 , n35926 , n35931 );
buf ( n35933 , n7117 );
buf ( n35934 , n35933 );
nand ( n7120 , n7110 , n35934 );
buf ( n35936 , n7120 );
xor ( n7122 , n7105 , n35936 );
buf ( n35938 , n6772 );
not ( n7124 , n35938 );
buf ( n35940 , n2668 );
not ( n7126 , n35940 );
or ( n7127 , n7124 , n7126 );
buf ( n35943 , n2591 );
buf ( n35944 , n513 );
buf ( n35945 , n493 );
xor ( n7131 , n35944 , n35945 );
buf ( n35947 , n7131 );
buf ( n35948 , n35947 );
nand ( n7134 , n35943 , n35948 );
buf ( n35950 , n7134 );
buf ( n35951 , n35950 );
nand ( n7137 , n7127 , n35951 );
buf ( n35953 , n7137 );
xor ( n7139 , n7122 , n35953 );
buf ( n35955 , n7139 );
xor ( n7141 , n35481 , n35486 );
and ( n7142 , n7141 , n35501 );
and ( n7143 , n35481 , n35486 );
or ( n7144 , n7142 , n7143 );
buf ( n35960 , n7144 );
buf ( n35961 , n35960 );
not ( n7147 , n6712 );
not ( n7148 , n35585 );
or ( n7149 , n7147 , n7148 );
buf ( n35965 , n35585 );
buf ( n35966 , n6712 );
nor ( n7152 , n35965 , n35966 );
buf ( n35968 , n7152 );
or ( n7154 , n35968 , n35524 );
nand ( n7155 , n7149 , n7154 );
buf ( n35971 , n7155 );
xor ( n7157 , n35961 , n35971 );
buf ( n35973 , n35623 );
buf ( n35974 , n6774 );
or ( n7160 , n35973 , n35974 );
buf ( n35976 , n35638 );
nand ( n7162 , n7160 , n35976 );
buf ( n35978 , n7162 );
buf ( n35979 , n35978 );
buf ( n35980 , n35623 );
buf ( n35981 , n6774 );
nand ( n7167 , n35980 , n35981 );
buf ( n35983 , n7167 );
buf ( n35984 , n35983 );
nand ( n35985 , n35979 , n35984 );
buf ( n35986 , n35985 );
buf ( n35987 , n35986 );
xor ( n7173 , n7157 , n35987 );
buf ( n35989 , n7173 );
buf ( n35990 , n35989 );
xor ( n35991 , n35955 , n35990 );
xor ( n7180 , n35504 , n35592 );
and ( n7181 , n7180 , n35640 );
and ( n35994 , n35504 , n35592 );
or ( n7186 , n7181 , n35994 );
buf ( n35996 , n7186 );
buf ( n35997 , n35996 );
xor ( n7189 , n35991 , n35997 );
buf ( n35999 , n7189 );
buf ( n36000 , n35999 );
xor ( n7192 , n7095 , n36000 );
buf ( n36002 , n7192 );
nor ( n7194 , n35818 , n36002 );
xor ( n7195 , n35643 , n35714 );
xor ( n7196 , n7195 , n35814 );
buf ( n36006 , n7196 );
xor ( n7198 , n33637 , n33681 );
and ( n7199 , n7198 , n33688 );
and ( n7200 , n33637 , n33681 );
or ( n7201 , n7199 , n7200 );
buf ( n36011 , n7201 );
not ( n7203 , n36011 );
not ( n7204 , n7203 );
not ( n7205 , n7204 );
xor ( n7206 , n35793 , n6980 );
xor ( n7207 , n7206 , n35807 );
not ( n7208 , n7207 );
nand ( n7209 , n7205 , n7208 );
not ( n7210 , n7209 );
xor ( n7211 , n35649 , n35702 );
xor ( n7212 , n7211 , n35709 );
buf ( n36022 , n7212 );
not ( n7214 , n36022 );
or ( n7215 , n7210 , n7214 );
not ( n7216 , n7208 );
nand ( n7217 , n7204 , n7216 );
nand ( n7218 , n7215 , n7217 );
nor ( n7219 , n36006 , n7218 );
nor ( n7220 , n7194 , n7219 );
not ( n7221 , n7220 );
not ( n7222 , n4616 );
not ( n7223 , n4612 );
or ( n7224 , n7222 , n7223 );
xor ( n7225 , n33607 , n33691 );
and ( n7226 , n7225 , n33697 );
and ( n7227 , n33607 , n33691 );
or ( n7228 , n7226 , n7227 );
buf ( n36038 , n7228 );
not ( n7230 , n36038 );
xor ( n36040 , n7207 , n36011 );
xnor ( n7232 , n36040 , n36022 );
nand ( n7233 , n7230 , n7232 );
nand ( n7234 , n33710 , n7233 );
not ( n7235 , n4592 );
not ( n7236 , n4600 );
nand ( n7237 , n7235 , n7236 );
nor ( n7238 , n7234 , n7237 );
nand ( n7239 , n7224 , n7238 );
not ( n7240 , n7234 );
and ( n7241 , n7240 , n4623 );
not ( n7242 , n4796 );
not ( n7243 , n7233 );
or ( n7244 , n7242 , n7243 );
not ( n7245 , n36022 );
not ( n7246 , n7203 );
not ( n7247 , n7216 );
or ( n7248 , n7246 , n7247 );
nand ( n7249 , n7208 , n36011 );
nand ( n7250 , n7248 , n7249 );
not ( n7251 , n7250 );
not ( n7252 , n7251 );
or ( n7253 , n7245 , n7252 );
not ( n7254 , n36022 );
nand ( n7255 , n7254 , n7250 );
nand ( n7256 , n7253 , n7255 );
not ( n7257 , n7230 );
nand ( n7258 , n7256 , n7257 );
nand ( n7259 , n7244 , n7258 );
nor ( n7260 , n7241 , n7259 );
nand ( n7261 , n7239 , n7260 );
not ( n7262 , n7261 );
or ( n7263 , n7221 , n7262 );
not ( n7264 , n7194 );
nand ( n7265 , n36002 , n35818 );
nand ( n7266 , n36006 , n7218 );
nand ( n36076 , n7265 , n7266 );
nand ( n36077 , n7264 , n36076 );
nand ( n7269 , n7263 , n36077 );
buf ( n36079 , n518 );
buf ( n36080 , n489 );
and ( n7275 , n36079 , n36080 );
buf ( n36082 , n7275 );
buf ( n36083 , n36082 );
not ( n7278 , n1999 );
not ( n36085 , n35883 );
or ( n7283 , n7278 , n36085 );
buf ( n36087 , n1865 );
xor ( n7285 , n499 , n506 );
buf ( n36089 , n7285 );
nand ( n7287 , n36087 , n36089 );
buf ( n36091 , n7287 );
nand ( n7289 , n7283 , n36091 );
buf ( n36093 , n7289 );
xor ( n7291 , n36083 , n36093 );
buf ( n36095 , n7044 );
not ( n7293 , n36095 );
buf ( n36097 , n33373 );
not ( n7295 , n36097 );
or ( n7296 , n7293 , n7295 );
buf ( n36100 , n31271 );
buf ( n36101 , n510 );
buf ( n36102 , n495 );
xor ( n7300 , n36101 , n36102 );
buf ( n36104 , n7300 );
buf ( n36105 , n36104 );
nand ( n7303 , n36100 , n36105 );
buf ( n36107 , n7303 );
buf ( n36108 , n36107 );
nand ( n7306 , n7296 , n36108 );
buf ( n36110 , n7306 );
buf ( n36111 , n36110 );
xor ( n7309 , n7291 , n36111 );
buf ( n36113 , n7309 );
buf ( n36114 , n36113 );
not ( n7312 , n35837 );
not ( n7313 , n6703 );
not ( n7314 , n4626 );
nand ( n7315 , n7313 , n7314 );
not ( n7316 , n7315 );
not ( n7317 , n7316 );
or ( n7318 , n7312 , n7317 );
buf ( n36122 , n4626 );
buf ( n36123 , n516 );
buf ( n36124 , n489 );
xor ( n7322 , n36123 , n36124 );
buf ( n36126 , n7322 );
buf ( n36127 , n36126 );
nand ( n7325 , n36122 , n36127 );
buf ( n36129 , n7325 );
nand ( n7327 , n7318 , n36129 );
xor ( n7328 , n7104 , n7327 );
not ( n7329 , n501 );
not ( n7330 , n1915 );
or ( n7331 , n7329 , n7330 );
nand ( n7332 , n35849 , n2160 );
nand ( n7333 , n7331 , n7332 );
not ( n7334 , n7333 );
xor ( n7335 , n7328 , n7334 );
buf ( n36139 , n7335 );
xor ( n7337 , n36114 , n36139 );
xor ( n7338 , n35961 , n35971 );
and ( n7339 , n7338 , n35987 );
and ( n7340 , n35961 , n35971 );
or ( n7341 , n7339 , n7340 );
buf ( n36145 , n7341 );
buf ( n36146 , n36145 );
xor ( n7344 , n7337 , n36146 );
buf ( n36148 , n7344 );
buf ( n36149 , n36148 );
xor ( n7347 , n35955 , n35990 );
and ( n7348 , n7347 , n35997 );
and ( n7349 , n35955 , n35990 );
or ( n7350 , n7348 , n7349 );
buf ( n36154 , n7350 );
buf ( n36155 , n36154 );
xor ( n7353 , n36149 , n36155 );
xor ( n36157 , n7105 , n35936 );
and ( n7355 , n36157 , n35953 );
and ( n36159 , n7105 , n35936 );
or ( n7360 , n7355 , n36159 );
xor ( n36161 , n35823 , n35824 );
and ( n7362 , n36161 , n35842 );
and ( n7363 , n35823 , n35824 );
or ( n36164 , n7362 , n7363 );
buf ( n36165 , n36164 );
not ( n7369 , n35947 );
not ( n7370 , n6769 );
or ( n7371 , n7369 , n7370 );
and ( n7372 , n512 , n493 );
not ( n7373 , n512 );
not ( n7374 , n493 );
and ( n7375 , n7373 , n7374 );
nor ( n7376 , n7372 , n7375 );
nand ( n7377 , n2591 , n7376 );
nand ( n7378 , n7371 , n7377 );
buf ( n36176 , n7378 );
not ( n7380 , n6669 );
not ( n7381 , n35915 );
or ( n7382 , n7380 , n7381 );
buf ( n36180 , n2081 );
buf ( n36181 , n508 );
buf ( n36182 , n497 );
xor ( n7386 , n36181 , n36182 );
buf ( n36184 , n7386 );
buf ( n36185 , n36184 );
nand ( n7389 , n36180 , n36185 );
buf ( n36187 , n7389 );
nand ( n7391 , n7382 , n36187 );
buf ( n36189 , n7391 );
xor ( n7393 , n36176 , n36189 );
buf ( n36191 , n35930 );
not ( n7395 , n36191 );
buf ( n36193 , n6779 );
not ( n7397 , n36193 );
or ( n7398 , n7395 , n7397 );
buf ( n36196 , n4286 );
buf ( n36197 , n514 );
buf ( n36198 , n491 );
xor ( n7402 , n36197 , n36198 );
buf ( n36200 , n7402 );
buf ( n36201 , n36200 );
nand ( n7405 , n36196 , n36201 );
buf ( n36203 , n7405 );
buf ( n36204 , n36203 );
nand ( n7408 , n7398 , n36204 );
buf ( n36206 , n7408 );
buf ( n36207 , n36206 );
xor ( n7411 , n7393 , n36207 );
buf ( n36209 , n7411 );
xor ( n7413 , n36165 , n36209 );
xor ( n7414 , n35855 , n35872 );
and ( n7415 , n7414 , n35890 );
and ( n7416 , n35855 , n35872 );
or ( n7417 , n7415 , n7416 );
buf ( n36215 , n7417 );
xor ( n7419 , n7413 , n36215 );
xor ( n7420 , n7360 , n7419 );
xor ( n7421 , n35845 , n35893 );
and ( n7422 , n7421 , n35900 );
and ( n7423 , n35845 , n35893 );
or ( n7424 , n7422 , n7423 );
buf ( n36222 , n7424 );
xor ( n7426 , n7420 , n36222 );
buf ( n36224 , n7426 );
xor ( n7428 , n7353 , n36224 );
buf ( n36226 , n7428 );
xor ( n7433 , n35903 , n35909 );
and ( n36228 , n7433 , n36000 );
and ( n7435 , n35903 , n35909 );
or ( n7436 , n36228 , n7435 );
buf ( n36231 , n7436 );
nor ( n7441 , n36226 , n36231 );
not ( n7442 , n7441 );
nand ( n7443 , n36226 , n36231 );
nand ( n7444 , n7442 , n7443 );
not ( n7445 , n7444 );
and ( n7446 , n7269 , n7445 );
not ( n7447 , n7269 );
and ( n7448 , n7447 , n7444 );
nor ( n7449 , n7446 , n7448 );
nand ( n7450 , n7449 , n2815 );
not ( n7451 , n7450 );
nand ( n7452 , n1488 , n489 );
not ( n7453 , n7452 );
xor ( n7454 , n503 , n7453 );
buf ( n7455 , n5328 );
not ( n7456 , n7455 );
not ( n7457 , n489 );
not ( n7458 , n29797 );
or ( n7459 , n7457 , n7458 );
buf ( n36251 , n712 );
not ( n7461 , n489 );
buf ( n36253 , n7461 );
nand ( n7463 , n36251 , n36253 );
buf ( n36255 , n7463 );
nand ( n7465 , n7459 , n36255 );
not ( n7466 , n7465 );
or ( n7467 , n7456 , n7466 );
not ( n7468 , n489 );
not ( n7469 , n827 );
or ( n7470 , n7468 , n7469 );
or ( n7471 , n827 , n489 );
nand ( n36263 , n7470 , n7471 );
xnor ( n7473 , n490 , n489 );
nor ( n7474 , n5328 , n7473 );
nand ( n7475 , n36263 , n7474 );
nand ( n7476 , n7467 , n7475 );
xnor ( n7477 , n7454 , n7476 );
buf ( n36269 , n7477 );
not ( n7479 , n29737 );
not ( n7480 , n501 );
not ( n7481 , n456 );
not ( n7482 , n473 );
nand ( n7483 , n7481 , n7482 );
not ( n7484 , n457 );
nand ( n7485 , n7484 , n456 );
nand ( n7486 , n7483 , n7485 );
not ( n7487 , n7486 );
or ( n7488 , n7480 , n7487 );
not ( n7489 , n501 );
nand ( n7490 , n7485 , n7489 , n7483 );
nand ( n7491 , n7488 , n7490 );
not ( n36283 , n7491 );
or ( n7496 , n7479 , n36283 );
buf ( n36285 , n501 );
not ( n7498 , n36285 );
and ( n7499 , n456 , n458 );
not ( n36288 , n456 );
and ( n7504 , n36288 , n474 );
nor ( n7505 , n7499 , n7504 );
buf ( n36291 , n7505 );
not ( n7507 , n36291 );
or ( n7508 , n7498 , n7507 );
nand ( n7509 , n456 , n458 );
not ( n7510 , n7509 );
not ( n7511 , n456 );
nand ( n7512 , n7511 , n474 );
not ( n7513 , n7512 );
or ( n7514 , n7510 , n7513 );
nand ( n7515 , n7514 , n29635 );
buf ( n36301 , n7515 );
nand ( n7517 , n7508 , n36301 );
buf ( n36303 , n7517 );
buf ( n36304 , n36303 );
buf ( n36305 , n693 );
nand ( n7521 , n36304 , n36305 );
buf ( n36307 , n7521 );
nand ( n7523 , n7496 , n36307 );
not ( n7524 , n29873 );
buf ( n36310 , n495 );
not ( n7526 , n36310 );
buf ( n36312 , n29505 );
not ( n7528 , n36312 );
buf ( n36314 , n7528 );
buf ( n36315 , n36314 );
not ( n7531 , n36315 );
or ( n7532 , n7526 , n7531 );
buf ( n36318 , n29505 );
buf ( n36319 , n29716 );
nand ( n7535 , n36318 , n36319 );
buf ( n36321 , n7535 );
buf ( n36322 , n36321 );
nand ( n7538 , n7532 , n36322 );
buf ( n36324 , n7538 );
not ( n7540 , n36324 );
or ( n7541 , n7524 , n7540 );
buf ( n36327 , n29844 );
buf ( n36328 , n495 );
not ( n7547 , n36328 );
buf ( n36330 , n4966 );
not ( n7549 , n36330 );
or ( n7550 , n7547 , n7549 );
or ( n36333 , n456 , n480 );
not ( n7555 , n464 );
nand ( n7556 , n7555 , n456 );
nand ( n7557 , n36333 , n29716 , n7556 );
buf ( n36337 , n7557 );
nand ( n7559 , n7550 , n36337 );
buf ( n36339 , n7559 );
buf ( n36340 , n36339 );
nand ( n7562 , n36327 , n36340 );
buf ( n36342 , n7562 );
nand ( n7564 , n7541 , n36342 );
xor ( n7565 , n7523 , n7564 );
not ( n7566 , n29596 );
not ( n7567 , n4906 );
not ( n7568 , n7567 );
or ( n7569 , n7566 , n7568 );
and ( n7570 , n456 , n460 );
not ( n7571 , n456 );
and ( n7572 , n7571 , n476 );
nor ( n7573 , n7570 , n7572 );
nand ( n7574 , n7573 , n499 );
nand ( n7575 , n7569 , n7574 );
not ( n36355 , n7575 );
not ( n7577 , n29624 );
or ( n7578 , n36355 , n7577 );
and ( n36358 , n456 , n459 );
not ( n7583 , n456 );
and ( n7584 , n7583 , n475 );
nor ( n7585 , n36358 , n7584 );
not ( n7586 , n7585 );
not ( n7587 , n499 );
or ( n7588 , n7586 , n7587 );
not ( n7589 , n499 );
nand ( n7590 , n7511 , n5060 );
not ( n7591 , n459 );
nand ( n7592 , n7591 , n456 );
nand ( n7593 , n7589 , n7590 , n7592 );
nand ( n7594 , n7588 , n7593 );
buf ( n36371 , n7594 );
buf ( n36372 , n29583 );
nand ( n7597 , n36371 , n36372 );
buf ( n36374 , n7597 );
nand ( n7602 , n7578 , n36374 );
xor ( n7603 , n7565 , n7602 );
buf ( n36377 , n7603 );
xor ( n7605 , n36269 , n36377 );
buf ( n36379 , n490 );
not ( n7610 , n36379 );
buf ( n36381 , n29551 );
nand ( n36382 , n7610 , n36381 );
buf ( n36383 , n36382 );
buf ( n36384 , n36383 );
buf ( n36385 , n491 );
and ( n7619 , n36384 , n36385 );
buf ( n36387 , n490 );
not ( n36388 , n36387 );
buf ( n36389 , n777 );
not ( n7623 , n36389 );
or ( n36391 , n36388 , n7623 );
buf ( n36392 , n489 );
nand ( n7629 , n36391 , n36392 );
buf ( n36394 , n7629 );
buf ( n36395 , n36394 );
nor ( n7632 , n7619 , n36395 );
buf ( n36397 , n7632 );
buf ( n36398 , n36397 );
buf ( n36399 , n504 );
not ( n36400 , n36399 );
nand ( n7640 , n7483 , n7485 );
not ( n7641 , n503 );
xor ( n36403 , n7640 , n7641 );
buf ( n36404 , n36403 );
not ( n36405 , n36404 );
or ( n36406 , n36400 , n36405 );
nand ( n36407 , n5343 , n4911 );
buf ( n36408 , n36407 );
nand ( n36409 , n36406 , n36408 );
buf ( n36410 , n36409 );
buf ( n36411 , n36410 );
and ( n36412 , n36398 , n36411 );
buf ( n36413 , n36412 );
buf ( n36414 , n36413 );
not ( n36415 , n29668 );
not ( n36416 , n7489 );
not ( n36417 , n5062 );
or ( n36418 , n36416 , n36417 );
nand ( n36419 , n7585 , n501 );
nand ( n36420 , n36418 , n36419 );
not ( n36421 , n36420 );
or ( n36422 , n36415 , n36421 );
not ( n36423 , n5352 );
not ( n36424 , n5359 );
or ( n36425 , n36423 , n36424 );
nand ( n36426 , n36425 , n693 );
nand ( n36427 , n36422 , n36426 );
buf ( n36428 , n36427 );
not ( n36429 , n36428 );
buf ( n36430 , n36429 );
buf ( n36431 , n36430 );
not ( n36432 , n36431 );
buf ( n36433 , n489 );
not ( n36434 , n36433 );
buf ( n36435 , n36434 );
or ( n36436 , n795 , n36435 );
not ( n36437 , n487 );
nand ( n36438 , n36437 , n7511 );
not ( n36439 , n471 );
nand ( n36440 , n36439 , n456 );
nand ( n36441 , n36438 , n36440 , n7461 );
nand ( n36442 , n36436 , n36441 );
not ( n36443 , n36442 );
not ( n36444 , n7455 );
or ( n36445 , n36443 , n36444 );
not ( n36446 , n7461 );
and ( n36447 , n456 , n472 );
not ( n36448 , n456 );
and ( n36449 , n36448 , n488 );
nor ( n36450 , n36447 , n36449 );
not ( n36451 , n36450 );
not ( n36452 , n36451 );
or ( n36453 , n36446 , n36452 );
or ( n36454 , n36451 , n36435 );
nand ( n36455 , n36453 , n36454 );
nor ( n36456 , n7473 , n5328 );
nand ( n36457 , n36455 , n36456 );
nand ( n36458 , n36445 , n36457 );
buf ( n36459 , n36458 );
not ( n36460 , n36459 );
buf ( n36461 , n36460 );
buf ( n36462 , n36461 );
not ( n36463 , n36462 );
or ( n36464 , n36432 , n36463 );
buf ( n36465 , n29829 );
not ( n36466 , n36465 );
not ( n36467 , n497 );
not ( n36468 , n34073 );
or ( n36469 , n36467 , n36468 );
buf ( n36470 , n29505 );
buf ( n36471 , n706 );
nand ( n36472 , n36470 , n36471 );
buf ( n36473 , n36472 );
nand ( n36474 , n36469 , n36473 );
buf ( n36475 , n36474 );
not ( n36476 , n36475 );
or ( n36477 , n36466 , n36476 );
buf ( n36478 , n835 );
buf ( n36479 , n34355 );
nand ( n36480 , n36478 , n36479 );
buf ( n36481 , n36480 );
buf ( n36482 , n36481 );
nand ( n36483 , n36477 , n36482 );
buf ( n36484 , n36483 );
buf ( n36485 , n36484 );
nand ( n36486 , n36464 , n36485 );
buf ( n36487 , n36486 );
buf ( n36488 , n36487 );
nand ( n36489 , n36427 , n36458 );
buf ( n36490 , n36489 );
nand ( n36491 , n36488 , n36490 );
buf ( n36492 , n36491 );
buf ( n36493 , n36492 );
xor ( n36494 , n36414 , n36493 );
not ( n36495 , n29522 );
and ( n36496 , n1204 , n29537 );
not ( n36497 , n1204 );
and ( n36498 , n36497 , n493 );
or ( n36499 , n36496 , n36498 );
not ( n36500 , n36499 );
or ( n36501 , n36495 , n36500 );
nand ( n36502 , n5443 , n29576 );
nand ( n36503 , n36501 , n36502 );
not ( n36504 , n30072 );
not ( n36505 , n34383 );
or ( n36506 , n36504 , n36505 );
not ( n36507 , n495 );
not ( n36508 , n1147 );
or ( n36509 , n36507 , n36508 );
not ( n36510 , n1155 );
nand ( n36511 , n7511 , n481 );
not ( n36512 , n36511 );
or ( n36513 , n36510 , n36512 );
nand ( n36514 , n36513 , n29716 );
nand ( n36515 , n36509 , n36514 );
buf ( n36516 , n36515 );
buf ( n36517 , n29873 );
nand ( n36518 , n36516 , n36517 );
buf ( n36519 , n36518 );
nand ( n36520 , n36506 , n36519 );
xor ( n36521 , n36503 , n36520 );
not ( n36522 , n29624 );
not ( n36523 , n5521 );
or ( n36524 , n36522 , n36523 );
not ( n36525 , n499 );
not ( n36526 , n29511 );
not ( n36527 , n36526 );
or ( n36528 , n36525 , n36527 );
buf ( n36529 , n29511 );
buf ( n36530 , n29596 );
nand ( n36531 , n36529 , n36530 );
buf ( n36532 , n36531 );
nand ( n36533 , n36528 , n36532 );
buf ( n36534 , n36533 );
buf ( n36535 , n29583 );
nand ( n36536 , n36534 , n36535 );
buf ( n36537 , n36536 );
nand ( n36538 , n36524 , n36537 );
and ( n36539 , n36521 , n36538 );
and ( n36540 , n36503 , n36520 );
or ( n36541 , n36539 , n36540 );
buf ( n36542 , n36541 );
and ( n36543 , n36494 , n36542 );
and ( n36544 , n36414 , n36493 );
or ( n36545 , n36543 , n36544 );
buf ( n36546 , n36545 );
buf ( n36547 , n36546 );
xor ( n36548 , n7605 , n36547 );
buf ( n36549 , n36548 );
buf ( n36550 , n29576 );
not ( n36551 , n36550 );
not ( n36552 , n493 );
not ( n36553 , n1260 );
or ( n36554 , n36552 , n36553 );
or ( n36555 , n1260 , n493 );
nand ( n36556 , n36554 , n36555 );
buf ( n36557 , n36556 );
not ( n36558 , n36557 );
or ( n36559 , n36551 , n36558 );
buf ( n36560 , n493 );
not ( n36561 , n36560 );
buf ( n36562 , n29591 );
not ( n36563 , n36562 );
or ( n36564 , n36561 , n36563 );
buf ( n36565 , n29742 );
not ( n36566 , n36565 );
buf ( n36567 , n29537 );
nand ( n36568 , n36566 , n36567 );
buf ( n36569 , n36568 );
buf ( n36570 , n36569 );
nand ( n36571 , n36564 , n36570 );
buf ( n36572 , n36571 );
buf ( n36573 , n36572 );
buf ( n36574 , n29522 );
nand ( n36575 , n36573 , n36574 );
buf ( n36576 , n36575 );
buf ( n36577 , n36576 );
nand ( n36578 , n36559 , n36577 );
buf ( n36579 , n36578 );
buf ( n36580 , n36579 );
buf ( n36581 , n34031 );
not ( n36582 , n36581 );
not ( n36583 , n491 );
and ( n36584 , n456 , n468 );
not ( n36585 , n456 );
and ( n36586 , n36585 , n484 );
or ( n36587 , n36584 , n36586 );
or ( n36588 , n36583 , n36587 );
nand ( n36589 , n33936 , n36587 );
nand ( n36590 , n36588 , n36589 );
buf ( n36591 , n36590 );
not ( n36592 , n36591 );
or ( n36593 , n36582 , n36592 );
and ( n36594 , n1204 , n33936 );
not ( n36595 , n1204 );
and ( n36596 , n36595 , n491 );
or ( n36597 , n36594 , n36596 );
buf ( n36598 , n36597 );
buf ( n36599 , n4821 );
nand ( n36600 , n36598 , n36599 );
buf ( n36601 , n36600 );
buf ( n36602 , n36601 );
nand ( n36603 , n36593 , n36602 );
buf ( n36604 , n36603 );
buf ( n36605 , n36604 );
xor ( n36606 , n36580 , n36605 );
not ( n36607 , n835 );
not ( n36608 , n706 );
not ( n36609 , n5519 );
or ( n36610 , n36608 , n36609 );
not ( n36611 , n925 );
not ( n36612 , n36611 );
nand ( n36613 , n36612 , n497 );
nand ( n36614 , n36610 , n36613 );
not ( n36615 , n36614 );
or ( n36616 , n36607 , n36615 );
buf ( n36617 , n497 );
not ( n36618 , n36617 );
buf ( n36619 , n29510 );
not ( n36620 , n36619 );
or ( n36621 , n36618 , n36620 );
buf ( n36622 , n29511 );
buf ( n36623 , n706 );
nand ( n36624 , n36622 , n36623 );
buf ( n36625 , n36624 );
buf ( n36626 , n36625 );
nand ( n36627 , n36621 , n36626 );
buf ( n36628 , n36627 );
buf ( n36629 , n36628 );
buf ( n36630 , n29829 );
nand ( n36631 , n36629 , n36630 );
buf ( n36632 , n36631 );
nand ( n36633 , n36616 , n36632 );
buf ( n36634 , n36633 );
not ( n36635 , n36634 );
buf ( n36636 , n36635 );
buf ( n36637 , n36636 );
xor ( n36638 , n36606 , n36637 );
buf ( n36639 , n36638 );
buf ( n36640 , n36639 );
buf ( n36641 , n29678 );
buf ( n36642 , n489 );
and ( n36643 , n36641 , n36642 );
buf ( n36644 , n36643 );
buf ( n36645 , n36644 );
and ( n36646 , n456 , n457 );
not ( n36647 , n456 );
and ( n36648 , n36647 , n473 );
nor ( n36649 , n36646 , n36648 );
and ( n36650 , n847 , n36649 );
and ( n36651 , n504 , n503 );
nor ( n36652 , n36650 , n36651 );
nand ( n36653 , C1 , n36652 );
buf ( n36654 , n36653 );
xor ( n36655 , n36645 , n36654 );
buf ( n36656 , n693 );
not ( n36657 , n36656 );
buf ( n36658 , n36420 );
not ( n36659 , n36658 );
or ( n36660 , n36657 , n36659 );
buf ( n36661 , n36303 );
buf ( n36662 , n29737 );
nand ( n36663 , n36661 , n36662 );
buf ( n36664 , n36663 );
buf ( n36665 , n36664 );
nand ( n36666 , n36660 , n36665 );
buf ( n36667 , n36666 );
buf ( n36668 , n36667 );
and ( n36669 , n36655 , n36668 );
and ( n36670 , n36645 , n36654 );
or ( n36671 , n36669 , n36670 );
buf ( n36672 , n36671 );
buf ( n36673 , n36672 );
not ( n36674 , n29522 );
not ( n36675 , n36556 );
or ( n36676 , n36674 , n36675 );
not ( n36677 , n493 );
not ( n36678 , n29569 );
or ( n36679 , n36677 , n36678 );
nand ( n36680 , n36679 , n29574 );
not ( n36681 , n36680 );
nand ( n36682 , n36499 , n36681 );
nand ( n36683 , n36676 , n36682 );
buf ( n36684 , n36683 );
not ( n36685 , n36684 );
not ( n36686 , n4821 );
not ( n36687 , n36590 );
or ( n36688 , n36686 , n36687 );
and ( n36689 , n712 , n33936 );
not ( n36690 , n712 );
and ( n36691 , n36690 , n491 );
or ( n36692 , n36689 , n36691 );
buf ( n36693 , n36692 );
buf ( n36694 , n33725 );
buf ( n36695 , n5134 );
nor ( n36696 , n36694 , n36695 );
buf ( n36697 , n36696 );
nand ( n36698 , n36693 , n36697 );
buf ( n36699 , n36698 );
nand ( n36700 , n36688 , n36699 );
buf ( n36701 , n36700 );
not ( n36702 , n36701 );
or ( n36703 , n36685 , n36702 );
buf ( n36704 , n36700 );
buf ( n36705 , n36683 );
or ( n36706 , n36704 , n36705 );
not ( n36707 , n1627 );
not ( n36708 , n7575 );
or ( n36709 , n36707 , n36708 );
nor ( n36710 , n29581 , n29622 );
nand ( n36711 , n36533 , n36710 );
nand ( n36712 , n36709 , n36711 );
buf ( n36713 , n36712 );
nand ( n36714 , n36706 , n36713 );
buf ( n36715 , n36714 );
buf ( n36716 , n36715 );
nand ( n36717 , n36703 , n36716 );
buf ( n36718 , n36717 );
buf ( n36719 , n36718 );
xor ( n36720 , n36673 , n36719 );
not ( n36721 , n36456 );
not ( n36722 , n36442 );
or ( n36723 , n36721 , n36722 );
not ( n36724 , n490 );
not ( n36725 , n36583 );
or ( n36726 , n36724 , n36725 );
not ( n36727 , n490 );
nand ( n36728 , n36727 , n491 );
nand ( n36729 , n36726 , n36728 );
nand ( n36730 , n36729 , n36263 );
nand ( n36731 , n36723 , n36730 );
buf ( n36732 , n36731 );
not ( n36733 , n29873 );
not ( n36734 , n36339 );
or ( n36735 , n36733 , n36734 );
nand ( n36736 , n36515 , n29844 );
nand ( n36737 , n36735 , n36736 );
buf ( n36738 , n36737 );
xor ( n36739 , n36732 , n36738 );
not ( n36740 , n835 );
not ( n36741 , n36474 );
or ( n36742 , n36740 , n36741 );
and ( n36743 , n497 , n36611 );
not ( n36744 , n29829 );
nor ( n36745 , n36743 , n36744 );
or ( n36746 , n5519 , n497 );
nand ( n36747 , n36745 , n36746 );
nand ( n36748 , n36742 , n36747 );
buf ( n36749 , n36748 );
and ( n36750 , n36739 , n36749 );
and ( n36751 , n36732 , n36738 );
or ( n36752 , n36750 , n36751 );
buf ( n36753 , n36752 );
buf ( n36754 , n36753 );
xor ( n36755 , n36720 , n36754 );
buf ( n36756 , n36755 );
buf ( n36757 , n36756 );
xor ( n36758 , n36640 , n36757 );
xor ( n36759 , n36645 , n36654 );
xor ( n36760 , n36759 , n36668 );
buf ( n36761 , n36760 );
buf ( n36762 , n36761 );
xor ( n36763 , n36732 , n36738 );
xor ( n36764 , n36763 , n36749 );
buf ( n36765 , n36764 );
buf ( n36766 , n36765 );
xor ( n36767 , n36762 , n36766 );
buf ( n36768 , n36700 );
buf ( n36769 , n36683 );
xor ( n36770 , n36768 , n36769 );
buf ( n36771 , n36770 );
buf ( n36772 , n36771 );
buf ( n36773 , n36712 );
xor ( n36774 , n36772 , n36773 );
buf ( n36775 , n36774 );
buf ( n36776 , n36775 );
and ( n36777 , n36767 , n36776 );
and ( n36778 , n36762 , n36766 );
or ( n36779 , n36777 , n36778 );
buf ( n36780 , n36779 );
buf ( n36781 , n36780 );
xor ( n36782 , n36758 , n36781 );
buf ( n36783 , n36782 );
xor ( n36784 , n36549 , n36783 );
buf ( n36785 , n34031 );
not ( n36786 , n36785 );
buf ( n36787 , n34300 );
not ( n36788 , n36787 );
or ( n36789 , n36786 , n36788 );
buf ( n36790 , n36692 );
buf ( n36791 , n4821 );
nand ( n36792 , n36790 , n36791 );
buf ( n36793 , n36792 );
buf ( n36794 , n36793 );
nand ( n36795 , n36789 , n36794 );
buf ( n36796 , n36795 );
buf ( n36797 , n36796 );
xor ( n36798 , n36398 , n36411 );
buf ( n36799 , n36798 );
buf ( n36800 , n36799 );
xor ( n36801 , n36797 , n36800 );
not ( n36802 , n504 );
not ( n36803 , n5343 );
or ( n36804 , n36802 , n36803 );
nand ( n36805 , n5333 , n4911 );
nand ( n36806 , n36804 , n36805 );
or ( n36807 , n36806 , n34218 );
nand ( n36808 , n36807 , n34252 );
buf ( n36809 , n36808 );
nand ( n36810 , n36806 , n34218 );
buf ( n36811 , n36810 );
nand ( n36812 , n36809 , n36811 );
buf ( n36813 , n36812 );
buf ( n36814 , n36813 );
and ( n36815 , n36801 , n36814 );
and ( n36816 , n36797 , n36800 );
or ( n36817 , n36815 , n36816 );
buf ( n36818 , n36817 );
xor ( n36819 , n36414 , n36493 );
xor ( n36820 , n36819 , n36542 );
buf ( n36821 , n36820 );
xor ( n36822 , n36818 , n36821 );
buf ( n36823 , n5523 );
buf ( n36824 , n34366 );
buf ( n36825 , n34390 );
nor ( n36826 , n36824 , n36825 );
buf ( n36827 , n36826 );
buf ( n36828 , n36827 );
or ( n36829 , n36823 , n36828 );
buf ( n36830 , n34366 );
buf ( n36831 , n34390 );
nand ( n36832 , n36830 , n36831 );
buf ( n36833 , n36832 );
buf ( n36834 , n36833 );
nand ( n36835 , n36829 , n36834 );
buf ( n36836 , n36835 );
buf ( n36837 , n36836 );
buf ( n36838 , n36484 );
not ( n36839 , n36838 );
buf ( n36840 , n36839 );
buf ( n36841 , n36840 );
not ( n36842 , n36841 );
buf ( n36843 , n36458 );
not ( n36844 , n36843 );
buf ( n36845 , n36430 );
not ( n36846 , n36845 );
or ( n36847 , n36844 , n36846 );
buf ( n36848 , n36430 );
buf ( n36849 , n36458 );
or ( n36850 , n36848 , n36849 );
nand ( n36851 , n36847 , n36850 );
buf ( n36852 , n36851 );
buf ( n36853 , n36852 );
not ( n36854 , n36853 );
or ( n36855 , n36842 , n36854 );
buf ( n36856 , n36852 );
buf ( n36857 , n36840 );
or ( n36858 , n36856 , n36857 );
nand ( n36859 , n36855 , n36858 );
buf ( n36860 , n36859 );
buf ( n36861 , n36860 );
xor ( n36862 , n36837 , n36861 );
xor ( n36863 , n36503 , n36520 );
xor ( n36864 , n36863 , n36538 );
buf ( n36865 , n36864 );
and ( n36866 , n36862 , n36865 );
and ( n36867 , n36837 , n36861 );
or ( n36868 , n36866 , n36867 );
buf ( n36869 , n36868 );
and ( n36870 , n36822 , n36869 );
and ( n36871 , n36818 , n36821 );
or ( n36872 , n36870 , n36871 );
xor ( n36873 , n36784 , n36872 );
not ( n36874 , n36873 );
xor ( n36875 , n34311 , n34330 );
and ( n36876 , n36875 , n34338 );
and ( n36877 , n34311 , n34330 );
or ( n36878 , n36876 , n36877 );
buf ( n36879 , n36878 );
buf ( n36880 , n36879 );
xor ( n36881 , n36797 , n36800 );
xor ( n36882 , n36881 , n36814 );
buf ( n36883 , n36882 );
buf ( n36884 , n36883 );
xor ( n36885 , n36880 , n36884 );
buf ( n36886 , n34256 );
not ( n36887 , n36886 );
buf ( n36888 , n5324 );
not ( n36889 , n36888 );
buf ( n36890 , n36889 );
buf ( n36891 , n36890 );
not ( n36892 , n36891 );
or ( n36893 , n36887 , n36892 );
buf ( n36894 , n34253 );
not ( n36895 , n36894 );
buf ( n36896 , n5324 );
not ( n36897 , n36896 );
or ( n36898 , n36895 , n36897 );
buf ( n36899 , n34270 );
nand ( n36900 , n36898 , n36899 );
buf ( n36901 , n36900 );
buf ( n36902 , n36901 );
nand ( n36903 , n36893 , n36902 );
buf ( n36904 , n36903 );
buf ( n36905 , n36904 );
and ( n36906 , n36885 , n36905 );
and ( n36907 , n36880 , n36884 );
or ( n36908 , n36906 , n36907 );
buf ( n36909 , n36908 );
not ( n36910 , n36909 );
xor ( n36911 , n36762 , n36766 );
xor ( n36912 , n36911 , n36776 );
buf ( n36913 , n36912 );
not ( n36914 , n36913 );
nand ( n36915 , n36910 , n36914 );
not ( n36916 , n36915 );
xor ( n36917 , n36818 , n36821 );
xor ( n36918 , n36917 , n36869 );
not ( n36919 , n36918 );
or ( n36920 , n36916 , n36919 );
nand ( n36921 , n36913 , n36909 );
nand ( n36922 , n36920 , n36921 );
not ( n36923 , n36922 );
and ( n36924 , n36874 , n36923 );
xor ( n36925 , n36837 , n36861 );
xor ( n36926 , n36925 , n36865 );
buf ( n36927 , n36926 );
buf ( n36928 , n36927 );
xor ( n36929 , n34341 , n34408 );
and ( n36930 , n36929 , n34415 );
and ( n36931 , n34341 , n34408 );
or ( n36932 , n36930 , n36931 );
buf ( n36933 , n36932 );
buf ( n36934 , n36933 );
xor ( n36935 , n36928 , n36934 );
xor ( n36936 , n36880 , n36884 );
xor ( n36937 , n36936 , n36905 );
buf ( n36938 , n36937 );
buf ( n36939 , n36938 );
and ( n36940 , n36935 , n36939 );
and ( n36941 , n36928 , n36934 );
or ( n36942 , n36940 , n36941 );
buf ( n36943 , n36942 );
not ( n36944 , n36918 );
not ( n36945 , n36909 );
and ( n36946 , n36914 , n36945 );
not ( n36947 , n36914 );
and ( n36948 , n36947 , n36909 );
nor ( n36949 , n36946 , n36948 );
not ( n36950 , n36949 );
not ( n36951 , n36950 );
or ( n36952 , n36944 , n36951 );
not ( n36953 , n36918 );
nand ( n36954 , n36953 , n36949 );
nand ( n36955 , n36952 , n36954 );
nor ( n36956 , n36943 , n36955 );
nor ( n36957 , n36924 , n36956 );
not ( n36958 , n36957 );
not ( n36959 , n5537 );
not ( n36960 , n5542 );
and ( n36961 , n36959 , n36960 );
xor ( n36962 , n36928 , n36934 );
xor ( n36963 , n36962 , n36939 );
buf ( n36964 , n36963 );
not ( n36965 , n36964 );
xor ( n36966 , n34280 , n34285 );
and ( n36967 , n36966 , n34417 );
and ( n36968 , n34280 , n34285 );
or ( n36969 , n36967 , n36968 );
not ( n36970 , n36969 );
and ( n36971 , n36965 , n36970 );
nor ( n36972 , n36961 , n36971 );
nand ( n36973 , n5299 , n36972 , n5287 );
not ( n36974 , n5310 );
and ( n36975 , n36974 , n36972 );
not ( n36976 , n5544 );
nand ( n36977 , n36965 , n36970 );
not ( n36978 , n36977 );
or ( n36979 , n36976 , n36978 );
buf ( n36980 , n36964 );
nand ( n36981 , n36980 , n36969 );
nand ( n36982 , n36979 , n36981 );
nor ( n36983 , n36975 , n36982 );
nand ( n36984 , n36973 , n36983 );
not ( n36985 , n36984 );
or ( n36986 , n36958 , n36985 );
nand ( n36987 , n36873 , n36922 );
nand ( n36988 , n36955 , n36943 );
nand ( n36989 , n36987 , n36988 );
not ( n36990 , n36873 );
not ( n36991 , n36922 );
nand ( n36992 , n36990 , n36991 );
nand ( n36993 , n36989 , n36992 );
buf ( n36994 , n36993 );
nand ( n36995 , n36986 , n36994 );
not ( n36996 , n1627 );
buf ( n36997 , n499 );
not ( n36998 , n36997 );
buf ( n36999 , n29498 );
not ( n37000 , n36999 );
or ( n37001 , n36998 , n37000 );
or ( n37002 , n456 , n474 );
not ( n37003 , n458 );
nand ( n37004 , n37003 , n456 );
nand ( n37005 , n29596 , n37002 , n37004 );
buf ( n37006 , n37005 );
nand ( n37007 , n37001 , n37006 );
buf ( n37008 , n37007 );
not ( n37009 , n37008 );
or ( n37010 , n36996 , n37009 );
nand ( n37011 , n7594 , n36710 );
nand ( n37012 , n37010 , n37011 );
buf ( n37013 , n37012 );
buf ( n37014 , n1332 );
not ( n37015 , n37014 );
buf ( n37016 , n489 );
nand ( n37017 , n37015 , n37016 );
buf ( n37018 , n37017 );
buf ( n37019 , n37018 );
not ( n37020 , n37019 );
buf ( n37021 , n37020 );
buf ( n37022 , n37021 );
and ( n37023 , n37013 , n37022 );
not ( n37024 , n37013 );
buf ( n37025 , n37018 );
and ( n37026 , n37024 , n37025 );
nor ( n37027 , n37023 , n37026 );
buf ( n37028 , n37027 );
buf ( n37029 , n37028 );
not ( n37030 , n29873 );
not ( n37031 , n36611 );
not ( n37032 , n29716 );
or ( n37033 , n37031 , n37032 );
and ( n37034 , n456 , n462 );
not ( n37035 , n456 );
and ( n37036 , n37035 , n478 );
nor ( n37037 , n37034 , n37036 );
nand ( n37038 , n37037 , n495 );
nand ( n37039 , n37033 , n37038 );
not ( n37040 , n37039 );
or ( n37041 , n37030 , n37040 );
not ( n37042 , n36321 );
nand ( n37043 , n495 , n36314 );
not ( n37044 , n37043 );
or ( n37045 , n37042 , n37044 );
nand ( n37046 , n37045 , n30072 );
nand ( n37047 , n37041 , n37046 );
buf ( n37048 , n37047 );
and ( n37049 , n37029 , n37048 );
not ( n37050 , n37029 );
buf ( n37051 , n37047 );
not ( n37052 , n37051 );
buf ( n37053 , n37052 );
buf ( n37054 , n37053 );
and ( n37055 , n37050 , n37054 );
nor ( n37056 , n37049 , n37055 );
buf ( n37057 , n37056 );
buf ( n37058 , n37057 );
not ( n37059 , n693 );
not ( n37060 , n7491 );
or ( n37061 , n37059 , n37060 );
buf ( n37062 , n29635 );
not ( n37063 , n37062 );
buf ( n37064 , n29647 );
nand ( n37065 , n37063 , n37064 );
buf ( n37066 , n37065 );
nand ( n37067 , n37061 , n37066 );
not ( n37068 , n37067 );
buf ( n37069 , n37068 );
nor ( n37070 , n5328 , n7473 );
buf ( n37071 , n37070 );
not ( n37072 , n37071 );
not ( n37073 , n7465 );
or ( n37074 , n37072 , n37073 );
buf ( n37075 , n489 );
not ( n37076 , n37075 );
buf ( n37077 , n734 );
not ( n37078 , n37077 );
or ( n37079 , n37076 , n37078 );
buf ( n37080 , n29493 );
buf ( n37081 , n7461 );
nand ( n37082 , n37080 , n37081 );
buf ( n37083 , n37082 );
buf ( n37084 , n37083 );
nand ( n37085 , n37079 , n37084 );
buf ( n37086 , n37085 );
buf ( n37087 , n37086 );
buf ( n37088 , n7455 );
nand ( n37089 , n37087 , n37088 );
buf ( n37090 , n37089 );
nand ( n37091 , n37074 , n37090 );
buf ( n37092 , n37091 );
xor ( n37093 , n37069 , n37092 );
buf ( n37094 , n36633 );
xor ( n37095 , n37093 , n37094 );
buf ( n37096 , n37095 );
buf ( n37097 , n37096 );
xor ( n37098 , n37058 , n37097 );
xor ( n37099 , n36673 , n36719 );
and ( n37100 , n37099 , n36754 );
and ( n37101 , n36673 , n36719 );
or ( n37102 , n37100 , n37101 );
buf ( n37103 , n37102 );
buf ( n37104 , n37103 );
xor ( n37105 , n37098 , n37104 );
buf ( n37106 , n37105 );
buf ( n37107 , n37106 );
xor ( n37108 , n36640 , n36757 );
and ( n37109 , n37108 , n36781 );
and ( n37110 , n36640 , n36757 );
or ( n37111 , n37109 , n37110 );
buf ( n37112 , n37111 );
buf ( n37113 , n37112 );
xor ( n37114 , n37107 , n37113 );
xor ( n37115 , n36580 , n36605 );
and ( n37116 , n37115 , n36637 );
and ( n37117 , n36580 , n36605 );
or ( n37118 , n37116 , n37117 );
buf ( n37119 , n37118 );
buf ( n37120 , n37119 );
not ( n37121 , n863 );
not ( n37122 , n7453 );
or ( n37123 , n37121 , n37122 );
not ( n37124 , n503 );
not ( n37125 , n7452 );
or ( n37126 , n37124 , n37125 );
nand ( n37127 , n37126 , n7476 );
nand ( n37128 , n37123 , n37127 );
xor ( n37129 , n7523 , n7564 );
and ( n37130 , n37129 , n7602 );
and ( n37131 , n7523 , n7564 );
or ( n37132 , n37130 , n37131 );
xor ( n37133 , n37128 , n37132 );
not ( n37134 , n36696 );
not ( n37135 , n36597 );
or ( n37136 , n37134 , n37135 );
or ( n37137 , n1261 , n36583 );
nand ( n37138 , n1261 , n33936 );
nand ( n37139 , n37137 , n37138 );
nand ( n37140 , n37139 , n4821 );
nand ( n37141 , n37136 , n37140 );
buf ( n37142 , n37141 );
buf ( n37143 , n29829 );
not ( n37144 , n37143 );
buf ( n37145 , n497 );
not ( n37146 , n37145 );
buf ( n37147 , n7573 );
not ( n37148 , n37147 );
or ( n37149 , n37146 , n37148 );
buf ( n37150 , n7567 );
buf ( n37151 , n706 );
nand ( n37152 , n37150 , n37151 );
buf ( n37153 , n37152 );
buf ( n37154 , n37153 );
nand ( n37155 , n37149 , n37154 );
buf ( n37156 , n37155 );
buf ( n37157 , n37156 );
not ( n37158 , n37157 );
or ( n37159 , n37144 , n37158 );
nand ( n37160 , n36628 , n29786 );
buf ( n37161 , n37160 );
nand ( n37162 , n37159 , n37161 );
buf ( n37163 , n37162 );
buf ( n37164 , n37163 );
xor ( n37165 , n37142 , n37164 );
buf ( n37166 , n29576 );
not ( n37167 , n37166 );
buf ( n37168 , n36572 );
not ( n37169 , n37168 );
or ( n37170 , n37167 , n37169 );
not ( n37171 , n493 );
not ( n37172 , n29658 );
or ( n37173 , n37171 , n37172 );
or ( n37174 , n493 , n29658 );
nand ( n37175 , n37173 , n37174 );
not ( n37176 , n37175 );
nand ( n37177 , n37176 , n29522 );
buf ( n37178 , n37177 );
nand ( n37179 , n37170 , n37178 );
buf ( n37180 , n37179 );
buf ( n37181 , n37180 );
xor ( n37182 , n37165 , n37181 );
buf ( n37183 , n37182 );
xor ( n37184 , n37133 , n37183 );
buf ( n37185 , n37184 );
xor ( n37186 , n37120 , n37185 );
xor ( n37187 , n36269 , n36377 );
and ( n37188 , n37187 , n36547 );
and ( n37189 , n36269 , n36377 );
or ( n37190 , n37188 , n37189 );
buf ( n37191 , n37190 );
buf ( n37192 , n37191 );
xor ( n37193 , n37186 , n37192 );
buf ( n37194 , n37193 );
buf ( n37195 , n37194 );
xor ( n37196 , n37114 , n37195 );
buf ( n37197 , n37196 );
xor ( n37198 , n36549 , n36783 );
and ( n37199 , n37198 , n36872 );
and ( n37200 , n36549 , n36783 );
or ( n37201 , n37199 , n37200 );
nor ( n37202 , n37197 , n37201 );
not ( n37203 , n37202 );
and ( n37204 , n37197 , n37201 );
not ( n37205 , n37204 );
and ( n37206 , n37203 , n37205 );
or ( n37207 , n36995 , n37206 );
nand ( n37208 , n36995 , n37206 );
nand ( n37209 , n37207 , n37208 , n455 );
not ( n37210 , n37209 );
or ( n37211 , n7451 , n37210 );
nand ( n37212 , n37211 , n454 );
not ( n37213 , n37212 );
or ( n37214 , n6637 , n37213 );
not ( n37215 , n3138 );
xor ( n37216 , n6103 , n35138 );
xor ( n37217 , n37216 , n35244 );
not ( n37218 , n37217 );
or ( n37219 , n37215 , n37218 );
nand ( n37220 , n454 , n538 );
nand ( n37221 , n37219 , n37220 );
not ( n37222 , n37221 );
not ( n37223 , n7194 );
buf ( n37224 , n7265 );
nand ( n37225 , n37223 , n37224 );
not ( n37226 , n37225 );
not ( n37227 , n7219 );
not ( n37228 , n37227 );
not ( n37229 , n7261 );
or ( n37230 , n37228 , n37229 );
buf ( n37231 , n7266 );
nand ( n37232 , n37230 , n37231 );
not ( n37233 , n37232 );
or ( n37234 , n37226 , n37233 );
or ( n37235 , n37232 , n37225 );
nand ( n37236 , n37234 , n37235 );
nand ( n37237 , n37236 , n5774 );
nand ( n37238 , n36987 , n36992 );
buf ( n37239 , n36988 );
buf ( n37240 , n37239 );
not ( n37241 , n36983 );
not ( n37242 , n36973 );
or ( n37243 , n37241 , n37242 );
or ( n37244 , n36955 , n36943 );
nand ( n37245 , n37243 , n37244 );
and ( n37246 , n37238 , n37240 , n37245 );
nand ( n37247 , n454 , n455 );
nor ( n37248 , n37246 , n37247 );
not ( n37249 , n37240 );
not ( n37250 , n37245 );
or ( n37251 , n37249 , n37250 );
not ( n37252 , n37238 );
nand ( n37253 , n37251 , n37252 );
nand ( n37254 , n37248 , n37253 );
xor ( n37255 , n35163 , n35169 );
xor ( n37256 , n37255 , n35174 );
buf ( n37257 , n37256 );
nor ( n37258 , n6293 , n6297 );
not ( n37259 , n6293 );
nor ( n37260 , n37259 , n35147 );
or ( n37261 , n37258 , n37260 );
not ( n37262 , n6307 );
nand ( n37263 , n37261 , n37262 );
not ( n37264 , n6298 );
nand ( n37265 , n37264 , n6307 );
nand ( n37266 , n6307 , n35147 , n6293 );
nand ( n37267 , n37263 , n37265 , n37266 );
xor ( n37268 , n35110 , n35118 );
xor ( n37269 , n37268 , n35127 );
and ( n37270 , n37267 , n37269 );
xor ( n37271 , n34453 , n34488 );
and ( n37272 , n37271 , n34495 );
and ( n37273 , n34453 , n34488 );
or ( n37274 , n37272 , n37273 );
buf ( n37275 , n37274 );
xor ( n37276 , n35110 , n35118 );
xor ( n37277 , n37276 , n35127 );
and ( n37278 , n37275 , n37277 );
and ( n37279 , n37267 , n37275 );
or ( n37280 , n37270 , n37278 , n37279 );
xor ( n37281 , n37257 , n37280 );
xor ( n37282 , n35000 , n35055 );
xor ( n37283 , n37282 , n35134 );
buf ( n37284 , n37283 );
and ( n37285 , n37281 , n37284 );
and ( n37286 , n37257 , n37280 );
or ( n37287 , n37285 , n37286 );
nand ( n37288 , n37287 , n3138 );
nand ( n37289 , n37222 , n37237 , n37254 , n37288 );
nand ( n37290 , n37214 , n37289 );
not ( n37291 , n37290 );
not ( n37292 , n454 );
not ( n37293 , n2815 );
nand ( n37294 , n37227 , n37231 );
not ( n37295 , n37294 );
and ( n37296 , n7261 , n37295 );
not ( n37297 , n7261 );
and ( n37298 , n37297 , n37294 );
nor ( n37299 , n37296 , n37298 );
not ( n37300 , n37299 );
or ( n37301 , n37293 , n37300 );
nand ( n37302 , n37244 , n37239 );
nand ( n37303 , n36984 , n37302 );
not ( n37304 , n37303 );
not ( n37305 , n36984 );
not ( n37306 , n37302 );
nand ( n37307 , n37305 , n37306 );
not ( n37308 , n37307 );
or ( n37309 , n37304 , n37308 );
nand ( n37310 , n37309 , n455 );
nand ( n37311 , n37301 , n37310 );
not ( n37312 , n37311 );
or ( n37313 , n37292 , n37312 );
xor ( n37314 , n5635 , n34527 );
xor ( n37315 , n37314 , n34544 );
and ( n37316 , n34601 , n37315 );
xor ( n37317 , n5635 , n34527 );
xor ( n37318 , n37317 , n34544 );
and ( n37319 , n34606 , n37318 );
and ( n37320 , n34601 , n34606 );
or ( n37321 , n37316 , n37319 , n37320 );
buf ( n37322 , n37321 );
xor ( n37323 , n34966 , n34989 );
xor ( n37324 , n37323 , n34995 );
buf ( n37325 , n37324 );
buf ( n37326 , n37325 );
xor ( n37327 , n37322 , n37326 );
xor ( n37328 , n35110 , n35118 );
xor ( n37329 , n37328 , n35127 );
xor ( n37330 , n37267 , n37275 );
xor ( n37331 , n37329 , n37330 );
buf ( n37332 , n37331 );
and ( n37333 , n37327 , n37332 );
and ( n37334 , n37322 , n37326 );
or ( n37335 , n37333 , n37334 );
buf ( n37336 , n37335 );
buf ( n37337 , n37336 );
buf ( n37338 , n3138 );
nand ( n37339 , n37337 , n37338 );
buf ( n37340 , n37339 );
nand ( n37341 , n37313 , n37340 );
buf ( n37342 , n539 );
not ( n37343 , n37342 );
buf ( n37344 , n454 );
not ( n37345 , n37344 );
or ( n37346 , n37343 , n37345 );
xor ( n37347 , n37257 , n37280 );
xor ( n37348 , n37347 , n37284 );
buf ( n37349 , n37348 );
buf ( n37350 , n3360 );
nand ( n37351 , n37349 , n37350 );
buf ( n37352 , n37351 );
buf ( n37353 , n37352 );
nand ( n37354 , n37346 , n37353 );
buf ( n37355 , n37354 );
buf ( n37356 , n37355 );
or ( n37357 , n37341 , n37356 );
not ( n37358 , n5547 );
not ( n37359 , n5312 );
or ( n37360 , n37358 , n37359 );
nand ( n37361 , n37360 , n5545 );
buf ( n37362 , n36977 );
and ( n37363 , n37362 , n36981 );
and ( n37364 , n37361 , n37363 );
not ( n37365 , n37361 );
not ( n37366 , n37363 );
and ( n37367 , n37365 , n37366 );
nor ( n37368 , n37364 , n37367 );
nand ( n37369 , n37368 , n3648 );
xor ( n37370 , n34447 , n34498 );
and ( n37371 , n37370 , n34609 );
and ( n37372 , n34447 , n34498 );
or ( n37373 , n37371 , n37372 );
buf ( n37374 , n37373 );
and ( n37375 , n37374 , n3138 );
not ( n37376 , n5847 );
xor ( n37377 , n37322 , n37326 );
xor ( n37378 , n37377 , n37332 );
buf ( n37379 , n37378 );
not ( n37380 , n37379 );
or ( n37381 , n37376 , n37380 );
nand ( n37382 , n454 , n540 );
nand ( n37383 , n37381 , n37382 );
nor ( n37384 , n37375 , n37383 );
not ( n37385 , n33710 );
not ( n37386 , n4625 );
or ( n37387 , n37385 , n37386 );
nand ( n37388 , n37387 , n33708 );
not ( n37389 , n7257 );
not ( n37390 , n7256 );
or ( n37391 , n37389 , n37390 );
nand ( n37392 , n37391 , n7233 );
and ( n37393 , n2815 , n37392 );
and ( n37394 , n37388 , n37393 );
not ( n37395 , n37388 );
not ( n37396 , n2815 );
nor ( n37397 , n37396 , n37392 );
and ( n37398 , n37395 , n37397 );
or ( n37399 , n37394 , n37398 );
nand ( n37400 , n37399 , n454 );
nand ( n37401 , n37369 , n37384 , n37400 );
nand ( n37402 , n37357 , n37401 );
not ( n37403 , n37402 );
nand ( n37404 , n5892 , n37291 , n37403 );
buf ( n37405 , n37311 );
nand ( n37406 , n37405 , n454 );
not ( n37407 , n37340 );
nor ( n37408 , n37407 , n37355 );
nand ( n37409 , n37406 , n37408 );
not ( n37410 , n454 );
not ( n37411 , n37399 );
or ( n37412 , n37410 , n37411 );
and ( n37413 , n37368 , n3648 );
nor ( n37414 , n37413 , n37375 );
nand ( n37415 , n37412 , n37414 );
nand ( n37416 , n37415 , n37383 );
not ( n37417 , n37416 );
nand ( n37418 , n37409 , n37417 );
not ( n37419 , n454 );
not ( n37420 , n37311 );
or ( n37421 , n37419 , n37420 );
nand ( n37422 , n37421 , n37340 );
nand ( n37423 , n37356 , n37422 );
not ( n37424 , n37253 );
nand ( n37425 , n37245 , n37240 );
or ( n37426 , n37425 , n37252 );
not ( n37427 , n37247 );
nand ( n37428 , n37426 , n37427 );
or ( n37429 , n37424 , n37428 );
nand ( n37430 , n37429 , n37288 );
not ( n37431 , n37237 );
or ( n37432 , n37430 , n37431 );
nand ( n37433 , n37432 , n37221 );
nand ( n37434 , n37418 , n37423 , n37433 );
nand ( n37435 , n37434 , n37291 );
not ( n37436 , n6400 );
not ( n37437 , n37212 );
or ( n37438 , n37436 , n37437 );
nand ( n37439 , n37438 , n6635 );
nand ( n37440 , n37404 , n37435 , n37439 );
buf ( n37441 , n37440 );
xor ( n37442 , n35256 , n35433 );
and ( n37443 , n37442 , n35468 );
and ( n37444 , n35256 , n35433 );
or ( n37445 , n37443 , n37444 );
buf ( n37446 , n37445 );
nand ( n37447 , n37446 , n3138 );
not ( n37448 , n37447 );
xor ( n37449 , n6599 , n6603 );
xor ( n37450 , n37449 , n35448 );
and ( n37451 , n6618 , n37450 );
xor ( n37452 , n6599 , n6603 );
xor ( n37453 , n37452 , n35448 );
and ( n37454 , n6626 , n37453 );
and ( n37455 , n6618 , n6626 );
or ( n37456 , n37451 , n37454 , n37455 );
buf ( n37457 , n37456 );
buf ( n37458 , n5636 );
buf ( n37459 , n35268 );
or ( n37460 , n37458 , n37459 );
buf ( n37461 , n4040 );
buf ( n37462 , n32981 );
buf ( n37463 , n528 );
and ( n37464 , n37462 , n37463 );
buf ( n37465 , n32183 );
buf ( n37466 , n543 );
and ( n37467 , n37465 , n37466 );
nor ( n37468 , n37464 , n37467 );
buf ( n37469 , n37468 );
buf ( n37470 , n37469 );
or ( n37471 , n37461 , n37470 );
nand ( n37472 , n37460 , n37471 );
buf ( n37473 , n37472 );
buf ( n37474 , n3020 );
buf ( n37475 , n35422 );
or ( n37476 , n37474 , n37475 );
buf ( n37477 , n31978 );
buf ( n37478 , n547 );
buf ( n37479 , n34779 );
and ( n37480 , n37478 , n37479 );
not ( n37481 , n37478 );
buf ( n37482 , n524 );
and ( n37483 , n37481 , n37482 );
nor ( n37484 , n37480 , n37483 );
buf ( n37485 , n37484 );
buf ( n37486 , n37485 );
or ( n37487 , n37477 , n37486 );
nand ( n37488 , n37476 , n37487 );
buf ( n37489 , n37488 );
not ( n37490 , n37489 );
not ( n37491 , n37490 );
nand ( n37492 , n35335 , n457 );
not ( n37493 , n37492 );
nand ( n37494 , n37473 , n37491 , n37493 );
not ( n37495 , n37473 );
nor ( n37496 , n37491 , n37492 );
nand ( n37497 , n37495 , n37496 );
nand ( n37498 , n37495 , n37491 , n37492 );
and ( n37499 , n37490 , n37492 );
nand ( n37500 , n37499 , n37473 );
nand ( n37501 , n37494 , n37497 , n37498 , n37500 );
not ( n37502 , n37501 );
buf ( n37503 , n3045 );
buf ( n37504 , n35312 );
or ( n37505 , n37503 , n37504 );
buf ( n37506 , n2918 );
buf ( n37507 , n31868 );
buf ( n37508 , n522 );
and ( n37509 , n37507 , n37508 );
buf ( n37510 , n35199 );
buf ( n37511 , n549 );
and ( n37512 , n37510 , n37511 );
nor ( n37513 , n37509 , n37512 );
buf ( n37514 , n37513 );
buf ( n37515 , n37514 );
or ( n37516 , n37506 , n37515 );
nand ( n37517 , n37505 , n37516 );
buf ( n37518 , n37517 );
buf ( n37519 , n37518 );
not ( n37520 , n6548 );
not ( n37521 , n6559 );
not ( n37522 , n37521 );
or ( n37523 , n37520 , n37522 );
buf ( n37524 , n537 );
buf ( n37525 , n32008 );
and ( n37526 , n37524 , n37525 );
not ( n37527 , n37524 );
buf ( n37528 , n534 );
and ( n37529 , n37527 , n37528 );
nor ( n37530 , n37526 , n37529 );
buf ( n37531 , n37530 );
or ( n37532 , n6337 , n37531 );
nand ( n37533 , n37523 , n37532 );
buf ( n37534 , n37533 );
xor ( n37535 , n37519 , n37534 );
not ( n37536 , n6305 );
buf ( n37537 , n6519 );
not ( n37538 , n37537 );
buf ( n37539 , n37538 );
not ( n37540 , n37539 );
or ( n37541 , n37536 , n37540 );
buf ( n37542 , n526 );
buf ( n37543 , n32053 );
and ( n37544 , n37542 , n37543 );
not ( n37545 , n37542 );
buf ( n37546 , n545 );
and ( n37547 , n37545 , n37546 );
nor ( n37548 , n37544 , n37547 );
buf ( n37549 , n37548 );
or ( n37550 , n37549 , n3087 );
nand ( n37551 , n37541 , n37550 );
buf ( n37552 , n37551 );
xor ( n37553 , n37535 , n37552 );
buf ( n37554 , n37553 );
not ( n37555 , n37554 );
nor ( n37556 , n37502 , n37555 );
not ( n37557 , n6016 );
buf ( n37558 , n37557 );
buf ( n37559 , n35381 );
or ( n37560 , n37558 , n37559 );
buf ( n37561 , n6010 );
buf ( n37562 , n6001 );
buf ( n37563 , n532 );
and ( n37564 , n37562 , n37563 );
buf ( n37565 , n31908 );
buf ( n37566 , n539 );
and ( n37567 , n37565 , n37566 );
nor ( n37568 , n37564 , n37567 );
buf ( n37569 , n37568 );
buf ( n37570 , n37569 );
or ( n37571 , n37561 , n37570 );
nand ( n37572 , n37560 , n37571 );
buf ( n37573 , n37572 );
buf ( n37574 , n37573 );
buf ( n37575 , n5582 );
buf ( n37576 , n35291 );
or ( n37577 , n37575 , n37576 );
buf ( n37578 , n33118 );
buf ( n37579 , n541 );
buf ( n37580 , n31853 );
and ( n37581 , n37579 , n37580 );
not ( n37582 , n37579 );
buf ( n37583 , n530 );
and ( n37584 , n37582 , n37583 );
nor ( n37585 , n37581 , n37584 );
buf ( n37586 , n37585 );
buf ( n37587 , n37586 );
or ( n37588 , n37578 , n37587 );
nand ( n37589 , n37577 , n37588 );
buf ( n37590 , n37589 );
buf ( n37591 , n37590 );
xor ( n37592 , n37574 , n37591 );
buf ( n37593 , n536 );
buf ( n37594 , n537 );
and ( n37595 , n37593 , n37594 );
buf ( n37596 , n37595 );
buf ( n37597 , n37596 );
buf ( n37598 , n2962 );
buf ( n37599 , n35350 );
or ( n37600 , n37598 , n37599 );
buf ( n37601 , n2848 );
buf ( n37602 , n2845 );
or ( n37603 , n37601 , n37602 );
nand ( n37604 , n37600 , n37603 );
buf ( n37605 , n37604 );
buf ( n37606 , n37605 );
xor ( n37607 , n37597 , n37606 );
buf ( n37608 , n37607 );
buf ( n37609 , n37608 );
xor ( n37610 , n37592 , n37609 );
buf ( n37611 , n37610 );
nand ( n37612 , n37556 , n37611 );
nand ( n37613 , n37502 , n37555 , n37611 );
not ( n37614 , n37611 );
nand ( n37615 , n37501 , n37614 , n37555 );
nand ( n37616 , n37502 , n37554 , n37614 );
nand ( n37617 , n37612 , n37613 , n37615 , n37616 );
buf ( n37618 , n37617 );
xor ( n37619 , n37457 , n37618 );
xor ( n37620 , n35320 , n35368 );
and ( n37621 , n37620 , n35430 );
and ( n37622 , n35320 , n35368 );
or ( n37623 , n37621 , n37622 );
buf ( n37624 , n37623 );
buf ( n37625 , n37624 );
xor ( n37626 , n6599 , n6603 );
and ( n37627 , n37626 , n35448 );
and ( n37628 , n6599 , n6603 );
or ( n37629 , n37627 , n37628 );
buf ( n37630 , n37629 );
xor ( n37631 , n37625 , n37630 );
xor ( n37632 , n35273 , n35296 );
and ( n37633 , n37632 , n35317 );
and ( n37634 , n35273 , n35296 );
or ( n37635 , n37633 , n37634 );
buf ( n37636 , n37635 );
buf ( n37637 , n37636 );
not ( n37638 , n6491 );
nand ( n37639 , n37638 , n6513 );
not ( n37640 , n37639 );
not ( n37641 , n6521 );
or ( n37642 , n37640 , n37641 );
nand ( n37643 , n35355 , n6491 );
nand ( n37644 , n37642 , n37643 );
buf ( n37645 , n37644 );
xor ( n37646 , n37637 , n37645 );
xor ( n37647 , n35384 , n35409 );
and ( n37648 , n37647 , n35427 );
and ( n37649 , n35384 , n35409 );
or ( n37650 , n37648 , n37649 );
buf ( n37651 , n37650 );
buf ( n37652 , n37651 );
xor ( n37653 , n37646 , n37652 );
buf ( n37654 , n37653 );
buf ( n37655 , n37654 );
xor ( n37656 , n37631 , n37655 );
buf ( n37657 , n37656 );
buf ( n37658 , n37657 );
xor ( n37659 , n37619 , n37658 );
buf ( n37660 , n37659 );
not ( n37661 , n37660 );
nor ( n37662 , n37661 , n454 );
nor ( n37663 , n37448 , n37662 );
not ( n37664 , n7443 );
nand ( n37665 , n7269 , n7442 );
not ( n37666 , n37665 );
or ( n37667 , n37664 , n37666 );
buf ( n37668 , n517 );
buf ( n37669 , n489 );
and ( n37670 , n37668 , n37669 );
buf ( n37671 , n37670 );
not ( n37672 , n6769 );
not ( n37673 , n7376 );
or ( n37674 , n37672 , n37673 );
not ( n37675 , n511 );
nand ( n37676 , n37675 , n493 );
not ( n37677 , n37676 );
not ( n37678 , n493 );
nand ( n37679 , n37678 , n511 );
not ( n37680 , n37679 );
or ( n37681 , n37677 , n37680 );
nand ( n37682 , n37681 , n2591 );
nand ( n37683 , n37674 , n37682 );
xor ( n37684 , n37671 , n37683 );
buf ( n37685 , n36184 );
not ( n37686 , n37685 );
buf ( n37687 , n2213 );
not ( n37688 , n37687 );
or ( n37689 , n37686 , n37688 );
buf ( n37690 , n2081 );
buf ( n37691 , n507 );
buf ( n37692 , n497 );
xor ( n37693 , n37691 , n37692 );
buf ( n37694 , n37693 );
buf ( n37695 , n37694 );
nand ( n37696 , n37690 , n37695 );
buf ( n37697 , n37696 );
buf ( n37698 , n37697 );
nand ( n37699 , n37689 , n37698 );
buf ( n37700 , n37699 );
xor ( n37701 , n37684 , n37700 );
buf ( n37702 , n37701 );
xor ( n37703 , n7104 , n7327 );
and ( n37704 , n37703 , n7334 );
and ( n37705 , n7104 , n7327 );
or ( n37706 , n37704 , n37705 );
buf ( n37707 , n37706 );
xor ( n37708 , n37702 , n37707 );
and ( n37709 , n513 , n491 );
not ( n37710 , n513 );
and ( n37711 , n37710 , n36583 );
nor ( n37712 , n37709 , n37711 );
not ( n37713 , n37712 );
not ( n37714 , n4519 );
or ( n37715 , n37713 , n37714 );
nand ( n37716 , n4512 , n36200 );
nand ( n37717 , n37715 , n37716 );
not ( n37718 , n36126 );
not ( n37719 , n7316 );
or ( n37720 , n37718 , n37719 );
buf ( n37721 , n4626 );
buf ( n37722 , n489 );
buf ( n37723 , n515 );
xor ( n37724 , n37722 , n37723 );
buf ( n37725 , n37724 );
buf ( n37726 , n37725 );
nand ( n37727 , n37721 , n37726 );
buf ( n37728 , n37727 );
nand ( n37729 , n37720 , n37728 );
and ( n37730 , n37717 , n37729 );
not ( n37731 , n37717 );
not ( n37732 , n37729 );
and ( n37733 , n37731 , n37732 );
nor ( n37734 , n37730 , n37733 );
and ( n37735 , n37734 , n7333 );
not ( n37736 , n37734 );
and ( n37737 , n37736 , n7334 );
nor ( n37738 , n37735 , n37737 );
buf ( n37739 , n37738 );
xor ( n37740 , n37708 , n37739 );
buf ( n37741 , n37740 );
xor ( n37742 , n7360 , n7419 );
and ( n37743 , n37742 , n36222 );
and ( n37744 , n7360 , n7419 );
or ( n37745 , n37743 , n37744 );
xor ( n37746 , n37741 , n37745 );
xor ( n37747 , n36165 , n36209 );
and ( n37748 , n37747 , n36215 );
and ( n37749 , n36165 , n36209 );
or ( n37750 , n37748 , n37749 );
xor ( n37751 , n36083 , n36093 );
and ( n37752 , n37751 , n36111 );
and ( n37753 , n36083 , n36093 );
or ( n37754 , n37752 , n37753 );
buf ( n37755 , n37754 );
buf ( n37756 , n37755 );
xor ( n37757 , n36176 , n36189 );
and ( n37758 , n37757 , n36207 );
and ( n37759 , n36176 , n36189 );
or ( n37760 , n37758 , n37759 );
buf ( n37761 , n37760 );
buf ( n37762 , n37761 );
xor ( n37763 , n37756 , n37762 );
not ( n37764 , n36104 );
not ( n37765 , n33373 );
or ( n37766 , n37764 , n37765 );
buf ( n37767 , n35574 );
buf ( n37768 , n509 );
buf ( n37769 , n495 );
xor ( n37770 , n37768 , n37769 );
buf ( n37771 , n37770 );
buf ( n37772 , n37771 );
nand ( n37773 , n37767 , n37772 );
buf ( n37774 , n37773 );
nand ( n37775 , n37766 , n37774 );
not ( n37776 , n37775 );
not ( n37777 , n37776 );
not ( n37778 , n1908 );
not ( n37779 , n1909 );
or ( n37780 , n37778 , n37779 );
nand ( n37781 , n37780 , n501 );
not ( n37782 , n37781 );
not ( n37783 , n37782 );
or ( n37784 , n37777 , n37783 );
nand ( n37785 , n37781 , n37775 );
nand ( n37786 , n37784 , n37785 );
not ( n37787 , n31011 );
buf ( n37788 , n505 );
buf ( n37789 , n499 );
xor ( n37790 , n37788 , n37789 );
buf ( n37791 , n37790 );
not ( n37792 , n37791 );
or ( n37793 , n37787 , n37792 );
nand ( n37794 , n2001 , n7285 );
nand ( n37795 , n37793 , n37794 );
not ( n37796 , n37795 );
and ( n37797 , n37786 , n37796 );
not ( n37798 , n37786 );
and ( n37799 , n37798 , n37795 );
nor ( n37800 , n37797 , n37799 );
buf ( n37801 , n37800 );
xor ( n37802 , n37763 , n37801 );
buf ( n37803 , n37802 );
xor ( n37804 , n37750 , n37803 );
xor ( n37805 , n36114 , n36139 );
and ( n37806 , n37805 , n36146 );
and ( n37807 , n36114 , n36139 );
or ( n37808 , n37806 , n37807 );
buf ( n37809 , n37808 );
xor ( n37810 , n37804 , n37809 );
xor ( n37811 , n37746 , n37810 );
not ( n37812 , n37811 );
xor ( n37813 , n36149 , n36155 );
and ( n37814 , n37813 , n36224 );
and ( n37815 , n36149 , n36155 );
or ( n37816 , n37814 , n37815 );
buf ( n37817 , n37816 );
not ( n37818 , n37817 );
nand ( n37819 , n37812 , n37818 );
buf ( n37820 , n37819 );
not ( n37821 , n37818 );
buf ( n37822 , n37811 );
nand ( n37823 , n37821 , n37822 );
nand ( n37824 , n37820 , n37823 );
and ( n37825 , n37824 , n2815 );
nand ( n37826 , n37667 , n37825 );
buf ( n37827 , n37067 );
buf ( n37828 , n4821 );
not ( n37829 , n37828 );
not ( n37830 , n491 );
not ( n37831 , n29742 );
or ( n37832 , n37830 , n37831 );
nand ( n37833 , n29749 , n33936 );
nand ( n37834 , n37832 , n37833 );
buf ( n37835 , n37834 );
not ( n37836 , n37835 );
or ( n37837 , n37829 , n37836 );
buf ( n37838 , n37139 );
buf ( n37839 , n34031 );
nand ( n37840 , n37838 , n37839 );
buf ( n37841 , n37840 );
buf ( n37842 , n37841 );
nand ( n37843 , n37837 , n37842 );
buf ( n37844 , n37843 );
buf ( n37845 , n37844 );
xor ( n37846 , n37827 , n37845 );
buf ( n37847 , n7455 );
not ( n37848 , n37847 );
buf ( n37849 , n489 );
not ( n37850 , n37849 );
buf ( n37851 , n971 );
not ( n37852 , n37851 );
or ( n37853 , n37850 , n37852 );
buf ( n37854 , n1204 );
buf ( n37855 , n7461 );
nand ( n37856 , n37854 , n37855 );
buf ( n37857 , n37856 );
buf ( n37858 , n37857 );
nand ( n37859 , n37853 , n37858 );
buf ( n37860 , n37859 );
buf ( n37861 , n37860 );
not ( n37862 , n37861 );
or ( n37863 , n37848 , n37862 );
buf ( n37864 , n37086 );
buf ( n37865 , n7474 );
nand ( n37866 , n37864 , n37865 );
buf ( n37867 , n37866 );
buf ( n37868 , n37867 );
nand ( n37869 , n37863 , n37868 );
buf ( n37870 , n37869 );
buf ( n37871 , n37870 );
xor ( n37872 , n37846 , n37871 );
buf ( n37873 , n37872 );
buf ( n37874 , n37873 );
xor ( n37875 , n37069 , n37092 );
and ( n37876 , n37875 , n37094 );
and ( n37877 , n37069 , n37092 );
or ( n37878 , n37876 , n37877 );
buf ( n37879 , n37878 );
buf ( n37880 , n37879 );
xor ( n37881 , n37874 , n37880 );
buf ( n37882 , n29829 );
not ( n37883 , n37882 );
buf ( n37884 , n497 );
not ( n37885 , n37884 );
buf ( n37886 , n7585 );
not ( n37887 , n37886 );
or ( n37888 , n37885 , n37887 );
buf ( n37889 , n706 );
buf ( n37890 , n5062 );
nand ( n37891 , n37889 , n37890 );
buf ( n37892 , n37891 );
buf ( n37893 , n37892 );
nand ( n37894 , n37888 , n37893 );
buf ( n37895 , n37894 );
buf ( n37896 , n37895 );
not ( n37897 , n37896 );
or ( n37898 , n37883 , n37897 );
buf ( n37899 , n37156 );
buf ( n37900 , n835 );
nand ( n37901 , n37899 , n37900 );
buf ( n37902 , n37901 );
buf ( n37903 , n37902 );
nand ( n37904 , n37898 , n37903 );
buf ( n37905 , n37904 );
buf ( n37906 , n1405 );
buf ( n37907 , n489 );
nand ( n37908 , n37906 , n37907 );
buf ( n37909 , n37908 );
buf ( n37910 , n37909 );
not ( n37911 , n37910 );
buf ( n37912 , n37911 );
xor ( n37913 , n37905 , n37912 );
not ( n37914 , n37175 );
not ( n37915 , n29575 );
and ( n37916 , n37914 , n37915 );
nand ( n37917 , n456 , n463 );
not ( n37918 , n456 );
nand ( n37919 , n37918 , n479 );
nand ( n37920 , n37917 , n37919 , n493 );
nand ( n37921 , n29505 , n7374 );
and ( n37922 , n37920 , n37921 );
not ( n37923 , n29522 );
nor ( n37924 , n37922 , n37923 );
nor ( n37925 , n37916 , n37924 );
not ( n37926 , n37925 );
xor ( n37927 , n37913 , n37926 );
buf ( n37928 , n37927 );
xor ( n37929 , n37881 , n37928 );
buf ( n37930 , n37929 );
buf ( n37931 , n37930 );
xor ( n37932 , n37120 , n37185 );
and ( n37933 , n37932 , n37192 );
and ( n37934 , n37120 , n37185 );
or ( n37935 , n37933 , n37934 );
buf ( n37936 , n37935 );
buf ( n37937 , n37936 );
xor ( n37938 , n37931 , n37937 );
xor ( n37939 , n37128 , n37132 );
and ( n37940 , n37939 , n37183 );
and ( n37941 , n37128 , n37132 );
or ( n37942 , n37940 , n37941 );
buf ( n37943 , n37942 );
buf ( n37944 , n37021 );
not ( n37945 , n37944 );
buf ( n37946 , n37047 );
not ( n37947 , n37946 );
or ( n37948 , n37945 , n37947 );
not ( n37949 , n29873 );
not ( n37950 , n37039 );
or ( n37951 , n37949 , n37950 );
nand ( n37952 , n37951 , n37018 );
not ( n37953 , n37046 );
or ( n37954 , n37952 , n37953 );
nand ( n37955 , n37954 , n37012 );
buf ( n37956 , n37955 );
nand ( n37957 , n37948 , n37956 );
buf ( n37958 , n37957 );
buf ( n37959 , n37958 );
xor ( n37960 , n37142 , n37164 );
and ( n37961 , n37960 , n37181 );
and ( n37962 , n37142 , n37164 );
or ( n37963 , n37961 , n37962 );
buf ( n37964 , n37963 );
buf ( n37965 , n37964 );
xor ( n37966 , n37959 , n37965 );
buf ( n37967 , n29669 );
not ( n37968 , n37967 );
buf ( n37969 , n29670 );
not ( n37970 , n37969 );
or ( n37971 , n37968 , n37970 );
buf ( n37972 , n501 );
nand ( n37973 , n37971 , n37972 );
buf ( n37974 , n37973 );
buf ( n37975 , n37974 );
buf ( n37976 , n29873 );
not ( n37977 , n37976 );
buf ( n37978 , n495 );
not ( n37979 , n37978 );
buf ( n37980 , n29510 );
not ( n37981 , n37980 );
or ( n37982 , n37979 , n37981 );
buf ( n37983 , n29511 );
buf ( n37984 , n29716 );
nand ( n37985 , n37983 , n37984 );
buf ( n37986 , n37985 );
buf ( n37987 , n37986 );
nand ( n37988 , n37982 , n37987 );
buf ( n37989 , n37988 );
buf ( n37990 , n37989 );
not ( n37991 , n37990 );
or ( n37992 , n37977 , n37991 );
buf ( n37993 , n37039 );
buf ( n37994 , n30072 );
nand ( n37995 , n37993 , n37994 );
buf ( n37996 , n37995 );
buf ( n37997 , n37996 );
nand ( n37998 , n37992 , n37997 );
buf ( n37999 , n37998 );
buf ( n38000 , n37999 );
xor ( n38001 , n37975 , n38000 );
buf ( n38002 , n29583 );
not ( n38003 , n38002 );
buf ( n38004 , n499 );
not ( n38005 , n38004 );
and ( n38006 , n456 , n457 );
not ( n38007 , n456 );
and ( n38008 , n38007 , n473 );
nor ( n38009 , n38006 , n38008 );
buf ( n38010 , n38009 );
not ( n38011 , n38010 );
or ( n38012 , n38005 , n38011 );
not ( n38013 , n36649 );
buf ( n38014 , n38013 );
buf ( n38015 , n29596 );
nand ( n38016 , n38014 , n38015 );
buf ( n38017 , n38016 );
buf ( n38018 , n38017 );
nand ( n38019 , n38012 , n38018 );
buf ( n38020 , n38019 );
buf ( n38021 , n38020 );
not ( n38022 , n38021 );
or ( n38023 , n38003 , n38022 );
buf ( n38024 , n37008 );
buf ( n38025 , n29624 );
nand ( n38026 , n38024 , n38025 );
buf ( n38027 , n38026 );
buf ( n38028 , n38027 );
nand ( n38029 , n38023 , n38028 );
buf ( n38030 , n38029 );
buf ( n38031 , n38030 );
xor ( n38032 , n38001 , n38031 );
buf ( n38033 , n38032 );
buf ( n38034 , n38033 );
xor ( n38035 , n37966 , n38034 );
buf ( n38036 , n38035 );
buf ( n38037 , n38036 );
xor ( n38038 , n37943 , n38037 );
xor ( n38039 , n37058 , n37097 );
and ( n38040 , n38039 , n37104 );
and ( n38041 , n37058 , n37097 );
or ( n38042 , n38040 , n38041 );
buf ( n38043 , n38042 );
buf ( n38044 , n38043 );
xor ( n38045 , n38038 , n38044 );
buf ( n38046 , n38045 );
buf ( n38047 , n38046 );
xor ( n38048 , n37938 , n38047 );
buf ( n38049 , n38048 );
xor ( n38050 , n37107 , n37113 );
and ( n38051 , n38050 , n37195 );
and ( n38052 , n37107 , n37113 );
or ( n38053 , n38051 , n38052 );
buf ( n38054 , n38053 );
nand ( n38055 , n38049 , n38054 );
buf ( n38056 , n38055 );
not ( n38057 , n38049 );
not ( n38058 , n38054 );
nand ( n38059 , n38057 , n38058 );
nand ( n38060 , n38056 , n38059 );
nand ( n38061 , n455 , n38060 );
not ( n38062 , n38061 );
buf ( n38063 , n37203 );
nand ( n38064 , n36995 , n38063 );
nand ( n38065 , n38064 , n37205 );
nand ( n38066 , n38062 , n38065 );
nand ( n38067 , n37826 , n38066 );
not ( n38068 , n38064 );
nand ( n38069 , n37205 , n455 );
nor ( n38070 , n38060 , n38069 );
not ( n38071 , n38070 );
or ( n38072 , n38068 , n38071 );
not ( n38073 , n7443 );
nor ( n38074 , n37824 , n38073 , n455 );
nand ( n38075 , n37665 , n38074 );
nand ( n38076 , n38072 , n38075 );
or ( n38077 , n38067 , n38076 );
nand ( n38078 , n38077 , n454 );
nand ( n38079 , n37663 , n38078 );
not ( n38080 , n38079 );
not ( n38081 , n38080 );
and ( n38082 , n36957 , n38059 , n37203 );
not ( n38083 , n38082 );
not ( n38084 , n36984 );
or ( n38085 , n38083 , n38084 );
nand ( n38086 , n36992 , n37203 );
nand ( n38087 , n36989 , n38059 );
nor ( n38088 , n38086 , n38087 );
nand ( n38089 , n38057 , n38058 );
not ( n38090 , n38089 );
not ( n38091 , n37204 );
or ( n38092 , n38090 , n38091 );
nand ( n38093 , n38092 , n38056 );
nor ( n38094 , n38088 , n38093 );
nand ( n38095 , n38085 , n38094 );
xor ( n38096 , n37874 , n37880 );
and ( n38097 , n38096 , n37928 );
and ( n38098 , n37874 , n37880 );
or ( n38099 , n38097 , n38098 );
buf ( n38100 , n38099 );
xor ( n38101 , n37943 , n38037 );
and ( n38102 , n38101 , n38044 );
and ( n38103 , n37943 , n38037 );
or ( n38104 , n38102 , n38103 );
buf ( n38105 , n38104 );
xor ( n38106 , n38100 , n38105 );
and ( n38107 , n38020 , n29624 );
and ( n38108 , n29581 , n499 );
nor ( n38109 , n38107 , n38108 );
not ( n38110 , n37926 );
not ( n38111 , n37912 );
or ( n38112 , n38110 , n38111 );
not ( n38113 , n37909 );
not ( n38114 , n37925 );
or ( n38115 , n38113 , n38114 );
nand ( n38116 , n38115 , n37905 );
nand ( n38117 , n38112 , n38116 );
xor ( n38118 , n38109 , n38117 );
xor ( n38119 , n37975 , n38000 );
and ( n38120 , n38119 , n38031 );
and ( n38121 , n37975 , n38000 );
or ( n38122 , n38120 , n38121 );
buf ( n38123 , n38122 );
xor ( n38124 , n38118 , n38123 );
buf ( n38125 , n38124 );
xor ( n38126 , n37959 , n37965 );
and ( n38127 , n38126 , n38034 );
and ( n38128 , n37959 , n37965 );
or ( n38129 , n38127 , n38128 );
buf ( n38130 , n38129 );
buf ( n38131 , n38130 );
xor ( n38132 , n38125 , n38131 );
xor ( n38133 , n37827 , n37845 );
and ( n38134 , n38133 , n37871 );
and ( n38135 , n37827 , n37845 );
or ( n38136 , n38134 , n38135 );
buf ( n38137 , n38136 );
buf ( n38138 , n38137 );
buf ( n38139 , n29493 );
buf ( n38140 , n489 );
and ( n38141 , n38139 , n38140 );
buf ( n38142 , n38141 );
buf ( n38143 , n38142 );
buf ( n38144 , n30072 );
not ( n38145 , n38144 );
buf ( n38146 , n37989 );
not ( n38147 , n38146 );
or ( n38148 , n38145 , n38147 );
buf ( n38149 , n495 );
not ( n38150 , n38149 );
buf ( n38151 , n7573 );
not ( n38152 , n38151 );
or ( n38153 , n38150 , n38152 );
buf ( n38154 , n7567 );
buf ( n38155 , n29716 );
nand ( n38156 , n38154 , n38155 );
buf ( n38157 , n38156 );
buf ( n38158 , n38157 );
nand ( n38159 , n38153 , n38158 );
buf ( n38160 , n38159 );
buf ( n38161 , n38160 );
buf ( n38162 , n29873 );
nand ( n38163 , n38161 , n38162 );
buf ( n38164 , n38163 );
buf ( n38165 , n38164 );
nand ( n38166 , n38148 , n38165 );
buf ( n38167 , n38166 );
buf ( n38168 , n38167 );
xor ( n38169 , n38143 , n38168 );
buf ( n38170 , n37071 );
not ( n38171 , n38170 );
buf ( n38172 , n37860 );
not ( n38173 , n38172 );
or ( n38174 , n38171 , n38173 );
buf ( n38175 , n489 );
buf ( n38176 , n29613 );
xor ( n38177 , n38175 , n38176 );
buf ( n38178 , n38177 );
buf ( n38179 , n38178 );
buf ( n38180 , n7455 );
nand ( n38181 , n38179 , n38180 );
buf ( n38182 , n38181 );
buf ( n38183 , n38182 );
nand ( n38184 , n38174 , n38183 );
buf ( n38185 , n38184 );
buf ( n38186 , n38185 );
xor ( n38187 , n38169 , n38186 );
buf ( n38188 , n38187 );
buf ( n38189 , n38188 );
xor ( n38190 , n38138 , n38189 );
not ( n38191 , n29522 );
not ( n38192 , n36611 );
not ( n38193 , n29537 );
or ( n38194 , n38192 , n38193 );
nand ( n38195 , n37037 , n493 );
nand ( n38196 , n38194 , n38195 );
not ( n38197 , n38196 );
or ( n38198 , n38191 , n38197 );
not ( n38199 , n37920 );
not ( n38200 , n37921 );
or ( n38201 , n38199 , n38200 );
nand ( n38202 , n38201 , n29576 );
nand ( n38203 , n38198 , n38202 );
not ( n38204 , n36694 );
not ( n38205 , n855 );
not ( n38206 , n491 );
or ( n38207 , n38205 , n38206 );
not ( n38208 , n29654 );
nand ( n38209 , n38208 , n33936 );
nand ( n38210 , n38207 , n38209 );
not ( n38211 , n38210 );
or ( n38212 , n38204 , n38211 );
nand ( n38213 , n37834 , n34031 );
nand ( n38214 , n38212 , n38213 );
xor ( n38215 , n38203 , n38214 );
not ( n38216 , n37895 );
not ( n38217 , n835 );
or ( n38218 , n38216 , n38217 );
buf ( n38219 , n497 );
not ( n38220 , n38219 );
buf ( n38221 , n29498 );
not ( n38222 , n38221 );
or ( n38223 , n38220 , n38222 );
and ( n38224 , n456 , n458 );
not ( n38225 , n456 );
and ( n38226 , n38225 , n474 );
nor ( n38227 , n38224 , n38226 );
not ( n38228 , n38227 );
buf ( n38229 , n38228 );
buf ( n38230 , n706 );
nand ( n38231 , n38229 , n38230 );
buf ( n38232 , n38231 );
buf ( n38233 , n38232 );
nand ( n38234 , n38223 , n38233 );
buf ( n38235 , n38234 );
buf ( n38236 , n38235 );
buf ( n38237 , n29829 );
nand ( n38238 , n38236 , n38237 );
buf ( n38239 , n38238 );
nand ( n38240 , n38218 , n38239 );
and ( n38241 , n38215 , n38240 );
not ( n38242 , n38215 );
not ( n38243 , n38240 );
and ( n38244 , n38242 , n38243 );
nor ( n38245 , n38241 , n38244 );
buf ( n38246 , n38245 );
xor ( n38247 , n38190 , n38246 );
buf ( n38248 , n38247 );
buf ( n38249 , n38248 );
xor ( n38250 , n38132 , n38249 );
buf ( n38251 , n38250 );
xor ( n38252 , n38106 , n38251 );
not ( n38253 , n38252 );
xor ( n38254 , n37931 , n37937 );
and ( n38255 , n38254 , n38047 );
and ( n38256 , n37931 , n37937 );
or ( n38257 , n38255 , n38256 );
buf ( n38258 , n38257 );
not ( n38259 , n38258 );
nand ( n38260 , n38253 , n38259 );
buf ( n38261 , n38260 );
nand ( n38262 , n38252 , n38258 );
buf ( n38263 , n38262 );
and ( n38264 , n38261 , n38263 );
and ( n38265 , n38095 , n38264 );
not ( n38266 , n38095 );
not ( n38267 , n38264 );
and ( n38268 , n38266 , n38267 );
nor ( n38269 , n38265 , n38268 );
nand ( n38270 , n38269 , n455 );
not ( n38271 , n38270 );
nand ( n38272 , n7239 , n7260 );
not ( n38273 , n38272 );
nor ( n38274 , n7194 , n7219 );
and ( n38275 , n37820 , n7442 , n38274 );
not ( n38276 , n38275 );
or ( n38277 , n38273 , n38276 );
not ( n38278 , n7266 );
not ( n38279 , n7265 );
or ( n38280 , n38278 , n38279 );
nor ( n38281 , n36002 , n35818 );
nor ( n38282 , n38281 , n7441 );
nand ( n38283 , n38280 , n38282 );
not ( n38284 , n37819 );
nor ( n38285 , n38283 , n38284 );
not ( n38286 , n38073 );
not ( n38287 , n37819 );
or ( n38288 , n38286 , n38287 );
nand ( n38289 , n38288 , n37823 );
nor ( n38290 , n38285 , n38289 );
nand ( n38291 , n38277 , n38290 );
xor ( n38292 , n37741 , n37745 );
and ( n38293 , n38292 , n37810 );
and ( n38294 , n37741 , n37745 );
or ( n38295 , n38293 , n38294 );
xor ( n38296 , n37702 , n37707 );
and ( n38297 , n38296 , n37739 );
and ( n38298 , n37702 , n37707 );
or ( n38299 , n38297 , n38298 );
buf ( n38300 , n38299 );
xor ( n38301 , n37750 , n37803 );
and ( n38302 , n38301 , n37809 );
and ( n38303 , n37750 , n37803 );
or ( n38304 , n38302 , n38303 );
xor ( n38305 , n38300 , n38304 );
not ( n38306 , n37791 );
not ( n38307 , n2001 );
or ( n38308 , n38306 , n38307 );
buf ( n38309 , n30884 );
buf ( n38310 , n499 );
nand ( n38311 , n38309 , n38310 );
buf ( n38312 , n38311 );
nand ( n38313 , n38308 , n38312 );
not ( n38314 , n38313 );
buf ( n38315 , n38314 );
xor ( n38316 , n37671 , n37683 );
and ( n38317 , n38316 , n37700 );
and ( n38318 , n37671 , n37683 );
or ( n38319 , n38317 , n38318 );
buf ( n38320 , n38319 );
xor ( n38321 , n38315 , n38320 );
or ( n38322 , n37795 , n37775 );
nand ( n38323 , n38322 , n37781 );
nand ( n38324 , n37795 , n37775 );
nand ( n38325 , n38323 , n38324 );
buf ( n38326 , n38325 );
xor ( n38327 , n38321 , n38326 );
buf ( n38328 , n38327 );
buf ( n38329 , n38328 );
xor ( n38330 , n37756 , n37762 );
and ( n38331 , n38330 , n37801 );
and ( n38332 , n37756 , n37762 );
or ( n38333 , n38331 , n38332 );
buf ( n38334 , n38333 );
buf ( n38335 , n38334 );
xor ( n38336 , n38329 , n38335 );
not ( n38337 , n7333 );
not ( n38338 , n37729 );
or ( n38339 , n38337 , n38338 );
not ( n38340 , n7334 );
not ( n38341 , n37732 );
or ( n38342 , n38340 , n38341 );
nand ( n38343 , n38342 , n37717 );
nand ( n38344 , n38339 , n38343 );
buf ( n38345 , n38344 );
not ( n38346 , n37694 );
not ( n38347 , n6669 );
or ( n38348 , n38346 , n38347 );
xor ( n38349 , n506 , n497 );
nand ( n38350 , n2081 , n38349 );
nand ( n38351 , n38348 , n38350 );
buf ( n38352 , n37712 );
not ( n38353 , n38352 );
buf ( n38354 , n4512 );
not ( n38355 , n38354 );
or ( n38356 , n38353 , n38355 );
buf ( n38357 , n4286 );
buf ( n38358 , n512 );
buf ( n38359 , n491 );
xor ( n38360 , n38358 , n38359 );
buf ( n38361 , n38360 );
buf ( n38362 , n38361 );
nand ( n38363 , n38357 , n38362 );
buf ( n38364 , n38363 );
buf ( n38365 , n38364 );
nand ( n38366 , n38356 , n38365 );
buf ( n38367 , n38366 );
xor ( n38368 , n38351 , n38367 );
nand ( n38369 , n37679 , n37676 );
not ( n38370 , n38369 );
not ( n38371 , n2668 );
or ( n38372 , n38370 , n38371 );
buf ( n38373 , n2591 );
buf ( n38374 , n510 );
buf ( n38375 , n493 );
xor ( n38376 , n38374 , n38375 );
buf ( n38377 , n38376 );
buf ( n38378 , n38377 );
nand ( n38379 , n38373 , n38378 );
buf ( n38380 , n38379 );
nand ( n38381 , n38372 , n38380 );
xor ( n38382 , n38368 , n38381 );
buf ( n38383 , n38382 );
xor ( n38384 , n38345 , n38383 );
buf ( n38385 , n516 );
buf ( n38386 , n489 );
and ( n38387 , n38385 , n38386 );
buf ( n38388 , n38387 );
buf ( n38389 , n38388 );
buf ( n38390 , n37771 );
not ( n38391 , n38390 );
buf ( n38392 , n35567 );
not ( n38393 , n38392 );
or ( n38394 , n38391 , n38393 );
buf ( n38395 , n508 );
buf ( n38396 , n495 );
xor ( n38397 , n38395 , n38396 );
buf ( n38398 , n38397 );
buf ( n38399 , n38398 );
buf ( n38400 , n35574 );
nand ( n38401 , n38399 , n38400 );
buf ( n38402 , n38401 );
buf ( n38403 , n38402 );
nand ( n38404 , n38394 , n38403 );
buf ( n38405 , n38404 );
buf ( n38406 , n38405 );
xor ( n38407 , n38389 , n38406 );
buf ( n38408 , n37725 );
not ( n38409 , n38408 );
not ( n38410 , n7315 );
buf ( n38411 , n38410 );
not ( n38412 , n38411 );
or ( n38413 , n38409 , n38412 );
buf ( n38414 , n35832 );
buf ( n38415 , n489 );
buf ( n38416 , n514 );
xor ( n38417 , n38415 , n38416 );
buf ( n38418 , n38417 );
buf ( n38419 , n38418 );
nand ( n38420 , n38414 , n38419 );
buf ( n38421 , n38420 );
buf ( n38422 , n38421 );
nand ( n38423 , n38413 , n38422 );
buf ( n38424 , n38423 );
buf ( n38425 , n38424 );
xor ( n38426 , n38407 , n38425 );
buf ( n38427 , n38426 );
buf ( n38428 , n38427 );
xor ( n38429 , n38384 , n38428 );
buf ( n38430 , n38429 );
buf ( n38431 , n38430 );
xor ( n38432 , n38336 , n38431 );
buf ( n38433 , n38432 );
xor ( n38434 , n38305 , n38433 );
nand ( n38435 , n38295 , n38434 );
not ( n38436 , n38435 );
nor ( n38437 , n38434 , n38295 );
nor ( n38438 , n38436 , n38437 );
and ( n38439 , n38291 , n38438 );
not ( n38440 , n38291 );
not ( n38441 , n38438 );
and ( n38442 , n38440 , n38441 );
nor ( n38443 , n38439 , n38442 );
nand ( n38444 , n38443 , n2815 );
not ( n38445 , n38444 );
or ( n38446 , n38271 , n38445 );
nand ( n38447 , n38446 , n454 );
xor ( n38448 , n37574 , n37591 );
and ( n38449 , n38448 , n37609 );
and ( n38450 , n37574 , n37591 );
or ( n38451 , n38449 , n38450 );
buf ( n38452 , n38451 );
buf ( n38453 , n38452 );
buf ( n38454 , n3045 );
buf ( n38455 , n37514 );
or ( n38456 , n38454 , n38455 );
buf ( n38457 , n2918 );
buf ( n38458 , n31868 );
buf ( n38459 , n521 );
and ( n38460 , n38458 , n38459 );
buf ( n38461 , n35343 );
buf ( n38462 , n549 );
and ( n38463 , n38461 , n38462 );
nor ( n38464 , n38460 , n38463 );
buf ( n38465 , n38464 );
buf ( n38466 , n38465 );
or ( n38467 , n38457 , n38466 );
nand ( n38468 , n38456 , n38467 );
buf ( n38469 , n38468 );
buf ( n38470 , n38469 );
buf ( n38471 , n5582 );
buf ( n38472 , n37586 );
or ( n38473 , n38471 , n38472 );
buf ( n38474 , n33118 );
buf ( n38475 , n541 );
buf ( n38476 , n2969 );
and ( n38477 , n38475 , n38476 );
not ( n38478 , n38475 );
buf ( n38479 , n529 );
and ( n38480 , n38478 , n38479 );
nor ( n38481 , n38477 , n38480 );
buf ( n38482 , n38481 );
buf ( n38483 , n38482 );
or ( n38484 , n38474 , n38483 );
nand ( n38485 , n38473 , n38484 );
buf ( n38486 , n38485 );
buf ( n38487 , n38486 );
xor ( n38488 , n38470 , n38487 );
buf ( n38489 , n3020 );
buf ( n38490 , n37485 );
or ( n38491 , n38489 , n38490 );
buf ( n38492 , n31978 );
buf ( n38493 , n547 );
buf ( n38494 , n523 );
xnor ( n38495 , n38493 , n38494 );
buf ( n38496 , n38495 );
buf ( n38497 , n38496 );
or ( n38498 , n38492 , n38497 );
nand ( n38499 , n38491 , n38498 );
buf ( n38500 , n38499 );
buf ( n38501 , n38500 );
xor ( n38502 , n38488 , n38501 );
buf ( n38503 , n38502 );
buf ( n38504 , n38503 );
xor ( n38505 , n38453 , n38504 );
xor ( n38506 , n37637 , n37645 );
and ( n38507 , n38506 , n37652 );
and ( n38508 , n37637 , n37645 );
or ( n38509 , n38507 , n38508 );
buf ( n38510 , n38509 );
buf ( n38511 , n38510 );
xor ( n38512 , n38505 , n38511 );
buf ( n38513 , n38512 );
buf ( n38514 , n38513 );
xor ( n38515 , n37625 , n37630 );
and ( n38516 , n38515 , n37655 );
and ( n38517 , n37625 , n37630 );
or ( n38518 , n38516 , n38517 );
buf ( n38519 , n38518 );
buf ( n38520 , n38519 );
xor ( n38521 , n38514 , n38520 );
and ( n38522 , n37597 , n37606 );
buf ( n38523 , n38522 );
buf ( n38524 , n38523 );
buf ( n38525 , n37557 );
buf ( n38526 , n37569 );
or ( n38527 , n38525 , n38526 );
buf ( n38528 , n6010 );
buf ( n38529 , n6001 );
buf ( n38530 , n531 );
and ( n38531 , n38529 , n38530 );
buf ( n38532 , n31840 );
buf ( n38533 , n539 );
and ( n38534 , n38532 , n38533 );
nor ( n38535 , n38531 , n38534 );
buf ( n38536 , n38535 );
buf ( n38537 , n38536 );
or ( n38538 , n38528 , n38537 );
nand ( n38539 , n38527 , n38538 );
buf ( n38540 , n38539 );
buf ( n38541 , n38540 );
xor ( n38542 , n38524 , n38541 );
or ( n38543 , n37495 , n37499 );
nand ( n38544 , n37491 , n37493 );
nand ( n38545 , n38543 , n38544 );
buf ( n38546 , n38545 );
xor ( n38547 , n38542 , n38546 );
buf ( n38548 , n38547 );
not ( n38549 , n37611 );
nand ( n38550 , n37555 , n37502 );
not ( n38551 , n38550 );
or ( n38552 , n38549 , n38551 );
nand ( n38553 , n37554 , n37501 );
nand ( n38554 , n38552 , n38553 );
xor ( n38555 , n38548 , n38554 );
buf ( n38556 , n6559 );
buf ( n38557 , n37531 );
or ( n38558 , n38556 , n38557 );
buf ( n38559 , n6337 );
buf ( n38560 , n537 );
buf ( n38561 , n31874 );
and ( n38562 , n38560 , n38561 );
not ( n38563 , n38560 );
buf ( n38564 , n533 );
and ( n38565 , n38563 , n38564 );
nor ( n38566 , n38562 , n38565 );
buf ( n38567 , n38566 );
buf ( n38568 , n38567 );
or ( n38569 , n38559 , n38568 );
nand ( n38570 , n38558 , n38569 );
buf ( n38571 , n38570 );
buf ( n38572 , n38571 );
buf ( n38573 , n535 );
buf ( n38574 , n537 );
and ( n38575 , n38573 , n38574 );
buf ( n38576 , n38575 );
buf ( n38577 , n38576 );
xor ( n38578 , n38572 , n38577 );
buf ( n38579 , n545 );
buf ( n38580 , n525 );
and ( n38581 , n38579 , n38580 );
not ( n38582 , n38579 );
buf ( n38583 , n34557 );
and ( n38584 , n38582 , n38583 );
nor ( n38585 , n38581 , n38584 );
buf ( n38586 , n38585 );
buf ( n38587 , n38586 );
not ( n38588 , n38587 );
buf ( n38589 , n3063 );
not ( n38590 , n38589 );
or ( n38591 , n38588 , n38590 );
buf ( n38592 , n3069 );
buf ( n38593 , n37549 );
or ( n38594 , n38592 , n38593 );
nand ( n38595 , n38591 , n38594 );
buf ( n38596 , n38595 );
buf ( n38597 , n38596 );
xor ( n38598 , n38578 , n38597 );
buf ( n38599 , n38598 );
buf ( n38600 , n38599 );
buf ( n38601 , n2848 );
not ( n38602 , n38601 );
buf ( n38603 , n5636 );
buf ( n38604 , n37469 );
or ( n38605 , n38603 , n38604 );
buf ( n38606 , n35070 );
buf ( n38607 , n32981 );
buf ( n38608 , n527 );
and ( n38609 , n38607 , n38608 );
buf ( n38610 , n33009 );
buf ( n38611 , n543 );
and ( n38612 , n38610 , n38611 );
nor ( n38613 , n38609 , n38612 );
buf ( n38614 , n38613 );
buf ( n38615 , n38614 );
or ( n38616 , n38606 , n38615 );
nand ( n38617 , n38605 , n38616 );
buf ( n38618 , n38617 );
buf ( n38619 , n38618 );
not ( n38620 , n38619 );
or ( n38621 , n38602 , n38620 );
buf ( n38622 , n38618 );
buf ( n38623 , n2848 );
or ( n38624 , n38622 , n38623 );
buf ( n38625 , n38624 );
buf ( n38626 , n38625 );
nand ( n38627 , n38621 , n38626 );
buf ( n38628 , n38627 );
buf ( n38629 , n38628 );
xor ( n38630 , n38600 , n38629 );
xor ( n38631 , n37519 , n37534 );
and ( n38632 , n38631 , n37552 );
and ( n38633 , n37519 , n37534 );
or ( n38634 , n38632 , n38633 );
buf ( n38635 , n38634 );
buf ( n38636 , n38635 );
xor ( n38637 , n38630 , n38636 );
buf ( n38638 , n38637 );
xor ( n38639 , n38555 , n38638 );
buf ( n38640 , n38639 );
xor ( n38641 , n38521 , n38640 );
buf ( n38642 , n38641 );
buf ( n38643 , n38642 );
buf ( n38644 , n3360 );
and ( n38645 , n38643 , n38644 );
buf ( n38646 , n38645 );
xor ( n38647 , n37457 , n37618 );
and ( n38648 , n38647 , n37658 );
and ( n38649 , n37457 , n37618 );
or ( n38650 , n38648 , n38649 );
buf ( n38651 , n38650 );
and ( n38652 , n38651 , n3138 );
nor ( n38653 , n38646 , n38652 );
nand ( n38654 , n38447 , n38653 );
not ( n38655 , n38654 );
not ( n38656 , n38655 );
nand ( n38657 , n38081 , n38656 );
buf ( n38658 , n38625 );
buf ( n38659 , n6559 );
buf ( n38660 , n38567 );
or ( n38661 , n38659 , n38660 );
buf ( n38662 , n6337 );
buf ( n38663 , n6541 );
buf ( n38664 , n532 );
and ( n38665 , n38663 , n38664 );
buf ( n38666 , n31908 );
buf ( n38667 , n537 );
and ( n38668 , n38666 , n38667 );
nor ( n38669 , n38665 , n38668 );
buf ( n38670 , n38669 );
buf ( n38671 , n38670 );
or ( n38672 , n38662 , n38671 );
nand ( n38673 , n38661 , n38672 );
buf ( n38674 , n38673 );
buf ( n38675 , n38674 );
xor ( n38676 , n38658 , n38675 );
xor ( n38677 , n38572 , n38577 );
and ( n38678 , n38677 , n38597 );
and ( n38679 , n38572 , n38577 );
or ( n38680 , n38678 , n38679 );
buf ( n38681 , n38680 );
buf ( n38682 , n38681 );
and ( n38683 , n38676 , n38682 );
and ( n38684 , n38658 , n38675 );
or ( n38685 , n38683 , n38684 );
buf ( n38686 , n38685 );
buf ( n38687 , n38686 );
buf ( n38688 , n5582 );
buf ( n38689 , n541 );
buf ( n38690 , n32183 );
and ( n38691 , n38689 , n38690 );
not ( n38692 , n38689 );
buf ( n38693 , n528 );
and ( n38694 , n38692 , n38693 );
nor ( n38695 , n38691 , n38694 );
buf ( n38696 , n38695 );
buf ( n38697 , n38696 );
or ( n38698 , n38688 , n38697 );
buf ( n38699 , n33118 );
buf ( n38700 , n541 );
buf ( n38701 , n33009 );
and ( n38702 , n38700 , n38701 );
not ( n38703 , n38700 );
buf ( n38704 , n527 );
and ( n38705 , n38703 , n38704 );
nor ( n38706 , n38702 , n38705 );
buf ( n38707 , n38706 );
buf ( n38708 , n38707 );
or ( n38709 , n38699 , n38708 );
nand ( n38710 , n38698 , n38709 );
buf ( n38711 , n38710 );
buf ( n38712 , n38711 );
buf ( n38713 , n533 );
buf ( n38714 , n537 );
and ( n38715 , n38713 , n38714 );
buf ( n38716 , n38715 );
buf ( n38717 , n38716 );
xor ( n38718 , n38712 , n38717 );
buf ( n38719 , n3069 );
buf ( n38720 , n32053 );
buf ( n38721 , n524 );
and ( n38722 , n38720 , n38721 );
buf ( n38723 , n34779 );
buf ( n38724 , n545 );
and ( n38725 , n38723 , n38724 );
nor ( n38726 , n38722 , n38725 );
buf ( n38727 , n38726 );
buf ( n38728 , n38727 );
or ( n38729 , n38719 , n38728 );
buf ( n38730 , n3087 );
buf ( n38731 , n523 );
buf ( n38732 , n32053 );
and ( n38733 , n38731 , n38732 );
not ( n38734 , n38731 );
buf ( n38735 , n545 );
and ( n38736 , n38734 , n38735 );
nor ( n38737 , n38733 , n38736 );
buf ( n38738 , n38737 );
buf ( n38739 , n38738 );
or ( n38740 , n38730 , n38739 );
nand ( n38741 , n38729 , n38740 );
buf ( n38742 , n38741 );
buf ( n38743 , n38742 );
xor ( n38744 , n38718 , n38743 );
buf ( n38745 , n38744 );
buf ( n38746 , n38745 );
xor ( n38747 , n38687 , n38746 );
buf ( n38748 , n37557 );
buf ( n38749 , n6001 );
buf ( n38750 , n530 );
and ( n38751 , n38749 , n38750 );
buf ( n38752 , n31853 );
buf ( n38753 , n539 );
and ( n38754 , n38752 , n38753 );
nor ( n38755 , n38751 , n38754 );
buf ( n38756 , n38755 );
buf ( n38757 , n38756 );
or ( n38758 , n38748 , n38757 );
buf ( n38759 , n6010 );
buf ( n38760 , n6001 );
buf ( n38761 , n529 );
and ( n38762 , n38760 , n38761 );
buf ( n38763 , n2969 );
buf ( n38764 , n539 );
and ( n38765 , n38763 , n38764 );
nor ( n38766 , n38762 , n38765 );
buf ( n38767 , n38766 );
buf ( n38768 , n38767 );
or ( n38769 , n38759 , n38768 );
nand ( n38770 , n38758 , n38769 );
buf ( n38771 , n38770 );
buf ( n38772 , n38771 );
nand ( n38773 , n35397 , n6337 );
buf ( n38774 , n38773 );
buf ( n38775 , n38670 );
or ( n38776 , n38774 , n38775 );
buf ( n38777 , n6337 );
buf ( n38778 , n6541 );
buf ( n38779 , n531 );
and ( n38780 , n38778 , n38779 );
buf ( n38781 , n31840 );
buf ( n38782 , n537 );
and ( n38783 , n38781 , n38782 );
nor ( n38784 , n38780 , n38783 );
buf ( n38785 , n38784 );
buf ( n38786 , n38785 );
or ( n38787 , n38777 , n38786 );
nand ( n38788 , n38776 , n38787 );
buf ( n38789 , n38788 );
buf ( n38790 , n38789 );
xor ( n38791 , n38772 , n38790 );
not ( n38792 , n38586 );
not ( n38793 , n6305 );
or ( n38794 , n38792 , n38793 );
or ( n38795 , n38727 , n3087 );
nand ( n38796 , n38794 , n38795 );
buf ( n38797 , n38796 );
buf ( n38798 , n6015 );
buf ( n38799 , n38536 );
or ( n38800 , n38798 , n38799 );
buf ( n38801 , n6010 );
buf ( n38802 , n38756 );
or ( n38803 , n38801 , n38802 );
nand ( n38804 , n38800 , n38803 );
buf ( n38805 , n38804 );
buf ( n38806 , n38805 );
and ( n38807 , n38797 , n38806 );
buf ( n38808 , n38807 );
buf ( n38809 , n38808 );
xor ( n38810 , n38791 , n38809 );
buf ( n38811 , n38810 );
buf ( n38812 , n38811 );
xor ( n38813 , n38747 , n38812 );
buf ( n38814 , n38813 );
buf ( n38815 , n38814 );
buf ( n38816 , n3045 );
buf ( n38817 , n38465 );
or ( n38818 , n38816 , n38817 );
buf ( n38819 , n2918 );
buf ( n38820 , n31868 );
or ( n38821 , n38819 , n38820 );
nand ( n38822 , n38818 , n38821 );
buf ( n38823 , n38822 );
buf ( n38824 , n38823 );
not ( n38825 , n38824 );
buf ( n38826 , n3020 );
buf ( n38827 , n38496 );
or ( n38828 , n38826 , n38827 );
buf ( n38829 , n31978 );
buf ( n38830 , n547 );
buf ( n38831 , n35199 );
and ( n38832 , n38830 , n38831 );
not ( n38833 , n38830 );
buf ( n38834 , n522 );
and ( n38835 , n38833 , n38834 );
nor ( n38836 , n38832 , n38835 );
buf ( n38837 , n38836 );
buf ( n38838 , n38837 );
or ( n38839 , n38829 , n38838 );
nand ( n38840 , n38828 , n38839 );
buf ( n38841 , n38840 );
buf ( n38842 , n38841 );
not ( n38843 , n38842 );
or ( n38844 , n38825 , n38843 );
buf ( n38845 , n38841 );
buf ( n38846 , n38823 );
or ( n38847 , n38845 , n38846 );
buf ( n38848 , n38847 );
buf ( n38849 , n38848 );
nand ( n38850 , n38844 , n38849 );
buf ( n38851 , n38850 );
buf ( n38852 , n38851 );
xor ( n38853 , n38797 , n38806 );
buf ( n38854 , n38853 );
buf ( n38855 , n38854 );
xor ( n38856 , n38852 , n38855 );
xor ( n38857 , n38470 , n38487 );
and ( n38858 , n38857 , n38501 );
and ( n38859 , n38470 , n38487 );
or ( n38860 , n38858 , n38859 );
buf ( n38861 , n38860 );
buf ( n38862 , n38861 );
xor ( n38863 , n38856 , n38862 );
buf ( n38864 , n38863 );
buf ( n38865 , n38864 );
xor ( n38866 , n38600 , n38629 );
and ( n38867 , n38866 , n38636 );
and ( n38868 , n38600 , n38629 );
or ( n38869 , n38867 , n38868 );
buf ( n38870 , n38869 );
buf ( n38871 , n38870 );
xor ( n38872 , n38865 , n38871 );
xor ( n38873 , n38453 , n38504 );
and ( n38874 , n38873 , n38511 );
and ( n38875 , n38453 , n38504 );
or ( n38876 , n38874 , n38875 );
buf ( n38877 , n38876 );
buf ( n38878 , n38877 );
and ( n38879 , n38872 , n38878 );
and ( n38880 , n38865 , n38871 );
or ( n38881 , n38879 , n38880 );
buf ( n38882 , n38881 );
buf ( n38883 , n38882 );
xor ( n38884 , n38815 , n38883 );
buf ( n38885 , n5582 );
buf ( n38886 , n38482 );
or ( n38887 , n38885 , n38886 );
buf ( n38888 , n33118 );
buf ( n38889 , n38696 );
or ( n38890 , n38888 , n38889 );
nand ( n38891 , n38887 , n38890 );
buf ( n38892 , n38891 );
buf ( n38893 , n38892 );
buf ( n38894 , n534 );
buf ( n38895 , n537 );
and ( n38896 , n38894 , n38895 );
buf ( n38897 , n38896 );
buf ( n38898 , n38897 );
xor ( n38899 , n38893 , n38898 );
buf ( n38900 , n4030 );
buf ( n38901 , n38614 );
or ( n38902 , n38900 , n38901 );
buf ( n38903 , n4040 );
buf ( n38904 , n526 );
buf ( n38905 , n32981 );
and ( n38906 , n38904 , n38905 );
not ( n38907 , n38904 );
buf ( n38908 , n543 );
and ( n38909 , n38907 , n38908 );
nor ( n38910 , n38906 , n38909 );
buf ( n38911 , n38910 );
buf ( n38912 , n38911 );
or ( n38913 , n38903 , n38912 );
nand ( n38914 , n38902 , n38913 );
buf ( n38915 , n38914 );
buf ( n38916 , n38915 );
and ( n38917 , n38899 , n38916 );
and ( n38918 , n38893 , n38898 );
or ( n38919 , n38917 , n38918 );
buf ( n38920 , n38919 );
buf ( n38921 , n38920 );
buf ( n38922 , n38848 );
xor ( n38923 , n38921 , n38922 );
not ( n38924 , n2918 );
not ( n38925 , n2911 );
or ( n38926 , n38924 , n38925 );
nand ( n38927 , n38926 , n549 );
buf ( n38928 , n38927 );
buf ( n38929 , n5636 );
buf ( n38930 , n38911 );
or ( n38931 , n38929 , n38930 );
buf ( n38932 , n4040 );
buf ( n38933 , n32981 );
buf ( n38934 , n525 );
and ( n38935 , n38933 , n38934 );
buf ( n38936 , n34557 );
buf ( n38937 , n543 );
and ( n38938 , n38936 , n38937 );
nor ( n38939 , n38935 , n38938 );
buf ( n38940 , n38939 );
buf ( n38941 , n38940 );
or ( n38942 , n38932 , n38941 );
nand ( n38943 , n38931 , n38942 );
buf ( n38944 , n38943 );
buf ( n38945 , n38944 );
xor ( n38946 , n38928 , n38945 );
buf ( n38947 , n3020 );
buf ( n38948 , n38837 );
or ( n38949 , n38947 , n38948 );
buf ( n38950 , n31978 );
buf ( n38951 , n547 );
buf ( n38952 , n35343 );
and ( n38953 , n38951 , n38952 );
not ( n38954 , n38951 );
buf ( n38955 , n521 );
and ( n38956 , n38954 , n38955 );
nor ( n38957 , n38953 , n38956 );
buf ( n38958 , n38957 );
buf ( n38959 , n38958 );
or ( n38960 , n38950 , n38959 );
nand ( n38961 , n38949 , n38960 );
buf ( n38962 , n38961 );
buf ( n38963 , n38962 );
xor ( n38964 , n38946 , n38963 );
buf ( n38965 , n38964 );
buf ( n38966 , n38965 );
xor ( n38967 , n38923 , n38966 );
buf ( n38968 , n38967 );
buf ( n38969 , n38968 );
xor ( n38970 , n38852 , n38855 );
and ( n38971 , n38970 , n38862 );
and ( n38972 , n38852 , n38855 );
or ( n38973 , n38971 , n38972 );
buf ( n38974 , n38973 );
buf ( n38975 , n38974 );
xor ( n38976 , n38969 , n38975 );
xor ( n38977 , n38524 , n38541 );
and ( n38978 , n38977 , n38546 );
and ( n38979 , n38524 , n38541 );
or ( n38980 , n38978 , n38979 );
buf ( n38981 , n38980 );
buf ( n38982 , n38981 );
xor ( n38983 , n38893 , n38898 );
xor ( n38984 , n38983 , n38916 );
buf ( n38985 , n38984 );
buf ( n38986 , n38985 );
xor ( n38987 , n38982 , n38986 );
xor ( n38988 , n38658 , n38675 );
xor ( n38989 , n38988 , n38682 );
buf ( n38990 , n38989 );
buf ( n38991 , n38990 );
and ( n38992 , n38987 , n38991 );
and ( n38993 , n38982 , n38986 );
or ( n38994 , n38992 , n38993 );
buf ( n38995 , n38994 );
buf ( n38996 , n38995 );
xor ( n38997 , n38976 , n38996 );
buf ( n38998 , n38997 );
buf ( n38999 , n38998 );
xor ( n39000 , n38884 , n38999 );
buf ( n39001 , n39000 );
nand ( n39002 , n39001 , n3360 );
xor ( n39003 , n38982 , n38986 );
xor ( n39004 , n39003 , n38991 );
buf ( n39005 , n39004 );
xor ( n39006 , n38548 , n38554 );
and ( n39007 , n39006 , n38638 );
and ( n39008 , n38548 , n38554 );
or ( n39009 , n39007 , n39008 );
xor ( n39010 , n39005 , n39009 );
xor ( n39011 , n38865 , n38871 );
xor ( n39012 , n39011 , n38878 );
buf ( n39013 , n39012 );
and ( n39014 , n39010 , n39013 );
and ( n39015 , n39005 , n39009 );
or ( n39016 , n39014 , n39015 );
nand ( n39017 , n3138 , n39016 );
and ( n39018 , n39002 , n39017 );
not ( n39019 , n39018 );
buf ( n39020 , n29873 );
not ( n39021 , n39020 );
buf ( n39022 , n495 );
not ( n39023 , n39022 );
and ( n39024 , n456 , n459 );
not ( n39025 , n456 );
and ( n39026 , n39025 , n475 );
nor ( n39027 , n39024 , n39026 );
buf ( n39028 , n39027 );
not ( n39029 , n39028 );
or ( n39030 , n39023 , n39029 );
buf ( n39031 , n5062 );
buf ( n39032 , n29716 );
nand ( n39033 , n39031 , n39032 );
buf ( n39034 , n39033 );
buf ( n39035 , n39034 );
nand ( n39036 , n39030 , n39035 );
buf ( n39037 , n39036 );
buf ( n39038 , n39037 );
not ( n39039 , n39038 );
or ( n39040 , n39021 , n39039 );
buf ( n39041 , n30072 );
buf ( n39042 , n38160 );
nand ( n39043 , n39041 , n39042 );
buf ( n39044 , n39043 );
buf ( n39045 , n39044 );
nand ( n39046 , n39040 , n39045 );
buf ( n39047 , n39046 );
buf ( n39048 , n39047 );
buf ( n39049 , n37071 );
not ( n39050 , n39049 );
buf ( n39051 , n38178 );
not ( n39052 , n39051 );
or ( n39053 , n39050 , n39052 );
not ( n39054 , n7461 );
not ( n39055 , n30193 );
or ( n39056 , n39054 , n39055 );
nand ( n39057 , n489 , n29748 );
nand ( n39058 , n39056 , n39057 );
buf ( n39059 , n39058 );
buf ( n39060 , n7455 );
nand ( n39061 , n39059 , n39060 );
buf ( n39062 , n39061 );
buf ( n39063 , n39062 );
nand ( n39064 , n39053 , n39063 );
buf ( n39065 , n39064 );
buf ( n39066 , n39065 );
xor ( n39067 , n39048 , n39066 );
not ( n39068 , n34031 );
not ( n39069 , n38210 );
or ( n39070 , n39068 , n39069 );
buf ( n39071 , n491 );
not ( n39072 , n39071 );
buf ( n39073 , n34073 );
not ( n39074 , n39073 );
or ( n39075 , n39072 , n39074 );
buf ( n39076 , n33936 );
buf ( n39077 , n29505 );
nand ( n39078 , n39076 , n39077 );
buf ( n39079 , n39078 );
buf ( n39080 , n39079 );
nand ( n39081 , n39075 , n39080 );
buf ( n39082 , n39081 );
buf ( n39083 , n39082 );
buf ( n39084 , n4821 );
nand ( n39085 , n39083 , n39084 );
buf ( n39086 , n39085 );
nand ( n39087 , n39070 , n39086 );
buf ( n39088 , n39087 );
and ( n39089 , n39067 , n39088 );
and ( n39090 , n39048 , n39066 );
or ( n39091 , n39089 , n39090 );
buf ( n39092 , n39091 );
buf ( n39093 , n39092 );
not ( n39094 , n29582 );
not ( n39095 , n29623 );
not ( n39096 , n39095 );
or ( n39097 , n39094 , n39096 );
nand ( n39098 , n39097 , n499 );
buf ( n39099 , n39098 );
buf ( n39100 , n835 );
not ( n39101 , n39100 );
buf ( n39102 , n38235 );
not ( n39103 , n39102 );
or ( n39104 , n39101 , n39103 );
buf ( n39105 , n497 );
not ( n39106 , n39105 );
buf ( n39107 , n38009 );
not ( n39108 , n39107 );
or ( n39109 , n39106 , n39108 );
buf ( n39110 , n38013 );
buf ( n39111 , n706 );
nand ( n39112 , n39110 , n39111 );
buf ( n39113 , n39112 );
buf ( n39114 , n39113 );
nand ( n39115 , n39109 , n39114 );
buf ( n39116 , n39115 );
buf ( n39117 , n39116 );
buf ( n39118 , n29829 );
nand ( n39119 , n39117 , n39118 );
buf ( n39120 , n39119 );
buf ( n39121 , n39120 );
nand ( n39122 , n39104 , n39121 );
buf ( n39123 , n39122 );
buf ( n39124 , n39123 );
xor ( n39125 , n39099 , n39124 );
buf ( n39126 , n29522 );
not ( n39127 , n39126 );
buf ( n39128 , n493 );
not ( n39129 , n39128 );
buf ( n39130 , n36526 );
not ( n39131 , n39130 );
or ( n39132 , n39129 , n39131 );
not ( n39133 , n5226 );
nand ( n39134 , n39133 , n29537 );
buf ( n39135 , n39134 );
nand ( n39136 , n39132 , n39135 );
buf ( n39137 , n39136 );
buf ( n39138 , n39137 );
not ( n39139 , n39138 );
or ( n39140 , n39127 , n39139 );
nand ( n39141 , n38196 , n29576 );
buf ( n39142 , n39141 );
nand ( n39143 , n39140 , n39142 );
buf ( n39144 , n39143 );
buf ( n39145 , n39144 );
and ( n39146 , n39125 , n39145 );
and ( n39147 , n39099 , n39124 );
or ( n39148 , n39146 , n39147 );
buf ( n39149 , n39148 );
buf ( n39150 , n39149 );
xor ( n39151 , n39093 , n39150 );
buf ( n39152 , n34031 );
not ( n39153 , n39152 );
buf ( n39154 , n39082 );
not ( n39155 , n39154 );
or ( n39156 , n39153 , n39155 );
not ( n39157 , n33936 );
not ( n39158 , n36611 );
or ( n39159 , n39157 , n39158 );
nand ( n39160 , n37037 , n491 );
nand ( n39161 , n39159 , n39160 );
buf ( n39162 , n39161 );
buf ( n39163 , n4821 );
nand ( n39164 , n39162 , n39163 );
buf ( n39165 , n39164 );
buf ( n39166 , n39165 );
nand ( n39167 , n39156 , n39166 );
buf ( n39168 , n39167 );
buf ( n39169 , n39168 );
buf ( n39170 , n835 );
not ( n39171 , n39170 );
buf ( n39172 , n39116 );
not ( n39173 , n39172 );
or ( n39174 , n39171 , n39173 );
buf ( n39175 , n706 );
not ( n39176 , n39175 );
buf ( n39177 , n29829 );
nand ( n39178 , n39176 , n39177 );
buf ( n39179 , n39178 );
buf ( n39180 , n39179 );
nand ( n39181 , n39174 , n39180 );
buf ( n39182 , n39181 );
buf ( n39183 , n39182 );
xor ( n39184 , n39169 , n39183 );
buf ( n39185 , n39184 );
buf ( n39186 , n39185 );
not ( n39187 , n37071 );
not ( n39188 , n39058 );
or ( n39189 , n39187 , n39188 );
not ( n39190 , n489 );
not ( n39191 , n855 );
or ( n39192 , n39190 , n39191 );
not ( n39193 , n4966 );
nand ( n39194 , n39193 , n7461 );
nand ( n39195 , n39192 , n39194 );
nand ( n39196 , n39195 , n5328 );
nand ( n39197 , n39189 , n39196 );
buf ( n39198 , n39197 );
and ( n39199 , n39186 , n39198 );
not ( n39200 , n39186 );
buf ( n39201 , n39197 );
not ( n39202 , n39201 );
buf ( n39203 , n39202 );
buf ( n39204 , n39203 );
and ( n39205 , n39200 , n39204 );
nor ( n39206 , n39199 , n39205 );
buf ( n39207 , n39206 );
buf ( n39208 , n39207 );
xor ( n39209 , n39151 , n39208 );
buf ( n39210 , n39209 );
buf ( n39211 , n39210 );
xor ( n39212 , n38109 , n38117 );
and ( n39213 , n39212 , n38123 );
and ( n39214 , n38109 , n38117 );
or ( n39215 , n39213 , n39214 );
buf ( n39216 , n39215 );
buf ( n39217 , n489 );
not ( n39218 , n39217 );
buf ( n39219 , n971 );
nor ( n39220 , n39218 , n39219 );
buf ( n39221 , n39220 );
not ( n39222 , n38109 );
xor ( n39223 , n39221 , n39222 );
or ( n39224 , n38214 , n38203 );
nand ( n39225 , n39224 , n38240 );
nand ( n39226 , n38214 , n38203 );
nand ( n39227 , n39225 , n39226 );
xor ( n39228 , n39223 , n39227 );
buf ( n39229 , n39228 );
xor ( n39230 , n39216 , n39229 );
xor ( n39231 , n38138 , n38189 );
and ( n39232 , n39231 , n38246 );
and ( n39233 , n38138 , n38189 );
or ( n39234 , n39232 , n39233 );
buf ( n39235 , n39234 );
buf ( n39236 , n39235 );
and ( n39237 , n39230 , n39236 );
and ( n39238 , n39216 , n39229 );
or ( n39239 , n39237 , n39238 );
buf ( n39240 , n39239 );
buf ( n39241 , n39240 );
xor ( n39242 , n39211 , n39241 );
and ( n39243 , n38175 , n38176 );
buf ( n39244 , n39243 );
buf ( n39245 , n39244 );
buf ( n39246 , n29873 );
not ( n39247 , n39246 );
buf ( n39248 , n495 );
not ( n39249 , n39248 );
buf ( n39250 , n38227 );
not ( n39251 , n39250 );
or ( n39252 , n39249 , n39251 );
buf ( n39253 , n38228 );
buf ( n39254 , n29716 );
nand ( n39255 , n39253 , n39254 );
buf ( n39256 , n39255 );
buf ( n39257 , n39256 );
nand ( n39258 , n39252 , n39257 );
buf ( n39259 , n39258 );
buf ( n39260 , n39259 );
not ( n39261 , n39260 );
or ( n39262 , n39247 , n39261 );
buf ( n39263 , n39037 );
buf ( n39264 , n30072 );
nand ( n39265 , n39263 , n39264 );
buf ( n39266 , n39265 );
buf ( n39267 , n39266 );
nand ( n39268 , n39262 , n39267 );
buf ( n39269 , n39268 );
buf ( n39270 , n39269 );
not ( n39271 , n39270 );
buf ( n39272 , n39271 );
buf ( n39273 , n39272 );
xor ( n39274 , n39245 , n39273 );
buf ( n39275 , n29576 );
buf ( n39276 , n39275 );
buf ( n39277 , n39276 );
buf ( n39278 , n39277 );
not ( n39279 , n39278 );
buf ( n39280 , n39137 );
not ( n39281 , n39280 );
or ( n39282 , n39279 , n39281 );
buf ( n39283 , n493 );
not ( n39284 , n39283 );
buf ( n39285 , n7573 );
not ( n39286 , n39285 );
or ( n39287 , n39284 , n39286 );
and ( n39288 , n456 , n5355 );
not ( n39289 , n456 );
not ( n39290 , n476 );
and ( n39291 , n39289 , n39290 );
nor ( n39292 , n39288 , n39291 );
nand ( n39293 , n39292 , n29537 );
buf ( n39294 , n39293 );
nand ( n39295 , n39287 , n39294 );
buf ( n39296 , n39295 );
buf ( n39297 , n39296 );
buf ( n39298 , n29522 );
nand ( n39299 , n39297 , n39298 );
buf ( n39300 , n39299 );
buf ( n39301 , n39300 );
nand ( n39302 , n39282 , n39301 );
buf ( n39303 , n39302 );
buf ( n39304 , n39303 );
xor ( n39305 , n39274 , n39304 );
buf ( n39306 , n39305 );
buf ( n39307 , n39306 );
xor ( n39308 , n39221 , n39222 );
and ( n39309 , n39308 , n39227 );
and ( n39310 , n39221 , n39222 );
or ( n39311 , n39309 , n39310 );
buf ( n39312 , n39311 );
xor ( n39313 , n39307 , n39312 );
xor ( n39314 , n38143 , n38168 );
and ( n39315 , n39314 , n38186 );
and ( n39316 , n38143 , n38168 );
or ( n39317 , n39315 , n39316 );
buf ( n39318 , n39317 );
buf ( n39319 , n39318 );
xor ( n39320 , n39099 , n39124 );
xor ( n39321 , n39320 , n39145 );
buf ( n39322 , n39321 );
buf ( n39323 , n39322 );
xor ( n39324 , n39319 , n39323 );
xor ( n39325 , n39048 , n39066 );
xor ( n39326 , n39325 , n39088 );
buf ( n39327 , n39326 );
buf ( n39328 , n39327 );
and ( n39329 , n39324 , n39328 );
and ( n39330 , n39319 , n39323 );
or ( n39331 , n39329 , n39330 );
buf ( n39332 , n39331 );
buf ( n39333 , n39332 );
xor ( n39334 , n39313 , n39333 );
buf ( n39335 , n39334 );
buf ( n39336 , n39335 );
xor ( n39337 , n39242 , n39336 );
buf ( n39338 , n39337 );
not ( n39339 , n39338 );
xor ( n39340 , n39319 , n39323 );
xor ( n39341 , n39340 , n39328 );
buf ( n39342 , n39341 );
buf ( n39343 , n39342 );
xor ( n39344 , n39216 , n39229 );
xor ( n39345 , n39344 , n39236 );
buf ( n39346 , n39345 );
buf ( n39347 , n39346 );
xor ( n39348 , n39343 , n39347 );
xor ( n39349 , n38125 , n38131 );
and ( n39350 , n39349 , n38249 );
and ( n39351 , n38125 , n38131 );
or ( n39352 , n39350 , n39351 );
buf ( n39353 , n39352 );
buf ( n39354 , n39353 );
and ( n39355 , n39348 , n39354 );
and ( n39356 , n39343 , n39347 );
or ( n39357 , n39355 , n39356 );
buf ( n39358 , n39357 );
not ( n39359 , n39358 );
nand ( n39360 , n39339 , n39359 );
buf ( n39361 , n39360 );
nand ( n39362 , n39338 , n39358 );
buf ( n39363 , n39362 );
nand ( n39364 , n39361 , n39363 );
not ( n39365 , n39364 );
nand ( n39366 , n39365 , n455 );
xor ( n39367 , n38100 , n38105 );
and ( n39368 , n39367 , n38251 );
and ( n39369 , n38100 , n38105 );
or ( n39370 , n39368 , n39369 );
xor ( n39371 , n39343 , n39347 );
xor ( n39372 , n39371 , n39354 );
buf ( n39373 , n39372 );
nor ( n39374 , n39370 , n39373 );
nor ( n39375 , n39374 , n38262 );
not ( n39376 , n39375 );
nand ( n39377 , n39370 , n39373 );
not ( n39378 , n39377 );
not ( n39379 , n39378 );
nand ( n39380 , n39376 , n39379 );
nor ( n39381 , n39366 , n39380 );
not ( n39382 , n39381 );
not ( n39383 , n39374 );
nand ( n39384 , n39383 , n38260 );
buf ( n39385 , n39384 );
not ( n39386 , n39385 );
nand ( n39387 , n38095 , n39386 );
not ( n39388 , n39387 );
or ( n39389 , n39382 , n39388 );
and ( n39390 , n39364 , n455 );
nand ( n39391 , n39380 , n39390 );
nand ( n39392 , n39389 , n39391 );
not ( n39393 , n39392 );
not ( n39394 , n39387 );
nand ( n39395 , n39394 , n39390 );
nand ( n39396 , n39393 , n39395 );
xor ( n39397 , n38300 , n38304 );
and ( n39398 , n39397 , n38433 );
and ( n39399 , n38300 , n38304 );
or ( n39400 , n39398 , n39399 );
not ( n39401 , n39400 );
not ( n39402 , n39401 );
xor ( n39403 , n38389 , n38406 );
and ( n39404 , n39403 , n38425 );
and ( n39405 , n38389 , n38406 );
or ( n39406 , n39404 , n39405 );
buf ( n39407 , n39406 );
buf ( n39408 , n39407 );
not ( n39409 , n38349 );
not ( n39410 , n2213 );
or ( n39411 , n39409 , n39410 );
buf ( n39412 , n2081 );
buf ( n39413 , n505 );
buf ( n39414 , n497 );
xor ( n39415 , n39413 , n39414 );
buf ( n39416 , n39415 );
buf ( n39417 , n39416 );
nand ( n39418 , n39412 , n39417 );
buf ( n39419 , n39418 );
nand ( n39420 , n39411 , n39419 );
buf ( n39421 , n39420 );
not ( n39422 , n30881 );
not ( n39423 , n2000 );
or ( n39424 , n39422 , n39423 );
nand ( n39425 , n39424 , n499 );
buf ( n39426 , n39425 );
xor ( n39427 , n39421 , n39426 );
buf ( n39428 , n38377 );
not ( n39429 , n39428 );
buf ( n39430 , n2668 );
not ( n39431 , n39430 );
or ( n39432 , n39429 , n39431 );
buf ( n39433 , n2591 );
buf ( n39434 , n509 );
buf ( n39435 , n493 );
xor ( n39436 , n39434 , n39435 );
buf ( n39437 , n39436 );
buf ( n39438 , n39437 );
nand ( n39439 , n39433 , n39438 );
buf ( n39440 , n39439 );
buf ( n39441 , n39440 );
nand ( n39442 , n39432 , n39441 );
buf ( n39443 , n39442 );
buf ( n39444 , n39443 );
xor ( n39445 , n39427 , n39444 );
buf ( n39446 , n39445 );
buf ( n39447 , n39446 );
xor ( n39448 , n39408 , n39447 );
buf ( n39449 , n38418 );
not ( n39450 , n39449 );
buf ( n39451 , n38410 );
not ( n39452 , n39451 );
or ( n39453 , n39450 , n39452 );
buf ( n39454 , n35832 );
buf ( n39455 , n489 );
buf ( n39456 , n513 );
xor ( n39457 , n39455 , n39456 );
buf ( n39458 , n39457 );
buf ( n39459 , n39458 );
nand ( n39460 , n39454 , n39459 );
buf ( n39461 , n39460 );
buf ( n39462 , n39461 );
nand ( n39463 , n39453 , n39462 );
buf ( n39464 , n39463 );
buf ( n39465 , n39464 );
buf ( n39466 , n38361 );
not ( n39467 , n39466 );
buf ( n39468 , n4512 );
not ( n39469 , n39468 );
or ( n39470 , n39467 , n39469 );
buf ( n39471 , n4519 );
buf ( n39472 , n511 );
buf ( n39473 , n491 );
xor ( n39474 , n39472 , n39473 );
buf ( n39475 , n39474 );
buf ( n39476 , n39475 );
nand ( n39477 , n39471 , n39476 );
buf ( n39478 , n39477 );
buf ( n39479 , n39478 );
nand ( n39480 , n39470 , n39479 );
buf ( n39481 , n39480 );
buf ( n39482 , n39481 );
xor ( n39483 , n39465 , n39482 );
buf ( n39484 , n38398 );
not ( n39485 , n39484 );
buf ( n39486 , n2412 );
not ( n39487 , n39486 );
or ( n39488 , n39485 , n39487 );
buf ( n39489 , n507 );
buf ( n39490 , n495 );
xnor ( n39491 , n39489 , n39490 );
buf ( n39492 , n39491 );
buf ( n39493 , n39492 );
not ( n39494 , n39493 );
buf ( n39495 , n31271 );
nand ( n39496 , n39494 , n39495 );
buf ( n39497 , n39496 );
buf ( n39498 , n39497 );
nand ( n39499 , n39488 , n39498 );
buf ( n39500 , n39499 );
buf ( n39501 , n39500 );
xor ( n39502 , n39483 , n39501 );
buf ( n39503 , n39502 );
buf ( n39504 , n39503 );
xor ( n39505 , n39448 , n39504 );
buf ( n39506 , n39505 );
not ( n39507 , n38351 );
not ( n39508 , n38367 );
nand ( n39509 , n39507 , n39508 );
not ( n39510 , n39509 );
not ( n39511 , n38381 );
or ( n39512 , n39510 , n39511 );
nand ( n39513 , n38351 , n38367 );
nand ( n39514 , n39512 , n39513 );
not ( n39515 , n39514 );
and ( n39516 , n37722 , n37723 );
buf ( n39517 , n39516 );
not ( n39518 , n39517 );
not ( n39519 , n38313 );
or ( n39520 , n39518 , n39519 );
or ( n39521 , n38313 , n39517 );
nand ( n39522 , n39520 , n39521 );
not ( n39523 , n39522 );
or ( n39524 , n39515 , n39523 );
or ( n39525 , n39522 , n39514 );
nand ( n39526 , n39524 , n39525 );
xor ( n39527 , n38315 , n38320 );
and ( n39528 , n39527 , n38326 );
and ( n39529 , n38315 , n38320 );
or ( n39530 , n39528 , n39529 );
buf ( n39531 , n39530 );
xor ( n39532 , n39526 , n39531 );
xor ( n39533 , n38345 , n38383 );
and ( n39534 , n39533 , n38428 );
and ( n39535 , n38345 , n38383 );
or ( n39536 , n39534 , n39535 );
buf ( n39537 , n39536 );
xor ( n39538 , n39532 , n39537 );
xor ( n39539 , n39506 , n39538 );
xor ( n39540 , n38329 , n38335 );
and ( n39541 , n39540 , n38431 );
and ( n39542 , n38329 , n38335 );
or ( n39543 , n39541 , n39542 );
buf ( n39544 , n39543 );
xor ( n39545 , n39539 , n39544 );
not ( n39546 , n39545 );
not ( n39547 , n39546 );
or ( n39548 , n39402 , n39547 );
not ( n39549 , n38434 );
not ( n39550 , n38295 );
nand ( n39551 , n39549 , n39550 );
nand ( n39552 , n39548 , n39551 );
not ( n39553 , n39552 );
not ( n39554 , n39553 );
not ( n39555 , n38291 );
or ( n39556 , n39554 , n39555 );
nor ( n39557 , n39545 , n39400 );
nor ( n39558 , n39557 , n38435 );
not ( n39559 , n39558 );
nand ( n39560 , n39545 , n39400 );
buf ( n39561 , n39560 );
nand ( n39562 , n39559 , n39561 );
not ( n39563 , n39562 );
nand ( n39564 , n39556 , n39563 );
xor ( n39565 , n39421 , n39426 );
and ( n39566 , n39565 , n39444 );
and ( n39567 , n39421 , n39426 );
or ( n39568 , n39566 , n39567 );
buf ( n39569 , n39568 );
buf ( n39570 , n39569 );
buf ( n39571 , n39416 );
not ( n39572 , n39571 );
buf ( n39573 , n2213 );
not ( n39574 , n39573 );
or ( n39575 , n39572 , n39574 );
buf ( n39576 , n497 );
buf ( n39577 , n2081 );
nand ( n39578 , n39576 , n39577 );
buf ( n39579 , n39578 );
buf ( n39580 , n39579 );
nand ( n39581 , n39575 , n39580 );
buf ( n39582 , n39581 );
not ( n39583 , n39458 );
not ( n39584 , n38410 );
or ( n39585 , n39583 , n39584 );
buf ( n39586 , n35832 );
buf ( n39587 , n489 );
buf ( n39588 , n512 );
xor ( n39589 , n39587 , n39588 );
buf ( n39590 , n39589 );
buf ( n39591 , n39590 );
nand ( n39592 , n39586 , n39591 );
buf ( n39593 , n39592 );
nand ( n39594 , n39585 , n39593 );
xor ( n39595 , n39582 , n39594 );
buf ( n39596 , n39475 );
not ( n39597 , n39596 );
buf ( n39598 , n33438 );
not ( n39599 , n39598 );
or ( n39600 , n39597 , n39599 );
buf ( n39601 , n4519 );
buf ( n39602 , n510 );
buf ( n39603 , n491 );
xor ( n39604 , n39602 , n39603 );
buf ( n39605 , n39604 );
buf ( n39606 , n39605 );
nand ( n39607 , n39601 , n39606 );
buf ( n39608 , n39607 );
buf ( n39609 , n39608 );
nand ( n39610 , n39600 , n39609 );
buf ( n39611 , n39610 );
xor ( n39612 , n39595 , n39611 );
buf ( n39613 , n39612 );
xor ( n39614 , n39570 , n39613 );
xor ( n39615 , n39465 , n39482 );
and ( n39616 , n39615 , n39501 );
and ( n39617 , n39465 , n39482 );
or ( n39618 , n39616 , n39617 );
buf ( n39619 , n39618 );
buf ( n39620 , n39619 );
xor ( n39621 , n39614 , n39620 );
buf ( n39622 , n39621 );
xor ( n39623 , n39526 , n39531 );
and ( n39624 , n39623 , n39537 );
and ( n39625 , n39526 , n39531 );
or ( n39626 , n39624 , n39625 );
xor ( n39627 , n39622 , n39626 );
and ( n39628 , n38415 , n38416 );
buf ( n39629 , n39628 );
buf ( n39630 , n39629 );
buf ( n39631 , n39437 );
not ( n39632 , n39631 );
buf ( n39633 , n31660 );
not ( n39634 , n39633 );
or ( n39635 , n39632 , n39634 );
buf ( n39636 , n2591 );
buf ( n39637 , n508 );
buf ( n39638 , n493 );
xor ( n39639 , n39637 , n39638 );
buf ( n39640 , n39639 );
buf ( n39641 , n39640 );
nand ( n39642 , n39636 , n39641 );
buf ( n39643 , n39642 );
buf ( n39644 , n39643 );
nand ( n39645 , n39635 , n39644 );
buf ( n39646 , n39645 );
buf ( n39647 , n39646 );
xor ( n39648 , n39630 , n39647 );
buf ( n39649 , n31271 );
not ( n39650 , n39649 );
buf ( n39651 , n506 );
buf ( n39652 , n495 );
xor ( n39653 , n39651 , n39652 );
buf ( n39654 , n39653 );
buf ( n39655 , n39654 );
not ( n39656 , n39655 );
or ( n39657 , n39650 , n39656 );
buf ( n39658 , n2411 );
buf ( n39659 , n39492 );
or ( n39660 , n39658 , n39659 );
nand ( n39661 , n39657 , n39660 );
buf ( n39662 , n39661 );
buf ( n39663 , n39662 );
not ( n39664 , n39663 );
buf ( n39665 , n39664 );
buf ( n39666 , n39665 );
xor ( n39667 , n39648 , n39666 );
buf ( n39668 , n39667 );
not ( n39669 , n39517 );
not ( n39670 , n38313 );
or ( n39671 , n39669 , n39670 );
or ( n39672 , n38313 , n39517 );
nand ( n39673 , n39672 , n39514 );
nand ( n39674 , n39671 , n39673 );
xor ( n39675 , n39668 , n39674 );
xor ( n39676 , n39408 , n39447 );
and ( n39677 , n39676 , n39504 );
and ( n39678 , n39408 , n39447 );
or ( n39679 , n39677 , n39678 );
buf ( n39680 , n39679 );
xor ( n39681 , n39675 , n39680 );
xor ( n39682 , n39627 , n39681 );
not ( n39683 , n39682 );
xor ( n39684 , n39506 , n39538 );
and ( n39685 , n39684 , n39544 );
and ( n39686 , n39506 , n39538 );
or ( n39687 , n39685 , n39686 );
not ( n39688 , n39687 );
nand ( n39689 , n39683 , n39688 );
buf ( n39690 , n39689 );
not ( n39691 , n39690 );
nand ( n39692 , n39687 , n39682 );
not ( n39693 , n39692 );
nor ( n39694 , n39691 , n39693 );
or ( n39695 , n39694 , n455 );
and ( n39696 , n39564 , n39695 );
not ( n39697 , n39564 );
nand ( n39698 , n39690 , n39692 , n2815 );
and ( n39699 , n39697 , n39698 );
nor ( n39700 , n39696 , n39699 );
or ( n39701 , n39396 , n39700 );
nand ( n39702 , n39701 , n454 );
not ( n39703 , n39702 );
or ( n39704 , n39019 , n39703 );
not ( n39705 , n38261 );
not ( n39706 , n38095 );
or ( n39707 , n39705 , n39706 );
nand ( n39708 , n39707 , n38263 );
not ( n39709 , n39708 );
not ( n39710 , n39709 );
nand ( n39711 , n39383 , n39379 );
nand ( n39712 , n39711 , n455 );
not ( n39713 , n39712 );
and ( n39714 , n39710 , n39713 );
not ( n39715 , n39708 );
not ( n39716 , n39711 );
and ( n39717 , n39716 , n455 );
and ( n39718 , n39715 , n39717 );
nor ( n39719 , n39714 , n39718 );
not ( n39720 , n39551 );
not ( n39721 , n38291 );
or ( n39722 , n39720 , n39721 );
nand ( n39723 , n39722 , n38435 );
not ( n39724 , n39723 );
not ( n39725 , n39557 );
nand ( n39726 , n39725 , n39561 );
not ( n39727 , n39726 );
nand ( n39728 , n39727 , n29516 );
not ( n39729 , n39728 );
and ( n39730 , n39724 , n39729 );
and ( n39731 , n39726 , n29516 );
and ( n39732 , n39723 , n39731 );
nor ( n39733 , n39730 , n39732 );
nand ( n39734 , n39719 , n39733 );
and ( n39735 , n39734 , n454 );
xor ( n39736 , n38514 , n38520 );
and ( n39737 , n39736 , n38640 );
and ( n39738 , n38514 , n38520 );
or ( n39739 , n39737 , n39738 );
buf ( n39740 , n39739 );
nand ( n39741 , n39740 , n3138 );
xor ( n39742 , n39005 , n39009 );
xor ( n39743 , n39742 , n39013 );
nand ( n39744 , n39743 , n3360 );
nand ( n39745 , n39741 , n39744 );
nor ( n39746 , n39735 , n39745 );
not ( n39747 , n39746 );
nand ( n39748 , n39704 , n39747 );
nor ( n39749 , n38657 , n39748 );
xor ( n39750 , n39622 , n39626 );
and ( n39751 , n39750 , n39681 );
and ( n39752 , n39622 , n39626 );
or ( n39753 , n39751 , n39752 );
xor ( n39754 , n39570 , n39613 );
and ( n39755 , n39754 , n39620 );
and ( n39756 , n39570 , n39613 );
or ( n39757 , n39755 , n39756 );
buf ( n39758 , n39757 );
buf ( n39759 , n39758 );
xor ( n39760 , n39668 , n39674 );
and ( n39761 , n39760 , n39680 );
and ( n39762 , n39668 , n39674 );
or ( n39763 , n39761 , n39762 );
buf ( n39764 , n39763 );
xor ( n39765 , n39759 , n39764 );
xor ( n39766 , n39630 , n39647 );
and ( n39767 , n39766 , n39666 );
and ( n39768 , n39630 , n39647 );
or ( n39769 , n39767 , n39768 );
buf ( n39770 , n39769 );
buf ( n39771 , n39770 );
buf ( n39772 , n31286 );
not ( n39773 , n39772 );
buf ( n39774 , n31280 );
not ( n39775 , n39774 );
or ( n39776 , n39773 , n39775 );
buf ( n39777 , n497 );
nand ( n39778 , n39776 , n39777 );
buf ( n39779 , n39778 );
buf ( n39780 , n39779 );
buf ( n39781 , n39605 );
not ( n39782 , n39781 );
buf ( n39783 , n33438 );
not ( n39784 , n39783 );
or ( n39785 , n39782 , n39784 );
buf ( n39786 , n4519 );
buf ( n39787 , n491 );
buf ( n39788 , n509 );
xor ( n39789 , n39787 , n39788 );
buf ( n39790 , n39789 );
buf ( n39791 , n39790 );
nand ( n39792 , n39786 , n39791 );
buf ( n39793 , n39792 );
buf ( n39794 , n39793 );
nand ( n39795 , n39785 , n39794 );
buf ( n39796 , n39795 );
buf ( n39797 , n39796 );
xor ( n39798 , n39780 , n39797 );
buf ( n39799 , n39654 );
not ( n39800 , n39799 );
buf ( n39801 , n2412 );
not ( n39802 , n39801 );
or ( n39803 , n39800 , n39802 );
buf ( n39804 , n495 );
buf ( n39805 , n505 );
xnor ( n39806 , n39804 , n39805 );
buf ( n39807 , n39806 );
buf ( n39808 , n39807 );
not ( n39809 , n39808 );
buf ( n39810 , n31271 );
nand ( n39811 , n39809 , n39810 );
buf ( n39812 , n39811 );
buf ( n39813 , n39812 );
nand ( n39814 , n39803 , n39813 );
buf ( n39815 , n39814 );
buf ( n39816 , n39815 );
xor ( n39817 , n39798 , n39816 );
buf ( n39818 , n39817 );
buf ( n39819 , n39818 );
xor ( n39820 , n39771 , n39819 );
buf ( n39821 , n39662 );
buf ( n39822 , n39594 );
not ( n39823 , n39822 );
buf ( n39824 , n39582 );
not ( n39825 , n39824 );
or ( n39826 , n39823 , n39825 );
buf ( n39827 , n39594 );
buf ( n39828 , n39582 );
or ( n39829 , n39827 , n39828 );
buf ( n39830 , n39611 );
nand ( n39831 , n39829 , n39830 );
buf ( n39832 , n39831 );
buf ( n39833 , n39832 );
nand ( n39834 , n39826 , n39833 );
buf ( n39835 , n39834 );
buf ( n39836 , n39835 );
xor ( n39837 , n39821 , n39836 );
and ( n39838 , n39455 , n39456 );
buf ( n39839 , n39838 );
buf ( n39840 , n39839 );
buf ( n39841 , n39590 );
not ( n39842 , n39841 );
buf ( n39843 , n38410 );
not ( n39844 , n39843 );
or ( n39845 , n39842 , n39844 );
buf ( n39846 , n35832 );
buf ( n39847 , n489 );
buf ( n39848 , n511 );
xor ( n39849 , n39847 , n39848 );
buf ( n39850 , n39849 );
buf ( n39851 , n39850 );
nand ( n39852 , n39846 , n39851 );
buf ( n39853 , n39852 );
buf ( n39854 , n39853 );
nand ( n39855 , n39845 , n39854 );
buf ( n39856 , n39855 );
buf ( n39857 , n39856 );
xor ( n39858 , n39840 , n39857 );
buf ( n39859 , n39640 );
not ( n39860 , n39859 );
buf ( n39861 , n2668 );
not ( n39862 , n39861 );
or ( n39863 , n39860 , n39862 );
buf ( n39864 , n2591 );
buf ( n39865 , n507 );
buf ( n39866 , n493 );
xor ( n39867 , n39865 , n39866 );
buf ( n39868 , n39867 );
buf ( n39869 , n39868 );
nand ( n39870 , n39864 , n39869 );
buf ( n39871 , n39870 );
buf ( n39872 , n39871 );
nand ( n39873 , n39863 , n39872 );
buf ( n39874 , n39873 );
buf ( n39875 , n39874 );
xor ( n39876 , n39858 , n39875 );
buf ( n39877 , n39876 );
buf ( n39878 , n39877 );
xor ( n39879 , n39837 , n39878 );
buf ( n39880 , n39879 );
buf ( n39881 , n39880 );
xor ( n39882 , n39820 , n39881 );
buf ( n39883 , n39882 );
buf ( n39884 , n39883 );
xor ( n39885 , n39765 , n39884 );
buf ( n39886 , n39885 );
nand ( n39887 , n39753 , n39886 );
nor ( n39888 , n39753 , n39886 );
not ( n39889 , n39888 );
nand ( n39890 , n39887 , n39889 );
and ( n39891 , n39890 , n2815 , n454 );
not ( n39892 , n39891 );
nand ( n39893 , n39553 , n39690 );
not ( n39894 , n39893 );
not ( n39895 , n39894 );
not ( n39896 , n38291 );
or ( n39897 , n39895 , n39896 );
and ( n39898 , n39562 , n39690 );
nor ( n39899 , n39898 , n39693 );
nand ( n39900 , n39897 , n39899 );
not ( n39901 , n39900 );
or ( n39902 , n39892 , n39901 );
xor ( n39903 , n38815 , n38883 );
and ( n39904 , n39903 , n38999 );
and ( n39905 , n38815 , n38883 );
or ( n39906 , n39904 , n39905 );
buf ( n39907 , n39906 );
buf ( n39908 , n39907 );
buf ( n39909 , n3138 );
nand ( n39910 , n39908 , n39909 );
buf ( n39911 , n39910 );
nand ( n39912 , n39902 , n39911 );
not ( n39913 , n39912 );
not ( n39914 , n39900 );
not ( n39915 , n454 );
not ( n39916 , n39890 );
nand ( n39917 , n39916 , n2815 );
nor ( n39918 , n39915 , n39917 );
nand ( n39919 , n39914 , n39918 );
not ( n39920 , n39361 );
nor ( n39921 , n39385 , n39920 );
not ( n39922 , n39921 );
not ( n39923 , n38095 );
or ( n39924 , n39922 , n39923 );
and ( n39925 , n39361 , n39380 );
not ( n39926 , n39363 );
nor ( n39927 , n39925 , n39926 );
nand ( n39928 , n39924 , n39927 );
not ( n39929 , n39928 );
xor ( n39930 , n39093 , n39150 );
and ( n39931 , n39930 , n39208 );
and ( n39932 , n39093 , n39150 );
or ( n39933 , n39931 , n39932 );
buf ( n39934 , n39933 );
buf ( n39935 , n39934 );
xor ( n39936 , n39245 , n39273 );
and ( n39937 , n39936 , n39304 );
and ( n39938 , n39245 , n39273 );
or ( n39939 , n39937 , n39938 );
buf ( n39940 , n39939 );
buf ( n39941 , n39940 );
buf ( n39942 , n36744 );
not ( n39943 , n39942 );
buf ( n39944 , n834 );
not ( n39945 , n39944 );
or ( n39946 , n39943 , n39945 );
buf ( n39947 , n497 );
nand ( n39948 , n39946 , n39947 );
buf ( n39949 , n39948 );
buf ( n39950 , n39949 );
buf ( n39951 , n30072 );
not ( n39952 , n39951 );
buf ( n39953 , n39259 );
not ( n39954 , n39953 );
or ( n39955 , n39952 , n39954 );
buf ( n39956 , n495 );
not ( n39957 , n39956 );
buf ( n39958 , n38009 );
not ( n39959 , n39958 );
or ( n39960 , n39957 , n39959 );
buf ( n39961 , n38013 );
buf ( n39962 , n29716 );
nand ( n39963 , n39961 , n39962 );
buf ( n39964 , n39963 );
buf ( n39965 , n39964 );
nand ( n39966 , n39960 , n39965 );
buf ( n39967 , n39966 );
buf ( n39968 , n39967 );
buf ( n39969 , n29873 );
nand ( n39970 , n39968 , n39969 );
buf ( n39971 , n39970 );
buf ( n39972 , n39971 );
nand ( n39973 , n39955 , n39972 );
buf ( n39974 , n39973 );
buf ( n39975 , n39974 );
xor ( n39976 , n39950 , n39975 );
buf ( n39977 , n34031 );
not ( n39978 , n39977 );
buf ( n39979 , n39161 );
not ( n39980 , n39979 );
or ( n39981 , n39978 , n39980 );
buf ( n39982 , n491 );
not ( n39983 , n39982 );
buf ( n39984 , n36526 );
not ( n39985 , n39984 );
or ( n39986 , n39983 , n39985 );
buf ( n39987 , n39133 );
buf ( n39988 , n33936 );
nand ( n39989 , n39987 , n39988 );
buf ( n39990 , n39989 );
buf ( n39991 , n39990 );
nand ( n39992 , n39986 , n39991 );
buf ( n39993 , n39992 );
buf ( n39994 , n39993 );
buf ( n39995 , n4821 );
nand ( n39996 , n39994 , n39995 );
buf ( n39997 , n39996 );
buf ( n39998 , n39997 );
nand ( n39999 , n39981 , n39998 );
buf ( n40000 , n39999 );
buf ( n40001 , n40000 );
xor ( n40002 , n39976 , n40001 );
buf ( n40003 , n40002 );
buf ( n40004 , n40003 );
xor ( n40005 , n39941 , n40004 );
buf ( n40006 , n39269 );
buf ( n40007 , n39197 );
buf ( n40008 , n39168 );
or ( n40009 , n40007 , n40008 );
buf ( n40010 , n39182 );
nand ( n40011 , n40009 , n40010 );
buf ( n40012 , n40011 );
buf ( n40013 , n40012 );
buf ( n40014 , n39197 );
buf ( n40015 , n39168 );
nand ( n40016 , n40014 , n40015 );
buf ( n40017 , n40016 );
buf ( n40018 , n40017 );
nand ( n40019 , n40013 , n40018 );
buf ( n40020 , n40019 );
buf ( n40021 , n40020 );
xor ( n40022 , n40006 , n40021 );
buf ( n40023 , n489 );
not ( n40024 , n40023 );
buf ( n40025 , n29591 );
nor ( n40026 , n40024 , n40025 );
buf ( n40027 , n40026 );
buf ( n40028 , n40027 );
buf ( n40029 , n29576 );
not ( n40030 , n40029 );
buf ( n40031 , n39296 );
not ( n40032 , n40031 );
or ( n40033 , n40030 , n40032 );
buf ( n40034 , n493 );
not ( n40035 , n40034 );
buf ( n40036 , n39027 );
not ( n40037 , n40036 );
or ( n40038 , n40035 , n40037 );
nand ( n40039 , n29537 , n5062 );
buf ( n40040 , n40039 );
nand ( n40041 , n40038 , n40040 );
buf ( n40042 , n40041 );
buf ( n40043 , n40042 );
buf ( n40044 , n29522 );
nand ( n40045 , n40043 , n40044 );
buf ( n40046 , n40045 );
buf ( n40047 , n40046 );
nand ( n40048 , n40033 , n40047 );
buf ( n40049 , n40048 );
buf ( n40050 , n40049 );
xor ( n40051 , n40028 , n40050 );
buf ( n40052 , n37071 );
not ( n40053 , n40052 );
buf ( n40054 , n39195 );
not ( n40055 , n40054 );
or ( n40056 , n40053 , n40055 );
buf ( n40057 , n34073 );
not ( n40058 , n40057 );
buf ( n40059 , n40058 );
xor ( n40060 , n489 , n40059 );
nand ( n40061 , n40060 , n7455 );
buf ( n40062 , n40061 );
nand ( n40063 , n40056 , n40062 );
buf ( n40064 , n40063 );
buf ( n40065 , n40064 );
xor ( n40066 , n40051 , n40065 );
buf ( n40067 , n40066 );
buf ( n40068 , n40067 );
xor ( n40069 , n40022 , n40068 );
buf ( n40070 , n40069 );
buf ( n40071 , n40070 );
xor ( n40072 , n40005 , n40071 );
buf ( n40073 , n40072 );
buf ( n40074 , n40073 );
xor ( n40075 , n39935 , n40074 );
xor ( n40076 , n39307 , n39312 );
and ( n40077 , n40076 , n39333 );
and ( n40078 , n39307 , n39312 );
or ( n40079 , n40077 , n40078 );
buf ( n40080 , n40079 );
buf ( n40081 , n40080 );
xor ( n40082 , n40075 , n40081 );
buf ( n40083 , n40082 );
xor ( n40084 , n39211 , n39241 );
and ( n40085 , n40084 , n39336 );
and ( n40086 , n39211 , n39241 );
or ( n40087 , n40085 , n40086 );
buf ( n40088 , n40087 );
or ( n40089 , n40083 , n40088 );
nand ( n40090 , n40083 , n40088 );
nand ( n40091 , n40089 , n40090 );
not ( n40092 , n5847 );
nand ( n40093 , n40092 , n455 );
nor ( n40094 , n40091 , n40093 );
nand ( n40095 , n39929 , n40094 );
and ( n40096 , n40091 , n455 );
nand ( n40097 , n39928 , n40096 , n454 );
nand ( n40098 , n39913 , n39919 , n40095 , n40097 );
buf ( n40099 , n6015 );
buf ( n40100 , n38767 );
or ( n40101 , n40099 , n40100 );
buf ( n40102 , n6010 );
buf ( n40103 , n6001 );
buf ( n40104 , n528 );
and ( n40105 , n40103 , n40104 );
buf ( n40106 , n32183 );
buf ( n40107 , n539 );
and ( n40108 , n40106 , n40107 );
nor ( n40109 , n40105 , n40108 );
buf ( n40110 , n40109 );
buf ( n40111 , n40110 );
or ( n40112 , n40102 , n40111 );
nand ( n40113 , n40101 , n40112 );
buf ( n40114 , n40113 );
buf ( n40115 , n5582 );
buf ( n40116 , n38707 );
or ( n40117 , n40115 , n40116 );
buf ( n40118 , n33118 );
buf ( n40119 , n541 );
buf ( n40120 , n526 );
not ( n40121 , n40120 );
buf ( n40122 , n40121 );
buf ( n40123 , n40122 );
and ( n40124 , n40119 , n40123 );
not ( n40125 , n40119 );
buf ( n40126 , n526 );
and ( n40127 , n40125 , n40126 );
nor ( n40128 , n40124 , n40127 );
buf ( n40129 , n40128 );
buf ( n40130 , n40129 );
or ( n40131 , n40118 , n40130 );
nand ( n40132 , n40117 , n40131 );
buf ( n40133 , n40132 );
xor ( n40134 , n40114 , n40133 );
buf ( n40135 , n3069 );
buf ( n40136 , n38738 );
or ( n40137 , n40135 , n40136 );
buf ( n40138 , n3087 );
buf ( n40139 , n32053 );
buf ( n40140 , n522 );
and ( n40141 , n40139 , n40140 );
buf ( n40142 , n35199 );
buf ( n40143 , n545 );
and ( n40144 , n40142 , n40143 );
nor ( n40145 , n40141 , n40144 );
buf ( n40146 , n40145 );
buf ( n40147 , n40146 );
or ( n40148 , n40138 , n40147 );
nand ( n40149 , n40137 , n40148 );
buf ( n40150 , n40149 );
xor ( n40151 , n40134 , n40150 );
buf ( n40152 , n6559 );
buf ( n40153 , n38785 );
or ( n40154 , n40152 , n40153 );
buf ( n40155 , n6337 );
buf ( n40156 , n6541 );
buf ( n40157 , n530 );
and ( n40158 , n40156 , n40157 );
buf ( n40159 , n31853 );
buf ( n40160 , n537 );
and ( n40161 , n40159 , n40160 );
nor ( n40162 , n40158 , n40161 );
buf ( n40163 , n40162 );
buf ( n40164 , n40163 );
or ( n40165 , n40155 , n40164 );
nand ( n40166 , n40154 , n40165 );
buf ( n40167 , n40166 );
buf ( n40168 , n40167 );
buf ( n40169 , n532 );
buf ( n40170 , n537 );
and ( n40171 , n40169 , n40170 );
buf ( n40172 , n40171 );
buf ( n40173 , n40172 );
xor ( n40174 , n40168 , n40173 );
buf ( n40175 , n5636 );
buf ( n40176 , n38940 );
or ( n40177 , n40175 , n40176 );
buf ( n40178 , n35070 );
buf ( n40179 , n32981 );
buf ( n40180 , n524 );
and ( n40181 , n40179 , n40180 );
buf ( n40182 , n34779 );
buf ( n40183 , n543 );
and ( n40184 , n40182 , n40183 );
nor ( n40185 , n40181 , n40184 );
buf ( n40186 , n40185 );
buf ( n40187 , n40186 );
or ( n40188 , n40178 , n40187 );
nand ( n40189 , n40177 , n40188 );
buf ( n40190 , n40189 );
buf ( n40191 , n40190 );
xor ( n40192 , n40174 , n40191 );
buf ( n40193 , n40192 );
xor ( n40194 , n38772 , n38790 );
and ( n40195 , n40194 , n38809 );
and ( n40196 , n38772 , n38790 );
or ( n40197 , n40195 , n40196 );
buf ( n40198 , n40197 );
xor ( n40199 , n40193 , n40198 );
xor ( n40200 , n40151 , n40199 );
buf ( n40201 , n40200 );
xor ( n40202 , n38969 , n38975 );
and ( n40203 , n40202 , n38996 );
and ( n40204 , n38969 , n38975 );
or ( n40205 , n40203 , n40204 );
buf ( n40206 , n40205 );
buf ( n40207 , n40206 );
xor ( n40208 , n40201 , n40207 );
xor ( n40209 , n38921 , n38922 );
and ( n40210 , n40209 , n38966 );
and ( n40211 , n38921 , n38922 );
or ( n40212 , n40210 , n40211 );
buf ( n40213 , n40212 );
buf ( n40214 , n40213 );
xor ( n40215 , n38712 , n38717 );
and ( n40216 , n40215 , n38743 );
and ( n40217 , n38712 , n38717 );
or ( n40218 , n40216 , n40217 );
buf ( n40219 , n40218 );
buf ( n40220 , n40219 );
buf ( n40221 , n3020 );
buf ( n40222 , n38958 );
or ( n40223 , n40221 , n40222 );
buf ( n40224 , n31978 );
buf ( n40225 , n547 );
not ( n40226 , n40225 );
buf ( n40227 , n40226 );
buf ( n40228 , n40227 );
or ( n40229 , n40224 , n40228 );
nand ( n40230 , n40223 , n40229 );
buf ( n40231 , n40230 );
buf ( n40232 , n40231 );
not ( n40233 , n40232 );
buf ( n40234 , n40233 );
buf ( n40235 , n40234 );
xor ( n40236 , n40220 , n40235 );
xor ( n40237 , n38928 , n38945 );
and ( n40238 , n40237 , n38963 );
and ( n40239 , n38928 , n38945 );
or ( n40240 , n40238 , n40239 );
buf ( n40241 , n40240 );
buf ( n40242 , n40241 );
xor ( n40243 , n40236 , n40242 );
buf ( n40244 , n40243 );
buf ( n40245 , n40244 );
xor ( n40246 , n40214 , n40245 );
xor ( n40247 , n38687 , n38746 );
and ( n40248 , n40247 , n38812 );
and ( n40249 , n38687 , n38746 );
or ( n40250 , n40248 , n40249 );
buf ( n40251 , n40250 );
buf ( n40252 , n40251 );
xor ( n40253 , n40246 , n40252 );
buf ( n40254 , n40253 );
buf ( n40255 , n40254 );
xor ( n40256 , n40208 , n40255 );
buf ( n40257 , n40256 );
and ( n40258 , n40257 , n3360 );
or ( n40259 , n40098 , n40258 );
nand ( n40260 , n37441 , n39749 , n40259 );
nand ( n40261 , n39700 , n454 );
nand ( n40262 , n39392 , n454 );
and ( n40263 , n39390 , n454 );
and ( n40264 , n39394 , n40263 );
not ( n40265 , n454 );
and ( n40266 , n39016 , n40265 );
nor ( n40267 , n40264 , n40266 );
and ( n40268 , n40261 , n40262 , n40267 , n39002 );
nor ( n40269 , n39746 , n40268 );
not ( n40270 , n40269 );
not ( n40271 , n37447 );
not ( n40272 , n38078 );
or ( n40273 , n40271 , n40272 );
nand ( n40274 , n40273 , n37662 );
not ( n40275 , n38654 );
or ( n40276 , n40274 , n40275 );
not ( n40277 , n38652 );
not ( n40278 , n40277 );
not ( n40279 , n38447 );
or ( n40280 , n40278 , n40279 );
nand ( n40281 , n40280 , n38646 );
nand ( n40282 , n40276 , n40281 );
not ( n40283 , n40282 );
or ( n40284 , n40270 , n40283 );
not ( n40285 , n39716 );
nand ( n40286 , n40285 , n39709 );
nand ( n40287 , n39716 , n39708 );
nand ( n40288 , n40286 , n40287 , n455 );
not ( n40289 , n40288 );
not ( n40290 , n39723 );
nand ( n40291 , n40290 , n39726 );
nand ( n40292 , n39723 , n39727 );
and ( n40293 , n40291 , n40292 , n29516 );
not ( n40294 , n39741 );
nor ( n40295 , n40293 , n40294 );
not ( n40296 , n40295 );
or ( n40297 , n40289 , n40296 );
not ( n40298 , n39744 );
nand ( n40299 , n39741 , n5847 );
and ( n40300 , n40298 , n40299 );
nand ( n40301 , n40297 , n40300 );
not ( n40302 , n40301 );
nand ( n40303 , n39018 , n39702 );
and ( n40304 , n40302 , n40303 );
nand ( n40305 , n40262 , n40267 );
not ( n40306 , n40261 );
or ( n40307 , n40305 , n40306 );
not ( n40308 , n39002 );
nand ( n40309 , n40307 , n40308 );
not ( n40310 , n40309 );
nor ( n40311 , n40304 , n40310 );
nand ( n40312 , n40284 , n40311 );
nand ( n40313 , n40259 , n40312 );
and ( n40314 , n40098 , n40258 );
buf ( n40315 , n40314 );
not ( n40316 , n40315 );
nand ( n40317 , n40260 , n40313 , n40316 );
not ( n40318 , n454 );
not ( n40319 , n455 );
nand ( n40320 , n39362 , n40090 );
nor ( n40321 , n39378 , n40320 );
and ( n40322 , n39384 , n40321 );
or ( n40323 , n40320 , n39360 );
nand ( n40324 , n40323 , n40089 );
nor ( n40325 , n40322 , n40324 );
not ( n40326 , n40325 );
nor ( n40327 , n39375 , n40320 );
not ( n40328 , n37197 );
not ( n40329 , n37201 );
and ( n40330 , n40328 , n40329 );
and ( n40331 , n36990 , n36991 );
nor ( n40332 , n40330 , n40331 );
nand ( n40333 , n40332 , n38089 , n36989 );
and ( n40334 , n39377 , n38055 );
nand ( n40335 , n37204 , n38089 );
nand ( n40336 , n40327 , n40333 , n40334 , n40335 );
not ( n40337 , n40336 );
or ( n40338 , n40326 , n40337 );
nand ( n40339 , n39360 , n40089 );
nor ( n40340 , n39384 , n40339 );
nand ( n40341 , n40340 , n36984 , n38082 );
nand ( n40342 , n40338 , n40341 );
xor ( n40343 , n39935 , n40074 );
and ( n40344 , n40343 , n40081 );
and ( n40345 , n39935 , n40074 );
or ( n40346 , n40344 , n40345 );
buf ( n40347 , n40346 );
xor ( n40348 , n40006 , n40021 );
and ( n40349 , n40348 , n40068 );
and ( n40350 , n40006 , n40021 );
or ( n40351 , n40349 , n40350 );
buf ( n40352 , n40351 );
buf ( n40353 , n40352 );
buf ( n40354 , n39193 );
buf ( n40355 , n489 );
and ( n40356 , n40354 , n40355 );
buf ( n40357 , n40356 );
buf ( n40358 , n40357 );
buf ( n40359 , n30072 );
not ( n40360 , n40359 );
buf ( n40361 , n39967 );
not ( n40362 , n40361 );
or ( n40363 , n40360 , n40362 );
buf ( n40364 , n29873 );
buf ( n40365 , n495 );
nand ( n40366 , n40364 , n40365 );
buf ( n40367 , n40366 );
buf ( n40368 , n40367 );
nand ( n40369 , n40363 , n40368 );
buf ( n40370 , n40369 );
buf ( n40371 , n40370 );
xor ( n40372 , n40358 , n40371 );
not ( n40373 , n37071 );
not ( n40374 , n40060 );
or ( n40375 , n40373 , n40374 );
buf ( n40376 , n489 );
not ( n40377 , n4835 );
buf ( n40378 , n40377 );
xor ( n40379 , n40376 , n40378 );
buf ( n40380 , n40379 );
buf ( n40381 , n40380 );
buf ( n40382 , n7455 );
nand ( n40383 , n40381 , n40382 );
buf ( n40384 , n40383 );
nand ( n40385 , n40375 , n40384 );
buf ( n40386 , n40385 );
xor ( n40387 , n40372 , n40386 );
buf ( n40388 , n40387 );
buf ( n40389 , n40388 );
xor ( n40390 , n39950 , n39975 );
and ( n40391 , n40390 , n40001 );
and ( n40392 , n39950 , n39975 );
or ( n40393 , n40391 , n40392 );
buf ( n40394 , n40393 );
buf ( n40395 , n40394 );
xor ( n40396 , n40389 , n40395 );
buf ( n40397 , n4821 );
not ( n40398 , n40397 );
buf ( n40399 , n491 );
not ( n40400 , n40399 );
buf ( n40401 , n7573 );
not ( n40402 , n40401 );
or ( n40403 , n40400 , n40402 );
nand ( n40404 , n39292 , n33936 );
buf ( n40405 , n40404 );
nand ( n40406 , n40403 , n40405 );
buf ( n40407 , n40406 );
buf ( n40408 , n40407 );
not ( n40409 , n40408 );
or ( n40410 , n40398 , n40409 );
buf ( n40411 , n39993 );
buf ( n40412 , n34031 );
nand ( n40413 , n40411 , n40412 );
buf ( n40414 , n40413 );
buf ( n40415 , n40414 );
nand ( n40416 , n40410 , n40415 );
buf ( n40417 , n40416 );
buf ( n40418 , n40417 );
buf ( n40419 , n29522 );
not ( n40420 , n40419 );
buf ( n40421 , n493 );
not ( n40422 , n40421 );
buf ( n40423 , n38227 );
not ( n40424 , n40423 );
or ( n40425 , n40422 , n40424 );
buf ( n40426 , n38228 );
buf ( n40427 , n29537 );
nand ( n40428 , n40426 , n40427 );
buf ( n40429 , n40428 );
buf ( n40430 , n40429 );
nand ( n40431 , n40425 , n40430 );
buf ( n40432 , n40431 );
buf ( n40433 , n40432 );
not ( n40434 , n40433 );
or ( n40435 , n40420 , n40434 );
buf ( n40436 , n40042 );
buf ( n40437 , n39277 );
nand ( n40438 , n40436 , n40437 );
buf ( n40439 , n40438 );
buf ( n40440 , n40439 );
nand ( n40441 , n40435 , n40440 );
buf ( n40442 , n40441 );
buf ( n40443 , n40442 );
not ( n40444 , n40443 );
buf ( n40445 , n40444 );
buf ( n40446 , n40445 );
xor ( n40447 , n40418 , n40446 );
xor ( n40448 , n40028 , n40050 );
and ( n40449 , n40448 , n40065 );
and ( n40450 , n40028 , n40050 );
or ( n40451 , n40449 , n40450 );
buf ( n40452 , n40451 );
buf ( n40453 , n40452 );
xor ( n40454 , n40447 , n40453 );
buf ( n40455 , n40454 );
buf ( n40456 , n40455 );
xor ( n40457 , n40396 , n40456 );
buf ( n40458 , n40457 );
buf ( n40459 , n40458 );
xor ( n40460 , n40353 , n40459 );
xor ( n40461 , n39941 , n40004 );
and ( n40462 , n40461 , n40071 );
and ( n40463 , n39941 , n40004 );
or ( n40464 , n40462 , n40463 );
buf ( n40465 , n40464 );
buf ( n40466 , n40465 );
xor ( n40467 , n40460 , n40466 );
buf ( n40468 , n40467 );
nor ( n40469 , n40347 , n40468 );
not ( n40470 , n40469 );
nand ( n40471 , n40347 , n40468 );
nand ( n40472 , n40470 , n40471 );
not ( n40473 , n40472 );
and ( n40474 , n40342 , n40473 );
not ( n40475 , n40342 );
and ( n40476 , n40475 , n40472 );
nor ( n40477 , n40474 , n40476 );
not ( n40478 , n40477 );
or ( n40479 , n40319 , n40478 );
not ( n40480 , n38272 );
not ( n40481 , n38284 );
nand ( n40482 , n40481 , n39889 , n38274 , n7442 );
nor ( n40483 , n39893 , n40482 );
not ( n40484 , n40483 );
or ( n40485 , n40480 , n40484 );
not ( n40486 , n39560 );
not ( n40487 , n39682 );
not ( n40488 , n39687 );
or ( n40489 , n40487 , n40488 );
nand ( n40490 , n40489 , n39887 );
nor ( n40491 , n40486 , n40490 );
not ( n40492 , n40491 );
nor ( n40493 , n40492 , n39558 );
not ( n40494 , n40493 );
not ( n40495 , n38290 );
or ( n40496 , n40494 , n40495 );
not ( n40497 , n40491 );
not ( n40498 , n39552 );
or ( n40499 , n40497 , n40498 );
not ( n40500 , n40490 );
not ( n40501 , n39689 );
and ( n40502 , n40500 , n40501 );
buf ( n40503 , n39888 );
nor ( n40504 , n40502 , n40503 );
nand ( n40505 , n40499 , n40504 );
not ( n40506 , n40505 );
nand ( n40507 , n40496 , n40506 );
nand ( n40508 , n40485 , n40507 );
xor ( n40509 , n39759 , n39764 );
and ( n40510 , n40509 , n39884 );
and ( n40511 , n39759 , n39764 );
or ( n40512 , n40510 , n40511 );
buf ( n40513 , n40512 );
buf ( n40514 , n40513 );
xor ( n40515 , n39821 , n39836 );
and ( n40516 , n40515 , n39878 );
and ( n40517 , n39821 , n39836 );
or ( n40518 , n40516 , n40517 );
buf ( n40519 , n40518 );
buf ( n40520 , n40519 );
xor ( n40521 , n39771 , n39819 );
and ( n40522 , n40521 , n39881 );
and ( n40523 , n39771 , n39819 );
or ( n40524 , n40522 , n40523 );
buf ( n40525 , n40524 );
buf ( n40526 , n40525 );
xor ( n40527 , n40520 , n40526 );
and ( n40528 , n39587 , n39588 );
buf ( n40529 , n40528 );
buf ( n40530 , n40529 );
buf ( n40531 , n495 );
not ( n40532 , n40531 );
buf ( n40533 , n31271 );
not ( n40534 , n40533 );
or ( n40535 , n40532 , n40534 );
buf ( n40536 , n2411 );
buf ( n40537 , n39807 );
or ( n40538 , n40536 , n40537 );
nand ( n40539 , n40535 , n40538 );
buf ( n40540 , n40539 );
buf ( n40541 , n40540 );
xor ( n40542 , n40530 , n40541 );
buf ( n40543 , n39850 );
not ( n40544 , n40543 );
buf ( n40545 , n38410 );
not ( n40546 , n40545 );
or ( n40547 , n40544 , n40546 );
buf ( n40548 , n35832 );
buf ( n40549 , n489 );
buf ( n40550 , n510 );
xor ( n40551 , n40549 , n40550 );
buf ( n40552 , n40551 );
buf ( n40553 , n40552 );
nand ( n40554 , n40548 , n40553 );
buf ( n40555 , n40554 );
buf ( n40556 , n40555 );
nand ( n40557 , n40547 , n40556 );
buf ( n40558 , n40557 );
buf ( n40559 , n40558 );
xor ( n40560 , n40542 , n40559 );
buf ( n40561 , n40560 );
buf ( n40562 , n40561 );
xor ( n40563 , n39780 , n39797 );
and ( n40564 , n40563 , n39816 );
and ( n40565 , n39780 , n39797 );
or ( n40566 , n40564 , n40565 );
buf ( n40567 , n40566 );
buf ( n40568 , n40567 );
xor ( n40569 , n40562 , n40568 );
buf ( n40570 , n39790 );
not ( n40571 , n40570 );
buf ( n40572 , n33438 );
not ( n40573 , n40572 );
or ( n40574 , n40571 , n40573 );
buf ( n40575 , n4519 );
buf ( n40576 , n508 );
buf ( n40577 , n491 );
xor ( n40578 , n40576 , n40577 );
buf ( n40579 , n40578 );
buf ( n40580 , n40579 );
nand ( n40581 , n40575 , n40580 );
buf ( n40582 , n40581 );
buf ( n40583 , n40582 );
nand ( n40584 , n40574 , n40583 );
buf ( n40585 , n40584 );
buf ( n40586 , n40585 );
buf ( n40587 , n39868 );
not ( n40588 , n40587 );
buf ( n40589 , n31660 );
not ( n40590 , n40589 );
or ( n40591 , n40588 , n40590 );
buf ( n40592 , n2591 );
buf ( n40593 , n493 );
buf ( n40594 , n506 );
xor ( n40595 , n40593 , n40594 );
buf ( n40596 , n40595 );
buf ( n40597 , n40596 );
nand ( n40598 , n40592 , n40597 );
buf ( n40599 , n40598 );
buf ( n40600 , n40599 );
nand ( n40601 , n40591 , n40600 );
buf ( n40602 , n40601 );
buf ( n40603 , n40602 );
not ( n40604 , n40603 );
buf ( n40605 , n40604 );
buf ( n40606 , n40605 );
xor ( n40607 , n40586 , n40606 );
xor ( n40608 , n39840 , n39857 );
and ( n40609 , n40608 , n39875 );
and ( n40610 , n39840 , n39857 );
or ( n40611 , n40609 , n40610 );
buf ( n40612 , n40611 );
buf ( n40613 , n40612 );
xor ( n40614 , n40607 , n40613 );
buf ( n40615 , n40614 );
buf ( n40616 , n40615 );
xor ( n40617 , n40569 , n40616 );
buf ( n40618 , n40617 );
buf ( n40619 , n40618 );
xor ( n40620 , n40527 , n40619 );
buf ( n40621 , n40620 );
nor ( n40622 , n40514 , n40621 );
not ( n40623 , n40622 );
nand ( n40624 , n40513 , n40621 );
nand ( n40625 , n40623 , n40624 );
not ( n40626 , n40625 );
and ( n40627 , n40508 , n40626 );
not ( n40628 , n40508 );
and ( n40629 , n40628 , n40625 );
nor ( n40630 , n40627 , n40629 );
nand ( n40631 , n40630 , n2815 );
nand ( n40632 , n40479 , n40631 );
not ( n40633 , n40632 );
or ( n40634 , n40318 , n40633 );
xor ( n40635 , n40214 , n40245 );
and ( n40636 , n40635 , n40252 );
and ( n40637 , n40214 , n40245 );
or ( n40638 , n40636 , n40637 );
buf ( n40639 , n40638 );
not ( n40640 , n40639 );
xor ( n40641 , n40114 , n40133 );
xor ( n40642 , n40641 , n40150 );
and ( n40643 , n40193 , n40642 );
xor ( n40644 , n40114 , n40133 );
xor ( n40645 , n40644 , n40150 );
and ( n40646 , n40198 , n40645 );
and ( n40647 , n40193 , n40198 );
or ( n40648 , n40643 , n40646 , n40647 );
not ( n40649 , n40648 );
xor ( n40650 , n40220 , n40235 );
and ( n40651 , n40650 , n40242 );
and ( n40652 , n40220 , n40235 );
or ( n40653 , n40651 , n40652 );
buf ( n40654 , n40653 );
buf ( n40655 , n40654 );
buf ( n40656 , n40231 );
buf ( n40657 , n6541 );
buf ( n40658 , n31840 );
nor ( n40659 , n40657 , n40658 );
buf ( n40660 , n40659 );
buf ( n40661 , n40660 );
xor ( n40662 , n40656 , n40661 );
xor ( n40663 , n40114 , n40133 );
and ( n40664 , n40663 , n40150 );
and ( n40665 , n40114 , n40133 );
or ( n40666 , n40664 , n40665 );
buf ( n40667 , n40666 );
xor ( n40668 , n40662 , n40667 );
buf ( n40669 , n40668 );
buf ( n40670 , n40669 );
xor ( n40671 , n40655 , n40670 );
buf ( n40672 , n6015 );
buf ( n40673 , n40110 );
or ( n40674 , n40672 , n40673 );
buf ( n40675 , n6010 );
buf ( n40676 , n6001 );
buf ( n40677 , n527 );
and ( n40678 , n40676 , n40677 );
buf ( n40679 , n33009 );
buf ( n40680 , n539 );
and ( n40681 , n40679 , n40680 );
nor ( n40682 , n40678 , n40681 );
buf ( n40683 , n40682 );
buf ( n40684 , n40683 );
or ( n40685 , n40675 , n40684 );
nand ( n40686 , n40674 , n40685 );
buf ( n40687 , n40686 );
buf ( n40688 , n40687 );
buf ( n40689 , n4030 );
buf ( n40690 , n40186 );
or ( n40691 , n40689 , n40690 );
buf ( n40692 , n4040 );
buf ( n40693 , n523 );
buf ( n40694 , n32981 );
and ( n40695 , n40693 , n40694 );
not ( n40696 , n40693 );
buf ( n40697 , n543 );
and ( n40698 , n40696 , n40697 );
nor ( n40699 , n40695 , n40698 );
buf ( n40700 , n40699 );
buf ( n40701 , n40700 );
or ( n40702 , n40692 , n40701 );
nand ( n40703 , n40691 , n40702 );
buf ( n40704 , n40703 );
buf ( n40705 , n40704 );
xor ( n40706 , n40688 , n40705 );
buf ( n40707 , n38773 );
buf ( n40708 , n40163 );
or ( n40709 , n40707 , n40708 );
buf ( n40710 , n6337 );
buf ( n40711 , n6541 );
buf ( n40712 , n529 );
and ( n40713 , n40711 , n40712 );
buf ( n40714 , n2969 );
buf ( n40715 , n537 );
and ( n40716 , n40714 , n40715 );
nor ( n40717 , n40713 , n40716 );
buf ( n40718 , n40717 );
buf ( n40719 , n40718 );
or ( n40720 , n40710 , n40719 );
nand ( n40721 , n40709 , n40720 );
buf ( n40722 , n40721 );
buf ( n40723 , n40722 );
xor ( n40724 , n40706 , n40723 );
buf ( n40725 , n40724 );
buf ( n40726 , n40725 );
xor ( n40727 , n40168 , n40173 );
and ( n40728 , n40727 , n40191 );
and ( n40729 , n40168 , n40173 );
or ( n40730 , n40728 , n40729 );
buf ( n40731 , n40730 );
buf ( n40732 , n40731 );
xor ( n40733 , n40726 , n40732 );
buf ( n40734 , n31978 );
not ( n40735 , n40734 );
buf ( n40736 , n3020 );
not ( n40737 , n40736 );
or ( n40738 , n40735 , n40737 );
buf ( n40739 , n547 );
nand ( n40740 , n40738 , n40739 );
buf ( n40741 , n40740 );
buf ( n40742 , n40741 );
buf ( n40743 , n5582 );
buf ( n40744 , n40129 );
or ( n40745 , n40743 , n40744 );
buf ( n40746 , n33118 );
buf ( n40747 , n541 );
buf ( n40748 , n34557 );
and ( n40749 , n40747 , n40748 );
not ( n40750 , n40747 );
buf ( n40751 , n525 );
and ( n40752 , n40750 , n40751 );
nor ( n40753 , n40749 , n40752 );
buf ( n40754 , n40753 );
buf ( n40755 , n40754 );
or ( n40756 , n40746 , n40755 );
nand ( n40757 , n40745 , n40756 );
buf ( n40758 , n40757 );
buf ( n40759 , n40758 );
xor ( n40760 , n40742 , n40759 );
buf ( n40761 , n3069 );
buf ( n40762 , n40146 );
or ( n40763 , n40761 , n40762 );
buf ( n40764 , n3087 );
buf ( n40765 , n32053 );
buf ( n40766 , n521 );
and ( n40767 , n40765 , n40766 );
buf ( n40768 , n35343 );
buf ( n40769 , n545 );
and ( n40770 , n40768 , n40769 );
nor ( n40771 , n40767 , n40770 );
buf ( n40772 , n40771 );
buf ( n40773 , n40772 );
or ( n40774 , n40764 , n40773 );
nand ( n40775 , n40763 , n40774 );
buf ( n40776 , n40775 );
buf ( n40777 , n40776 );
xor ( n40778 , n40760 , n40777 );
buf ( n40779 , n40778 );
buf ( n40780 , n40779 );
xor ( n40781 , n40733 , n40780 );
buf ( n40782 , n40781 );
buf ( n40783 , n40782 );
xor ( n40784 , n40671 , n40783 );
buf ( n40785 , n40784 );
not ( n40786 , n40785 );
not ( n40787 , n40786 );
and ( n40788 , n40649 , n40787 );
not ( n40789 , n40649 );
and ( n40790 , n40789 , n40786 );
nor ( n40791 , n40788 , n40790 );
nand ( n40792 , n40640 , n40791 );
not ( n40793 , n40791 );
nand ( n40794 , n40793 , n40639 );
nand ( n40795 , n40792 , n40794 , n3138 );
not ( n40796 , n40795 );
xor ( n40797 , n40201 , n40207 );
and ( n40798 , n40797 , n40255 );
and ( n40799 , n40201 , n40207 );
or ( n40800 , n40798 , n40799 );
buf ( n40801 , n40800 );
and ( n40802 , n40801 , n3360 );
nor ( n40803 , n40796 , n40802 );
nand ( n40804 , n40634 , n40803 );
not ( n40805 , n40795 );
not ( n40806 , n40805 );
not ( n40807 , n40806 );
nand ( n40808 , n40632 , n454 );
not ( n40809 , n40808 );
or ( n40810 , n40807 , n40809 );
nand ( n40811 , n40810 , n40802 );
nand ( n40812 , n40804 , n40811 );
and ( n40813 , n40317 , n40812 );
not ( n40814 , n40317 );
not ( n40815 , n40812 );
and ( n40816 , n40814 , n40815 );
nor ( n40817 , n40813 , n40816 );
not ( n40818 , n37402 );
buf ( n40819 , n5860 );
buf ( n40820 , n3827 );
nand ( n40821 , n40818 , n40819 , n40820 );
nand ( n40822 , n5889 , n5880 , n5886 );
or ( n40823 , n37355 , n37341 );
or ( n40824 , n37383 , n37415 );
nand ( n40825 , n40822 , n40823 , n40824 );
not ( n40826 , n37417 );
not ( n40827 , n37409 );
or ( n40828 , n40826 , n40827 );
nand ( n40829 , n40828 , n37423 );
not ( n40830 , n40829 );
nand ( n40831 , n40821 , n40825 , n40830 );
not ( n40832 , n37430 );
nand ( n40833 , n5774 , n37236 );
not ( n40834 , n37221 );
nand ( n40835 , n40832 , n40833 , n40834 );
nand ( n40836 , n40835 , n37433 );
not ( n40837 , n40836 );
and ( n40838 , n40831 , n40837 );
not ( n40839 , n40831 );
and ( n40840 , n40839 , n40836 );
nor ( n40841 , n40838 , n40840 );
nor ( n40842 , n37341 , n37355 );
not ( n40843 , n40842 );
nand ( n40844 , n40843 , n37423 );
not ( n40845 , n40844 );
nor ( n40846 , n37415 , n37383 );
not ( n40847 , n40846 );
buf ( n40848 , n5890 );
nand ( n40849 , n40847 , n40848 );
nor ( n40850 , n40846 , n3830 );
nand ( n40851 , n40819 , n40850 );
not ( n40852 , n37417 );
nand ( n40853 , n40849 , n40851 , n40852 );
not ( n40854 , n40853 );
or ( n40855 , n40845 , n40854 );
buf ( n40856 , n37417 );
nor ( n40857 , n40856 , n40844 );
nand ( n40858 , n40849 , n40857 , n40851 );
nand ( n40859 , n40855 , n40858 );
nand ( n40860 , n40841 , n40859 );
not ( n40861 , n40860 );
nand ( n40862 , n37212 , n6636 );
nand ( n40863 , n37439 , n40862 );
not ( n40864 , n40863 );
and ( n40865 , n37403 , n40835 );
nand ( n40866 , n40865 , n40819 , n40820 );
not ( n40867 , n40835 );
not ( n40868 , n40829 );
or ( n40869 , n40867 , n40868 );
buf ( n40870 , n37433 );
nand ( n40871 , n40869 , n40870 );
not ( n40872 , n40871 );
nand ( n40873 , n40865 , n40848 );
nand ( n40874 , n40866 , n40872 , n40873 );
not ( n40875 , n40874 );
or ( n40876 , n40864 , n40875 );
not ( n40877 , n40863 );
nand ( n40878 , n40866 , n40873 , n40872 , n40877 );
nand ( n40879 , n40876 , n40878 );
nand ( n40880 , n40861 , n40879 );
nand ( n40881 , n3891 , n3833 , n3860 );
nand ( n40882 , n3899 , n3833 );
nand ( n40883 , n40881 , n40882 , n3834 );
not ( n40884 , n5859 );
not ( n40885 , n3827 );
or ( n40886 , n40884 , n40885 );
buf ( n40887 , n5879 );
not ( n40888 , n40887 );
nand ( n40889 , n40886 , n40888 );
nand ( n40890 , n5815 , n5884 );
not ( n40891 , n40890 );
and ( n40892 , n40889 , n40891 );
not ( n40893 , n40889 );
and ( n40894 , n40893 , n40890 );
nor ( n40895 , n40892 , n40894 );
not ( n40896 , n3249 );
not ( n40897 , n3827 );
or ( n40898 , n40896 , n40897 );
buf ( n40899 , n3251 );
nand ( n40900 , n40898 , n40899 );
nand ( n40901 , n5878 , n5857 );
not ( n40902 , n40901 );
and ( n40903 , n40900 , n40902 );
not ( n40904 , n40900 );
and ( n40905 , n40904 , n40901 );
nor ( n40906 , n40903 , n40905 );
nand ( n40907 , n40895 , n40906 );
not ( n40908 , n40907 );
nor ( n40909 , n40846 , n37417 );
not ( n40910 , n40909 );
not ( n40911 , n5892 );
not ( n40912 , n40911 );
or ( n40913 , n40910 , n40912 );
not ( n40914 , n40909 );
not ( n40915 , n40911 );
nand ( n40916 , n40914 , n40915 );
nand ( n40917 , n40913 , n40916 );
and ( n40918 , n5815 , n5859 );
not ( n40919 , n40918 );
not ( n40920 , n3827 );
or ( n40921 , n40919 , n40920 );
buf ( n40922 , n5815 );
and ( n40923 , n40887 , n40922 );
nor ( n40924 , n40923 , n5885 );
nand ( n40925 , n40921 , n40924 );
nand ( n40926 , n5743 , n5889 );
not ( n40927 , n40926 );
and ( n40928 , n40925 , n40927 );
not ( n40929 , n40925 );
and ( n40930 , n40929 , n40926 );
nor ( n40931 , n40928 , n40930 );
not ( n40932 , n40931 );
not ( n40933 , n40932 );
nand ( n40934 , n40883 , n40908 , n40917 , n40933 );
nor ( n40935 , n40880 , n40934 );
not ( n40936 , n37441 );
not ( n40937 , n40936 );
not ( n40938 , n38080 );
buf ( n40939 , n40274 );
nand ( n40940 , n40938 , n40939 );
not ( n40941 , n40940 );
not ( n40942 , n40941 );
or ( n40943 , n40937 , n40942 );
nand ( n40944 , n40940 , n37441 );
nand ( n40945 , n40943 , n40944 );
nand ( n40946 , n40935 , n40945 );
not ( n40947 , n454 );
not ( n40948 , n39734 );
or ( n40949 , n40947 , n40948 );
not ( n40950 , n39745 );
nand ( n40951 , n40949 , n40950 );
nand ( n40952 , n40938 , n40951 , n38656 );
not ( n40953 , n40952 );
not ( n40954 , n37289 );
not ( n40955 , n40862 );
or ( n40956 , n40954 , n40955 );
nand ( n40957 , n40956 , n37439 );
and ( n40958 , n40957 , n40303 );
not ( n40959 , n37403 );
not ( n40960 , n5892 );
or ( n40961 , n40959 , n40960 );
not ( n40962 , n37439 );
nand ( n40963 , n37418 , n37433 , n37423 );
nor ( n40964 , n40962 , n40963 );
nand ( n40965 , n40961 , n40964 );
nand ( n40966 , n40953 , n40958 , n40965 );
not ( n40967 , n40269 );
not ( n40968 , n40282 );
or ( n40969 , n40967 , n40968 );
nand ( n40970 , n40969 , n40311 );
not ( n40971 , n40970 );
nand ( n40972 , n40966 , n40971 );
not ( n40973 , n40315 );
nand ( n40974 , n40973 , n40259 );
not ( n40975 , n40974 );
and ( n40976 , n40972 , n40975 );
not ( n40977 , n40972 );
and ( n40978 , n40977 , n40974 );
nor ( n40979 , n40976 , n40978 );
not ( n40980 , n40310 );
nand ( n40981 , n40980 , n40303 );
not ( n40982 , n40981 );
not ( n40983 , n40952 );
buf ( n40984 , n40957 );
nand ( n40985 , n40983 , n40965 , n40984 );
not ( n40986 , n40282 );
not ( n40987 , n40951 );
or ( n40988 , n40986 , n40987 );
buf ( n40989 , n40301 );
nand ( n40990 , n40988 , n40989 );
not ( n40991 , n40990 );
nand ( n40992 , n40985 , n40991 );
not ( n40993 , n40992 );
or ( n40994 , n40982 , n40993 );
not ( n40995 , n40981 );
nand ( n40996 , n40985 , n40995 , n40991 );
nand ( n40997 , n40994 , n40996 );
nor ( n40998 , n38655 , n38080 );
and ( n40999 , n40998 , n40957 );
not ( n41000 , n40999 );
not ( n41001 , n40965 );
or ( n41002 , n41000 , n41001 );
or ( n41003 , n40274 , n40275 );
nand ( n41004 , n41003 , n40281 );
not ( n41005 , n41004 );
nand ( n41006 , n41002 , n41005 );
nand ( n41007 , n40301 , n40951 );
not ( n41008 , n41007 );
and ( n41009 , n41006 , n41008 );
not ( n41010 , n41006 );
and ( n41011 , n41010 , n41007 );
nor ( n41012 , n41009 , n41011 );
not ( n41013 , n40939 );
not ( n41014 , n40275 );
nand ( n41015 , n41014 , n40281 );
nor ( n41016 , n41013 , n41015 );
not ( n41017 , n41016 );
and ( n41018 , n40957 , n40938 );
nand ( n41019 , n41018 , n40965 );
not ( n41020 , n41019 );
or ( n41021 , n41017 , n41020 );
not ( n41022 , n40939 );
not ( n41023 , n41019 );
or ( n41024 , n41022 , n41023 );
not ( n41025 , n41015 );
not ( n41026 , n41025 );
nand ( n41027 , n41024 , n41026 );
nand ( n41028 , n41021 , n41027 );
nand ( n41029 , n40979 , n40997 , n41012 , n41028 );
nor ( n41030 , n40946 , n41029 );
buf ( n41031 , n41030 );
not ( n41032 , n41031 );
and ( n41033 , n40817 , n41032 );
not ( n41034 , n40817 );
not ( n41035 , n41032 );
and ( n41036 , n41034 , n41035 );
nor ( n41037 , n41033 , n41036 );
not ( n41038 , n41037 );
or ( n41039 , n3997 , n41038 );
not ( n41040 , n29512 );
and ( n41041 , n497 , n41040 );
not ( n41042 , n497 );
and ( n41043 , n41042 , n29512 );
nor ( n41044 , n41041 , n41043 );
not ( n41045 , n29506 );
not ( n41046 , n41045 );
not ( n41047 , n40377 );
and ( n41048 , n41046 , n41047 );
not ( n41049 , n29506 );
and ( n41050 , n41049 , n40377 );
nor ( n41051 , n41048 , n41050 );
not ( n41052 , n41051 );
not ( n41053 , n41052 );
or ( n41054 , n41044 , n41053 );
not ( n41055 , n29512 );
and ( n41056 , n498 , n41055 );
not ( n41057 , n498 );
and ( n41058 , n41057 , n29512 );
nor ( n41059 , n41056 , n41058 );
not ( n41060 , n41059 );
and ( n41061 , n40377 , n41055 );
not ( n41062 , n40377 );
and ( n41063 , n41062 , n29512 );
or ( n41064 , n41061 , n41063 );
nand ( n41065 , n41051 , n41064 );
not ( n41066 , n41065 );
nand ( n41067 , n41060 , n41066 );
nand ( n41068 , n41054 , n41067 );
not ( n41069 , n1147 );
not ( n41070 , n41069 );
and ( n41071 , n494 , n41070 );
not ( n41072 , n494 );
not ( n41073 , n41070 );
and ( n41074 , n41072 , n41073 );
nor ( n41075 , n41071 , n41074 );
not ( n41076 , n41075 );
not ( n41077 , n41076 );
buf ( n41078 , n1261 );
and ( n41079 , n41078 , n41070 );
not ( n41080 , n41078 );
not ( n41081 , n1147 );
and ( n41082 , n41080 , n41081 );
or ( n41083 , n41079 , n41082 );
xnor ( n41084 , n1261 , n3916 );
nand ( n41085 , n41083 , n41084 );
not ( n41086 , n41085 );
not ( n41087 , n41086 );
or ( n41088 , n41077 , n41087 );
not ( n41089 , n493 );
and ( n41090 , n41073 , n41089 );
and ( n41091 , n41070 , n493 );
nor ( n41092 , n41090 , n41091 );
not ( n41093 , n41084 );
not ( n41094 , n41093 );
or ( n41095 , n41092 , n41094 );
nand ( n41096 , n41088 , n41095 );
xor ( n41097 , n41068 , n41096 );
and ( n41098 , n456 , n459 );
not ( n41099 , n456 );
and ( n41100 , n41099 , n475 );
nor ( n41101 , n41098 , n41100 );
not ( n41102 , n41101 );
not ( n41103 , n41102 );
and ( n41104 , n499 , n41103 );
not ( n41105 , n499 );
and ( n41106 , n41105 , n41102 );
nor ( n41107 , n41104 , n41106 );
not ( n41108 , n5358 );
not ( n41109 , n29512 );
or ( n41110 , n41108 , n41109 );
not ( n41111 , n5358 );
not ( n41112 , n41111 );
or ( n41113 , n29512 , n41112 );
nand ( n41114 , n41110 , n41113 );
buf ( n41115 , n41114 );
or ( n41116 , n41107 , n41115 );
and ( n41117 , n41103 , n500 );
not ( n41118 , n500 );
and ( n41119 , n41102 , n41118 );
nor ( n41120 , n41117 , n41119 );
not ( n41121 , n41120 );
or ( n41122 , n41102 , n41111 );
nand ( n41123 , n41102 , n41111 );
nand ( n41124 , n41122 , n41123 );
nand ( n41125 , n41115 , n41124 );
not ( n41126 , n41125 );
nand ( n41127 , n41121 , n41126 );
nand ( n41128 , n41116 , n41127 );
and ( n41129 , n41097 , n41128 );
and ( n41130 , n41068 , n41096 );
or ( n41131 , n41129 , n41130 );
not ( n41132 , n41086 );
or ( n41133 , n41132 , n41092 );
not ( n41134 , n492 );
buf ( n41135 , n41081 );
and ( n41136 , n41134 , n41135 );
not ( n41137 , n41134 );
not ( n41138 , n41135 );
and ( n41139 , n41137 , n41138 );
nor ( n41140 , n41136 , n41139 );
or ( n41141 , n41140 , n41094 );
nand ( n41142 , n41133 , n41141 );
or ( n41143 , n41125 , n41107 );
and ( n41144 , n498 , n41101 );
not ( n41145 , n498 );
and ( n41146 , n41145 , n41102 );
nor ( n41147 , n41144 , n41146 );
or ( n41148 , n41115 , n41147 );
nand ( n41149 , n41143 , n41148 );
xor ( n41150 , n41142 , n41149 );
xor ( n41151 , n29500 , n41101 );
not ( n41152 , n29500 );
and ( n41153 , n456 , n457 );
not ( n41154 , n456 );
and ( n41155 , n41154 , n473 );
nor ( n41156 , n41153 , n41155 );
not ( n41157 , n41156 );
not ( n41158 , n41157 );
and ( n41159 , n41152 , n41158 );
and ( n41160 , n41157 , n29500 );
nor ( n41161 , n41159 , n41160 );
nand ( n41162 , n41151 , n41161 );
not ( n41163 , n41162 );
not ( n41164 , n41163 );
buf ( n41165 , n41157 );
and ( n41166 , n41165 , n3959 );
not ( n41167 , n41157 );
and ( n41168 , n41167 , n501 );
nor ( n41169 , n41166 , n41168 );
or ( n41170 , n41164 , n41169 );
not ( n41171 , n41151 );
not ( n41172 , n41171 );
and ( n41173 , n41165 , n41118 );
and ( n41174 , n41167 , n500 );
nor ( n41175 , n41173 , n41174 );
or ( n41176 , n41172 , n41175 );
nand ( n41177 , n41170 , n41176 );
xor ( n41178 , n41150 , n41177 );
xor ( n41179 , n41131 , n41178 );
buf ( n41180 , n29658 );
nand ( n41181 , n41180 , n41049 );
not ( n41182 , n41181 );
not ( n41183 , n41180 );
not ( n41184 , n41045 );
nand ( n41185 , n41183 , n41184 );
not ( n41186 , n41185 );
or ( n41187 , n41182 , n41186 );
xnor ( n41188 , n41081 , n41180 );
nand ( n41189 , n41187 , n41188 );
and ( n41190 , n495 , n41049 );
not ( n41191 , n495 );
not ( n41192 , n41049 );
and ( n41193 , n41191 , n41192 );
nor ( n41194 , n41190 , n41193 );
or ( n41195 , n41189 , n41194 );
not ( n41196 , n494 );
and ( n41197 , n41192 , n41196 );
and ( n41198 , n41049 , n494 );
nor ( n41199 , n41197 , n41198 );
not ( n41200 , n41188 );
not ( n41201 , n41200 );
or ( n41202 , n41199 , n41201 );
nand ( n41203 , n41195 , n41202 );
and ( n41204 , n41157 , n502 );
xor ( n41205 , n41203 , n41204 );
not ( n41206 , n41066 );
or ( n41207 , n41206 , n41044 );
not ( n41208 , n496 );
and ( n41209 , n29512 , n41208 );
and ( n41210 , n41040 , n496 );
nor ( n41211 , n41209 , n41210 );
or ( n41212 , n41211 , n41053 );
nand ( n41213 , n41207 , n41212 );
xor ( n41214 , n41205 , n41213 );
xor ( n41215 , n41179 , n41214 );
and ( n41216 , n489 , n3931 );
not ( n41217 , n489 );
and ( n41218 , n41217 , n32891 );
nor ( n41219 , n41216 , n41218 );
not ( n41220 , n3946 );
or ( n41221 , n41219 , n41220 );
not ( n41222 , n32891 );
or ( n41223 , n41222 , n3945 );
nand ( n41224 , n41221 , n41223 );
and ( n41225 , n491 , n3921 );
not ( n41226 , n491 );
and ( n41227 , n41226 , n3916 );
nor ( n41228 , n41225 , n41227 );
or ( n41229 , n3920 , n41228 );
not ( n41230 , n3980 );
and ( n41231 , n36727 , n3916 );
not ( n41232 , n36727 );
and ( n41233 , n41232 , n3921 );
nor ( n41234 , n41231 , n41233 );
or ( n41235 , n41230 , n41234 );
nand ( n41236 , n41229 , n41235 );
xor ( n41237 , n41224 , n41236 );
and ( n41238 , n41134 , n3916 );
not ( n41239 , n41134 );
and ( n41240 , n456 , n467 );
not ( n41241 , n456 );
and ( n41242 , n41241 , n483 );
nor ( n41243 , n41240 , n41242 );
and ( n41244 , n41239 , n41243 );
nor ( n41245 , n41238 , n41244 );
or ( n41246 , n3920 , n41245 );
or ( n41247 , n41230 , n41228 );
nand ( n41248 , n41246 , n41247 );
and ( n41249 , n41157 , n503 );
xor ( n41250 , n41248 , n41249 );
not ( n41251 , n41189 );
not ( n41252 , n41251 );
and ( n41253 , n41208 , n41045 );
not ( n41254 , n41208 );
and ( n41255 , n41254 , n41184 );
nor ( n41256 , n41253 , n41255 );
not ( n41257 , n41256 );
or ( n41258 , n41252 , n41257 );
or ( n41259 , n41194 , n41201 );
nand ( n41260 , n41258 , n41259 );
and ( n41261 , n41250 , n41260 );
and ( n41262 , n41248 , n41249 );
or ( n41263 , n41261 , n41262 );
xor ( n41264 , n41237 , n41263 );
and ( n41265 , n41157 , n3951 );
and ( n41266 , n41156 , n502 );
nor ( n41267 , n41265 , n41266 );
or ( n41268 , n41164 , n41267 );
or ( n41269 , n41169 , n41172 );
nand ( n41270 , n41268 , n41269 );
and ( n41271 , n490 , n32891 );
not ( n41272 , n490 );
and ( n41273 , n41272 , n41222 );
nor ( n41274 , n41271 , n41273 );
not ( n41275 , n41274 );
or ( n41276 , n41275 , n41220 );
or ( n41277 , n41219 , n3945 );
nand ( n41278 , n41276 , n41277 );
xor ( n41279 , n41270 , n41278 );
not ( n41280 , n41165 );
not ( n41281 , n504 );
nor ( n41282 , n41280 , n41281 );
not ( n41283 , n3944 );
not ( n41284 , n41274 );
or ( n41285 , n41283 , n41284 );
and ( n41286 , n491 , n1405 );
not ( n41287 , n491 );
and ( n41288 , n41287 , n41222 );
nor ( n41289 , n41286 , n41288 );
nand ( n41290 , n41289 , n3946 );
nand ( n41291 , n41285 , n41290 );
xor ( n41292 , n41282 , n41291 );
and ( n41293 , n41089 , n3916 );
not ( n41294 , n41089 );
and ( n41295 , n41294 , n3921 );
nor ( n41296 , n41293 , n41295 );
or ( n41297 , n3920 , n41296 );
or ( n41298 , n41230 , n41245 );
nand ( n41299 , n41297 , n41298 );
and ( n41300 , n41292 , n41299 );
and ( n41301 , n41282 , n41291 );
or ( n41302 , n41300 , n41301 );
and ( n41303 , n41279 , n41302 );
and ( n41304 , n41270 , n41278 );
or ( n41305 , n41303 , n41304 );
xor ( n41306 , n41264 , n41305 );
and ( n41307 , n497 , n41192 );
not ( n41308 , n497 );
and ( n41309 , n41308 , n41045 );
nor ( n41310 , n41307 , n41309 );
not ( n41311 , n41310 );
and ( n41312 , n41181 , n41185 );
nor ( n41313 , n41312 , n41200 );
not ( n41314 , n41313 );
or ( n41315 , n41311 , n41314 );
nand ( n41316 , n41256 , n41200 );
nand ( n41317 , n41315 , n41316 );
not ( n41318 , n41065 );
not ( n41319 , n41318 );
and ( n41320 , n29596 , n29512 );
not ( n41321 , n29596 );
and ( n41322 , n41321 , n41040 );
nor ( n41323 , n41320 , n41322 );
or ( n41324 , n41319 , n41323 );
or ( n41325 , n41059 , n41053 );
nand ( n41326 , n41324 , n41325 );
xor ( n41327 , n41317 , n41326 );
not ( n41328 , n495 );
and ( n41329 , n41135 , n41328 );
and ( n41330 , n41070 , n495 );
nor ( n41331 , n41329 , n41330 );
or ( n41332 , n41132 , n41331 );
or ( n41333 , n41094 , n41075 );
nand ( n41334 , n41332 , n41333 );
and ( n41335 , n41327 , n41334 );
and ( n41336 , n41317 , n41326 );
or ( n41337 , n41335 , n41336 );
xor ( n41338 , n41068 , n41096 );
xor ( n41339 , n41338 , n41128 );
xor ( n41340 , n41337 , n41339 );
xor ( n41341 , n41248 , n41249 );
xor ( n41342 , n41341 , n41260 );
and ( n41343 , n41340 , n41342 );
and ( n41344 , n41337 , n41339 );
or ( n41345 , n41343 , n41344 );
xor ( n41346 , n41306 , n41345 );
xor ( n41347 , n41215 , n41346 );
not ( n41348 , n41126 );
and ( n41349 , n501 , n41103 );
not ( n41350 , n501 );
and ( n41351 , n41350 , n41102 );
nor ( n41352 , n41349 , n41351 );
not ( n41353 , n41352 );
not ( n41354 , n41353 );
or ( n41355 , n41348 , n41354 );
or ( n41356 , n41120 , n41115 );
nand ( n41357 , n41355 , n41356 );
and ( n41358 , n41157 , n32922 );
and ( n41359 , n41156 , n503 );
nor ( n41360 , n41358 , n41359 );
or ( n41361 , n41164 , n41360 );
or ( n41362 , n41267 , n41172 );
nand ( n41363 , n41361 , n41362 );
xor ( n41364 , n41357 , n41363 );
or ( n41365 , n41102 , n29500 );
nand ( n41366 , n41365 , n504 );
nand ( n41367 , n41102 , n29500 );
and ( n41368 , n41366 , n41367 , n41157 );
not ( n41369 , n3944 );
not ( n41370 , n41289 );
or ( n41371 , n41369 , n41370 );
not ( n41372 , n492 );
not ( n41373 , n3931 );
or ( n41374 , n41372 , n41373 );
nand ( n41375 , n32891 , n41134 );
nand ( n41376 , n41374 , n41375 );
nand ( n41377 , n3946 , n41376 );
nand ( n41378 , n41371 , n41377 );
and ( n41379 , n41368 , n41378 );
and ( n41380 , n41364 , n41379 );
and ( n41381 , n41357 , n41363 );
or ( n41382 , n41380 , n41381 );
xor ( n41383 , n41270 , n41278 );
xor ( n41384 , n41383 , n41302 );
xor ( n41385 , n41382 , n41384 );
not ( n41386 , n494 );
not ( n41387 , n3921 );
or ( n41388 , n41386 , n41387 );
not ( n41389 , n41243 );
nand ( n41390 , n41389 , n41196 );
nand ( n41391 , n41388 , n41390 );
not ( n41392 , n41391 );
or ( n41393 , n3920 , n41392 );
or ( n41394 , n41230 , n41296 );
nand ( n41395 , n41393 , n41394 );
and ( n41396 , n498 , n41045 );
not ( n41397 , n498 );
and ( n41398 , n41397 , n41192 );
nor ( n41399 , n41396 , n41398 );
or ( n41400 , n41252 , n41399 );
not ( n41401 , n41310 );
or ( n41402 , n41201 , n41401 );
nand ( n41403 , n41400 , n41402 );
xor ( n41404 , n41395 , n41403 );
and ( n41405 , n41118 , n41055 );
not ( n41406 , n41118 );
and ( n41407 , n41406 , n29512 );
nor ( n41408 , n41405 , n41407 );
not ( n41409 , n41408 );
or ( n41410 , n41206 , n41409 );
or ( n41411 , n41323 , n41053 );
nand ( n41412 , n41410 , n41411 );
and ( n41413 , n41404 , n41412 );
and ( n41414 , n41395 , n41403 );
or ( n41415 , n41413 , n41414 );
and ( n41416 , n41135 , n41208 );
and ( n41417 , n41070 , n496 );
nor ( n41418 , n41416 , n41417 );
or ( n41419 , n41132 , n41418 );
or ( n41420 , n41084 , n41331 );
nand ( n41421 , n41419 , n41420 );
and ( n41422 , n502 , n41101 );
not ( n41423 , n502 );
and ( n41424 , n41423 , n41102 );
nor ( n41425 , n41422 , n41424 );
or ( n41426 , n41125 , n41425 );
or ( n41427 , n41352 , n41115 );
nand ( n41428 , n41426 , n41427 );
xor ( n41429 , n41421 , n41428 );
and ( n41430 , n41157 , n41281 );
and ( n41431 , n41167 , n504 );
nor ( n41432 , n41430 , n41431 );
or ( n41433 , n41164 , n41432 );
or ( n41434 , n41360 , n41172 );
nand ( n41435 , n41433 , n41434 );
and ( n41436 , n41429 , n41435 );
and ( n41437 , n41421 , n41428 );
or ( n41438 , n41436 , n41437 );
xor ( n41439 , n41415 , n41438 );
xor ( n41440 , n41282 , n41291 );
xor ( n41441 , n41440 , n41299 );
and ( n41442 , n41439 , n41441 );
and ( n41443 , n41415 , n41438 );
or ( n41444 , n41442 , n41443 );
and ( n41445 , n41385 , n41444 );
and ( n41446 , n41382 , n41384 );
or ( n41447 , n41445 , n41446 );
xor ( n41448 , n41347 , n41447 );
xor ( n41449 , n41337 , n41339 );
xor ( n41450 , n41449 , n41342 );
xor ( n41451 , n41317 , n41326 );
xor ( n41452 , n41451 , n41334 );
xor ( n41453 , n41357 , n41363 );
xor ( n41454 , n41453 , n41379 );
xor ( n41455 , n41452 , n41454 );
xor ( n41456 , n41368 , n41378 );
and ( n41457 , n41171 , n504 );
and ( n41458 , n495 , n3916 );
not ( n41459 , n495 );
and ( n41460 , n41459 , n41243 );
nor ( n41461 , n41458 , n41460 );
not ( n41462 , n41461 );
and ( n41463 , n3908 , n3919 );
not ( n41464 , n41463 );
or ( n41465 , n41462 , n41464 );
nand ( n41466 , n41391 , n3980 );
nand ( n41467 , n41465 , n41466 );
xor ( n41468 , n41457 , n41467 );
and ( n41469 , n499 , n41049 );
not ( n41470 , n499 );
and ( n41471 , n41470 , n41192 );
nor ( n41472 , n41469 , n41471 );
or ( n41473 , n41252 , n41472 );
or ( n41474 , n41399 , n41201 );
nand ( n41475 , n41473 , n41474 );
and ( n41476 , n41468 , n41475 );
and ( n41477 , n41457 , n41467 );
or ( n41478 , n41476 , n41477 );
xor ( n41479 , n41456 , n41478 );
and ( n41480 , n3959 , n41055 );
not ( n41481 , n3959 );
and ( n41482 , n41481 , n29512 );
nor ( n41483 , n41480 , n41482 );
not ( n41484 , n41483 );
not ( n41485 , n41066 );
or ( n41486 , n41484 , n41485 );
nand ( n41487 , n41408 , n41052 );
nand ( n41488 , n41486 , n41487 );
not ( n41489 , n3946 );
xor ( n41490 , n41089 , n41222 );
not ( n41491 , n41490 );
or ( n41492 , n41489 , n41491 );
nand ( n41493 , n41376 , n3944 );
nand ( n41494 , n41492 , n41493 );
xor ( n41495 , n41488 , n41494 );
and ( n41496 , n41102 , n32922 );
not ( n41497 , n41102 );
and ( n41498 , n41497 , n503 );
nor ( n41499 , n41496 , n41498 );
or ( n41500 , n41125 , n41499 );
or ( n41501 , n41425 , n41115 );
nand ( n41502 , n41500 , n41501 );
and ( n41503 , n41495 , n41502 );
and ( n41504 , n41488 , n41494 );
or ( n41505 , n41503 , n41504 );
and ( n41506 , n41479 , n41505 );
and ( n41507 , n41456 , n41478 );
or ( n41508 , n41506 , n41507 );
and ( n41509 , n41455 , n41508 );
and ( n41510 , n41452 , n41454 );
or ( n41511 , n41509 , n41510 );
xor ( n41512 , n41450 , n41511 );
xor ( n41513 , n41382 , n41384 );
xor ( n41514 , n41513 , n41444 );
and ( n41515 , n41512 , n41514 );
and ( n41516 , n41450 , n41511 );
or ( n41517 , n41515 , n41516 );
nor ( n41518 , n41448 , n41517 );
and ( n41519 , n41448 , n41517 );
or ( n41520 , n41518 , n41519 );
not ( n41521 , n41520 );
xor ( n41522 , n41415 , n41438 );
xor ( n41523 , n41522 , n41441 );
xor ( n41524 , n41452 , n41454 );
xor ( n41525 , n41524 , n41508 );
xor ( n41526 , n41523 , n41525 );
xor ( n41527 , n41421 , n41428 );
xor ( n41528 , n41527 , n41435 );
xor ( n41529 , n41395 , n41403 );
xor ( n41530 , n41529 , n41412 );
xor ( n41531 , n41528 , n41530 );
not ( n41532 , n497 );
and ( n41533 , n41135 , n41532 );
and ( n41534 , n41138 , n497 );
nor ( n41535 , n41533 , n41534 );
or ( n41536 , n41535 , n41085 );
or ( n41537 , n41094 , n41418 );
nand ( n41538 , n41536 , n41537 );
or ( n41539 , n29512 , n41112 );
nand ( n41540 , n41539 , n504 );
nand ( n41541 , n29512 , n41112 );
and ( n41542 , n41540 , n41541 , n41102 );
and ( n41543 , n496 , n3916 );
not ( n41544 , n496 );
and ( n41545 , n41544 , n41243 );
nor ( n41546 , n41543 , n41545 );
not ( n41547 , n41546 );
not ( n41548 , n41463 );
or ( n41549 , n41547 , n41548 );
nand ( n41550 , n41461 , n3980 );
nand ( n41551 , n41549 , n41550 );
and ( n41552 , n41542 , n41551 );
xor ( n41553 , n41538 , n41552 );
and ( n41554 , n41118 , n41192 );
not ( n41555 , n41118 );
and ( n41556 , n41555 , n41049 );
nor ( n41557 , n41554 , n41556 );
or ( n41558 , n41189 , n41557 );
or ( n41559 , n41472 , n41188 );
nand ( n41560 , n41558 , n41559 );
and ( n41561 , n3951 , n29512 );
not ( n41562 , n3951 );
and ( n41563 , n41562 , n41040 );
nor ( n41564 , n41561 , n41563 );
or ( n41565 , n41319 , n41564 );
not ( n41566 , n41483 );
or ( n41567 , n41566 , n41053 );
nand ( n41568 , n41565 , n41567 );
xor ( n41569 , n41560 , n41568 );
not ( n41570 , n3944 );
not ( n41571 , n41490 );
or ( n41572 , n41570 , n41571 );
not ( n41573 , n32891 );
not ( n41574 , n41196 );
and ( n41575 , n41573 , n41574 );
and ( n41576 , n32891 , n41196 );
nor ( n41577 , n41575 , n41576 );
or ( n41578 , n41577 , n41220 );
nand ( n41579 , n41572 , n41578 );
and ( n41580 , n41569 , n41579 );
and ( n41581 , n41560 , n41568 );
or ( n41582 , n41580 , n41581 );
and ( n41583 , n41553 , n41582 );
and ( n41584 , n41538 , n41552 );
or ( n41585 , n41583 , n41584 );
and ( n41586 , n41531 , n41585 );
and ( n41587 , n41528 , n41530 );
or ( n41588 , n41586 , n41587 );
xor ( n41589 , n41526 , n41588 );
xor ( n41590 , n41456 , n41478 );
xor ( n41591 , n41590 , n41505 );
xor ( n41592 , n41488 , n41494 );
xor ( n41593 , n41592 , n41502 );
xor ( n41594 , n41457 , n41467 );
xor ( n41595 , n41594 , n41475 );
xor ( n41596 , n41593 , n41595 );
not ( n41597 , n41126 );
and ( n41598 , n41102 , n41281 );
and ( n41599 , n41103 , n504 );
nor ( n41600 , n41598 , n41599 );
or ( n41601 , n41597 , n41600 );
or ( n41602 , n41115 , n41499 );
nand ( n41603 , n41601 , n41602 );
and ( n41604 , n701 , n41073 );
not ( n41605 , n701 );
and ( n41606 , n41605 , n41070 );
nor ( n41607 , n41604 , n41606 );
or ( n41608 , n41085 , n41607 );
or ( n41609 , n41094 , n41535 );
nand ( n41610 , n41608 , n41609 );
xor ( n41611 , n41603 , n41610 );
xor ( n41612 , n41542 , n41551 );
and ( n41613 , n41611 , n41612 );
and ( n41614 , n41603 , n41610 );
or ( n41615 , n41613 , n41614 );
and ( n41616 , n41596 , n41615 );
and ( n41617 , n41593 , n41595 );
or ( n41618 , n41616 , n41617 );
xor ( n41619 , n41591 , n41618 );
xor ( n41620 , n41528 , n41530 );
xor ( n41621 , n41620 , n41585 );
and ( n41622 , n41619 , n41621 );
and ( n41623 , n41591 , n41618 );
or ( n41624 , n41622 , n41623 );
or ( n41625 , n41589 , n41624 );
xor ( n41626 , n41591 , n41618 );
xor ( n41627 , n41626 , n41621 );
xor ( n41628 , n41538 , n41552 );
xor ( n41629 , n41628 , n41582 );
not ( n41630 , n41115 );
and ( n41631 , n41630 , n504 );
or ( n41632 , n3921 , n497 );
or ( n41633 , n41389 , n41532 );
nand ( n41634 , n41632 , n41633 );
not ( n41635 , n41634 );
not ( n41636 , n41463 );
or ( n41637 , n41635 , n41636 );
nand ( n41638 , n41546 , n3980 );
nand ( n41639 , n41637 , n41638 );
xor ( n41640 , n41631 , n41639 );
and ( n41641 , n3959 , n41049 );
not ( n41642 , n3959 );
and ( n41643 , n41642 , n41192 );
nor ( n41644 , n41641 , n41643 );
not ( n41645 , n41644 );
or ( n41646 , n41189 , n41645 );
or ( n41647 , n41557 , n41201 );
nand ( n41648 , n41646 , n41647 );
and ( n41649 , n41640 , n41648 );
and ( n41650 , n41631 , n41639 );
or ( n41651 , n41649 , n41650 );
and ( n41652 , n503 , n41055 );
not ( n41653 , n503 );
and ( n41654 , n41653 , n29512 );
nor ( n41655 , n41652 , n41654 );
or ( n41656 , n41206 , n41655 );
or ( n41657 , n41564 , n41053 );
nand ( n41658 , n41656 , n41657 );
not ( n41659 , n3944 );
not ( n41660 , n41577 );
not ( n41661 , n41660 );
or ( n41662 , n41659 , n41661 );
and ( n41663 , n495 , n1404 );
not ( n41664 , n495 );
and ( n41665 , n41664 , n32891 );
nor ( n41666 , n41663 , n41665 );
or ( n41667 , n41666 , n41220 );
nand ( n41668 , n41662 , n41667 );
xor ( n41669 , n41658 , n41668 );
and ( n41670 , n41073 , n29596 );
and ( n41671 , n41070 , n499 );
nor ( n41672 , n41670 , n41671 );
or ( n41673 , n41085 , n41672 );
or ( n41674 , n41607 , n41094 );
nand ( n41675 , n41673 , n41674 );
and ( n41676 , n41669 , n41675 );
and ( n41677 , n41658 , n41668 );
or ( n41678 , n41676 , n41677 );
xor ( n41679 , n41651 , n41678 );
xor ( n41680 , n41560 , n41568 );
xor ( n41681 , n41680 , n41579 );
and ( n41682 , n41679 , n41681 );
and ( n41683 , n41651 , n41678 );
or ( n41684 , n41682 , n41683 );
xor ( n41685 , n41629 , n41684 );
xor ( n41686 , n41593 , n41595 );
xor ( n41687 , n41686 , n41615 );
and ( n41688 , n41685 , n41687 );
and ( n41689 , n41629 , n41684 );
or ( n41690 , n41688 , n41689 );
and ( n41691 , n41627 , n41690 );
and ( n41692 , n41625 , n41691 );
and ( n41693 , n41589 , n41624 );
nor ( n41694 , n41692 , n41693 );
not ( n41695 , n3946 );
and ( n41696 , n701 , n1405 );
not ( n41697 , n701 );
and ( n41698 , n41697 , n3931 );
or ( n41699 , n41696 , n41698 );
not ( n41700 , n41699 );
or ( n41701 , n41695 , n41700 );
not ( n41702 , n41532 );
not ( n41703 , n1405 );
or ( n41704 , n41702 , n41703 );
nand ( n41705 , n41222 , n497 );
nand ( n41706 , n41704 , n41705 );
nand ( n41707 , n41706 , n3944 );
nand ( n41708 , n41701 , n41707 );
or ( n41709 , n41073 , n41180 );
nand ( n41710 , n41709 , n504 );
nand ( n41711 , n41135 , n41180 );
and ( n41712 , n41710 , n41711 , n41192 );
xor ( n41713 , n41708 , n41712 );
and ( n41714 , n41200 , n504 );
not ( n41715 , n3944 );
not ( n41716 , n41699 );
or ( n41717 , n41715 , n41716 );
and ( n41718 , n29596 , n1405 );
not ( n41719 , n29596 );
and ( n41720 , n41719 , n41222 );
or ( n41721 , n41718 , n41720 );
nand ( n41722 , n41721 , n3946 );
nand ( n41723 , n41717 , n41722 );
xor ( n41724 , n41714 , n41723 );
and ( n41725 , n3959 , n3916 );
not ( n41726 , n3959 );
and ( n41727 , n41726 , n3921 );
nor ( n41728 , n41725 , n41727 );
or ( n41729 , n3920 , n41728 );
not ( n41730 , n3916 );
not ( n41731 , n41118 );
and ( n41732 , n41730 , n41731 );
and ( n41733 , n3916 , n41118 );
nor ( n41734 , n41732 , n41733 );
or ( n41735 , n41734 , n41230 );
nand ( n41736 , n41729 , n41735 );
and ( n41737 , n41724 , n41736 );
and ( n41738 , n41714 , n41723 );
or ( n41739 , n41737 , n41738 );
xor ( n41740 , n41713 , n41739 );
and ( n41741 , n504 , n41049 );
not ( n41742 , n504 );
and ( n41743 , n41742 , n41184 );
nor ( n41744 , n41741 , n41743 );
or ( n41745 , n41189 , n41744 );
and ( n41746 , n503 , n41049 );
not ( n41747 , n503 );
and ( n41748 , n41747 , n41184 );
nor ( n41749 , n41746 , n41748 );
or ( n41750 , n41749 , n41188 );
nand ( n41751 , n41745 , n41750 );
not ( n41752 , n41734 );
not ( n41753 , n41752 );
not ( n41754 , n41463 );
or ( n41755 , n41753 , n41754 );
and ( n41756 , n499 , n41389 );
not ( n41757 , n499 );
and ( n41758 , n41757 , n3921 );
nor ( n41759 , n41756 , n41758 );
nand ( n41760 , n41759 , n3980 );
nand ( n41761 , n41755 , n41760 );
xor ( n41762 , n41751 , n41761 );
and ( n41763 , n3951 , n41135 );
not ( n41764 , n3951 );
and ( n41765 , n41764 , n41138 );
nor ( n41766 , n41763 , n41765 );
or ( n41767 , n41085 , n41766 );
and ( n41768 , n501 , n41070 );
not ( n41769 , n501 );
and ( n41770 , n41769 , n41073 );
nor ( n41771 , n41768 , n41770 );
or ( n41772 , n41771 , n41084 );
nand ( n41773 , n41767 , n41772 );
xor ( n41774 , n41762 , n41773 );
and ( n41775 , n41740 , n41774 );
and ( n41776 , n41713 , n41739 );
or ( n41777 , n41775 , n41776 );
xor ( n41778 , n41751 , n41761 );
and ( n41779 , n41778 , n41773 );
and ( n41780 , n41751 , n41761 );
or ( n41781 , n41779 , n41780 );
and ( n41782 , n41052 , n504 );
not ( n41783 , n3944 );
and ( n41784 , n41208 , n3931 );
not ( n41785 , n41208 );
and ( n41786 , n41785 , n32891 );
nor ( n41787 , n41784 , n41786 );
not ( n41788 , n41787 );
or ( n41789 , n41783 , n41788 );
nand ( n41790 , n41706 , n3946 );
nand ( n41791 , n41789 , n41790 );
xor ( n41792 , n41782 , n41791 );
not ( n41793 , n41749 );
not ( n41794 , n41793 );
not ( n41795 , n41313 );
or ( n41796 , n41794 , n41795 );
and ( n41797 , n502 , n41184 );
not ( n41798 , n502 );
and ( n41799 , n41798 , n41049 );
nor ( n41800 , n41797 , n41799 );
nand ( n41801 , n41800 , n41200 );
nand ( n41802 , n41796 , n41801 );
xor ( n41803 , n41792 , n41802 );
xor ( n41804 , n41781 , n41803 );
not ( n41805 , n41759 );
or ( n41806 , n3920 , n41805 );
and ( n41807 , n701 , n3916 );
not ( n41808 , n701 );
and ( n41809 , n41808 , n3921 );
nor ( n41810 , n41807 , n41809 );
or ( n41811 , n41230 , n41810 );
nand ( n41812 , n41806 , n41811 );
or ( n41813 , n41132 , n41771 );
and ( n41814 , n41073 , n41118 );
and ( n41815 , n41070 , n500 );
nor ( n41816 , n41814 , n41815 );
or ( n41817 , n41816 , n41094 );
nand ( n41818 , n41813 , n41817 );
xor ( n41819 , n41812 , n41818 );
and ( n41820 , n41708 , n41712 );
xor ( n41821 , n41819 , n41820 );
xor ( n41822 , n41804 , n41821 );
xor ( n41823 , n41777 , n41822 );
and ( n41824 , n41093 , n504 );
and ( n41825 , n3951 , n3921 );
not ( n41826 , n3951 );
and ( n41827 , n41826 , n41389 );
nor ( n41828 , n41825 , n41827 );
not ( n41829 , n41828 );
not ( n41830 , n3980 );
or ( n41831 , n41829 , n41830 );
not ( n41832 , n3927 );
nand ( n41833 , n41832 , n41463 );
nand ( n41834 , n41831 , n41833 );
xor ( n41835 , n41824 , n41834 );
not ( n41836 , n3944 );
not ( n41837 , n500 );
not ( n41838 , n41222 );
or ( n41839 , n41837 , n41838 );
nand ( n41840 , n32891 , n41118 );
nand ( n41841 , n41839 , n41840 );
not ( n41842 , n41841 );
or ( n41843 , n41836 , n41842 );
not ( n41844 , n3961 );
or ( n41845 , n41844 , n41220 );
nand ( n41846 , n41843 , n41845 );
and ( n41847 , n41835 , n41846 );
and ( n41848 , n41824 , n41834 );
or ( n41849 , n41847 , n41848 );
not ( n41850 , n41828 );
or ( n41851 , n3920 , n41850 );
or ( n41852 , n41728 , n41230 );
nand ( n41853 , n41851 , n41852 );
and ( n41854 , n41073 , n41281 );
and ( n41855 , n41070 , n504 );
nor ( n41856 , n41854 , n41855 );
or ( n41857 , n41085 , n41856 );
and ( n41858 , n41135 , n32922 );
and ( n41859 , n41138 , n503 );
nor ( n41860 , n41858 , n41859 );
or ( n41861 , n41860 , n41084 );
nand ( n41862 , n41857 , n41861 );
xor ( n41863 , n41853 , n41862 );
or ( n41864 , n41389 , n41078 );
nand ( n41865 , n41864 , n504 );
nand ( n41866 , n3916 , n41078 );
and ( n41867 , n41865 , n41866 , n41073 );
not ( n41868 , n3944 );
not ( n41869 , n41721 );
or ( n41870 , n41868 , n41869 );
not ( n41871 , n41841 );
or ( n41872 , n41871 , n41220 );
nand ( n41873 , n41870 , n41872 );
xor ( n41874 , n41867 , n41873 );
xor ( n41875 , n41863 , n41874 );
xor ( n41876 , n41849 , n41875 );
and ( n41877 , n3943 , n3963 );
xor ( n41878 , n41824 , n41834 );
xor ( n41879 , n41878 , n41846 );
xor ( n41880 , n41877 , n41879 );
xor ( n41881 , n3929 , n3964 );
and ( n41882 , n41881 , n32940 );
and ( n41883 , n3929 , n3964 );
or ( n41884 , n41882 , n41883 );
and ( n41885 , n41880 , n41884 );
and ( n41886 , n41877 , n41879 );
or ( n41887 , n41885 , n41886 );
and ( n41888 , n41876 , n41887 );
and ( n41889 , n41849 , n41875 );
or ( n41890 , n41888 , n41889 );
or ( n41891 , n41132 , n41860 );
or ( n41892 , n41766 , n41094 );
nand ( n41893 , n41891 , n41892 );
and ( n41894 , n41867 , n41873 );
xor ( n41895 , n41893 , n41894 );
xor ( n41896 , n41714 , n41723 );
xor ( n41897 , n41896 , n41736 );
xor ( n41898 , n41895 , n41897 );
xor ( n41899 , n41853 , n41862 );
and ( n41900 , n41899 , n41874 );
and ( n41901 , n41853 , n41862 );
or ( n41902 , n41900 , n41901 );
or ( n41903 , n41898 , n41902 );
nand ( n41904 , n41890 , n41903 );
xor ( n41905 , n41713 , n41739 );
xor ( n41906 , n41905 , n41774 );
xor ( n41907 , n41893 , n41894 );
and ( n41908 , n41907 , n41897 );
and ( n41909 , n41893 , n41894 );
or ( n41910 , n41908 , n41909 );
nor ( n41911 , n41906 , n41910 );
or ( n41912 , n41904 , n41911 );
not ( n41913 , n41911 );
nand ( n41914 , n41898 , n41902 );
not ( n41915 , n41914 );
and ( n41916 , n41913 , n41915 );
and ( n41917 , n41906 , n41910 );
nor ( n41918 , n41916 , n41917 );
nand ( n41919 , n41912 , n41918 );
and ( n41920 , n41823 , n41919 );
and ( n41921 , n41777 , n41822 );
or ( n41922 , n41920 , n41921 );
not ( n41923 , n41922 );
xor ( n41924 , n41658 , n41668 );
xor ( n41925 , n41924 , n41675 );
or ( n41926 , n41132 , n41816 );
or ( n41927 , n41672 , n41094 );
nand ( n41928 , n41926 , n41927 );
or ( n41929 , n41192 , n40377 );
nand ( n41930 , n41929 , n504 );
nand ( n41931 , n41192 , n40377 );
and ( n41932 , n41930 , n41931 , n29512 );
not ( n41933 , n3980 );
not ( n41934 , n41634 );
or ( n41935 , n41933 , n41934 );
not ( n41936 , n41810 );
nand ( n41937 , n41936 , n41463 );
nand ( n41938 , n41935 , n41937 );
xor ( n41939 , n41932 , n41938 );
xor ( n41940 , n41928 , n41939 );
xor ( n41941 , n41782 , n41791 );
and ( n41942 , n41941 , n41802 );
and ( n41943 , n41782 , n41791 );
or ( n41944 , n41942 , n41943 );
and ( n41945 , n41940 , n41944 );
and ( n41946 , n41928 , n41939 );
or ( n41947 , n41945 , n41946 );
xor ( n41948 , n41925 , n41947 );
and ( n41949 , n41932 , n41938 );
not ( n41950 , n41800 );
not ( n41951 , n41313 );
or ( n41952 , n41950 , n41951 );
nand ( n41953 , n41644 , n41200 );
nand ( n41954 , n41952 , n41953 );
and ( n41955 , n41281 , n29512 );
and ( n41956 , n41055 , n504 );
nor ( n41957 , n41955 , n41956 );
or ( n41958 , n41206 , n41957 );
or ( n41959 , n41655 , n41053 );
nand ( n41960 , n41958 , n41959 );
xor ( n41961 , n41954 , n41960 );
not ( n41962 , n41787 );
or ( n41963 , n41962 , n41220 );
or ( n41964 , n41666 , n3945 );
nand ( n41965 , n41963 , n41964 );
and ( n41966 , n41961 , n41965 );
and ( n41967 , n41954 , n41960 );
or ( n41968 , n41966 , n41967 );
xor ( n41969 , n41949 , n41968 );
xor ( n41970 , n41631 , n41639 );
xor ( n41971 , n41970 , n41648 );
xor ( n41972 , n41969 , n41971 );
xor ( n41973 , n41948 , n41972 );
xor ( n41974 , n41954 , n41960 );
xor ( n41975 , n41974 , n41965 );
xor ( n41976 , n41812 , n41818 );
and ( n41977 , n41976 , n41820 );
and ( n41978 , n41812 , n41818 );
or ( n41979 , n41977 , n41978 );
xor ( n41980 , n41975 , n41979 );
xor ( n41981 , n41928 , n41939 );
xor ( n41982 , n41981 , n41944 );
and ( n41983 , n41980 , n41982 );
and ( n41984 , n41975 , n41979 );
or ( n41985 , n41983 , n41984 );
or ( n41986 , n41973 , n41985 );
xor ( n41987 , n41975 , n41979 );
xor ( n41988 , n41987 , n41982 );
xor ( n41989 , n41781 , n41803 );
and ( n41990 , n41989 , n41821 );
and ( n41991 , n41781 , n41803 );
or ( n41992 , n41990 , n41991 );
or ( n41993 , n41988 , n41992 );
and ( n41994 , n41986 , n41993 );
not ( n41995 , n41994 );
or ( n41996 , n41923 , n41995 );
nand ( n41997 , n41988 , n41992 );
not ( n41998 , n41997 );
nand ( n41999 , n41973 , n41985 );
not ( n42000 , n41999 );
or ( n42001 , n41998 , n42000 );
nand ( n42002 , n42001 , n41986 );
nand ( n42003 , n41996 , n42002 );
not ( n42004 , n42003 );
xor ( n42005 , n41603 , n41610 );
xor ( n42006 , n42005 , n41612 );
xor ( n42007 , n41651 , n41678 );
xor ( n42008 , n42007 , n41681 );
xor ( n42009 , n42006 , n42008 );
xor ( n42010 , n41949 , n41968 );
and ( n42011 , n42010 , n41971 );
and ( n42012 , n41949 , n41968 );
or ( n42013 , n42011 , n42012 );
xor ( n42014 , n42009 , n42013 );
xor ( n42015 , n41925 , n41947 );
and ( n42016 , n42015 , n41972 );
and ( n42017 , n41925 , n41947 );
or ( n42018 , n42016 , n42017 );
nor ( n42019 , n42014 , n42018 );
xor ( n42020 , n42006 , n42008 );
and ( n42021 , n42020 , n42013 );
and ( n42022 , n42006 , n42008 );
or ( n42023 , n42021 , n42022 );
not ( n42024 , n42023 );
not ( n42025 , n42024 );
xor ( n42026 , n41629 , n41684 );
xor ( n42027 , n42026 , n41687 );
nor ( n42028 , n42025 , n42027 );
nor ( n42029 , n42019 , n42028 );
not ( n42030 , n42029 );
or ( n42031 , n42004 , n42030 );
and ( n42032 , n42014 , n42018 );
not ( n42033 , n42028 );
and ( n42034 , n42032 , n42033 );
not ( n42035 , n42027 );
nor ( n42036 , n42035 , n42024 );
nor ( n42037 , n42034 , n42036 );
nand ( n42038 , n42031 , n42037 );
or ( n42039 , n41627 , n41690 );
nand ( n42040 , n42038 , n41625 , n42039 );
nand ( n42041 , n41694 , n42040 );
not ( n42042 , n42041 );
xor ( n42043 , n41450 , n41511 );
xor ( n42044 , n42043 , n41514 );
xor ( n42045 , n41523 , n41525 );
and ( n42046 , n42045 , n41588 );
and ( n42047 , n41523 , n41525 );
or ( n42048 , n42046 , n42047 );
nor ( n42049 , n42044 , n42048 );
or ( n42050 , n42042 , n42049 );
nand ( n42051 , n42044 , n42048 );
nand ( n42052 , n42050 , n42051 );
not ( n42053 , n42052 );
or ( n42054 , n41521 , n42053 );
or ( n42055 , n42052 , n41520 );
nand ( n42056 , n42054 , n42055 );
nand ( n42057 , n42056 , n29519 );
nand ( n42058 , n41039 , n42057 );
not ( n42059 , n29520 );
not ( n42060 , n40879 );
not ( n42061 , n42060 );
not ( n42062 , n42061 );
not ( n42063 , n40861 );
not ( n42064 , n42063 );
not ( n42065 , n40934 );
nand ( n42066 , n42064 , n42065 );
not ( n42067 , n42066 );
or ( n42068 , n42062 , n42067 );
or ( n42069 , n42061 , n42066 );
nand ( n42070 , n42068 , n42069 );
not ( n42071 , n42070 );
or ( n42072 , n42059 , n42071 );
nand ( n42073 , n41986 , n41999 );
not ( n42074 , n42073 );
not ( n42075 , n41993 );
not ( n42076 , n41922 );
or ( n42077 , n42075 , n42076 );
nand ( n42078 , n42077 , n41997 );
not ( n42079 , n42078 );
or ( n42080 , n42074 , n42079 );
or ( n42081 , n42078 , n42073 );
nand ( n42082 , n42080 , n42081 );
nand ( n42083 , n42082 , n29519 );
nand ( n42084 , n42072 , n42083 );
not ( n42085 , n29520 );
buf ( n42086 , n41012 );
not ( n42087 , n42086 );
nor ( n42088 , n42060 , n42063 );
buf ( n42089 , n40945 );
and ( n42090 , n42088 , n42089 );
not ( n42091 , n41028 );
not ( n42092 , n42091 );
and ( n42093 , n42065 , n42092 );
nand ( n42094 , n42090 , n42093 );
not ( n42095 , n42094 );
or ( n42096 , n42087 , n42095 );
or ( n42097 , n42086 , n42094 );
nand ( n42098 , n42096 , n42097 );
not ( n42099 , n42098 );
or ( n42100 , n42085 , n42099 );
not ( n42101 , n41691 );
nand ( n42102 , n42039 , n42101 );
not ( n42103 , n42102 );
buf ( n42104 , n42038 );
not ( n42105 , n42104 );
or ( n42106 , n42103 , n42105 );
or ( n42107 , n42104 , n42102 );
nand ( n42108 , n42106 , n42107 );
nand ( n42109 , n42108 , n29519 );
nand ( n42110 , n42100 , n42109 );
not ( n42111 , n29520 );
and ( n42112 , n42092 , n42086 , n42065 );
nand ( n42113 , n42112 , n42088 , n42089 );
buf ( n42114 , n40992 );
and ( n42115 , n42114 , n40995 );
not ( n42116 , n42114 );
and ( n42117 , n42116 , n40981 );
nor ( n42118 , n42115 , n42117 );
not ( n42119 , n42118 );
and ( n42120 , n42113 , n42119 );
not ( n42121 , n42113 );
and ( n42122 , n42121 , n42118 );
nor ( n42123 , n42120 , n42122 );
not ( n42124 , n42123 );
or ( n42125 , n42111 , n42124 );
not ( n42126 , n41693 );
nand ( n42127 , n42126 , n41625 );
not ( n42128 , n42127 );
not ( n42129 , n42039 );
not ( n42130 , n42104 );
or ( n42131 , n42129 , n42130 );
nand ( n42132 , n42131 , n42101 );
not ( n42133 , n42132 );
or ( n42134 , n42128 , n42133 );
or ( n42135 , n42132 , n42127 );
nand ( n42136 , n42134 , n42135 );
nand ( n42137 , n42136 , n29519 );
nand ( n42138 , n42125 , n42137 );
not ( n42139 , n29520 );
buf ( n42140 , n40841 );
not ( n42141 , n42140 );
buf ( n42142 , n40859 );
nand ( n42143 , n42142 , n42065 );
not ( n42144 , n42143 );
or ( n42145 , n42141 , n42144 );
or ( n42146 , n42140 , n42143 );
nand ( n42147 , n42145 , n42146 );
not ( n42148 , n42147 );
or ( n42149 , n42139 , n42148 );
nand ( n42150 , n41993 , n41997 );
not ( n42151 , n42150 );
not ( n42152 , n41922 );
or ( n42153 , n42151 , n42152 );
or ( n42154 , n41922 , n42150 );
nand ( n42155 , n42153 , n42154 );
nand ( n42156 , n42155 , n29519 );
nand ( n42157 , n42149 , n42156 );
nand ( n42158 , n41903 , n41914 );
xor ( n42159 , n41890 , n42158 );
and ( n42160 , n29519 , n42159 );
not ( n42161 , n29519 );
not ( n42162 , n40932 );
nand ( n42163 , n3834 , n40881 , n40882 );
nand ( n42164 , n42163 , n40908 );
not ( n42165 , n42164 );
or ( n42166 , n42162 , n42165 );
or ( n42167 , n40932 , n42164 );
nand ( n42168 , n42166 , n42167 );
and ( n42169 , n42161 , n42168 );
nor ( n42170 , n42160 , n42169 );
not ( n42171 , n29520 );
nand ( n42172 , n40883 , n40906 );
not ( n42173 , n42172 );
not ( n42174 , n40895 );
or ( n42175 , n42173 , n42174 );
or ( n42176 , n40895 , n42172 );
nand ( n42177 , n42175 , n42176 );
not ( n42178 , n42177 );
or ( n42179 , n42171 , n42178 );
xor ( n42180 , n41849 , n41875 );
xor ( n42181 , n42180 , n41887 );
nand ( n42182 , n42181 , n29519 );
nand ( n42183 , n42179 , n42182 );
or ( n42184 , n41163 , n41171 );
nand ( n42185 , n42184 , n41157 );
buf ( n42186 , n41156 );
nor ( n42187 , n42186 , n36435 );
xor ( n42188 , n42185 , n42187 );
nand ( n42189 , n41157 , n490 );
not ( n42190 , n42189 );
xor ( n42191 , n42188 , n42190 );
and ( n42192 , n41157 , n36435 );
and ( n42193 , n41167 , n489 );
nor ( n42194 , n42192 , n42193 );
or ( n42195 , n41164 , n42194 );
or ( n42196 , n41172 , n42186 );
nand ( n42197 , n42195 , n42196 );
xor ( n42198 , n42197 , n42189 );
not ( n42199 , n41115 );
not ( n42200 , n41597 );
or ( n42201 , n42199 , n42200 );
nand ( n42202 , n42201 , n41102 );
and ( n42203 , n41157 , n36727 );
and ( n42204 , n41167 , n490 );
nor ( n42205 , n42203 , n42204 );
or ( n42206 , n41164 , n42205 );
or ( n42207 , n42194 , n41172 );
nand ( n42208 , n42206 , n42207 );
xor ( n42209 , n42202 , n42208 );
nor ( n42210 , n42186 , n36583 );
and ( n42211 , n42209 , n42210 );
and ( n42212 , n42202 , n42208 );
or ( n42213 , n42211 , n42212 );
and ( n42214 , n42198 , n42213 );
and ( n42215 , n42197 , n42189 );
or ( n42216 , n42214 , n42215 );
xnor ( n42217 , n42191 , n42216 );
not ( n42218 , n42217 );
or ( n42219 , n41103 , n496 );
or ( n42220 , n41102 , n41208 );
nand ( n42221 , n42219 , n42220 );
not ( n42222 , n42221 );
not ( n42223 , n41126 );
or ( n42224 , n42222 , n42223 );
or ( n42225 , n41103 , n495 );
or ( n42226 , n41102 , n41328 );
nand ( n42227 , n42225 , n42226 );
nand ( n42228 , n42227 , n41630 );
nand ( n42229 , n42224 , n42228 );
and ( n42230 , n492 , n41045 );
not ( n42231 , n492 );
and ( n42232 , n42231 , n41192 );
nor ( n42233 , n42230 , n42232 );
or ( n42234 , n41252 , n42233 );
and ( n42235 , n491 , n41049 );
not ( n42236 , n491 );
and ( n42237 , n42236 , n41192 );
nor ( n42238 , n42235 , n42237 );
or ( n42239 , n41188 , n42238 );
nand ( n42240 , n42234 , n42239 );
xor ( n42241 , n42229 , n42240 );
and ( n42242 , n41165 , n701 );
and ( n42243 , n41167 , n498 );
nor ( n42244 , n42242 , n42243 );
or ( n42245 , n41164 , n42244 );
and ( n42246 , n41165 , n41532 );
and ( n42247 , n41167 , n497 );
nor ( n42248 , n42246 , n42247 );
or ( n42249 , n42248 , n41172 );
nand ( n42250 , n42245 , n42249 );
and ( n42251 , n42241 , n42250 );
and ( n42252 , n42229 , n42240 );
or ( n42253 , n42251 , n42252 );
or ( n42254 , n41463 , n3980 );
nand ( n42255 , n42254 , n3916 );
and ( n42256 , n490 , n41070 );
not ( n42257 , n490 );
and ( n42258 , n42257 , n41073 );
nor ( n42259 , n42256 , n42258 );
or ( n42260 , n41132 , n42259 );
and ( n42261 , n41135 , n36435 );
and ( n42262 , n41070 , n489 );
nor ( n42263 , n42261 , n42262 );
or ( n42264 , n41094 , n42263 );
nand ( n42265 , n42260 , n42264 );
xor ( n42266 , n42255 , n42265 );
and ( n42267 , n29512 , n41196 );
and ( n42268 , n41040 , n494 );
nor ( n42269 , n42267 , n42268 );
or ( n42270 , n41319 , n42269 );
and ( n42271 , n29512 , n41089 );
and ( n42272 , n41040 , n493 );
nor ( n42273 , n42271 , n42272 );
or ( n42274 , n41053 , n42273 );
nand ( n42275 , n42270 , n42274 );
and ( n42276 , n42266 , n42275 );
and ( n42277 , n42255 , n42265 );
or ( n42278 , n42276 , n42277 );
xor ( n42279 , n42253 , n42278 );
not ( n42280 , n42227 );
not ( n42281 , n41126 );
or ( n42282 , n42280 , n42281 );
or ( n42283 , n41103 , n494 );
or ( n42284 , n41102 , n41196 );
nand ( n42285 , n42283 , n42284 );
nand ( n42286 , n42285 , n41630 );
nand ( n42287 , n42282 , n42286 );
or ( n42288 , n41164 , n42248 );
not ( n42289 , n41157 );
not ( n42290 , n41208 );
and ( n42291 , n42289 , n42290 );
and ( n42292 , n41157 , n41208 );
nor ( n42293 , n42291 , n42292 );
or ( n42294 , n42293 , n41172 );
nand ( n42295 , n42288 , n42294 );
xor ( n42296 , n42287 , n42295 );
or ( n42297 , n41085 , n42263 );
or ( n42298 , n41094 , n41070 );
nand ( n42299 , n42297 , n42298 );
xor ( n42300 , n42296 , n42299 );
xor ( n42301 , n42279 , n42300 );
nor ( n42302 , n41280 , n701 );
or ( n42303 , n41319 , n42273 );
and ( n42304 , n41134 , n29512 );
not ( n42305 , n41134 );
and ( n42306 , n42305 , n41040 );
nor ( n42307 , n42304 , n42306 );
or ( n42308 , n41053 , n42307 );
nand ( n42309 , n42303 , n42308 );
xor ( n42310 , n42302 , n42309 );
or ( n42311 , n41189 , n42238 );
and ( n42312 , n41192 , n36727 );
and ( n42313 , n41049 , n490 );
nor ( n42314 , n42312 , n42313 );
or ( n42315 , n41201 , n42314 );
nand ( n42316 , n42311 , n42315 );
not ( n42317 , n42316 );
xor ( n42318 , n42310 , n42317 );
nor ( n42319 , n42186 , n29596 );
and ( n42320 , n3916 , n36435 );
and ( n42321 , n3921 , n489 );
nor ( n42322 , n42320 , n42321 );
or ( n42323 , n3920 , n42322 );
or ( n42324 , n41230 , n3921 );
nand ( n42325 , n42323 , n42324 );
xor ( n42326 , n42319 , n42325 );
and ( n42327 , n491 , n41073 );
not ( n42328 , n491 );
and ( n42329 , n42328 , n41070 );
nor ( n42330 , n42327 , n42329 );
not ( n42331 , n42330 );
or ( n42332 , n41085 , n42331 );
or ( n42333 , n41094 , n42259 );
nand ( n42334 , n42332 , n42333 );
and ( n42335 , n29512 , n41328 );
and ( n42336 , n41040 , n495 );
nor ( n42337 , n42335 , n42336 );
or ( n42338 , n41319 , n42337 );
or ( n42339 , n42269 , n41053 );
nand ( n42340 , n42338 , n42339 );
xor ( n42341 , n42334 , n42340 );
and ( n42342 , n41102 , n41532 );
and ( n42343 , n41103 , n497 );
nor ( n42344 , n42342 , n42343 );
or ( n42345 , n41597 , n42344 );
not ( n42346 , n42221 );
or ( n42347 , n42346 , n41115 );
nand ( n42348 , n42345 , n42347 );
and ( n42349 , n42341 , n42348 );
and ( n42350 , n42334 , n42340 );
or ( n42351 , n42349 , n42350 );
and ( n42352 , n42326 , n42351 );
and ( n42353 , n42319 , n42325 );
or ( n42354 , n42352 , n42353 );
xor ( n42355 , n42318 , n42354 );
and ( n42356 , n493 , n41045 );
not ( n42357 , n493 );
and ( n42358 , n42357 , n41192 );
nor ( n42359 , n42356 , n42358 );
or ( n42360 , n42359 , n41252 );
not ( n42361 , n42233 );
nand ( n42362 , n42361 , n41200 );
nand ( n42363 , n42360 , n42362 );
and ( n42364 , n41157 , n29596 );
and ( n42365 , n41156 , n499 );
nor ( n42366 , n42364 , n42365 );
not ( n42367 , n42366 );
not ( n42368 , n42367 );
not ( n42369 , n41163 );
or ( n42370 , n42368 , n42369 );
not ( n42371 , n42244 );
nand ( n42372 , n42371 , n41171 );
nand ( n42373 , n42370 , n42372 );
xor ( n42374 , n42363 , n42373 );
nor ( n42375 , n41167 , n41118 );
and ( n42376 , n42374 , n42375 );
and ( n42377 , n42363 , n42373 );
or ( n42378 , n42376 , n42377 );
xor ( n42379 , n42229 , n42240 );
xor ( n42380 , n42379 , n42250 );
xor ( n42381 , n42378 , n42380 );
xor ( n42382 , n42255 , n42265 );
xor ( n42383 , n42382 , n42275 );
and ( n42384 , n42381 , n42383 );
and ( n42385 , n42378 , n42380 );
or ( n42386 , n42384 , n42385 );
xor ( n42387 , n42355 , n42386 );
xor ( n42388 , n42301 , n42387 );
xor ( n42389 , n42319 , n42325 );
xor ( n42390 , n42389 , n42351 );
not ( n42391 , n42325 );
or ( n42392 , n3920 , n41234 );
or ( n42393 , n41230 , n42322 );
nand ( n42394 , n42392 , n42393 );
or ( n42395 , n3946 , n3944 );
nand ( n42396 , n42395 , n32891 );
or ( n42397 , n42394 , n42396 );
xor ( n42398 , n42391 , n42397 );
nor ( n42399 , n41167 , n3959 );
or ( n42400 , n41252 , n41199 );
or ( n42401 , n42359 , n41201 );
nand ( n42402 , n42400 , n42401 );
xor ( n42403 , n42399 , n42402 );
or ( n42404 , n41319 , n41211 );
or ( n42405 , n42337 , n41053 );
nand ( n42406 , n42404 , n42405 );
and ( n42407 , n42403 , n42406 );
and ( n42408 , n42399 , n42402 );
or ( n42409 , n42407 , n42408 );
and ( n42410 , n42398 , n42409 );
and ( n42411 , n42391 , n42397 );
or ( n42412 , n42410 , n42411 );
xor ( n42413 , n42390 , n42412 );
not ( n42414 , n41140 );
not ( n42415 , n42414 );
not ( n42416 , n41086 );
or ( n42417 , n42415 , n42416 );
nand ( n42418 , n42330 , n41093 );
nand ( n42419 , n42417 , n42418 );
not ( n42420 , n41630 );
not ( n42421 , n42344 );
not ( n42422 , n42421 );
or ( n42423 , n42420 , n42422 );
not ( n42424 , n41126 );
or ( n42425 , n42424 , n41147 );
nand ( n42426 , n42423 , n42425 );
xor ( n42427 , n42419 , n42426 );
or ( n42428 , n41164 , n41175 );
or ( n42429 , n42366 , n41172 );
nand ( n42430 , n42428 , n42429 );
and ( n42431 , n42427 , n42430 );
and ( n42432 , n42419 , n42426 );
or ( n42433 , n42431 , n42432 );
xor ( n42434 , n42363 , n42373 );
xor ( n42435 , n42434 , n42375 );
xor ( n42436 , n42433 , n42435 );
xor ( n42437 , n42334 , n42340 );
xor ( n42438 , n42437 , n42348 );
and ( n42439 , n42436 , n42438 );
and ( n42440 , n42433 , n42435 );
or ( n42441 , n42439 , n42440 );
and ( n42442 , n42413 , n42441 );
and ( n42443 , n42390 , n42412 );
or ( n42444 , n42442 , n42443 );
and ( n42445 , n42388 , n42444 );
and ( n42446 , n42301 , n42387 );
or ( n42447 , n42445 , n42446 );
xor ( n42448 , n42253 , n42278 );
and ( n42449 , n42448 , n42300 );
and ( n42450 , n42253 , n42278 );
or ( n42451 , n42449 , n42450 );
not ( n42452 , n41094 );
not ( n42453 , n41085 );
or ( n42454 , n42452 , n42453 );
nand ( n42455 , n42454 , n41073 );
or ( n42456 , n41252 , n42314 );
and ( n42457 , n41192 , n36435 );
and ( n42458 , n41049 , n489 );
nor ( n42459 , n42457 , n42458 );
or ( n42460 , n41201 , n42459 );
nand ( n42461 , n42456 , n42460 );
xor ( n42462 , n42455 , n42461 );
not ( n42463 , n42285 );
or ( n42464 , n42424 , n42463 );
and ( n42465 , n41102 , n41089 );
and ( n42466 , n41103 , n493 );
nor ( n42467 , n42465 , n42466 );
or ( n42468 , n41115 , n42467 );
nand ( n42469 , n42464 , n42468 );
xor ( n42470 , n42462 , n42469 );
xor ( n42471 , n42302 , n42309 );
and ( n42472 , n42471 , n42317 );
and ( n42473 , n42302 , n42309 );
or ( n42474 , n42472 , n42473 );
xor ( n42475 , n42470 , n42474 );
xor ( n42476 , n42287 , n42295 );
and ( n42477 , n42476 , n42299 );
and ( n42478 , n42287 , n42295 );
or ( n42479 , n42477 , n42478 );
xor ( n42480 , n42316 , n42479 );
not ( n42481 , n42293 );
not ( n42482 , n42481 );
not ( n42483 , n41163 );
or ( n42484 , n42482 , n42483 );
and ( n42485 , n495 , n41165 );
not ( n42486 , n495 );
and ( n42487 , n42486 , n41167 );
nor ( n42488 , n42485 , n42487 );
nand ( n42489 , n42488 , n41171 );
nand ( n42490 , n42484 , n42489 );
not ( n42491 , n42307 );
not ( n42492 , n42491 );
not ( n42493 , n41066 );
or ( n42494 , n42492 , n42493 );
and ( n42495 , n491 , n29512 );
not ( n42496 , n491 );
and ( n42497 , n42496 , n41040 );
nor ( n42498 , n42495 , n42497 );
nand ( n42499 , n41052 , n42498 );
nand ( n42500 , n42494 , n42499 );
xor ( n42501 , n42490 , n42500 );
nor ( n42502 , n41280 , n41532 );
xor ( n42503 , n42501 , n42502 );
xor ( n42504 , n42480 , n42503 );
xor ( n42505 , n42475 , n42504 );
xor ( n42506 , n42451 , n42505 );
xor ( n42507 , n42318 , n42354 );
and ( n42508 , n42507 , n42386 );
and ( n42509 , n42318 , n42354 );
or ( n42510 , n42508 , n42509 );
xor ( n42511 , n42506 , n42510 );
or ( n42512 , n42447 , n42511 );
xor ( n42513 , n42451 , n42505 );
and ( n42514 , n42513 , n42510 );
and ( n42515 , n42451 , n42505 );
or ( n42516 , n42514 , n42515 );
xor ( n42517 , n42316 , n42479 );
and ( n42518 , n42517 , n42503 );
and ( n42519 , n42316 , n42479 );
or ( n42520 , n42518 , n42519 );
xor ( n42521 , n42455 , n42461 );
and ( n42522 , n42521 , n42469 );
and ( n42523 , n42455 , n42461 );
or ( n42524 , n42522 , n42523 );
not ( n42525 , n42488 );
or ( n42526 , n41162 , n42525 );
and ( n42527 , n494 , n41167 );
not ( n42528 , n494 );
and ( n42529 , n42528 , n41157 );
nor ( n42530 , n42527 , n42529 );
or ( n42531 , n42530 , n41151 );
nand ( n42532 , n42526 , n42531 );
and ( n42533 , n41165 , n496 );
xor ( n42534 , n42532 , n42533 );
or ( n42535 , n41252 , n42459 );
or ( n42536 , n41201 , n41049 );
nand ( n42537 , n42535 , n42536 );
xor ( n42538 , n42534 , n42537 );
xor ( n42539 , n42524 , n42538 );
or ( n42540 , n41597 , n42467 );
and ( n42541 , n41102 , n41134 );
and ( n42542 , n41103 , n492 );
nor ( n42543 , n42541 , n42542 );
or ( n42544 , n41115 , n42543 );
nand ( n42545 , n42540 , n42544 );
not ( n42546 , n42498 );
or ( n42547 , n41319 , n42546 );
and ( n42548 , n36727 , n29512 );
not ( n42549 , n36727 );
and ( n42550 , n42549 , n41040 );
nor ( n42551 , n42548 , n42550 );
or ( n42552 , n41053 , n42551 );
nand ( n42553 , n42547 , n42552 );
not ( n42554 , n42553 );
xor ( n42555 , n42545 , n42554 );
xor ( n42556 , n42490 , n42500 );
and ( n42557 , n42556 , n42502 );
and ( n42558 , n42490 , n42500 );
or ( n42559 , n42557 , n42558 );
xor ( n42560 , n42555 , n42559 );
xor ( n42561 , n42539 , n42560 );
xor ( n42562 , n42520 , n42561 );
xor ( n42563 , n42470 , n42474 );
and ( n42564 , n42563 , n42504 );
and ( n42565 , n42470 , n42474 );
or ( n42566 , n42564 , n42565 );
xor ( n42567 , n42562 , n42566 );
nor ( n42568 , n42516 , n42567 );
not ( n42569 , n42568 );
xor ( n42570 , n42520 , n42561 );
and ( n42571 , n42570 , n42566 );
and ( n42572 , n42520 , n42561 );
or ( n42573 , n42571 , n42572 );
xor ( n42574 , n42545 , n42554 );
and ( n42575 , n42574 , n42559 );
and ( n42576 , n42545 , n42554 );
or ( n42577 , n42575 , n42576 );
xor ( n42578 , n42532 , n42533 );
and ( n42579 , n42578 , n42537 );
and ( n42580 , n42532 , n42533 );
or ( n42581 , n42579 , n42580 );
not ( n42582 , n41201 );
not ( n42583 , n41252 );
or ( n42584 , n42582 , n42583 );
nand ( n42585 , n42584 , n41192 );
or ( n42586 , n41319 , n42551 );
and ( n42587 , n489 , n41040 );
not ( n42588 , n489 );
and ( n42589 , n42588 , n29512 );
nor ( n42590 , n42587 , n42589 );
or ( n42591 , n41053 , n42590 );
nand ( n42592 , n42586 , n42591 );
xor ( n42593 , n42585 , n42592 );
or ( n42594 , n41164 , n42530 );
and ( n42595 , n41165 , n41089 );
and ( n42596 , n42186 , n493 );
nor ( n42597 , n42595 , n42596 );
or ( n42598 , n42597 , n41172 );
nand ( n42599 , n42594 , n42598 );
xor ( n42600 , n42593 , n42599 );
xor ( n42601 , n42581 , n42600 );
nor ( n42602 , n41167 , n41328 );
or ( n42603 , n41597 , n42543 );
and ( n42604 , n491 , n41103 );
not ( n42605 , n491 );
and ( n42606 , n42605 , n41102 );
nor ( n42607 , n42604 , n42606 );
or ( n42608 , n41115 , n42607 );
nand ( n42609 , n42603 , n42608 );
xor ( n42610 , n42602 , n42609 );
xor ( n42611 , n42610 , n42553 );
xor ( n42612 , n42601 , n42611 );
xor ( n42613 , n42577 , n42612 );
xor ( n42614 , n42524 , n42538 );
and ( n42615 , n42614 , n42560 );
and ( n42616 , n42524 , n42538 );
or ( n42617 , n42615 , n42616 );
xor ( n42618 , n42613 , n42617 );
or ( n42619 , n42573 , n42618 );
and ( n42620 , n42512 , n42569 , n42619 );
xor ( n42621 , n42577 , n42612 );
and ( n42622 , n42621 , n42617 );
and ( n42623 , n42577 , n42612 );
or ( n42624 , n42622 , n42623 );
xor ( n42625 , n42602 , n42609 );
and ( n42626 , n42625 , n42553 );
and ( n42627 , n42602 , n42609 );
or ( n42628 , n42626 , n42627 );
or ( n42629 , n41319 , n42590 );
or ( n42630 , n41053 , n41040 );
nand ( n42631 , n42629 , n42630 );
not ( n42632 , n42631 );
xor ( n42633 , n42585 , n42592 );
and ( n42634 , n42633 , n42599 );
and ( n42635 , n42585 , n42592 );
or ( n42636 , n42634 , n42635 );
xor ( n42637 , n42632 , n42636 );
nor ( n42638 , n41167 , n41196 );
not ( n42639 , n42607 );
not ( n42640 , n42639 );
not ( n42641 , n41126 );
or ( n42642 , n42640 , n42641 );
or ( n42643 , n41103 , n490 );
or ( n42644 , n41102 , n36727 );
nand ( n42645 , n42643 , n42644 );
nand ( n42646 , n42645 , n41630 );
nand ( n42647 , n42642 , n42646 );
xor ( n42648 , n42638 , n42647 );
or ( n42649 , n41164 , n42597 );
and ( n42650 , n41157 , n41134 );
and ( n42651 , n41280 , n492 );
nor ( n42652 , n42650 , n42651 );
or ( n42653 , n42652 , n41172 );
nand ( n42654 , n42649 , n42653 );
xor ( n42655 , n42648 , n42654 );
xor ( n42656 , n42637 , n42655 );
xor ( n42657 , n42628 , n42656 );
xor ( n42658 , n42581 , n42600 );
and ( n42659 , n42658 , n42611 );
and ( n42660 , n42581 , n42600 );
or ( n42661 , n42659 , n42660 );
xor ( n42662 , n42657 , n42661 );
or ( n42663 , n42624 , n42662 );
xor ( n42664 , n42628 , n42656 );
and ( n42665 , n42664 , n42661 );
and ( n42666 , n42628 , n42656 );
or ( n42667 , n42665 , n42666 );
not ( n42668 , n42667 );
or ( n42669 , n41066 , n41052 );
nand ( n42670 , n42669 , n29512 );
not ( n42671 , n42645 );
or ( n42672 , n41597 , n42671 );
and ( n42673 , n41102 , n36435 );
and ( n42674 , n41103 , n489 );
nor ( n42675 , n42673 , n42674 );
or ( n42676 , n42675 , n41115 );
nand ( n42677 , n42672 , n42676 );
xor ( n42678 , n42670 , n42677 );
nor ( n42679 , n42186 , n41089 );
xor ( n42680 , n42678 , n42679 );
or ( n42681 , n41164 , n42652 );
and ( n42682 , n41165 , n36583 );
and ( n42683 , n42186 , n491 );
nor ( n42684 , n42682 , n42683 );
or ( n42685 , n42684 , n41172 );
nand ( n42686 , n42681 , n42685 );
xor ( n42687 , n42686 , n42631 );
xor ( n42688 , n42638 , n42647 );
and ( n42689 , n42688 , n42654 );
and ( n42690 , n42638 , n42647 );
or ( n42691 , n42689 , n42690 );
xor ( n42692 , n42687 , n42691 );
xor ( n42693 , n42680 , n42692 );
xor ( n42694 , n42632 , n42636 );
and ( n42695 , n42694 , n42655 );
and ( n42696 , n42632 , n42636 );
or ( n42697 , n42695 , n42696 );
xor ( n42698 , n42693 , n42697 );
not ( n42699 , n42698 );
nand ( n42700 , n42668 , n42699 );
xor ( n42701 , n42680 , n42692 );
and ( n42702 , n42701 , n42697 );
and ( n42703 , n42680 , n42692 );
or ( n42704 , n42702 , n42703 );
xor ( n42705 , n42670 , n42677 );
and ( n42706 , n42705 , n42679 );
and ( n42707 , n42670 , n42677 );
or ( n42708 , n42706 , n42707 );
or ( n42709 , n41164 , n42684 );
or ( n42710 , n42205 , n41172 );
nand ( n42711 , n42709 , n42710 );
nor ( n42712 , n41167 , n41134 );
xor ( n42713 , n42711 , n42712 );
not ( n42714 , n42675 );
and ( n42715 , n41126 , n42714 );
and ( n42716 , n41630 , n41102 );
nor ( n42717 , n42715 , n42716 );
xor ( n42718 , n42713 , n42717 );
xor ( n42719 , n42708 , n42718 );
xor ( n42720 , n42686 , n42631 );
and ( n42721 , n42720 , n42691 );
and ( n42722 , n42686 , n42631 );
or ( n42723 , n42721 , n42722 );
xor ( n42724 , n42719 , n42723 );
nor ( n42725 , n42704 , n42724 );
xor ( n42726 , n42708 , n42718 );
and ( n42727 , n42726 , n42723 );
and ( n42728 , n42708 , n42718 );
or ( n42729 , n42727 , n42728 );
not ( n42730 , n42717 );
xor ( n42731 , n42202 , n42208 );
xor ( n42732 , n42731 , n42210 );
xor ( n42733 , n42730 , n42732 );
xor ( n42734 , n42711 , n42712 );
and ( n42735 , n42734 , n42717 );
and ( n42736 , n42711 , n42712 );
or ( n42737 , n42735 , n42736 );
xor ( n42738 , n42733 , n42737 );
nor ( n42739 , n42729 , n42738 );
nor ( n42740 , n42725 , n42739 );
xor ( n42741 , n42730 , n42732 );
and ( n42742 , n42741 , n42737 );
and ( n42743 , n42730 , n42732 );
or ( n42744 , n42742 , n42743 );
xor ( n42745 , n42197 , n42189 );
xor ( n42746 , n42745 , n42213 );
or ( n42747 , n42744 , n42746 );
and ( n42748 , n42663 , n42700 , n42740 , n42747 );
and ( n42749 , n42620 , n42748 );
not ( n42750 , n42749 );
xor ( n42751 , n42378 , n42380 );
xor ( n42752 , n42751 , n42383 );
xor ( n42753 , n42390 , n42412 );
xor ( n42754 , n42753 , n42441 );
xor ( n42755 , n42752 , n42754 );
and ( n42756 , n41224 , n41236 );
xor ( n42757 , n41203 , n41204 );
and ( n42758 , n42757 , n41213 );
and ( n42759 , n41203 , n41204 );
or ( n42760 , n42758 , n42759 );
xor ( n42761 , n42756 , n42760 );
xor ( n42762 , n41142 , n41149 );
and ( n42763 , n42762 , n41177 );
and ( n42764 , n41142 , n41149 );
or ( n42765 , n42763 , n42764 );
and ( n42766 , n42761 , n42765 );
and ( n42767 , n42756 , n42760 );
or ( n42768 , n42766 , n42767 );
xor ( n42769 , n42391 , n42397 );
xor ( n42770 , n42769 , n42409 );
xor ( n42771 , n42768 , n42770 );
xor ( n42772 , n42419 , n42426 );
xor ( n42773 , n42772 , n42430 );
not ( n42774 , n42396 );
not ( n42775 , n42394 );
or ( n42776 , n42774 , n42775 );
nand ( n42777 , n42776 , n42397 );
xor ( n42778 , n42773 , n42777 );
xor ( n42779 , n42399 , n42402 );
xor ( n42780 , n42779 , n42406 );
and ( n42781 , n42778 , n42780 );
and ( n42782 , n42773 , n42777 );
or ( n42783 , n42781 , n42782 );
and ( n42784 , n42771 , n42783 );
and ( n42785 , n42768 , n42770 );
or ( n42786 , n42784 , n42785 );
and ( n42787 , n42755 , n42786 );
and ( n42788 , n42752 , n42754 );
or ( n42789 , n42787 , n42788 );
not ( n42790 , n42789 );
xor ( n42791 , n42301 , n42387 );
xor ( n42792 , n42791 , n42444 );
not ( n42793 , n42792 );
nand ( n42794 , n42790 , n42793 );
xor ( n42795 , n42773 , n42777 );
xor ( n42796 , n42795 , n42780 );
xor ( n42797 , n41264 , n41305 );
and ( n42798 , n42797 , n41345 );
and ( n42799 , n41264 , n41305 );
or ( n42800 , n42798 , n42799 );
xor ( n42801 , n42796 , n42800 );
and ( n42802 , n41237 , n41263 );
xor ( n42803 , n42756 , n42760 );
xor ( n42804 , n42803 , n42765 );
xor ( n42805 , n42802 , n42804 );
xor ( n42806 , n41131 , n41178 );
and ( n42807 , n42806 , n41214 );
and ( n42808 , n41131 , n41178 );
or ( n42809 , n42807 , n42808 );
xor ( n42810 , n42805 , n42809 );
xor ( n42811 , n42801 , n42810 );
xor ( n42812 , n41215 , n41346 );
and ( n42813 , n42812 , n41447 );
and ( n42814 , n41215 , n41346 );
or ( n42815 , n42813 , n42814 );
nor ( n42816 , n42811 , n42815 );
xor ( n42817 , n42433 , n42435 );
xor ( n42818 , n42817 , n42438 );
xor ( n42819 , n42802 , n42804 );
and ( n42820 , n42819 , n42809 );
and ( n42821 , n42802 , n42804 );
or ( n42822 , n42820 , n42821 );
xor ( n42823 , n42818 , n42822 );
xor ( n42824 , n42768 , n42770 );
xor ( n42825 , n42824 , n42783 );
xor ( n42826 , n42823 , n42825 );
xor ( n42827 , n42796 , n42800 );
and ( n42828 , n42827 , n42810 );
and ( n42829 , n42796 , n42800 );
or ( n42830 , n42828 , n42829 );
nor ( n42831 , n42826 , n42830 );
nor ( n42832 , n42816 , n42831 );
xor ( n42833 , n42752 , n42754 );
xor ( n42834 , n42833 , n42786 );
xor ( n42835 , n42818 , n42822 );
and ( n42836 , n42835 , n42825 );
and ( n42837 , n42818 , n42822 );
or ( n42838 , n42836 , n42837 );
or ( n42839 , n42834 , n42838 );
and ( n42840 , n42794 , n42832 , n42839 );
not ( n42841 , n42840 );
nor ( n42842 , n41518 , n42049 );
not ( n42843 , n42842 );
not ( n42844 , n42041 );
or ( n42845 , n42843 , n42844 );
not ( n42846 , n41518 );
not ( n42847 , n42051 );
and ( n42848 , n42846 , n42847 );
nor ( n42849 , n42848 , n41519 );
nand ( n42850 , n42845 , n42849 );
not ( n42851 , n42850 );
or ( n42852 , n42841 , n42851 );
not ( n42853 , n42839 );
nand ( n42854 , n42815 , n42811 );
or ( n42855 , n42831 , n42854 );
nand ( n42856 , n42826 , n42830 );
nand ( n42857 , n42855 , n42856 );
not ( n42858 , n42857 );
or ( n42859 , n42853 , n42858 );
nand ( n42860 , n42834 , n42838 );
nand ( n42861 , n42859 , n42860 );
nand ( n42862 , n42793 , n42790 );
and ( n42863 , n42861 , n42862 );
nand ( n42864 , n42792 , n42789 );
not ( n42865 , n42864 );
nor ( n42866 , n42863 , n42865 );
nand ( n42867 , n42852 , n42866 );
buf ( n42868 , n42867 );
not ( n42869 , n42868 );
or ( n42870 , n42750 , n42869 );
not ( n42871 , n42619 );
nand ( n42872 , n42447 , n42511 );
or ( n42873 , n42872 , n42568 );
nand ( n42874 , n42516 , n42567 );
nand ( n42875 , n42873 , n42874 );
not ( n42876 , n42875 );
or ( n42877 , n42871 , n42876 );
nand ( n42878 , n42573 , n42618 );
nand ( n42879 , n42877 , n42878 );
and ( n42880 , n42748 , n42879 );
and ( n42881 , n42624 , n42662 );
and ( n42882 , n42881 , n42700 );
nor ( n42883 , n42668 , n42699 );
nor ( n42884 , n42882 , n42883 );
not ( n42885 , n42884 );
nand ( n42886 , n42885 , n42740 );
not ( n42887 , n42747 );
or ( n42888 , n42886 , n42887 );
nand ( n42889 , n42704 , n42724 );
not ( n42890 , n42889 );
not ( n42891 , n42739 );
and ( n42892 , n42890 , n42891 );
and ( n42893 , n42729 , n42738 );
nor ( n42894 , n42892 , n42893 );
or ( n42895 , n42894 , n42887 );
nand ( n42896 , n42744 , n42746 );
nand ( n42897 , n42888 , n42895 , n42896 );
nor ( n42898 , n42880 , n42897 );
nand ( n42899 , n42870 , n42898 );
not ( n42900 , n42899 );
or ( n42901 , n42218 , n42900 );
or ( n42902 , n42899 , n42217 );
nand ( n42903 , n42901 , n42902 );
and ( n42904 , n42903 , n29519 );
not ( n42905 , n32935 );
and ( n42906 , n29519 , n42905 );
not ( n42907 , n29519 );
xor ( n42908 , n3877 , n472 );
and ( n42909 , n42907 , n42908 );
or ( n42910 , n42906 , n42909 );
xor ( n42911 , n41777 , n41822 );
xor ( n42912 , n42911 , n41919 );
and ( n42913 , n29519 , n42912 );
not ( n42914 , n29519 );
xor ( n42915 , n42142 , n42065 );
and ( n42916 , n42914 , n42915 );
or ( n42917 , n42913 , n42916 );
or ( n42918 , n3987 , n3989 );
nand ( n42919 , n42918 , n3990 );
not ( n42920 , n42919 );
and ( n42921 , n29519 , n42920 );
not ( n42922 , n29519 );
xor ( n42923 , n471 , n3879 );
xor ( n42924 , n42923 , n3888 );
and ( n42925 , n42922 , n42924 );
or ( n42926 , n42921 , n42925 );
xor ( n42927 , n41877 , n41879 );
xor ( n42928 , n42927 , n41884 );
and ( n42929 , n29519 , n42928 );
not ( n42930 , n29519 );
xor ( n42931 , n42163 , n40906 );
and ( n42932 , n42930 , n42931 );
or ( n42933 , n42929 , n42932 );
nand ( n42934 , n3861 , n3900 );
not ( n42935 , n32848 );
and ( n42936 , n42934 , n42935 );
not ( n42937 , n42934 );
and ( n42938 , n42937 , n32848 );
nor ( n42939 , n42936 , n42938 );
not ( n42940 , n454 );
not ( n42941 , n2815 );
buf ( n42942 , n33438 );
not ( n42943 , n42942 );
buf ( n42944 , n42943 );
buf ( n42945 , n42944 );
not ( n42946 , n42945 );
buf ( n42947 , n36583 );
buf ( n42948 , n505 );
and ( n42949 , n42947 , n42948 );
buf ( n42950 , n505 );
not ( n42951 , n42950 );
buf ( n42952 , n42951 );
buf ( n42953 , n42952 );
buf ( n42954 , n491 );
and ( n42955 , n42953 , n42954 );
nor ( n42956 , n42949 , n42955 );
buf ( n42957 , n42956 );
buf ( n42958 , n42957 );
not ( n42959 , n42958 );
and ( n42960 , n42946 , n42959 );
buf ( n42961 , n4519 );
buf ( n42962 , n491 );
and ( n42963 , n42961 , n42962 );
nor ( n42964 , n42960 , n42963 );
buf ( n42965 , n42964 );
buf ( n42966 , n42965 );
not ( n42967 , n42966 );
buf ( n42968 , n42967 );
buf ( n42969 , n508 );
buf ( n42970 , n489 );
and ( n42971 , n42969 , n42970 );
buf ( n42972 , n42971 );
not ( n42973 , n42972 );
buf ( n42974 , n7008 );
not ( n42975 , n42974 );
not ( n42976 , n42975 );
and ( n42977 , n506 , n36435 );
not ( n42978 , n506 );
and ( n42979 , n42978 , n489 );
or ( n42980 , n42977 , n42979 );
not ( n42981 , n42980 );
or ( n42982 , n42976 , n42981 );
buf ( n42983 , n36435 );
buf ( n42984 , n507 );
and ( n42985 , n42983 , n42984 );
buf ( n42986 , n33214 );
buf ( n42987 , n489 );
and ( n42988 , n42986 , n42987 );
nor ( n42989 , n42985 , n42988 );
buf ( n42990 , n42989 );
not ( n42991 , n42990 );
not ( n42992 , n7315 );
nand ( n42993 , n42991 , n42992 );
nand ( n42994 , n42982 , n42993 );
not ( n42995 , n42994 );
or ( n42996 , n42973 , n42995 );
not ( n42997 , n42972 );
not ( n42998 , n42997 );
not ( n42999 , n42994 );
not ( n43000 , n42999 );
or ( n43001 , n42998 , n43000 );
nand ( n43002 , n43001 , n42965 );
nand ( n43003 , n42996 , n43002 );
xor ( n43004 , n42968 , n43003 );
not ( n43005 , n42992 );
not ( n43006 , n42980 );
or ( n43007 , n43005 , n43006 );
buf ( n43008 , n36435 );
buf ( n43009 , n505 );
and ( n43010 , n43008 , n43009 );
buf ( n43011 , n42952 );
buf ( n43012 , n489 );
and ( n43013 , n43011 , n43012 );
nor ( n43014 , n43010 , n43013 );
buf ( n43015 , n43014 );
not ( n43016 , n43015 );
nand ( n43017 , n43016 , n42975 );
nand ( n43018 , n43007 , n43017 );
buf ( n43019 , n43018 );
buf ( n43020 , n36435 );
buf ( n43021 , n33214 );
nor ( n43022 , n43020 , n43021 );
buf ( n43023 , n43022 );
buf ( n43024 , n43023 );
xor ( n43025 , n43019 , n43024 );
buf ( n43026 , n4519 );
not ( n43027 , n43026 );
buf ( n43028 , n43027 );
buf ( n43029 , n43028 );
not ( n43030 , n43029 );
buf ( n43031 , n42944 );
not ( n43032 , n43031 );
or ( n43033 , n43030 , n43032 );
buf ( n43034 , n491 );
nand ( n43035 , n43033 , n43034 );
buf ( n43036 , n43035 );
buf ( n43037 , n43036 );
xor ( n43038 , n43025 , n43037 );
buf ( n43039 , n43038 );
and ( n43040 , n43004 , n43039 );
and ( n43041 , n42968 , n43003 );
or ( n43042 , n43040 , n43041 );
not ( n43043 , n42992 );
or ( n43044 , n43015 , n43043 );
or ( n43045 , n42974 , n36435 );
nand ( n43046 , n43044 , n43045 );
buf ( n43047 , n43046 );
buf ( n43048 , n506 );
buf ( n43049 , n489 );
nand ( n43050 , n43048 , n43049 );
buf ( n43051 , n43050 );
buf ( n43052 , n43051 );
xor ( n43053 , n43047 , n43052 );
xor ( n43054 , n43019 , n43024 );
and ( n43055 , n43054 , n43037 );
and ( n43056 , n43019 , n43024 );
or ( n43057 , n43055 , n43056 );
buf ( n43058 , n43057 );
buf ( n43059 , n43058 );
xor ( n43060 , n43053 , n43059 );
buf ( n43061 , n43060 );
or ( n43062 , n43042 , n43061 );
not ( n43063 , n43062 );
xor ( n43064 , n40586 , n40606 );
and ( n43065 , n43064 , n40613 );
and ( n43066 , n40586 , n40606 );
or ( n43067 , n43065 , n43066 );
buf ( n43068 , n43067 );
buf ( n43069 , n43068 );
xor ( n43070 , n40530 , n40541 );
and ( n43071 , n43070 , n40559 );
and ( n43072 , n40530 , n40541 );
or ( n43073 , n43071 , n43072 );
buf ( n43074 , n43073 );
buf ( n43075 , n43074 );
and ( n43076 , n39847 , n39848 );
buf ( n43077 , n43076 );
buf ( n43078 , n43077 );
buf ( n43079 , n40602 );
xor ( n43080 , n43078 , n43079 );
buf ( n43081 , n40579 );
not ( n43082 , n43081 );
buf ( n43083 , n33438 );
not ( n43084 , n43083 );
or ( n43085 , n43082 , n43084 );
buf ( n43086 , n491 );
buf ( n43087 , n507 );
xnor ( n43088 , n43086 , n43087 );
buf ( n43089 , n43088 );
buf ( n43090 , n43089 );
not ( n43091 , n43090 );
buf ( n43092 , n4519 );
nand ( n43093 , n43091 , n43092 );
buf ( n43094 , n43093 );
buf ( n43095 , n43094 );
nand ( n43096 , n43085 , n43095 );
buf ( n43097 , n43096 );
buf ( n43098 , n43097 );
xor ( n43099 , n43080 , n43098 );
buf ( n43100 , n43099 );
buf ( n43101 , n43100 );
xor ( n43102 , n43075 , n43101 );
buf ( n43103 , n31271 );
not ( n43104 , n43103 );
buf ( n43105 , n43104 );
buf ( n43106 , n43105 );
not ( n43107 , n43106 );
buf ( n43108 , n2411 );
not ( n43109 , n43108 );
or ( n43110 , n43107 , n43109 );
buf ( n43111 , n495 );
nand ( n43112 , n43110 , n43111 );
buf ( n43113 , n43112 );
buf ( n43114 , n43113 );
buf ( n43115 , n40552 );
not ( n43116 , n43115 );
buf ( n43117 , n38410 );
not ( n43118 , n43117 );
or ( n43119 , n43116 , n43118 );
buf ( n43120 , n35832 );
buf ( n43121 , n489 );
buf ( n43122 , n509 );
xor ( n43123 , n43121 , n43122 );
buf ( n43124 , n43123 );
buf ( n43125 , n43124 );
nand ( n43126 , n43120 , n43125 );
buf ( n43127 , n43126 );
buf ( n43128 , n43127 );
nand ( n43129 , n43119 , n43128 );
buf ( n43130 , n43129 );
buf ( n43131 , n43130 );
xor ( n43132 , n43114 , n43131 );
buf ( n43133 , n40596 );
not ( n43134 , n43133 );
buf ( n43135 , n31660 );
not ( n43136 , n43135 );
or ( n43137 , n43134 , n43136 );
buf ( n43138 , n505 );
buf ( n43139 , n493 );
xnor ( n43140 , n43138 , n43139 );
buf ( n43141 , n43140 );
buf ( n43142 , n43141 );
not ( n43143 , n43142 );
buf ( n43144 , n2591 );
nand ( n43145 , n43143 , n43144 );
buf ( n43146 , n43145 );
buf ( n43147 , n43146 );
nand ( n43148 , n43137 , n43147 );
buf ( n43149 , n43148 );
buf ( n43150 , n43149 );
xor ( n43151 , n43132 , n43150 );
buf ( n43152 , n43151 );
buf ( n43153 , n43152 );
xor ( n43154 , n43102 , n43153 );
buf ( n43155 , n43154 );
buf ( n43156 , n43155 );
xor ( n43157 , n43069 , n43156 );
xor ( n43158 , n40562 , n40568 );
and ( n43159 , n43158 , n40616 );
and ( n43160 , n40562 , n40568 );
or ( n43161 , n43159 , n43160 );
buf ( n43162 , n43161 );
buf ( n43163 , n43162 );
xor ( n43164 , n43157 , n43163 );
buf ( n43165 , n43164 );
xor ( n43166 , n40520 , n40526 );
and ( n43167 , n43166 , n40619 );
and ( n43168 , n40520 , n40526 );
or ( n43169 , n43167 , n43168 );
buf ( n43170 , n43169 );
nor ( n43171 , n43165 , n43170 );
nor ( n43172 , n40622 , n43171 );
xor ( n43173 , n43078 , n43079 );
and ( n43174 , n43173 , n43098 );
and ( n43175 , n43078 , n43079 );
or ( n43176 , n43174 , n43175 );
buf ( n43177 , n43176 );
buf ( n43178 , n43177 );
buf ( n43179 , n31660 );
not ( n43180 , n43179 );
buf ( n43181 , n43180 );
buf ( n43182 , n43181 );
buf ( n43183 , n43141 );
or ( n43184 , n43182 , n43183 );
buf ( n43185 , n2591 );
not ( n43186 , n43185 );
buf ( n43187 , n43186 );
buf ( n43188 , n43187 );
buf ( n43189 , n493 );
not ( n43190 , n43189 );
buf ( n43191 , n43190 );
buf ( n43192 , n43191 );
or ( n43193 , n43188 , n43192 );
nand ( n43194 , n43184 , n43193 );
buf ( n43195 , n43194 );
buf ( n43196 , n43195 );
not ( n43197 , n43196 );
buf ( n43198 , n43197 );
buf ( n43199 , n43198 );
and ( n43200 , n40549 , n40550 );
buf ( n43201 , n43200 );
buf ( n43202 , n43201 );
buf ( n43203 , n43124 );
not ( n43204 , n43203 );
buf ( n43205 , n38410 );
not ( n43206 , n43205 );
or ( n43207 , n43204 , n43206 );
buf ( n43208 , n489 );
buf ( n43209 , n508 );
xnor ( n43210 , n43208 , n43209 );
buf ( n43211 , n43210 );
buf ( n43212 , n43211 );
not ( n43213 , n43212 );
buf ( n43214 , n35832 );
nand ( n43215 , n43213 , n43214 );
buf ( n43216 , n43215 );
buf ( n43217 , n43216 );
nand ( n43218 , n43207 , n43217 );
buf ( n43219 , n43218 );
buf ( n43220 , n43219 );
xor ( n43221 , n43202 , n43220 );
buf ( n43222 , n42944 );
buf ( n43223 , n43089 );
or ( n43224 , n43222 , n43223 );
buf ( n43225 , n43028 );
buf ( n43226 , n506 );
buf ( n43227 , n36583 );
and ( n43228 , n43226 , n43227 );
not ( n43229 , n43226 );
buf ( n43230 , n491 );
and ( n43231 , n43229 , n43230 );
nor ( n43232 , n43228 , n43231 );
buf ( n43233 , n43232 );
buf ( n43234 , n43233 );
or ( n43235 , n43225 , n43234 );
nand ( n43236 , n43224 , n43235 );
buf ( n43237 , n43236 );
buf ( n43238 , n43237 );
xor ( n43239 , n43221 , n43238 );
buf ( n43240 , n43239 );
buf ( n43241 , n43240 );
xor ( n43242 , n43199 , n43241 );
xor ( n43243 , n43114 , n43131 );
and ( n43244 , n43243 , n43150 );
and ( n43245 , n43114 , n43131 );
or ( n43246 , n43244 , n43245 );
buf ( n43247 , n43246 );
buf ( n43248 , n43247 );
xor ( n43249 , n43242 , n43248 );
buf ( n43250 , n43249 );
buf ( n43251 , n43250 );
xor ( n43252 , n43178 , n43251 );
xor ( n43253 , n43075 , n43101 );
and ( n43254 , n43253 , n43153 );
and ( n43255 , n43075 , n43101 );
or ( n43256 , n43254 , n43255 );
buf ( n43257 , n43256 );
buf ( n43258 , n43257 );
and ( n43259 , n43252 , n43258 );
and ( n43260 , n43178 , n43251 );
or ( n43261 , n43259 , n43260 );
buf ( n43262 , n43261 );
and ( n43263 , n43121 , n43122 );
buf ( n43264 , n43263 );
buf ( n43265 , n42944 );
buf ( n43266 , n43233 );
or ( n43267 , n43265 , n43266 );
buf ( n43268 , n43028 );
buf ( n43269 , n42957 );
or ( n43270 , n43268 , n43269 );
nand ( n43271 , n43267 , n43270 );
buf ( n43272 , n43271 );
not ( n43273 , n43272 );
xor ( n43274 , n43264 , n43273 );
buf ( n43275 , n43187 );
not ( n43276 , n43275 );
buf ( n43277 , n43181 );
not ( n43278 , n43277 );
or ( n43279 , n43276 , n43278 );
buf ( n43280 , n493 );
nand ( n43281 , n43279 , n43280 );
buf ( n43282 , n43281 );
xnor ( n43283 , n43274 , n43282 );
not ( n43284 , n42975 );
not ( n43285 , n42991 );
or ( n43286 , n43284 , n43285 );
not ( n43287 , n43211 );
nand ( n43288 , n43287 , n42992 );
nand ( n43289 , n43286 , n43288 );
buf ( n43290 , n43195 );
xor ( n43291 , n43289 , n43290 );
xor ( n43292 , n43202 , n43220 );
and ( n43293 , n43292 , n43238 );
and ( n43294 , n43202 , n43220 );
or ( n43295 , n43293 , n43294 );
buf ( n43296 , n43295 );
xor ( n43297 , n43291 , n43296 );
xor ( n43298 , n43283 , n43297 );
xor ( n43299 , n43199 , n43241 );
and ( n43300 , n43299 , n43248 );
and ( n43301 , n43199 , n43241 );
or ( n43302 , n43300 , n43301 );
buf ( n43303 , n43302 );
xor ( n43304 , n43298 , n43303 );
or ( n43305 , n43262 , n43304 );
xor ( n43306 , n43069 , n43156 );
and ( n43307 , n43306 , n43163 );
and ( n43308 , n43069 , n43156 );
or ( n43309 , n43307 , n43308 );
buf ( n43310 , n43309 );
xor ( n43311 , n43178 , n43251 );
xor ( n43312 , n43311 , n43258 );
buf ( n43313 , n43312 );
or ( n43314 , n43310 , n43313 );
nand ( n43315 , n43172 , n43305 , n43314 );
not ( n43316 , n43282 );
not ( n43317 , n43264 );
nand ( n43318 , n43317 , n43273 );
not ( n43319 , n43318 );
or ( n43320 , n43316 , n43319 );
nand ( n43321 , n43264 , n43272 );
nand ( n43322 , n43320 , n43321 );
not ( n43323 , n43289 );
not ( n43324 , n43323 );
not ( n43325 , n43324 );
not ( n43326 , n43290 );
or ( n43327 , n43325 , n43326 );
not ( n43328 , n43323 );
not ( n43329 , n43290 );
not ( n43330 , n43329 );
or ( n43331 , n43328 , n43330 );
nand ( n43332 , n43331 , n43296 );
nand ( n43333 , n43327 , n43332 );
xor ( n43334 , n43322 , n43333 );
xor ( n43335 , n42972 , n42999 );
xnor ( n43336 , n43335 , n42965 );
xor ( n43337 , n43334 , n43336 );
not ( n43338 , n43337 );
xor ( n43339 , n43283 , n43297 );
and ( n43340 , n43339 , n43303 );
and ( n43341 , n43283 , n43297 );
or ( n43342 , n43340 , n43341 );
not ( n43343 , n43342 );
nand ( n43344 , n43338 , n43343 );
xor ( n43345 , n42968 , n43003 );
xor ( n43346 , n43345 , n43039 );
not ( n43347 , n43346 );
not ( n43348 , n43336 );
nand ( n43349 , n43324 , n43290 );
nand ( n43350 , n43348 , n43332 , n43349 );
and ( n43351 , n43350 , n43322 );
nand ( n43352 , n43332 , n43349 );
and ( n43353 , n43336 , n43352 );
nor ( n43354 , n43351 , n43353 );
nand ( n43355 , n43347 , n43354 );
nand ( n43356 , n43344 , n43355 );
nor ( n43357 , n43315 , n43356 );
not ( n43358 , n43357 );
not ( n43359 , n40508 );
or ( n43360 , n43358 , n43359 );
not ( n43361 , n43347 );
not ( n43362 , n43354 );
and ( n43363 , n43361 , n43362 );
not ( n43364 , n43344 );
nand ( n43365 , n43262 , n43304 );
not ( n43366 , n43365 );
not ( n43367 , n43366 );
or ( n43368 , n43364 , n43367 );
not ( n43369 , n43343 );
nand ( n43370 , n43369 , n43337 );
nand ( n43371 , n43368 , n43370 );
not ( n43372 , n43371 );
nand ( n43373 , n43310 , n43313 );
not ( n43374 , n43373 );
or ( n43375 , n40624 , n43171 );
nand ( n43376 , n43165 , n43170 );
nand ( n43377 , n43375 , n43376 );
nand ( n43378 , n43314 , n43377 );
not ( n43379 , n43378 );
or ( n43380 , n43374 , n43379 );
and ( n43381 , n43305 , n43344 );
nand ( n43382 , n43380 , n43381 );
nand ( n43383 , n43372 , n43382 );
and ( n43384 , n43383 , n43355 );
nor ( n43385 , n43363 , n43384 );
nand ( n43386 , n43360 , n43385 );
not ( n43387 , n43386 );
or ( n43388 , n43063 , n43387 );
nand ( n43389 , n43042 , n43061 );
nand ( n43390 , n43388 , n43389 );
xor ( n43391 , n43047 , n43052 );
and ( n43392 , n43391 , n43059 );
and ( n43393 , n43047 , n43052 );
or ( n43394 , n43392 , n43393 );
buf ( n43395 , n43394 );
xor ( n43396 , n43395 , n43051 );
buf ( n43397 , n505 );
buf ( n43398 , n489 );
nand ( n43399 , n43397 , n43398 );
buf ( n43400 , n43399 );
buf ( n43401 , n43400 );
not ( n43402 , n43401 );
buf ( n43403 , n38410 );
buf ( n43404 , n35832 );
or ( n43405 , n43403 , n43404 );
buf ( n43406 , n489 );
nand ( n43407 , n43405 , n43406 );
buf ( n43408 , n43407 );
buf ( n43409 , n43408 );
not ( n43410 , n43409 );
or ( n43411 , n43402 , n43410 );
buf ( n43412 , n43408 );
buf ( n43413 , n43400 );
or ( n43414 , n43412 , n43413 );
nand ( n43415 , n43411 , n43414 );
buf ( n43416 , n43415 );
xnor ( n43417 , n43396 , n43416 );
and ( n43418 , n43390 , n43417 );
not ( n43419 , n43390 );
buf ( n43420 , n43051 );
not ( n43421 , n43420 );
buf ( n43422 , n43416 );
not ( n43423 , n43422 );
or ( n43424 , n43421 , n43423 );
buf ( n43425 , n43416 );
buf ( n43426 , n43051 );
or ( n43427 , n43425 , n43426 );
nand ( n43428 , n43424 , n43427 );
buf ( n43429 , n43428 );
xnor ( n43430 , n43395 , n43429 );
and ( n43431 , n43419 , n43430 );
nor ( n43432 , n43418 , n43431 );
not ( n43433 , n43432 );
or ( n43434 , n42941 , n43433 );
buf ( n43435 , n491 );
buf ( n43436 , n38013 );
and ( n43437 , n43435 , n43436 );
not ( n43438 , n43435 );
buf ( n43439 , n38013 );
not ( n43440 , n43439 );
buf ( n43441 , n43440 );
buf ( n43442 , n43441 );
and ( n43443 , n43438 , n43442 );
nor ( n43444 , n43437 , n43443 );
buf ( n43445 , n43444 );
buf ( n43446 , n43445 );
buf ( n43447 , n34031 );
and ( n43448 , n43446 , n43447 );
buf ( n43449 , n4821 );
buf ( n43450 , n491 );
and ( n43451 , n43449 , n43450 );
nor ( n43452 , n43448 , n43451 );
buf ( n43453 , n43452 );
buf ( n43454 , n43453 );
not ( n43455 , n43454 );
buf ( n43456 , n43455 );
buf ( n43457 , n43456 );
buf ( n43458 , n34031 );
buf ( n43459 , n4821 );
or ( n43460 , n43458 , n43459 );
buf ( n43461 , n491 );
nand ( n43462 , n43460 , n43461 );
buf ( n43463 , n43462 );
buf ( n43464 , n43463 );
buf ( n43465 , n489 );
not ( n43466 , n7585 );
buf ( n43467 , n43466 );
and ( n43468 , n43465 , n43467 );
buf ( n43469 , n43468 );
buf ( n43470 , n43469 );
xor ( n43471 , n43464 , n43470 );
buf ( n43472 , n37071 );
not ( n43473 , n43472 );
buf ( n43474 , n38228 );
buf ( n43475 , n7461 );
and ( n43476 , n43474 , n43475 );
buf ( n43477 , n38227 );
buf ( n43478 , n489 );
and ( n43479 , n43477 , n43478 );
nor ( n43480 , n43476 , n43479 );
buf ( n43481 , n43480 );
buf ( n43482 , n43481 );
not ( n43483 , n43482 );
buf ( n43484 , n43483 );
buf ( n43485 , n43484 );
not ( n43486 , n43485 );
or ( n43487 , n43473 , n43486 );
buf ( n43488 , n38013 );
buf ( n43489 , n7461 );
and ( n43490 , n43488 , n43489 );
buf ( n43491 , n43441 );
buf ( n43492 , n489 );
and ( n43493 , n43491 , n43492 );
nor ( n43494 , n43490 , n43493 );
buf ( n43495 , n43494 );
buf ( n43496 , n43495 );
buf ( n43497 , n7455 );
not ( n43498 , n43497 );
buf ( n43499 , n43498 );
buf ( n43500 , n43499 );
or ( n43501 , n43496 , n43500 );
nand ( n43502 , n43487 , n43501 );
buf ( n43503 , n43502 );
buf ( n43504 , n43503 );
xor ( n43505 , n43471 , n43504 );
buf ( n43506 , n43505 );
buf ( n43507 , n43506 );
xor ( n43508 , n43457 , n43507 );
buf ( n43509 , n43453 );
and ( n43510 , n489 , n39292 );
buf ( n43511 , n43510 );
xor ( n43512 , n43509 , n43511 );
buf ( n43513 , n37071 );
not ( n43514 , n43513 );
xor ( n43515 , n43465 , n43467 );
buf ( n43516 , n43515 );
buf ( n43517 , n43516 );
not ( n43518 , n43517 );
or ( n43519 , n43514 , n43518 );
buf ( n43520 , n43481 );
buf ( n43521 , n43499 );
or ( n43522 , n43520 , n43521 );
nand ( n43523 , n43519 , n43522 );
buf ( n43524 , n43523 );
buf ( n43525 , n43524 );
and ( n43526 , n43512 , n43525 );
and ( n43527 , n43509 , n43511 );
or ( n43528 , n43526 , n43527 );
buf ( n43529 , n43528 );
buf ( n43530 , n43529 );
and ( n43531 , n43508 , n43530 );
and ( n43532 , n43457 , n43507 );
or ( n43533 , n43531 , n43532 );
buf ( n43534 , n43533 );
buf ( n43535 , n43495 );
buf ( n43536 , n37071 );
not ( n43537 , n43536 );
buf ( n43538 , n43537 );
buf ( n43539 , n43538 );
or ( n43540 , n43535 , n43539 );
buf ( n43541 , n43499 );
buf ( n43542 , n7461 );
or ( n43543 , n43541 , n43542 );
nand ( n43544 , n43540 , n43543 );
buf ( n43545 , n43544 );
buf ( n43546 , n43545 );
buf ( n43547 , n38228 );
buf ( n43548 , n489 );
nand ( n43549 , n43547 , n43548 );
buf ( n43550 , n43549 );
buf ( n43551 , n43550 );
xor ( n43552 , n43546 , n43551 );
xor ( n43553 , n43464 , n43470 );
and ( n43554 , n43553 , n43504 );
and ( n43555 , n43464 , n43470 );
or ( n43556 , n43554 , n43555 );
buf ( n43557 , n43556 );
buf ( n43558 , n43557 );
xor ( n43559 , n43552 , n43558 );
buf ( n43560 , n43559 );
or ( n43561 , n43534 , n43560 );
not ( n43562 , n43561 );
xor ( n43563 , n40418 , n40446 );
and ( n43564 , n43563 , n40453 );
and ( n43565 , n40418 , n40446 );
or ( n43566 , n43564 , n43565 );
buf ( n43567 , n43566 );
buf ( n43568 , n43567 );
xor ( n43569 , n40358 , n40371 );
and ( n43570 , n43569 , n40386 );
and ( n43571 , n40358 , n40371 );
or ( n43572 , n43570 , n43571 );
buf ( n43573 , n43572 );
buf ( n43574 , n43573 );
buf ( n43575 , n29873 );
buf ( n43576 , n30072 );
or ( n43577 , n43575 , n43576 );
buf ( n43578 , n495 );
nand ( n43579 , n43577 , n43578 );
buf ( n43580 , n43579 );
buf ( n43581 , n43580 );
buf ( n43582 , n7455 );
not ( n43583 , n43582 );
buf ( n43584 , n489 );
buf ( n43585 , n39133 );
xor ( n43586 , n43584 , n43585 );
buf ( n43587 , n43586 );
buf ( n43588 , n43587 );
not ( n43589 , n43588 );
or ( n43590 , n43583 , n43589 );
buf ( n43591 , n40380 );
buf ( n43592 , n37071 );
nand ( n43593 , n43591 , n43592 );
buf ( n43594 , n43593 );
buf ( n43595 , n43594 );
nand ( n43596 , n43590 , n43595 );
buf ( n43597 , n43596 );
buf ( n43598 , n43597 );
xor ( n43599 , n43581 , n43598 );
buf ( n43600 , n39277 );
not ( n43601 , n43600 );
buf ( n43602 , n40432 );
not ( n43603 , n43602 );
or ( n43604 , n43601 , n43603 );
buf ( n43605 , n38013 );
buf ( n43606 , n29537 );
nand ( n43607 , n43605 , n43606 );
buf ( n43608 , n43607 );
nand ( n43609 , n38009 , n493 );
nand ( n43610 , n43608 , n43609 );
buf ( n43611 , n43610 );
buf ( n43612 , n29522 );
nand ( n43613 , n43611 , n43612 );
buf ( n43614 , n43613 );
buf ( n43615 , n43614 );
nand ( n43616 , n43604 , n43615 );
buf ( n43617 , n43616 );
buf ( n43618 , n43617 );
xor ( n43619 , n43599 , n43618 );
buf ( n43620 , n43619 );
buf ( n43621 , n43620 );
xor ( n43622 , n43574 , n43621 );
and ( n43623 , n489 , n40059 );
xor ( n43624 , n43623 , n40442 );
buf ( n43625 , n34031 );
not ( n43626 , n43625 );
buf ( n43627 , n40407 );
not ( n43628 , n43627 );
or ( n43629 , n43626 , n43628 );
buf ( n43630 , n491 );
not ( n43631 , n43630 );
buf ( n43632 , n7585 );
not ( n43633 , n43632 );
or ( n43634 , n43631 , n43633 );
buf ( n43635 , n43466 );
buf ( n43636 , n33936 );
nand ( n43637 , n43635 , n43636 );
buf ( n43638 , n43637 );
buf ( n43639 , n43638 );
nand ( n43640 , n43634 , n43639 );
buf ( n43641 , n43640 );
buf ( n43642 , n43641 );
buf ( n43643 , n4821 );
nand ( n43644 , n43642 , n43643 );
buf ( n43645 , n43644 );
buf ( n43646 , n43645 );
nand ( n43647 , n43629 , n43646 );
buf ( n43648 , n43647 );
xor ( n43649 , n43624 , n43648 );
buf ( n43650 , n43649 );
xor ( n43651 , n43622 , n43650 );
buf ( n43652 , n43651 );
buf ( n43653 , n43652 );
xor ( n43654 , n43568 , n43653 );
xor ( n43655 , n40389 , n40395 );
and ( n43656 , n43655 , n40456 );
and ( n43657 , n40389 , n40395 );
or ( n43658 , n43656 , n43657 );
buf ( n43659 , n43658 );
buf ( n43660 , n43659 );
and ( n43661 , n43654 , n43660 );
and ( n43662 , n43568 , n43653 );
or ( n43663 , n43661 , n43662 );
buf ( n43664 , n43663 );
xor ( n43665 , n43623 , n40442 );
and ( n43666 , n43665 , n43648 );
and ( n43667 , n43623 , n40442 );
or ( n43668 , n43666 , n43667 );
and ( n43669 , n39277 , n43610 );
and ( n43670 , n29522 , n493 );
nor ( n43671 , n43669 , n43670 );
buf ( n43672 , n43671 );
xor ( n43673 , n43581 , n43598 );
and ( n43674 , n43673 , n43618 );
and ( n43675 , n43581 , n43598 );
or ( n43676 , n43674 , n43675 );
buf ( n43677 , n43676 );
buf ( n43678 , n43677 );
xor ( n43679 , n43672 , n43678 );
and ( n43680 , n40376 , n40378 );
buf ( n43681 , n43680 );
buf ( n43682 , n43681 );
buf ( n43683 , n7455 );
not ( n43684 , n43683 );
xor ( n43685 , n489 , n39292 );
buf ( n43686 , n43685 );
not ( n43687 , n43686 );
or ( n43688 , n43684 , n43687 );
buf ( n43689 , n43587 );
buf ( n43690 , n37071 );
nand ( n43691 , n43689 , n43690 );
buf ( n43692 , n43691 );
buf ( n43693 , n43692 );
nand ( n43694 , n43688 , n43693 );
buf ( n43695 , n43694 );
buf ( n43696 , n43695 );
xor ( n43697 , n43682 , n43696 );
buf ( n43698 , n34031 );
not ( n43699 , n43698 );
buf ( n43700 , n43641 );
not ( n43701 , n43700 );
or ( n43702 , n43699 , n43701 );
and ( n43703 , n33936 , n38227 );
not ( n43704 , n33936 );
and ( n43705 , n43704 , n38228 );
nor ( n43706 , n43703 , n43705 );
buf ( n43707 , n43706 );
buf ( n43708 , n4821 );
nand ( n43709 , n43707 , n43708 );
buf ( n43710 , n43709 );
buf ( n43711 , n43710 );
nand ( n43712 , n43702 , n43711 );
buf ( n43713 , n43712 );
buf ( n43714 , n43713 );
xor ( n43715 , n43697 , n43714 );
buf ( n43716 , n43715 );
buf ( n43717 , n43716 );
xor ( n43718 , n43679 , n43717 );
buf ( n43719 , n43718 );
xor ( n43720 , n43668 , n43719 );
xor ( n43721 , n43574 , n43621 );
and ( n43722 , n43721 , n43650 );
and ( n43723 , n43574 , n43621 );
or ( n43724 , n43722 , n43723 );
buf ( n43725 , n43724 );
xor ( n43726 , n43720 , n43725 );
nor ( n43727 , n43664 , n43726 );
not ( n43728 , n43727 );
not ( n43729 , n40347 );
not ( n43730 , n40468 );
and ( n43731 , n43729 , n43730 );
xor ( n43732 , n43568 , n43653 );
xor ( n43733 , n43732 , n43660 );
buf ( n43734 , n43733 );
xor ( n43735 , n40353 , n40459 );
and ( n43736 , n43735 , n40466 );
and ( n43737 , n40353 , n40459 );
or ( n43738 , n43736 , n43737 );
buf ( n43739 , n43738 );
nor ( n43740 , n43734 , n43739 );
nor ( n43741 , n43731 , n43740 );
xor ( n43742 , n43672 , n43678 );
and ( n43743 , n43742 , n43717 );
and ( n43744 , n43672 , n43678 );
or ( n43745 , n43743 , n43744 );
buf ( n43746 , n43745 );
buf ( n43747 , n39277 );
buf ( n43748 , n29522 );
or ( n43749 , n43747 , n43748 );
buf ( n43750 , n493 );
nand ( n43751 , n43749 , n43750 );
buf ( n43752 , n43751 );
buf ( n43753 , n43752 );
and ( n43754 , n43584 , n43585 );
buf ( n43755 , n43754 );
buf ( n43756 , n43755 );
xor ( n43757 , n43753 , n43756 );
buf ( n43758 , n34031 );
not ( n43759 , n43758 );
buf ( n43760 , n43706 );
not ( n43761 , n43760 );
or ( n43762 , n43759 , n43761 );
buf ( n43763 , n43445 );
not ( n43764 , n43763 );
buf ( n43765 , n43764 );
buf ( n43766 , n43765 );
buf ( n43767 , n4821 );
not ( n43768 , n43767 );
buf ( n43769 , n43768 );
buf ( n43770 , n43769 );
or ( n43771 , n43766 , n43770 );
nand ( n43772 , n43762 , n43771 );
buf ( n43773 , n43772 );
buf ( n43774 , n43773 );
xor ( n43775 , n43757 , n43774 );
buf ( n43776 , n43775 );
xor ( n43777 , n43746 , n43776 );
buf ( n43778 , n43671 );
not ( n43779 , n43778 );
buf ( n43780 , n43779 );
buf ( n43781 , n43780 );
buf ( n43782 , n7455 );
not ( n43783 , n43782 );
buf ( n43784 , n43516 );
not ( n43785 , n43784 );
or ( n43786 , n43783 , n43785 );
buf ( n43787 , n43685 );
buf ( n43788 , n37071 );
nand ( n43789 , n43787 , n43788 );
buf ( n43790 , n43789 );
buf ( n43791 , n43790 );
nand ( n43792 , n43786 , n43791 );
buf ( n43793 , n43792 );
buf ( n43794 , n43793 );
xor ( n43795 , n43781 , n43794 );
xor ( n43796 , n43682 , n43696 );
and ( n43797 , n43796 , n43714 );
and ( n43798 , n43682 , n43696 );
or ( n43799 , n43797 , n43798 );
buf ( n43800 , n43799 );
buf ( n43801 , n43800 );
xor ( n43802 , n43795 , n43801 );
buf ( n43803 , n43802 );
xor ( n43804 , n43777 , n43803 );
xor ( n43805 , n43668 , n43719 );
and ( n43806 , n43805 , n43725 );
and ( n43807 , n43668 , n43719 );
or ( n43808 , n43806 , n43807 );
or ( n43809 , n43804 , n43808 );
nand ( n43810 , n43728 , n43741 , n43809 );
xor ( n43811 , n43746 , n43776 );
and ( n43812 , n43811 , n43803 );
and ( n43813 , n43746 , n43776 );
or ( n43814 , n43812 , n43813 );
not ( n43815 , n43814 );
xor ( n43816 , n43753 , n43756 );
and ( n43817 , n43816 , n43774 );
and ( n43818 , n43753 , n43756 );
or ( n43819 , n43817 , n43818 );
buf ( n43820 , n43819 );
xor ( n43821 , n43781 , n43794 );
and ( n43822 , n43821 , n43801 );
and ( n43823 , n43781 , n43794 );
or ( n43824 , n43822 , n43823 );
buf ( n43825 , n43824 );
xor ( n43826 , n43820 , n43825 );
xor ( n43827 , n43509 , n43511 );
xor ( n43828 , n43827 , n43525 );
buf ( n43829 , n43828 );
xnor ( n43830 , n43826 , n43829 );
nand ( n43831 , n43815 , n43830 );
xor ( n43832 , n43457 , n43507 );
xor ( n43833 , n43832 , n43530 );
buf ( n43834 , n43833 );
not ( n43835 , n43820 );
not ( n43836 , n43829 );
or ( n43837 , n43835 , n43836 );
or ( n43838 , n43829 , n43820 );
nand ( n43839 , n43838 , n43825 );
nand ( n43840 , n43837 , n43839 );
or ( n43841 , n43834 , n43840 );
nand ( n43842 , n43831 , n43841 );
nor ( n43843 , n43810 , n43842 );
not ( n43844 , n43843 );
not ( n43845 , n40325 );
not ( n43846 , n40336 );
or ( n43847 , n43845 , n43846 );
nand ( n43848 , n43847 , n40341 );
not ( n43849 , n43848 );
or ( n43850 , n43844 , n43849 );
not ( n43851 , n43727 );
not ( n43852 , n43851 );
or ( n43853 , n43740 , n40471 );
nand ( n43854 , n43734 , n43739 );
nand ( n43855 , n43853 , n43854 );
not ( n43856 , n43855 );
or ( n43857 , n43852 , n43856 );
nand ( n43858 , n43726 , n43664 );
nand ( n43859 , n43857 , n43858 );
nand ( n43860 , n43859 , n43809 , n43831 );
nand ( n43861 , n43804 , n43808 );
not ( n43862 , n43861 );
and ( n43863 , n43862 , n43831 );
not ( n43864 , n43830 );
nand ( n43865 , n43864 , n43814 );
not ( n43866 , n43865 );
nor ( n43867 , n43863 , n43866 );
nand ( n43868 , n43860 , n43867 );
and ( n43869 , n43868 , n43841 );
and ( n43870 , n43834 , n43840 );
nor ( n43871 , n43869 , n43870 );
nand ( n43872 , n43850 , n43871 );
not ( n43873 , n43872 );
or ( n43874 , n43562 , n43873 );
nand ( n43875 , n43534 , n43560 );
nand ( n43876 , n43874 , n43875 );
not ( n43877 , n43876 );
xor ( n43878 , n43546 , n43551 );
and ( n43879 , n43878 , n43558 );
and ( n43880 , n43546 , n43551 );
or ( n43881 , n43879 , n43880 );
buf ( n43882 , n43881 );
not ( n43883 , n43882 );
buf ( n43884 , n43550 );
not ( n43885 , n43884 );
buf ( n43886 , n38013 );
buf ( n43887 , n489 );
nand ( n43888 , n43886 , n43887 );
buf ( n43889 , n43888 );
buf ( n43890 , n43889 );
not ( n43891 , n43890 );
buf ( n43892 , n37071 );
buf ( n43893 , n7455 );
or ( n43894 , n43892 , n43893 );
buf ( n43895 , n489 );
nand ( n43896 , n43894 , n43895 );
buf ( n43897 , n43896 );
buf ( n43898 , n43897 );
not ( n43899 , n43898 );
or ( n43900 , n43891 , n43899 );
buf ( n43901 , n43897 );
buf ( n43902 , n43889 );
or ( n43903 , n43901 , n43902 );
nand ( n43904 , n43900 , n43903 );
buf ( n43905 , n43904 );
buf ( n43906 , n43905 );
not ( n43907 , n43906 );
or ( n43908 , n43885 , n43907 );
buf ( n43909 , n43905 );
buf ( n43910 , n43550 );
or ( n43911 , n43909 , n43910 );
nand ( n43912 , n43908 , n43911 );
buf ( n43913 , n43912 );
not ( n43914 , n43913 );
and ( n43915 , n43883 , n43914 );
and ( n43916 , n43882 , n43913 );
nor ( n43917 , n43915 , n43916 );
and ( n43918 , n455 , n43917 );
and ( n43919 , n43877 , n43918 );
not ( n43920 , n455 );
nor ( n43921 , n43920 , n43917 );
and ( n43922 , n43876 , n43921 );
nor ( n43923 , n43919 , n43922 );
nand ( n43924 , n43434 , n43923 );
not ( n43925 , n43924 );
or ( n43926 , n42940 , n43925 );
buf ( n43927 , n5582 );
not ( n43928 , n43927 );
buf ( n43929 , n43928 );
or ( n43930 , n43929 , n4173 );
nand ( n43931 , n43930 , n541 );
buf ( n43932 , n43931 );
buf ( n43933 , n6541 );
buf ( n43934 , n34557 );
nor ( n43935 , n43933 , n43934 );
buf ( n43936 , n43935 );
buf ( n43937 , n43936 );
xor ( n43938 , n43932 , n43937 );
buf ( n43939 , n6015 );
buf ( n43940 , n6001 );
buf ( n43941 , n522 );
and ( n43942 , n43940 , n43941 );
buf ( n43943 , n35199 );
buf ( n43944 , n539 );
and ( n43945 , n43943 , n43944 );
nor ( n43946 , n43942 , n43945 );
buf ( n43947 , n43946 );
buf ( n43948 , n43947 );
or ( n43949 , n43939 , n43948 );
buf ( n43950 , n6010 );
buf ( n43951 , n6001 );
buf ( n43952 , n521 );
and ( n43953 , n43951 , n43952 );
buf ( n43954 , n35343 );
buf ( n43955 , n539 );
and ( n43956 , n43954 , n43955 );
nor ( n43957 , n43953 , n43956 );
buf ( n43958 , n43957 );
buf ( n43959 , n43958 );
or ( n43960 , n43950 , n43959 );
nand ( n43961 , n43949 , n43960 );
buf ( n43962 , n43961 );
buf ( n43963 , n43962 );
xor ( n43964 , n43938 , n43963 );
buf ( n43965 , n43964 );
not ( n43966 , n43965 );
buf ( n43967 , n38773 );
buf ( n43968 , n6541 );
buf ( n43969 , n524 );
and ( n43970 , n43968 , n43969 );
buf ( n43971 , n34779 );
buf ( n43972 , n537 );
and ( n43973 , n43971 , n43972 );
nor ( n43974 , n43970 , n43973 );
buf ( n43975 , n43974 );
buf ( n43976 , n43975 );
or ( n43977 , n43967 , n43976 );
buf ( n43978 , n6337 );
buf ( n43979 , n6541 );
buf ( n43980 , n523 );
and ( n43981 , n43979 , n43980 );
buf ( n43982 , n35307 );
buf ( n43983 , n537 );
and ( n43984 , n43982 , n43983 );
nor ( n43985 , n43981 , n43984 );
buf ( n43986 , n43985 );
buf ( n43987 , n43986 );
or ( n43988 , n43978 , n43987 );
nand ( n43989 , n43977 , n43988 );
buf ( n43990 , n43989 );
buf ( n43991 , n43990 );
buf ( n43992 , n5582 );
buf ( n43993 , n541 );
buf ( n43994 , n35343 );
and ( n43995 , n43993 , n43994 );
not ( n43996 , n43993 );
buf ( n43997 , n521 );
and ( n43998 , n43996 , n43997 );
nor ( n43999 , n43995 , n43998 );
buf ( n44000 , n43999 );
buf ( n44001 , n44000 );
or ( n44002 , n43992 , n44001 );
buf ( n44003 , n33118 );
buf ( n44004 , n5578 );
or ( n44005 , n44003 , n44004 );
nand ( n44006 , n44002 , n44005 );
buf ( n44007 , n44006 );
buf ( n44008 , n44007 );
xor ( n44009 , n43991 , n44008 );
buf ( n44010 , n38773 );
buf ( n44011 , n6541 );
buf ( n44012 , n525 );
and ( n44013 , n44011 , n44012 );
buf ( n44014 , n34557 );
buf ( n44015 , n537 );
and ( n44016 , n44014 , n44015 );
nor ( n44017 , n44013 , n44016 );
buf ( n44018 , n44017 );
buf ( n44019 , n44018 );
or ( n44020 , n44010 , n44019 );
buf ( n44021 , n6337 );
buf ( n44022 , n43975 );
or ( n44023 , n44021 , n44022 );
nand ( n44024 , n44020 , n44023 );
buf ( n44025 , n44024 );
buf ( n44026 , n44025 );
buf ( n44027 , n526 );
not ( n44028 , n44027 );
buf ( n44029 , n6541 );
nor ( n44030 , n44028 , n44029 );
buf ( n44031 , n44030 );
buf ( n44032 , n44031 );
xor ( n44033 , n44026 , n44032 );
buf ( n44034 , n6015 );
buf ( n44035 , n523 );
buf ( n44036 , n6001 );
and ( n44037 , n44035 , n44036 );
not ( n44038 , n44035 );
buf ( n44039 , n539 );
and ( n44040 , n44038 , n44039 );
nor ( n44041 , n44037 , n44040 );
buf ( n44042 , n44041 );
buf ( n44043 , n44042 );
or ( n44044 , n44034 , n44043 );
buf ( n44045 , n6010 );
buf ( n44046 , n43947 );
or ( n44047 , n44045 , n44046 );
nand ( n44048 , n44044 , n44047 );
buf ( n44049 , n44048 );
buf ( n44050 , n44049 );
and ( n44051 , n44033 , n44050 );
and ( n44052 , n44026 , n44032 );
or ( n44053 , n44051 , n44052 );
buf ( n44054 , n44053 );
buf ( n44055 , n44054 );
xor ( n44056 , n44009 , n44055 );
buf ( n44057 , n44056 );
not ( n44058 , n44057 );
or ( n44059 , n43966 , n44058 );
or ( n44060 , n44057 , n43965 );
buf ( n44061 , n5582 );
buf ( n44062 , n541 );
buf ( n44063 , n35199 );
and ( n44064 , n44062 , n44063 );
not ( n44065 , n44062 );
buf ( n44066 , n522 );
and ( n44067 , n44065 , n44066 );
nor ( n44068 , n44064 , n44067 );
buf ( n44069 , n44068 );
buf ( n44070 , n44069 );
or ( n44071 , n44061 , n44070 );
buf ( n44072 , n33118 );
buf ( n44073 , n44000 );
or ( n44074 , n44072 , n44073 );
nand ( n44075 , n44071 , n44074 );
buf ( n44076 , n44075 );
buf ( n44077 , n44076 );
not ( n44078 , n4030 );
buf ( n44079 , n44078 );
buf ( n44080 , n32165 );
or ( n44081 , n44079 , n44080 );
buf ( n44082 , n543 );
nand ( n44083 , n44081 , n44082 );
buf ( n44084 , n44083 );
buf ( n44085 , n44084 );
xor ( n44086 , n44077 , n44085 );
buf ( n44087 , n38773 );
buf ( n44088 , n526 );
buf ( n44089 , n6541 );
and ( n44090 , n44088 , n44089 );
not ( n44091 , n44088 );
buf ( n44092 , n537 );
and ( n44093 , n44091 , n44092 );
nor ( n44094 , n44090 , n44093 );
buf ( n44095 , n44094 );
buf ( n44096 , n44095 );
or ( n44097 , n44087 , n44096 );
buf ( n44098 , n6337 );
buf ( n44099 , n44018 );
or ( n44100 , n44098 , n44099 );
nand ( n44101 , n44097 , n44100 );
buf ( n44102 , n44101 );
buf ( n44103 , n44102 );
and ( n44104 , n44086 , n44103 );
and ( n44105 , n44077 , n44085 );
or ( n44106 , n44104 , n44105 );
buf ( n44107 , n44106 );
buf ( n44108 , n44007 );
not ( n44109 , n44108 );
buf ( n44110 , n44109 );
xor ( n44111 , n44107 , n44110 );
xor ( n44112 , n44026 , n44032 );
xor ( n44113 , n44112 , n44050 );
buf ( n44114 , n44113 );
and ( n44115 , n44111 , n44114 );
and ( n44116 , n44107 , n44110 );
or ( n44117 , n44115 , n44116 );
nand ( n44118 , n44060 , n44117 );
nand ( n44119 , n44059 , n44118 );
nand ( n44120 , n44119 , n5847 );
buf ( n44121 , n38773 );
buf ( n44122 , n43986 );
or ( n44123 , n44121 , n44122 );
buf ( n44124 , n6337 );
buf ( n44125 , n6541 );
buf ( n44126 , n522 );
and ( n44127 , n44125 , n44126 );
buf ( n44128 , n35199 );
buf ( n44129 , n537 );
and ( n44130 , n44128 , n44129 );
nor ( n44131 , n44127 , n44130 );
buf ( n44132 , n44131 );
buf ( n44133 , n44132 );
or ( n44134 , n44124 , n44133 );
nand ( n44135 , n44123 , n44134 );
buf ( n44136 , n44135 );
buf ( n44137 , n44136 );
buf ( n44138 , n6541 );
buf ( n44139 , n34779 );
nor ( n44140 , n44138 , n44139 );
buf ( n44141 , n44140 );
buf ( n44142 , n44141 );
xor ( n44143 , n44137 , n44142 );
buf ( n44144 , n6016 );
buf ( n44145 , n43958 );
not ( n44146 , n44145 );
buf ( n44147 , n44146 );
buf ( n44148 , n44147 );
and ( n44149 , n44144 , n44148 );
buf ( n44150 , n6009 );
buf ( n44151 , n539 );
and ( n44152 , n44150 , n44151 );
nor ( n44153 , n44149 , n44152 );
buf ( n44154 , n44153 );
buf ( n44155 , n44154 );
xor ( n44156 , n44143 , n44155 );
buf ( n44157 , n44156 );
buf ( n44158 , n44157 );
xor ( n44159 , n43932 , n43937 );
and ( n44160 , n44159 , n43963 );
and ( n44161 , n43932 , n43937 );
or ( n44162 , n44160 , n44161 );
buf ( n44163 , n44162 );
buf ( n44164 , n44163 );
xor ( n44165 , n44158 , n44164 );
xor ( n44166 , n43991 , n44008 );
and ( n44167 , n44166 , n44055 );
and ( n44168 , n43991 , n44008 );
or ( n44169 , n44167 , n44168 );
buf ( n44170 , n44169 );
buf ( n44171 , n44170 );
xor ( n44172 , n44165 , n44171 );
buf ( n44173 , n44172 );
nand ( n44174 , n44173 , n3138 );
and ( n44175 , n44120 , n44174 );
nand ( n44176 , n43926 , n44175 );
not ( n44177 , n44176 );
xor ( n44178 , n44158 , n44164 );
and ( n44179 , n44178 , n44171 );
and ( n44180 , n44158 , n44164 );
or ( n44181 , n44179 , n44180 );
buf ( n44182 , n44181 );
nand ( n44183 , n44182 , n3360 );
xor ( n44184 , n44137 , n44142 );
and ( n44185 , n44184 , n44155 );
and ( n44186 , n44137 , n44142 );
or ( n44187 , n44185 , n44186 );
buf ( n44188 , n44187 );
buf ( n44189 , n44188 );
buf ( n44190 , n44154 );
not ( n44191 , n44190 );
buf ( n44192 , n44191 );
buf ( n44193 , n44192 );
xor ( n44194 , n44189 , n44193 );
buf ( n44195 , n38773 );
buf ( n44196 , n44132 );
or ( n44197 , n44195 , n44196 );
buf ( n44198 , n6337 );
buf ( n44199 , n6541 );
buf ( n44200 , n521 );
and ( n44201 , n44199 , n44200 );
buf ( n44202 , n35343 );
buf ( n44203 , n537 );
and ( n44204 , n44202 , n44203 );
nor ( n44205 , n44201 , n44204 );
buf ( n44206 , n44205 );
buf ( n44207 , n44206 );
or ( n44208 , n44198 , n44207 );
nand ( n44209 , n44197 , n44208 );
buf ( n44210 , n44209 );
buf ( n44211 , n44210 );
buf ( n44212 , n523 );
not ( n44213 , n44212 );
buf ( n44214 , n6541 );
nor ( n44215 , n44213 , n44214 );
buf ( n44216 , n44215 );
buf ( n44217 , n44216 );
xor ( n44218 , n44211 , n44217 );
buf ( n44219 , n6016 );
buf ( n44220 , n6009 );
or ( n44221 , n44219 , n44220 );
buf ( n44222 , n539 );
nand ( n44223 , n44221 , n44222 );
buf ( n44224 , n44223 );
buf ( n44225 , n44224 );
xor ( n44226 , n44218 , n44225 );
buf ( n44227 , n44226 );
buf ( n44228 , n44227 );
xor ( n44229 , n44194 , n44228 );
buf ( n44230 , n44229 );
nand ( n44231 , n44230 , n3138 );
and ( n44232 , n44183 , n44231 );
not ( n44233 , n44232 );
xor ( n44234 , n44189 , n44193 );
and ( n44235 , n44234 , n44228 );
and ( n44236 , n44189 , n44193 );
or ( n44237 , n44235 , n44236 );
buf ( n44238 , n44237 );
buf ( n44239 , n44238 );
buf ( n44240 , n3360 );
and ( n44241 , n44239 , n44240 );
buf ( n44242 , n44241 );
buf ( n44243 , n38773 );
buf ( n44244 , n44206 );
or ( n44245 , n44243 , n44244 );
buf ( n44246 , n6337 );
buf ( n44247 , n6541 );
or ( n44248 , n44246 , n44247 );
nand ( n44249 , n44245 , n44248 );
buf ( n44250 , n44249 );
buf ( n44251 , n44250 );
buf ( n44252 , n522 );
buf ( n44253 , n537 );
nand ( n44254 , n44252 , n44253 );
buf ( n44255 , n44254 );
buf ( n44256 , n44255 );
xor ( n44257 , n44251 , n44256 );
xor ( n44258 , n44211 , n44217 );
and ( n44259 , n44258 , n44225 );
and ( n44260 , n44211 , n44217 );
or ( n44261 , n44259 , n44260 );
buf ( n44262 , n44261 );
buf ( n44263 , n44262 );
xor ( n44264 , n44257 , n44263 );
buf ( n44265 , n44264 );
buf ( n44266 , n44265 );
buf ( n44267 , n3138 );
and ( n44268 , n44266 , n44267 );
buf ( n44269 , n44268 );
or ( n44270 , n44242 , n44269 );
nand ( n44271 , n44233 , n44270 );
nor ( n44272 , n44177 , n44271 );
buf ( n44273 , n4030 );
buf ( n44274 , n32981 );
buf ( n44275 , n522 );
and ( n44276 , n44274 , n44275 );
buf ( n44277 , n35199 );
buf ( n44278 , n543 );
and ( n44279 , n44277 , n44278 );
nor ( n44280 , n44276 , n44279 );
buf ( n44281 , n44280 );
buf ( n44282 , n44281 );
or ( n44283 , n44273 , n44282 );
buf ( n44284 , n4040 );
buf ( n44285 , n32981 );
buf ( n44286 , n521 );
and ( n44287 , n44285 , n44286 );
buf ( n44288 , n35343 );
buf ( n44289 , n543 );
and ( n44290 , n44288 , n44289 );
nor ( n44291 , n44287 , n44290 );
buf ( n44292 , n44291 );
buf ( n44293 , n44292 );
or ( n44294 , n44284 , n44293 );
nand ( n44295 , n44283 , n44294 );
buf ( n44296 , n44295 );
buf ( n44297 , n44296 );
not ( n44298 , n3064 );
not ( n44299 , n3069 );
or ( n44300 , n44298 , n44299 );
nand ( n44301 , n44300 , n545 );
buf ( n44302 , n44301 );
xor ( n44303 , n44297 , n44302 );
buf ( n44304 , n37557 );
buf ( n44305 , n6001 );
buf ( n44306 , n526 );
and ( n44307 , n44305 , n44306 );
buf ( n44308 , n40122 );
buf ( n44309 , n539 );
and ( n44310 , n44308 , n44309 );
nor ( n44311 , n44307 , n44310 );
buf ( n44312 , n44311 );
buf ( n44313 , n44312 );
or ( n44314 , n44304 , n44313 );
buf ( n44315 , n6010 );
buf ( n44316 , n6001 );
buf ( n44317 , n525 );
and ( n44318 , n44316 , n44317 );
buf ( n44319 , n34557 );
buf ( n44320 , n539 );
and ( n44321 , n44319 , n44320 );
nor ( n44322 , n44318 , n44321 );
buf ( n44323 , n44322 );
buf ( n44324 , n44323 );
or ( n44325 , n44315 , n44324 );
nand ( n44326 , n44314 , n44325 );
buf ( n44327 , n44326 );
buf ( n44328 , n44327 );
and ( n44329 , n44303 , n44328 );
and ( n44330 , n44297 , n44302 );
or ( n44331 , n44329 , n44330 );
buf ( n44332 , n44331 );
buf ( n44333 , n6559 );
buf ( n44334 , n6541 );
buf ( n44335 , n527 );
and ( n44336 , n44334 , n44335 );
buf ( n44337 , n33009 );
buf ( n44338 , n537 );
and ( n44339 , n44337 , n44338 );
nor ( n44340 , n44336 , n44339 );
buf ( n44341 , n44340 );
buf ( n44342 , n44341 );
or ( n44343 , n44333 , n44342 );
buf ( n44344 , n6337 );
buf ( n44345 , n44095 );
or ( n44346 , n44344 , n44345 );
nand ( n44347 , n44343 , n44346 );
buf ( n44348 , n44347 );
buf ( n44349 , n44348 );
buf ( n44350 , n6541 );
buf ( n44351 , n32183 );
nor ( n44352 , n44350 , n44351 );
buf ( n44353 , n44352 );
buf ( n44354 , n44353 );
xor ( n44355 , n44349 , n44354 );
buf ( n44356 , n543 );
not ( n44357 , n44356 );
buf ( n44358 , n32165 );
not ( n44359 , n44358 );
or ( n44360 , n44357 , n44359 );
buf ( n44361 , n5636 );
buf ( n44362 , n44292 );
or ( n44363 , n44361 , n44362 );
nand ( n44364 , n44360 , n44363 );
buf ( n44365 , n44364 );
buf ( n44366 , n44365 );
xor ( n44367 , n44355 , n44366 );
buf ( n44368 , n44367 );
xor ( n44369 , n44332 , n44368 );
buf ( n44370 , n6015 );
buf ( n44371 , n44323 );
or ( n44372 , n44370 , n44371 );
buf ( n44373 , n6010 );
buf ( n44374 , n6001 );
buf ( n44375 , n524 );
and ( n44376 , n44374 , n44375 );
buf ( n44377 , n34779 );
buf ( n44378 , n539 );
and ( n44379 , n44377 , n44378 );
nor ( n44380 , n44376 , n44379 );
buf ( n44381 , n44380 );
buf ( n44382 , n44381 );
or ( n44383 , n44373 , n44382 );
nand ( n44384 , n44372 , n44383 );
buf ( n44385 , n44384 );
buf ( n44386 , n44385 );
buf ( n44387 , n5582 );
buf ( n44388 , n541 );
buf ( n44389 , n35307 );
and ( n44390 , n44388 , n44389 );
not ( n44391 , n44388 );
buf ( n44392 , n523 );
and ( n44393 , n44391 , n44392 );
nor ( n44394 , n44390 , n44393 );
buf ( n44395 , n44394 );
buf ( n44396 , n44395 );
or ( n44397 , n44387 , n44396 );
buf ( n44398 , n33118 );
buf ( n44399 , n44069 );
or ( n44400 , n44398 , n44399 );
nand ( n44401 , n44397 , n44400 );
buf ( n44402 , n44401 );
buf ( n44403 , n44402 );
not ( n44404 , n44403 );
buf ( n44405 , n44404 );
buf ( n44406 , n44405 );
xor ( n44407 , n44386 , n44406 );
buf ( n44408 , n6559 );
buf ( n44409 , n6541 );
buf ( n44410 , n528 );
and ( n44411 , n44409 , n44410 );
buf ( n44412 , n32183 );
buf ( n44413 , n537 );
and ( n44414 , n44412 , n44413 );
nor ( n44415 , n44411 , n44414 );
buf ( n44416 , n44415 );
buf ( n44417 , n44416 );
or ( n44418 , n44408 , n44417 );
buf ( n44419 , n6337 );
buf ( n44420 , n44341 );
or ( n44421 , n44419 , n44420 );
nand ( n44422 , n44418 , n44421 );
buf ( n44423 , n44422 );
buf ( n44424 , n44423 );
buf ( n44425 , n529 );
buf ( n44426 , n537 );
and ( n44427 , n44425 , n44426 );
buf ( n44428 , n44427 );
buf ( n44429 , n44428 );
xor ( n44430 , n44424 , n44429 );
buf ( n44431 , n5582 );
buf ( n44432 , n541 );
buf ( n44433 , n34779 );
and ( n44434 , n44432 , n44433 );
not ( n44435 , n44432 );
buf ( n44436 , n524 );
and ( n44437 , n44435 , n44436 );
nor ( n44438 , n44434 , n44437 );
buf ( n44439 , n44438 );
buf ( n44440 , n44439 );
or ( n44441 , n44431 , n44440 );
buf ( n44442 , n33118 );
buf ( n44443 , n44395 );
or ( n44444 , n44442 , n44443 );
nand ( n44445 , n44441 , n44444 );
buf ( n44446 , n44445 );
buf ( n44447 , n44446 );
and ( n44448 , n44430 , n44447 );
and ( n44449 , n44424 , n44429 );
or ( n44450 , n44448 , n44449 );
buf ( n44451 , n44450 );
buf ( n44452 , n44451 );
xor ( n44453 , n44407 , n44452 );
buf ( n44454 , n44453 );
and ( n44455 , n44369 , n44454 );
and ( n44456 , n44332 , n44368 );
or ( n44457 , n44455 , n44456 );
buf ( n44458 , n44457 );
xor ( n44459 , n44386 , n44406 );
and ( n44460 , n44459 , n44452 );
and ( n44461 , n44386 , n44406 );
or ( n44462 , n44460 , n44461 );
buf ( n44463 , n44462 );
buf ( n44464 , n44463 );
xor ( n44465 , n44458 , n44464 );
buf ( n44466 , n6541 );
buf ( n44467 , n33009 );
nor ( n44468 , n44466 , n44467 );
buf ( n44469 , n44468 );
xor ( n44470 , n44402 , n44469 );
buf ( n44471 , n6015 );
buf ( n44472 , n44381 );
or ( n44473 , n44471 , n44472 );
buf ( n44474 , n6010 );
buf ( n44475 , n44042 );
or ( n44476 , n44474 , n44475 );
nand ( n44477 , n44473 , n44476 );
buf ( n44478 , n44477 );
xor ( n44479 , n44470 , n44478 );
xor ( n44480 , n44349 , n44354 );
and ( n44481 , n44480 , n44366 );
and ( n44482 , n44349 , n44354 );
or ( n44483 , n44481 , n44482 );
buf ( n44484 , n44483 );
xor ( n44485 , n44077 , n44085 );
xor ( n44486 , n44485 , n44103 );
buf ( n44487 , n44486 );
xor ( n44488 , n44484 , n44487 );
xor ( n44489 , n44479 , n44488 );
buf ( n44490 , n44489 );
and ( n44491 , n44465 , n44490 );
and ( n44492 , n44458 , n44464 );
or ( n44493 , n44491 , n44492 );
buf ( n44494 , n44493 );
buf ( n44495 , n44494 );
buf ( n44496 , n3360 );
and ( n44497 , n44495 , n44496 );
buf ( n44498 , n44497 );
xor ( n44499 , n44107 , n44110 );
xor ( n44500 , n44499 , n44114 );
xor ( n44501 , n44402 , n44469 );
and ( n44502 , n44501 , n44478 );
and ( n44503 , n44402 , n44469 );
or ( n44504 , n44502 , n44503 );
xor ( n44505 , n44402 , n44469 );
xor ( n44506 , n44505 , n44478 );
and ( n44507 , n44484 , n44506 );
xor ( n44508 , n44402 , n44469 );
xor ( n44509 , n44508 , n44478 );
and ( n44510 , n44487 , n44509 );
and ( n44511 , n44484 , n44487 );
or ( n44512 , n44507 , n44510 , n44511 );
xor ( n44513 , n44504 , n44512 );
xor ( n44514 , n44500 , n44513 );
and ( n44515 , n44514 , n3138 );
nor ( n44516 , n44498 , n44515 );
not ( n44517 , n44516 );
not ( n44518 , n43344 );
not ( n44519 , n43354 );
not ( n44520 , n43347 );
or ( n44521 , n44519 , n44520 );
or ( n44522 , n43347 , n43354 );
nand ( n44523 , n44521 , n44522 );
nor ( n44524 , n44518 , n44523 );
not ( n44525 , n44524 );
not ( n44526 , n44525 );
not ( n44527 , n40483 );
not ( n44528 , n38272 );
or ( n44529 , n44527 , n44528 );
nand ( n44530 , n44529 , n40507 );
not ( n44531 , n43315 );
nand ( n44532 , n44530 , n44531 );
not ( n44533 , n44532 );
and ( n44534 , n44526 , n44533 );
not ( n44535 , n43383 );
and ( n44536 , n44535 , n44523 );
and ( n44537 , n44532 , n44536 );
nor ( n44538 , n44534 , n44537 );
not ( n44539 , n44523 );
or ( n44540 , n44539 , n43344 );
nand ( n44541 , n44540 , n29516 );
not ( n44542 , n44541 );
not ( n44543 , n44542 );
not ( n44544 , n44535 );
or ( n44545 , n44543 , n44544 );
not ( n44546 , n29516 );
nor ( n44547 , n44546 , n44539 );
nand ( n44548 , n43383 , n44547 );
nand ( n44549 , n44545 , n44548 );
nand ( n44550 , n44538 , n44549 );
not ( n44551 , n43870 );
nand ( n44552 , n44551 , n43841 );
not ( n44553 , n44552 );
not ( n44554 , n43831 );
nor ( n44555 , n44554 , n43810 );
not ( n44556 , n44555 );
not ( n44557 , n43848 );
or ( n44558 , n44556 , n44557 );
not ( n44559 , n43868 );
nand ( n44560 , n44558 , n44559 );
not ( n44561 , n44560 );
not ( n44562 , n44561 );
or ( n44563 , n44553 , n44562 );
not ( n44564 , n44552 );
and ( n44565 , n44560 , n44564 );
nor ( n44566 , n44565 , n29516 );
nand ( n44567 , n44563 , n44566 );
nand ( n44568 , n44550 , n44567 );
nand ( n44569 , n44568 , n454 );
not ( n44570 , n44569 );
or ( n44571 , n44517 , n44570 );
not ( n44572 , n454 );
not ( n44573 , n2815 );
nand ( n44574 , n43062 , n43389 );
not ( n44575 , n44574 );
and ( n44576 , n43386 , n44575 );
not ( n44577 , n43386 );
and ( n44578 , n44577 , n44574 );
nor ( n44579 , n44576 , n44578 );
not ( n44580 , n44579 );
or ( n44581 , n44573 , n44580 );
nand ( n44582 , n43561 , n43875 );
and ( n44583 , n455 , n44582 );
and ( n44584 , n43872 , n44583 );
not ( n44585 , n43872 );
not ( n44586 , n455 );
nor ( n44587 , n44586 , n44582 );
and ( n44588 , n44585 , n44587 );
nor ( n44589 , n44584 , n44588 );
nand ( n44590 , n44581 , n44589 );
not ( n44591 , n44590 );
or ( n44592 , n44572 , n44591 );
xor ( n44593 , n43965 , n44057 );
xor ( n44594 , n44593 , n44117 );
nand ( n44595 , n44594 , n3138 );
xor ( n44596 , n44107 , n44110 );
xor ( n44597 , n44596 , n44114 );
and ( n44598 , n44504 , n44597 );
xor ( n44599 , n44107 , n44110 );
xor ( n44600 , n44599 , n44114 );
and ( n44601 , n44512 , n44600 );
and ( n44602 , n44504 , n44512 );
or ( n44603 , n44598 , n44601 , n44602 );
nand ( n44604 , n44603 , n3360 );
and ( n44605 , n44595 , n44604 );
nand ( n44606 , n44592 , n44605 );
nand ( n44607 , n44571 , n44606 );
not ( n44608 , n44607 );
nand ( n44609 , n44530 , n43172 );
not ( n44610 , n44609 );
not ( n44611 , n43365 );
not ( n44612 , n43305 );
or ( n44613 , n44611 , n44612 );
nand ( n44614 , n44613 , n29516 );
not ( n44615 , n44614 );
not ( n44616 , n44615 );
nand ( n44617 , n43378 , n43373 );
not ( n44618 , n44617 );
not ( n44619 , n44618 );
not ( n44620 , n44619 );
and ( n44621 , n44616 , n44620 );
not ( n44622 , n43314 );
and ( n44623 , n44622 , n44618 );
not ( n44624 , n44623 );
not ( n44625 , n44614 );
or ( n44626 , n44624 , n44625 );
not ( n44627 , n43304 );
not ( n44628 , n43262 );
or ( n44629 , n44627 , n44628 );
or ( n44630 , n43262 , n43304 );
nand ( n44631 , n44629 , n44630 );
or ( n44632 , n44631 , n455 );
nand ( n44633 , n44632 , n44619 );
nand ( n44634 , n44626 , n44633 );
nor ( n44635 , n44621 , n44634 );
not ( n44636 , n44635 );
or ( n44637 , n44610 , n44636 );
not ( n44638 , n44634 );
not ( n44639 , n44609 );
nand ( n44640 , n44632 , n43314 );
nand ( n44641 , n44638 , n44639 , n44640 );
nand ( n44642 , n44637 , n44641 );
not ( n44643 , n43859 );
nand ( n44644 , n43809 , n43861 );
nand ( n44645 , n44643 , n44644 , n455 );
not ( n44646 , n44645 );
nand ( n44647 , n43809 , n43861 , n455 );
not ( n44648 , n44647 );
and ( n44649 , n44648 , n43859 );
nor ( n44650 , n44649 , n5847 );
not ( n44651 , n44650 );
or ( n44652 , n44646 , n44651 );
not ( n44653 , n43851 );
nor ( n44654 , n44653 , n40469 , n43740 );
nand ( n44655 , n40342 , n44650 , n44654 );
nand ( n44656 , n44652 , n44655 );
not ( n44657 , n44654 );
nor ( n44658 , n44657 , n44647 );
nand ( n44659 , n40342 , n44658 );
nand ( n44660 , n44656 , n44659 );
or ( n44661 , n44642 , n44660 );
xor ( n44662 , n44297 , n44302 );
xor ( n44663 , n44662 , n44328 );
buf ( n44664 , n44663 );
buf ( n44665 , n44664 );
buf ( n44666 , n5582 );
buf ( n44667 , n40754 );
or ( n44668 , n44666 , n44667 );
buf ( n44669 , n33118 );
buf ( n44670 , n44439 );
or ( n44671 , n44669 , n44670 );
nand ( n44672 , n44668 , n44671 );
buf ( n44673 , n44672 );
buf ( n44674 , n44673 );
buf ( n44675 , n6541 );
buf ( n44676 , n31853 );
nor ( n44677 , n44675 , n44676 );
buf ( n44678 , n44677 );
buf ( n44679 , n44678 );
xor ( n44680 , n44674 , n44679 );
buf ( n44681 , n4030 );
buf ( n44682 , n40700 );
or ( n44683 , n44681 , n44682 );
buf ( n44684 , n35070 );
buf ( n44685 , n44281 );
or ( n44686 , n44684 , n44685 );
nand ( n44687 , n44683 , n44686 );
buf ( n44688 , n44687 );
buf ( n44689 , n44688 );
not ( n44690 , n44689 );
buf ( n44691 , n44690 );
buf ( n44692 , n44691 );
and ( n44693 , n44680 , n44692 );
and ( n44694 , n44674 , n44679 );
or ( n44695 , n44693 , n44694 );
buf ( n44696 , n44695 );
buf ( n44697 , n44696 );
xor ( n44698 , n44665 , n44697 );
buf ( n44699 , n6015 );
buf ( n44700 , n40683 );
or ( n44701 , n44699 , n44700 );
buf ( n44702 , n6010 );
buf ( n44703 , n44312 );
or ( n44704 , n44702 , n44703 );
nand ( n44705 , n44701 , n44704 );
buf ( n44706 , n44705 );
buf ( n44707 , n44706 );
buf ( n44708 , n6559 );
buf ( n44709 , n40718 );
or ( n44710 , n44708 , n44709 );
buf ( n44711 , n6337 );
buf ( n44712 , n44416 );
or ( n44713 , n44711 , n44712 );
nand ( n44714 , n44710 , n44713 );
buf ( n44715 , n44714 );
buf ( n44716 , n44715 );
xor ( n44717 , n44707 , n44716 );
buf ( n44718 , n545 );
not ( n44719 , n44718 );
buf ( n44720 , n3063 );
not ( n44721 , n44720 );
or ( n44722 , n44719 , n44721 );
buf ( n44723 , n3069 );
buf ( n44724 , n40772 );
or ( n44725 , n44723 , n44724 );
nand ( n44726 , n44722 , n44725 );
buf ( n44727 , n44726 );
buf ( n44728 , n44727 );
and ( n44729 , n44717 , n44728 );
and ( n44730 , n44707 , n44716 );
or ( n44731 , n44729 , n44730 );
buf ( n44732 , n44731 );
buf ( n44733 , n44732 );
buf ( n44734 , n44688 );
xor ( n44735 , n44733 , n44734 );
xor ( n44736 , n44424 , n44429 );
xor ( n44737 , n44736 , n44447 );
buf ( n44738 , n44737 );
buf ( n44739 , n44738 );
xor ( n44740 , n44735 , n44739 );
buf ( n44741 , n44740 );
buf ( n44742 , n44741 );
xor ( n44743 , n44698 , n44742 );
buf ( n44744 , n44743 );
buf ( n44745 , n44744 );
xor ( n44746 , n40688 , n40705 );
and ( n44747 , n44746 , n40723 );
and ( n44748 , n40688 , n40705 );
or ( n44749 , n44747 , n44748 );
buf ( n44750 , n44749 );
buf ( n44751 , n44750 );
xor ( n44752 , n44707 , n44716 );
xor ( n44753 , n44752 , n44728 );
buf ( n44754 , n44753 );
buf ( n44755 , n44754 );
xor ( n44756 , n44751 , n44755 );
xor ( n44757 , n40742 , n40759 );
and ( n44758 , n44757 , n40777 );
and ( n44759 , n40742 , n40759 );
or ( n44760 , n44758 , n44759 );
buf ( n44761 , n44760 );
buf ( n44762 , n44761 );
and ( n44763 , n44756 , n44762 );
and ( n44764 , n44751 , n44755 );
or ( n44765 , n44763 , n44764 );
buf ( n44766 , n44765 );
buf ( n44767 , n44766 );
xor ( n44768 , n44745 , n44767 );
xor ( n44769 , n40656 , n40661 );
and ( n44770 , n44769 , n40667 );
and ( n44771 , n40656 , n40661 );
or ( n44772 , n44770 , n44771 );
buf ( n44773 , n44772 );
xor ( n44774 , n44674 , n44679 );
xor ( n44775 , n44774 , n44692 );
buf ( n44776 , n44775 );
xor ( n44777 , n44773 , n44776 );
xor ( n44778 , n40726 , n40732 );
and ( n44779 , n44778 , n40780 );
and ( n44780 , n40726 , n40732 );
or ( n44781 , n44779 , n44780 );
buf ( n44782 , n44781 );
and ( n44783 , n44777 , n44782 );
and ( n44784 , n44773 , n44776 );
or ( n44785 , n44783 , n44784 );
buf ( n44786 , n44785 );
and ( n44787 , n44768 , n44786 );
and ( n44788 , n44745 , n44767 );
or ( n44789 , n44787 , n44788 );
buf ( n44790 , n44789 );
buf ( n44791 , n44790 );
buf ( n44792 , n3138 );
nand ( n44793 , n44791 , n44792 );
buf ( n44794 , n44793 );
nand ( n44795 , n44661 , n44794 );
not ( n44796 , n44795 );
xor ( n44797 , n44332 , n44368 );
xor ( n44798 , n44797 , n44454 );
xor ( n44799 , n44733 , n44734 );
and ( n44800 , n44799 , n44739 );
and ( n44801 , n44733 , n44734 );
or ( n44802 , n44800 , n44801 );
buf ( n44803 , n44802 );
xor ( n44804 , n44665 , n44697 );
and ( n44805 , n44804 , n44742 );
and ( n44806 , n44665 , n44697 );
or ( n44807 , n44805 , n44806 );
buf ( n44808 , n44807 );
xor ( n44809 , n44803 , n44808 );
xor ( n44810 , n44798 , n44809 );
buf ( n44811 , n44810 );
not ( n44812 , n44811 );
buf ( n44813 , n454 );
nor ( n44814 , n44812 , n44813 );
buf ( n44815 , n44814 );
not ( n44816 , n44815 );
and ( n44817 , n44796 , n44816 );
not ( n44818 , n43305 );
not ( n44819 , n44617 );
or ( n44820 , n44818 , n44819 );
nand ( n44821 , n44820 , n43365 );
not ( n44822 , n44821 );
nand ( n44823 , n44822 , n44532 );
nand ( n44824 , n43344 , n43370 );
and ( n44825 , n44823 , n44824 );
not ( n44826 , n44823 );
not ( n44827 , n44824 );
and ( n44828 , n44826 , n44827 );
nor ( n44829 , n44825 , n44828 );
and ( n44830 , n44829 , n2815 );
nor ( n44831 , n44830 , n5847 );
not ( n44832 , n43810 );
not ( n44833 , n44832 );
not ( n44834 , n40342 );
or ( n44835 , n44833 , n44834 );
not ( n44836 , n43809 );
not ( n44837 , n43859 );
or ( n44838 , n44836 , n44837 );
nand ( n44839 , n44838 , n43861 );
not ( n44840 , n44839 );
nand ( n44841 , n44835 , n44840 );
nand ( n44842 , n43831 , n43865 );
and ( n44843 , n44841 , n44842 );
not ( n44844 , n44841 );
not ( n44845 , n44842 );
and ( n44846 , n44844 , n44845 );
nor ( n44847 , n44843 , n44846 );
nand ( n44848 , n44847 , n455 );
nand ( n44849 , n44831 , n44848 );
xor ( n44850 , n44458 , n44464 );
xor ( n44851 , n44850 , n44490 );
buf ( n44852 , n44851 );
buf ( n44853 , n44852 );
buf ( n44854 , n3138 );
nand ( n44855 , n44853 , n44854 );
buf ( n44856 , n44855 );
not ( n44857 , n44856 );
xor ( n44858 , n44332 , n44368 );
xor ( n44859 , n44858 , n44454 );
and ( n44860 , n44803 , n44859 );
xor ( n44861 , n44332 , n44368 );
xor ( n44862 , n44861 , n44454 );
and ( n44863 , n44808 , n44862 );
and ( n44864 , n44803 , n44808 );
or ( n44865 , n44860 , n44863 , n44864 );
not ( n44866 , n44865 );
nor ( n44867 , n44866 , n454 );
nor ( n44868 , n44857 , n44867 );
and ( n44869 , n44849 , n44868 );
nor ( n44870 , n44817 , n44869 );
nand ( n44871 , n44608 , n44870 );
not ( n44872 , n44871 );
and ( n44873 , n44272 , n44872 );
not ( n44874 , n40098 );
not ( n44875 , n40258 );
and ( n44876 , n44874 , n44875 );
nor ( n44877 , n40802 , n40805 );
and ( n44878 , n40808 , n44877 );
nor ( n44879 , n44876 , n44878 );
not ( n44880 , n43740 );
nand ( n44881 , n44880 , n43854 );
and ( n44882 , n455 , n44881 , n454 );
not ( n44883 , n44882 );
not ( n44884 , n40470 );
not ( n44885 , n43848 );
or ( n44886 , n44884 , n44885 );
buf ( n44887 , n40471 );
nand ( n44888 , n44886 , n44887 );
not ( n44889 , n44888 );
or ( n44890 , n44883 , n44889 );
xor ( n44891 , n44773 , n44776 );
xor ( n44892 , n44891 , n44782 );
xor ( n44893 , n44751 , n44755 );
xor ( n44894 , n44893 , n44762 );
buf ( n44895 , n44894 );
xor ( n44896 , n40655 , n40670 );
and ( n44897 , n44896 , n40783 );
and ( n44898 , n40655 , n40670 );
or ( n44899 , n44897 , n44898 );
buf ( n44900 , n44899 );
xor ( n44901 , n44895 , n44900 );
xor ( n44902 , n44892 , n44901 );
nand ( n44903 , n44902 , n3138 );
nand ( n44904 , n44890 , n44903 );
nand ( n44905 , n40786 , n40649 );
not ( n44906 , n44905 );
not ( n44907 , n40639 );
or ( n44908 , n44906 , n44907 );
nand ( n44909 , n40787 , n40648 );
nand ( n44910 , n44908 , n44909 );
nand ( n44911 , n44910 , n3360 );
not ( n44912 , n44911 );
nor ( n44913 , n44904 , n44912 );
not ( n44914 , n2815 );
not ( n44915 , n43171 );
nand ( n44916 , n44915 , n43376 );
not ( n44917 , n40623 );
not ( n44918 , n44530 );
or ( n44919 , n44917 , n44918 );
nand ( n44920 , n44919 , n40624 );
nor ( n44921 , n44914 , n44916 , n44920 );
not ( n44922 , n44881 );
nand ( n44923 , n44922 , n455 );
not ( n44924 , n44923 );
not ( n44925 , n44924 );
not ( n44926 , n44888 );
not ( n44927 , n44926 );
or ( n44928 , n44925 , n44927 );
nand ( n44929 , n44920 , n44916 , n2815 );
nand ( n44930 , n44928 , n44929 );
or ( n44931 , n44921 , n44930 );
nand ( n44932 , n44931 , n454 );
nand ( n44933 , n44913 , n44932 );
not ( n44934 , n454 );
not ( n44935 , n43741 );
not ( n44936 , n43848 );
or ( n44937 , n44935 , n44936 );
not ( n44938 , n43855 );
nand ( n44939 , n44937 , n44938 );
nand ( n44940 , n43851 , n43858 );
and ( n44941 , n44940 , n455 );
and ( n44942 , n44939 , n44941 );
not ( n44943 , n44939 );
not ( n44944 , n455 );
nor ( n44945 , n44944 , n44940 );
and ( n44946 , n44943 , n44945 );
nor ( n44947 , n44942 , n44946 );
nand ( n44948 , n43314 , n43373 );
and ( n44949 , n44948 , n2815 );
buf ( n44950 , n43377 );
and ( n44951 , n44949 , n44950 );
nor ( n44952 , n44948 , n44950 , n455 );
nor ( n44953 , n44951 , n44952 );
not ( n44954 , n44953 );
not ( n44955 , n44609 );
or ( n44956 , n44954 , n44955 );
not ( n44957 , n44639 );
or ( n44958 , n44957 , n44949 );
nand ( n44959 , n44956 , n44958 );
nand ( n44960 , n44947 , n44959 );
not ( n44961 , n44960 );
or ( n44962 , n44934 , n44961 );
xor ( n44963 , n44745 , n44767 );
xor ( n44964 , n44963 , n44786 );
buf ( n44965 , n44964 );
not ( n44966 , n44965 );
nor ( n44967 , n44966 , n454 );
xor ( n44968 , n44773 , n44776 );
xor ( n44969 , n44968 , n44782 );
and ( n44970 , n44895 , n44969 );
xor ( n44971 , n44773 , n44776 );
xor ( n44972 , n44971 , n44782 );
and ( n44973 , n44900 , n44972 );
and ( n44974 , n44895 , n44900 );
or ( n44975 , n44970 , n44973 , n44974 );
nand ( n44976 , n44975 , n3138 );
not ( n44977 , n44976 );
nor ( n44978 , n44967 , n44977 );
nand ( n44979 , n44962 , n44978 );
and ( n44980 , n44879 , n44933 , n44979 );
nand ( n44981 , n39749 , n44980 );
not ( n44982 , n44981 );
not ( n44983 , n40936 );
nand ( n44984 , n44873 , n44982 , n44983 );
nand ( n44985 , n3710 , n3759 );
nand ( n44986 , n3754 , n44985 );
not ( n44987 , n44986 );
nand ( n44988 , n32766 , n3803 );
not ( n44989 , n44988 );
or ( n44990 , n44987 , n44989 );
or ( n44991 , n44986 , n44988 );
nand ( n44992 , n44990 , n44991 );
not ( n44993 , n3710 );
nand ( n44994 , n3759 , n3754 );
not ( n44995 , n44994 );
or ( n44996 , n44993 , n44995 );
or ( n44997 , n3710 , n44994 );
nand ( n44998 , n44996 , n44997 );
not ( n44999 , n44607 );
not ( n45000 , n44999 );
nand ( n45001 , n44815 , n44795 );
not ( n45002 , n45001 );
not ( n45003 , n45002 );
not ( n45004 , n44848 );
and ( n45005 , n44829 , n2815 );
nor ( n45006 , n45005 , n5847 );
not ( n45007 , n45006 );
or ( n45008 , n45004 , n45007 );
not ( n45009 , n44867 );
and ( n45010 , n45009 , n44856 );
nand ( n45011 , n45008 , n45010 );
not ( n45012 , n45011 );
or ( n45013 , n45003 , n45012 );
not ( n45014 , n44856 );
not ( n45015 , n44831 );
not ( n45016 , n45015 );
or ( n45017 , n45014 , n45016 );
and ( n45018 , n44847 , n44856 , n455 );
nor ( n45019 , n45018 , n45009 );
nand ( n45020 , n45017 , n45019 );
nand ( n45021 , n45013 , n45020 );
not ( n45022 , n45021 );
or ( n45023 , n45000 , n45022 );
not ( n45024 , n454 );
not ( n45025 , n44590 );
or ( n45026 , n45024 , n45025 );
and ( n45027 , n44604 , n44595 );
nand ( n45028 , n45026 , n45027 );
nand ( n45029 , n44514 , n3138 );
nand ( n45030 , n44550 , n44567 , n45029 );
not ( n45031 , n454 );
nand ( n45032 , n45031 , n45029 );
and ( n45033 , n45032 , n44498 );
nand ( n45034 , n45030 , n45033 );
not ( n45035 , n45034 );
and ( n45036 , n45028 , n45035 );
not ( n45037 , n454 );
not ( n45038 , n44590 );
or ( n45039 , n45037 , n45038 );
nand ( n45040 , n45039 , n44595 );
not ( n45041 , n44604 );
and ( n45042 , n45040 , n45041 );
nor ( n45043 , n45036 , n45042 );
nand ( n45044 , n45023 , n45043 );
not ( n45045 , n45044 );
not ( n45046 , n44270 );
xor ( n45047 , n44251 , n44256 );
and ( n45048 , n45047 , n44263 );
and ( n45049 , n44251 , n44256 );
or ( n45050 , n45048 , n45049 );
buf ( n45051 , n45050 );
buf ( n45052 , n45051 );
not ( n45053 , n45052 );
buf ( n45054 , n454 );
nor ( n45055 , n45053 , n45054 );
buf ( n45056 , n45055 );
buf ( n45057 , n6541 );
buf ( n45058 , n35343 );
nor ( n45059 , n45057 , n45058 );
buf ( n45060 , n45059 );
buf ( n45061 , n45060 );
buf ( n45062 , n44255 );
not ( n45063 , n45062 );
buf ( n45064 , n45063 );
buf ( n45065 , n45064 );
xor ( n45066 , n45061 , n45065 );
buf ( n45067 , n6337 );
not ( n45068 , n45067 );
buf ( n45069 , n38773 );
not ( n45070 , n45069 );
or ( n45071 , n45068 , n45070 );
buf ( n45072 , n537 );
nand ( n45073 , n45071 , n45072 );
buf ( n45074 , n45073 );
buf ( n45075 , n45074 );
xor ( n45076 , n45066 , n45075 );
buf ( n45077 , n45076 );
buf ( n45078 , n45077 );
buf ( n45079 , n3138 );
and ( n45080 , n45078 , n45079 );
buf ( n45081 , n45080 );
nor ( n45082 , n45056 , n45081 );
nor ( n45083 , n45046 , n45082 );
not ( n45084 , n45083 );
nor ( n45085 , n45084 , n44232 );
and ( n45086 , n44176 , n45085 );
not ( n45087 , n45086 );
or ( n45088 , n45045 , n45087 );
nor ( n45089 , n44120 , n44232 );
not ( n45090 , n45089 );
not ( n45091 , n454 );
not ( n45092 , n43924 );
or ( n45093 , n45091 , n45092 );
nand ( n45094 , n45093 , n44174 );
not ( n45095 , n45094 );
or ( n45096 , n45090 , n45095 );
or ( n45097 , n44183 , n44231 );
nand ( n45098 , n45096 , n45097 );
and ( n45099 , n45098 , n45083 );
nand ( n45100 , n44242 , n44269 );
or ( n45101 , n45100 , n45082 );
nand ( n45102 , n45056 , n45081 );
nand ( n45103 , n45101 , n45102 );
nor ( n45104 , n45099 , n45103 );
nand ( n45105 , n45088 , n45104 );
not ( n45106 , n45105 );
nor ( n45107 , n44515 , n44498 );
nand ( n45108 , n45107 , n44569 );
not ( n45109 , n45108 );
not ( n45110 , n45021 );
or ( n45111 , n45109 , n45110 );
buf ( n45112 , n45034 );
nand ( n45113 , n45111 , n45112 );
not ( n45114 , n45113 );
and ( n45115 , n45098 , n44270 );
not ( n45116 , n45100 );
nor ( n45117 , n45115 , n45116 );
not ( n45118 , n40804 );
not ( n45119 , n40314 );
or ( n45120 , n45118 , n45119 );
nand ( n45121 , n45120 , n40811 );
not ( n45122 , n45121 );
nand ( n45123 , n45108 , n45112 );
nand ( n45124 , n44960 , n454 );
nor ( n45125 , n44977 , n44967 );
nand ( n45126 , n45124 , n45125 );
nand ( n45127 , n44933 , n45126 );
not ( n45128 , n45127 );
buf ( n45129 , n45128 );
buf ( n45130 , n44870 );
not ( n45131 , n45130 );
xor ( n45132 , n32659 , n32667 );
buf ( n45133 , n45001 );
not ( n45134 , n44660 );
not ( n45135 , n44642 );
and ( n45136 , n45134 , n45135 );
not ( n45137 , n44794 );
or ( n45138 , n45137 , n44815 );
nor ( n45139 , n45136 , n45138 );
not ( n45140 , n45139 );
nor ( n45141 , n44903 , n44911 );
buf ( n45142 , n45141 );
not ( n45143 , n45142 );
xor ( n45144 , n45061 , n45065 );
and ( n45145 , n45144 , n45075 );
and ( n45146 , n45061 , n45065 );
or ( n45147 , n45145 , n45146 );
buf ( n45148 , n45147 );
not ( n45149 , n42620 );
not ( n45150 , n42867 );
or ( n45151 , n45149 , n45150 );
not ( n45152 , n42879 );
nand ( n45153 , n45151 , n45152 );
and ( n45154 , n45153 , n42663 );
or ( n45155 , n45154 , n42881 );
not ( n45156 , n42881 );
nand ( n45157 , n45156 , n42663 );
not ( n45158 , n45157 );
not ( n45159 , n45153 );
or ( n45160 , n45158 , n45159 );
or ( n45161 , n45153 , n45157 );
nand ( n45162 , n45160 , n45161 );
not ( n45163 , n42850 );
not ( n45164 , n42832 );
or ( n45165 , n45163 , n45164 );
not ( n45166 , n42857 );
nand ( n45167 , n45165 , n45166 );
and ( n45168 , n45167 , n42839 );
not ( n45169 , n42860 );
nor ( n45170 , n45168 , n45169 );
not ( n45171 , n42049 );
nand ( n45172 , n45171 , n42051 );
not ( n45173 , n45172 );
not ( n45174 , n42041 );
or ( n45175 , n45173 , n45174 );
or ( n45176 , n42041 , n45172 );
nand ( n45177 , n45175 , n45176 );
nand ( n45178 , n42839 , n42860 );
not ( n45179 , n42831 );
nand ( n45180 , n45179 , n42856 );
and ( n45181 , n42569 , n42874 );
nand ( n45182 , n42512 , n42872 );
and ( n45183 , n42794 , n42864 );
not ( n45184 , n42872 );
nand ( n45185 , n42619 , n42878 );
not ( n45186 , n42036 );
nand ( n45187 , n45186 , n42033 );
not ( n45188 , n45187 );
not ( n45189 , n42003 );
or ( n45190 , n45189 , n42019 );
not ( n45191 , n42032 );
nand ( n45192 , n45190 , n45191 );
not ( n45193 , n45192 );
or ( n45194 , n45188 , n45193 );
or ( n45195 , n45192 , n45187 );
nand ( n45196 , n45194 , n45195 );
nor ( n45197 , n42019 , n42032 );
not ( n45198 , n45197 );
not ( n45199 , n45189 );
or ( n45200 , n45198 , n45199 );
or ( n45201 , n45189 , n45197 );
nand ( n45202 , n45200 , n45201 );
not ( n45203 , n42883 );
nand ( n45204 , n45203 , n42700 );
not ( n45205 , n42725 );
nand ( n45206 , n45205 , n42889 );
or ( n45207 , n42739 , n42893 );
or ( n45208 , n41917 , n41911 );
not ( n45209 , n45208 );
nand ( n45210 , n41904 , n41914 );
not ( n45211 , n45210 );
or ( n45212 , n45209 , n45211 );
or ( n45213 , n45210 , n45208 );
nand ( n45214 , n45212 , n45213 );
not ( n45215 , n3990 );
not ( n45216 , n3992 );
nor ( n45217 , n45216 , n3982 );
not ( n45218 , n45217 );
or ( n45219 , n45215 , n45218 );
or ( n45220 , n45217 , n3990 );
nand ( n45221 , n45219 , n45220 );
and ( n45222 , n42867 , n42512 );
nor ( n45223 , n45222 , n45184 );
xor ( n45224 , n45181 , n45223 );
xor ( n45225 , n45178 , n45167 );
not ( n45226 , n42704 );
not ( n45227 , n42724 );
and ( n45228 , n45226 , n45227 );
nor ( n45229 , n45228 , n42739 );
not ( n45230 , n45040 );
nor ( n45231 , n45230 , n44604 );
not ( n45232 , n45231 );
nand ( n45233 , n45232 , n45028 );
not ( n45234 , n45233 );
and ( n45235 , n45108 , n45130 );
buf ( n45236 , n44879 );
buf ( n45237 , n44933 );
buf ( n45238 , n45126 );
not ( n45239 , n40268 );
nand ( n45240 , n45236 , n45237 , n45238 , n45239 );
not ( n45241 , n45240 );
not ( n45242 , n45241 );
not ( n45243 , n40951 );
not ( n45244 , n40282 );
or ( n45245 , n45243 , n45244 );
and ( n45246 , n40301 , n40309 );
nand ( n45247 , n45245 , n45246 );
not ( n45248 , n45247 );
or ( n45249 , n45242 , n45248 );
not ( n45250 , n45121 );
not ( n45251 , n45128 );
or ( n45252 , n45250 , n45251 );
not ( n45253 , n44976 );
not ( n45254 , n45124 );
or ( n45255 , n45253 , n45254 );
buf ( n45256 , n44967 );
nand ( n45257 , n45255 , n45256 );
not ( n45258 , n44978 );
not ( n45259 , n45124 );
or ( n45260 , n45258 , n45259 );
nand ( n45261 , n45260 , n45141 );
nand ( n45262 , n45257 , n45261 );
not ( n45263 , n45262 );
nand ( n45264 , n45252 , n45263 );
not ( n45265 , n45264 );
nand ( n45266 , n45249 , n45265 );
nand ( n45267 , n45235 , n45266 );
not ( n45268 , n40936 );
nand ( n45269 , n45235 , n44982 , n45268 );
nand ( n45270 , n45267 , n45269 , n45114 );
not ( n45271 , n45270 );
or ( n45272 , n45234 , n45271 );
not ( n45273 , n45233 );
and ( n45274 , n45273 , n45114 );
nand ( n45275 , n45274 , n45267 , n45269 );
nand ( n45276 , n45272 , n45275 );
buf ( n45277 , n45276 );
not ( n45278 , n45277 );
not ( n45279 , n44176 );
not ( n45280 , n45279 );
not ( n45281 , n45280 );
not ( n45282 , n44999 );
nand ( n45283 , n45040 , n45041 );
nand ( n45284 , n45035 , n45028 );
nand ( n45285 , n45282 , n45283 , n45284 );
not ( n45286 , n45285 );
or ( n45287 , n45281 , n45286 );
not ( n45288 , n44120 );
nand ( n45289 , n45288 , n45094 );
nand ( n45290 , n45287 , n45289 );
not ( n45291 , n45290 );
and ( n45292 , n39747 , n40998 , n40303 );
nand ( n45293 , n37441 , n45130 , n44980 , n45292 );
not ( n45294 , n45289 );
not ( n45295 , n45028 );
not ( n45296 , n45035 );
or ( n45297 , n45295 , n45296 );
nand ( n45298 , n45297 , n45283 );
not ( n45299 , n45011 );
not ( n45300 , n45002 );
or ( n45301 , n45299 , n45300 );
nand ( n45302 , n45301 , n45020 );
nor ( n45303 , n45294 , n45298 , n45302 );
nand ( n45304 , n45293 , n45303 );
not ( n45305 , n45304 );
or ( n45306 , n45291 , n45305 );
not ( n45307 , n44872 );
nor ( n45308 , n45307 , n45279 );
nand ( n45309 , n45308 , n45266 );
nand ( n45310 , n45306 , n45309 );
not ( n45311 , n40815 );
not ( n45312 , n45311 );
not ( n45313 , n40317 );
or ( n45314 , n45312 , n45313 );
nor ( n45315 , n40315 , n40812 );
nand ( n45316 , n40260 , n45315 , n40313 );
nand ( n45317 , n45314 , n45316 );
nand ( n45318 , n45237 , n45143 );
not ( n45319 , n45318 );
not ( n45320 , n39748 );
nand ( n45321 , n45320 , n45236 );
not ( n45322 , n45321 );
not ( n45323 , n38657 );
nand ( n45324 , n45322 , n37441 , n45323 );
nand ( n45325 , n40312 , n45236 );
nand ( n45326 , n45324 , n45325 , n45122 );
not ( n45327 , n45326 );
or ( n45328 , n45319 , n45327 );
not ( n45329 , n45122 );
nor ( n45330 , n45329 , n45318 );
nand ( n45331 , n45330 , n45324 , n45325 );
nand ( n45332 , n45328 , n45331 );
nand ( n45333 , n45317 , n45332 );
not ( n45334 , n44176 );
nor ( n45335 , n45334 , n44232 );
nand ( n45336 , n44872 , n45335 );
not ( n45337 , n45336 );
nand ( n45338 , n45337 , n44982 , n44983 );
nor ( n45339 , n40907 , n40932 );
and ( n45340 , n45236 , n45237 );
not ( n45341 , n45133 );
buf ( n45342 , n44979 );
buf ( n45343 , n45257 );
nand ( n45344 , n45342 , n45343 );
not ( n45345 , n45344 );
not ( n45346 , n45123 );
nor ( n45347 , n45121 , n45262 );
not ( n45348 , n45347 );
not ( n45349 , n45325 );
or ( n45350 , n45348 , n45349 );
not ( n45351 , n45262 );
not ( n45352 , n45129 );
and ( n45353 , n45351 , n45352 );
nor ( n45354 , n45353 , n45131 );
nand ( n45355 , n45350 , n45354 );
and ( n45356 , n37441 , n45130 );
nand ( n45357 , n45356 , n44982 );
not ( n45358 , n45002 );
not ( n45359 , n45011 );
or ( n45360 , n45358 , n45359 );
nand ( n45361 , n45360 , n45020 );
not ( n45362 , n45361 );
nand ( n45363 , n45355 , n45357 , n45362 );
not ( n45364 , n45363 );
or ( n45365 , n45346 , n45364 );
not ( n45366 , n45362 );
nor ( n45367 , n45366 , n45123 );
nand ( n45368 , n45367 , n45355 , n45357 );
nand ( n45369 , n45365 , n45368 );
buf ( n45370 , n45369 );
not ( n45371 , n45370 );
nor ( n45372 , n45371 , n29519 );
buf ( n45373 , n41031 );
and ( n45374 , n45011 , n45020 );
not ( n45375 , n45374 );
not ( n45376 , n45375 );
not ( n45377 , n40971 );
not ( n45378 , n40966 );
or ( n45379 , n45377 , n45378 );
not ( n45380 , n44980 );
nor ( n45381 , n45380 , n45139 );
nand ( n45382 , n45379 , n45381 );
not ( n45383 , n45128 );
not ( n45384 , n45121 );
or ( n45385 , n45383 , n45384 );
nand ( n45386 , n45385 , n45263 );
and ( n45387 , n45386 , n45140 );
nor ( n45388 , n45387 , n45341 );
nand ( n45389 , n45382 , n45388 );
not ( n45390 , n45389 );
or ( n45391 , n45376 , n45390 );
nand ( n45392 , n45382 , n45388 , n45374 );
nand ( n45393 , n45391 , n45392 );
buf ( n45394 , n45393 );
and ( n45395 , n45241 , n45247 );
nor ( n45396 , n45395 , n45264 );
not ( n45397 , n45396 );
nand ( n45398 , n44982 , n45268 );
not ( n45399 , n45398 );
or ( n45400 , n45397 , n45399 );
nand ( n45401 , n45140 , n45133 );
nand ( n45402 , n45400 , n45401 );
not ( n45403 , n45402 );
not ( n45404 , n45401 );
nand ( n45405 , n45398 , n45396 , n45404 );
not ( n45406 , n45405 );
or ( n45407 , n45403 , n45406 );
not ( n45408 , n45345 );
not ( n45409 , n45408 );
nand ( n45410 , n45340 , n45292 , n37441 );
nand ( n45411 , n40970 , n45236 , n45237 );
nand ( n45412 , n45237 , n45121 );
and ( n45413 , n45412 , n45143 );
nand ( n45414 , n45410 , n45411 , n45413 );
not ( n45415 , n45414 );
or ( n45416 , n45409 , n45415 );
not ( n45417 , n45344 );
nand ( n45418 , n45417 , n45410 , n45411 , n45413 );
nand ( n45419 , n45416 , n45418 );
nand ( n45420 , n45407 , n45419 );
nor ( n45421 , n45420 , n45333 );
nand ( n45422 , n45373 , n45394 , n45421 );
nand ( n45423 , n45372 , n45422 );
xor ( n45424 , n42868 , n45182 );
not ( n45425 , n45424 );
nand ( n45426 , n45425 , n29519 );
not ( n45427 , n29519 );
nand ( n45428 , n45427 , n45278 );
nor ( n45429 , n45278 , n29519 );
not ( n45430 , n45224 );
nand ( n45431 , n45430 , n29519 );
not ( n45432 , n45290 );
not ( n45433 , n45304 );
or ( n45434 , n45432 , n45433 );
nand ( n45435 , n45434 , n45309 );
not ( n45436 , n44232 );
nand ( n45437 , n45436 , n45097 );
not ( n45438 , n45437 );
and ( n45439 , n45435 , n45438 );
not ( n45440 , n45435 );
and ( n45441 , n45440 , n45437 );
nor ( n45442 , n45439 , n45441 );
and ( n45443 , n44270 , n45100 );
not ( n45444 , n45443 );
not ( n45445 , n45444 );
not ( n45446 , n45241 );
not ( n45447 , n45247 );
or ( n45448 , n45446 , n45447 );
nand ( n45449 , n45448 , n45265 );
not ( n45450 , n45336 );
nand ( n45451 , n45449 , n45450 );
not ( n45452 , n45335 );
not ( n45453 , n45044 );
or ( n45454 , n45452 , n45453 );
not ( n45455 , n45098 );
nand ( n45456 , n45454 , n45455 );
not ( n45457 , n45456 );
nand ( n45458 , n45451 , n45338 , n45457 );
not ( n45459 , n45458 );
or ( n45460 , n45445 , n45459 );
nand ( n45461 , n45451 , n45338 , n45457 , n45443 );
nand ( n45462 , n45460 , n45461 );
nand ( n45463 , n45442 , n45462 );
nor ( n45464 , n45463 , n41032 );
not ( n45465 , n45408 );
not ( n45466 , n45414 );
or ( n45467 , n45465 , n45466 );
nand ( n45468 , n45467 , n45418 );
nand ( n45469 , n45393 , n45468 );
not ( n45470 , n45469 );
nand ( n45471 , n45317 , n45332 );
not ( n45472 , n45471 );
nand ( n45473 , n45405 , n45402 );
nand ( n45474 , n45470 , n45472 , n45369 , n45473 );
nor ( n45475 , n45298 , n45361 );
not ( n45476 , n45475 );
not ( n45477 , n45293 );
or ( n45478 , n45476 , n45477 );
buf ( n45479 , n45285 );
nand ( n45480 , n45478 , n45479 );
not ( n45481 , n45307 );
nand ( n45482 , n45481 , n45449 );
and ( n45483 , n45280 , n45289 );
nand ( n45484 , n45480 , n45482 , n45483 );
not ( n45485 , n45484 );
not ( n45486 , n45482 );
not ( n45487 , n45480 );
or ( n45488 , n45486 , n45487 );
not ( n45489 , n45483 );
nand ( n45490 , n45488 , n45489 );
not ( n45491 , n45490 );
or ( n45492 , n45485 , n45491 );
nand ( n45493 , n45492 , n45276 );
nor ( n45494 , n45474 , n45493 );
nand ( n45495 , n45464 , n45494 );
not ( n45496 , n45495 );
not ( n45497 , n45082 );
nand ( n45498 , n45497 , n45102 );
not ( n45499 , n45498 );
not ( n45500 , n44272 );
not ( n45501 , n45044 );
or ( n45502 , n45500 , n45501 );
nand ( n45503 , n45502 , n45117 );
not ( n45504 , n45503 );
nand ( n45505 , n44873 , n45449 );
nand ( n45506 , n45504 , n45505 , n44984 );
not ( n45507 , n45506 );
not ( n45508 , n45507 );
or ( n45509 , n45499 , n45508 );
not ( n45510 , n45498 );
nand ( n45511 , n45506 , n45510 );
nand ( n45512 , n45509 , n45511 );
and ( n45513 , n45512 , n29518 );
nand ( n45514 , n45496 , n45513 );
and ( n45515 , n42663 , n42700 );
not ( n45516 , n45515 );
not ( n45517 , n45153 );
or ( n45518 , n45516 , n45517 );
nand ( n45519 , n45518 , n42884 );
xor ( n45520 , n45519 , n45206 );
not ( n45521 , n45520 );
nand ( n45522 , n45521 , n29519 );
not ( n45523 , n45511 );
nor ( n45524 , n45506 , n45510 );
nor ( n45525 , n45523 , n45524 );
and ( n45526 , n45525 , n29518 );
nand ( n45527 , n45495 , n45526 );
nand ( n45528 , n45514 , n45522 , n45527 );
buf ( n45529 , n29519 );
xnor ( n45530 , n45204 , n45155 );
not ( n45531 , n45207 );
buf ( n45532 , n45317 );
nand ( n45533 , n41031 , n45532 );
or ( n45534 , n45332 , n29519 );
or ( n45535 , n45533 , n45534 );
not ( n45536 , n45332 );
nor ( n45537 , n45536 , n29519 );
nand ( n45538 , n45533 , n45537 );
not ( n45539 , n42854 );
nor ( n45540 , n45539 , n42816 );
not ( n45541 , n45540 );
not ( n45542 , n45163 );
or ( n45543 , n45541 , n45542 );
or ( n45544 , n45163 , n45540 );
nand ( n45545 , n45543 , n45544 );
nand ( n45546 , n45545 , n29519 );
nand ( n45547 , n45535 , n45538 , n45546 );
not ( n45548 , n45442 );
and ( n45549 , n45310 , n45438 );
not ( n45550 , n45310 );
and ( n45551 , n45550 , n45437 );
nor ( n45552 , n45549 , n45551 );
not ( n45553 , n45233 );
not ( n45554 , n45270 );
or ( n45555 , n45553 , n45554 );
nand ( n45556 , n45555 , n45275 );
nand ( n45557 , n41031 , n45556 );
not ( n45558 , n45557 );
not ( n45559 , n45345 );
not ( n45560 , n45414 );
not ( n45561 , n45560 );
or ( n45562 , n45559 , n45561 );
nand ( n45563 , n45408 , n45414 );
nand ( n45564 , n45562 , n45563 );
nor ( n45565 , n45564 , n29519 );
nand ( n45566 , n45565 , n45373 , n45472 );
or ( n45567 , n45163 , n42816 );
nand ( n45568 , n45567 , n42854 );
xor ( n45569 , n45180 , n45568 );
not ( n45570 , n45569 );
nand ( n45571 , n45570 , n29519 );
not ( n45572 , n45472 );
not ( n45573 , n29519 );
nand ( n45574 , n45573 , n45564 );
not ( n45575 , n45574 );
and ( n45576 , n45572 , n45575 );
nor ( n45577 , n45574 , n41031 );
nor ( n45578 , n45576 , n45577 );
nand ( n45579 , n45566 , n45571 , n45578 );
not ( n45580 , n45564 );
not ( n45581 , n41031 );
nor ( n45582 , n45581 , n45548 );
nand ( n45583 , n45339 , n42163 );
not ( n45584 , n45420 );
not ( n45585 , n45333 );
nand ( n45586 , n45373 , n45584 , n45585 );
not ( n45587 , n45394 );
nor ( n45588 , n45587 , n29519 );
nand ( n45589 , n45586 , n45588 );
and ( n45590 , n45585 , n29518 );
nand ( n45591 , n45590 , n45584 , n45587 , n45373 );
not ( n45592 , n45183 );
not ( n45593 , n45170 );
or ( n45594 , n45592 , n45593 );
or ( n45595 , n45170 , n45183 );
nand ( n45596 , n45594 , n45595 );
nand ( n45597 , n45596 , n29519 );
nand ( n45598 , n45589 , n45591 , n45597 );
not ( n45599 , n45229 );
not ( n45600 , n45519 );
or ( n45601 , n45599 , n45600 );
nand ( n45602 , n45601 , n42894 );
nand ( n45603 , n42747 , n42896 );
not ( n45604 , n45603 );
and ( n45605 , n45602 , n45604 );
not ( n45606 , n45602 );
and ( n45607 , n45606 , n45603 );
nor ( n45608 , n45605 , n45607 );
and ( n45609 , n45148 , n3360 );
xor ( n45610 , n45609 , n3138 );
not ( n45611 , n29519 );
nand ( n45612 , n45611 , n45610 );
and ( n45613 , n45558 , n45421 );
not ( n45614 , n42874 );
nor ( n45615 , n45185 , n45614 );
not ( n45616 , n45185 );
buf ( n45617 , n42568 );
and ( n45618 , n45616 , n42874 , n45617 );
and ( n45619 , n45185 , n45614 );
nor ( n45620 , n45618 , n45619 );
not ( n45621 , n45473 );
nor ( n45622 , n45621 , n29519 );
not ( n45623 , n45580 );
nand ( n45624 , n45373 , n45623 , n45585 );
nand ( n45625 , n45622 , n45624 );
nor ( n45626 , n45580 , n29519 );
nand ( n45627 , n45621 , n45626 , n45585 , n45373 );
not ( n45628 , n45225 );
nand ( n45629 , n45628 , n29519 );
nand ( n45630 , n45625 , n45627 , n45629 );
buf ( n45631 , n40997 );
and ( n45632 , n45631 , n42065 );
buf ( n45633 , n45462 );
nor ( n45634 , n45633 , n45529 );
nand ( n45635 , n45363 , n45123 );
buf ( n45636 , n40979 );
not ( n45637 , n45368 );
not ( n45638 , n45635 );
or ( n45639 , n45637 , n45638 );
nand ( n45640 , n45639 , n45394 );
not ( n45641 , n45640 );
nand ( n45642 , n45373 , n45641 , n45421 );
nand ( n45643 , n45086 , n45481 , n45449 );
nand ( n45644 , n45086 , n45481 , n44983 , n44982 );
nand ( n45645 , n45610 , n45644 , n45106 , n45643 );
nand ( n45646 , C1 , n45645 );
nand ( n45647 , n45490 , n45484 );
buf ( n45648 , n45647 );
nor ( n45649 , n45648 , n29519 );
nand ( n45650 , n45207 , n42889 );
not ( n45651 , n42889 );
and ( n45652 , n45531 , n45651 );
or ( n45653 , n45205 , n45650 );
nand ( n45654 , n45653 , n29519 );
nor ( n45655 , n45652 , n45654 );
nand ( n45656 , n45584 , n45462 );
nand ( n45657 , n45552 , n45647 , n45556 , n45472 );
nor ( n45658 , n45656 , n45657 );
nor ( n45659 , n45512 , n45640 );
not ( n45660 , n45581 );
nand ( n45661 , n45658 , n45659 , n45660 );
not ( n45662 , n45612 );
nand ( n45663 , n45662 , n45106 , n45644 , n45643 );
nand ( n45664 , C1 , n45663 );
not ( n45665 , n45634 );
nand ( n45666 , n45530 , n45529 );
or ( n45667 , n45642 , n45428 );
nand ( n45668 , n45642 , n45429 );
nand ( n45669 , n45667 , n45668 , n45431 );
nand ( n45670 , n45162 , n29519 );
not ( n45671 , n3706 );
nand ( n45672 , n3709 , n3669 );
not ( n45673 , n45672 );
or ( n45674 , n45671 , n45673 );
and ( n45675 , n3651 , n3667 );
not ( n45676 , n3651 );
and ( n45677 , n45676 , n3668 );
nor ( n45678 , n45675 , n45677 );
or ( n45679 , n45678 , n3706 );
nand ( n45680 , n45674 , n45679 );
buf ( n45681 , n40935 );
nand ( n45682 , n45681 , n40945 );
and ( n45683 , n45682 , n42091 );
not ( n45684 , n45682 );
and ( n45685 , n45684 , n42092 );
nor ( n45686 , n45683 , n45685 );
not ( n45687 , n42086 );
nor ( n45688 , n45687 , n42091 );
nand ( n45689 , n45688 , n42090 , n45632 );
not ( n45690 , n45636 );
not ( n45691 , n29520 );
not ( n45692 , n45686 );
or ( n45693 , n45691 , n45692 );
nand ( n45694 , n45196 , n29519 );
nand ( n45695 , n45693 , n45694 );
not ( n45696 , n29520 );
not ( n45697 , n42939 );
or ( n45698 , n45696 , n45697 );
nand ( n45699 , n45221 , n29519 );
nand ( n45700 , n45698 , n45699 );
not ( n45701 , n45689 );
and ( n45702 , n45690 , n29520 );
nand ( n45703 , n45701 , n45702 );
not ( n45704 , n29520 );
nor ( n45705 , n45704 , n45690 );
nand ( n45706 , n45689 , n45705 );
nand ( n45707 , n45177 , n29519 );
nand ( n45708 , n45703 , n45706 , n45707 );
not ( n45709 , n45641 );
not ( n45710 , n45613 );
or ( n45711 , n45709 , n45710 );
not ( n45712 , n45648 );
nor ( n45713 , n45712 , n29519 );
nand ( n45714 , n45711 , n45713 );
nand ( n45715 , n45613 , n45649 , n45641 );
or ( n45716 , n45223 , n45616 , n45617 );
not ( n45717 , n45620 );
and ( n45718 , n45223 , n45615 );
nor ( n45719 , n45717 , n45718 );
nand ( n45720 , n45716 , n45719 );
nand ( n45721 , n45720 , n29519 );
nand ( n45722 , n45714 , n45715 , n45721 );
nand ( n45723 , n45661 , n45664 );
or ( n45724 , n45519 , n45650 );
nand ( n45725 , n45531 , n45205 , n45519 );
nand ( n45726 , n45724 , n45725 , n45655 );
nand ( n45727 , n29520 , n40945 );
or ( n45728 , n45727 , n45681 );
not ( n45729 , n40945 );
nand ( n45730 , n45729 , n45681 , n29520 );
nand ( n45731 , n45202 , n29519 );
nand ( n45732 , n45728 , n45730 , n45731 );
or ( n45733 , n45583 , n29519 , n40917 );
nand ( n45734 , n29520 , n40917 , n45583 );
nand ( n45735 , n45214 , n29519 );
nand ( n45736 , n45733 , n45734 , n45735 );
not ( n45737 , n41032 );
not ( n45738 , n45463 );
nand ( n45739 , n3865 , n3497 );
and ( n45740 , n45739 , n3808 );
not ( n45741 , n45739 );
and ( n45742 , n45741 , n32823 );
nor ( n45743 , n45740 , n45742 );
or ( n45744 , n45552 , n29519 );
nand ( n45745 , n45744 , n45670 );
not ( n45746 , n45370 );
and ( n45747 , n45394 , n29518 );
nand ( n45748 , n45746 , n45747 , n45373 , n45421 );
nand ( n45749 , n45748 , n45423 , n45426 );
nor ( n45750 , n45548 , n29519 );
not ( n45751 , n45745 );
nand ( n45752 , C1 , n45723 , n45726 );
nand ( n45753 , n29520 , n45737 , n45494 );
nand ( n45754 , n45738 , n45646 , n45525 );
or ( n45755 , n45753 , n45754 );
nand ( n45756 , n45608 , n29519 );
nand ( n45757 , n45755 , n45756 );
not ( n45758 , n45474 );
not ( n45759 , n45493 );
nand ( n45760 , n45758 , n45759 , n45660 );
not ( n45761 , n45670 );
nor ( n45762 , n45761 , n45750 );
and ( n45763 , n45760 , n45762 );
not ( n45764 , n45760 );
and ( n45765 , n45764 , n45751 );
nor ( n45766 , n45763 , n45765 );
not ( n45767 , n45633 );
nor ( n45768 , n45767 , n45529 );
nand ( n45769 , n45582 , n45494 );
or ( n45770 , n45665 , n45769 );
nand ( n45771 , n45769 , n45768 );
nand ( n45772 , n45770 , n45771 , n45666 );
not ( C0n , n0 );
and ( C0 , C0n , n0 );
not ( C1n , n0 );
or ( C1 , C1n , n0 );
endmodule
