module top ( g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 , g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 , g157 , g158 , g159 , g160 , g161 , g162 , g163 , g164 , g165 , g166 );
input g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 , g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 ;
output g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 , g157 , g158 , g159 , g160 , g161 , g162 , g163 , g164 , g165 , g166 ;

wire n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , 
     n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , 
     n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , 
     n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , 
     n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , 
     n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , 
     n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , 
     n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , 
     n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , 
     n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , 
     n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , 
     n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , 
     n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , 
     n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , 
     n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , 
     n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , 
     n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , 
     n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , 
     n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , 
     n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , 
     n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , 
     n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , 
     n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , 
     n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , 
     n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , 
     n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , 
     n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , 
     n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , 
     n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , 
     n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , 
     n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , 
     n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , 
     n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , 
     n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , 
     n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , 
     n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , 
     n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , 
     n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , 
     n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , 
     n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , 
     n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , 
     n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , 
     n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , 
     n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , 
     n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , 
     n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , 
     n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , 
     n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , 
     n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , 
     n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , 
     n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , 
     n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , 
     n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , 
     n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , 
     n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , 
     n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , 
     n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , 
     n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , 
     n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , 
     n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , 
     n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , 
     n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , 
     n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , 
     n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , 
     n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , 
     n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , 
     n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , 
     n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , 
     n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , 
     n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , 
     n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , 
     n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , 
     n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , 
     n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , 
     n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , 
     n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , 
     n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , 
     n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , 
     n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , 
     n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , 
     n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , 
     n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , 
     n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , 
     n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , 
     n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , 
     n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , 
     n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , 
     n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , 
     n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , 
     n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , 
     n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , 
     n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , 
     n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , 
     n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , 
     n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , 
     n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , 
     n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , 
     n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , 
     n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , 
     n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , 
     n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , 
     n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , 
     n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , 
     n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , 
     n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , 
     n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , 
     n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , 
     n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , 
     n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , 
     n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , 
     n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , 
     n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , 
     n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , 
     n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , 
     n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , 
     n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , 
     n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , 
     n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , 
     n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , 
     n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , 
     n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , 
     n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , 
     n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , 
     n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , 
     n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , 
     n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , 
     n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , 
     n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , 
     n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , 
     n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , 
     n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , 
     n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , 
     n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , 
     n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , 
     n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , 
     n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , 
     n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , 
     n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , 
     n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , 
     n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , 
     n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , 
     n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , 
     n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , 
     n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , 
     n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , 
     n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , 
     n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , 
     n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , 
     n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , 
     n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , 
     n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , 
     n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , 
     n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , 
     n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , 
     n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , 
     n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , 
     n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , 
     n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , 
     n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , 
     n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , 
     n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , 
     n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , 
     n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , 
     n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , 
     n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , 
     n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , 
     n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , 
     n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , 
     n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , 
     n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , 
     n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , 
     n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , 
     n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , 
     n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , 
     n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , 
     n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , 
     n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , 
     n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , 
     n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , 
     n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , 
     n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , 
     n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , 
     n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , 
     n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , 
     n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , 
     n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , 
     n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , 
     n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , 
     n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , 
     n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , 
     n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , 
     n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , 
     n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , 
     n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , 
     n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , 
     n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , 
     n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , 
     n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , 
     n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , 
     n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , 
     n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , 
     n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , 
     n2020 , n2021 , n2022 , n2023 ;
buf ( n1 , g0 );
buf ( n2 , g1 );
buf ( n3 , g2 );
buf ( n4 , g3 );
buf ( n5 , g4 );
buf ( n6 , g5 );
buf ( n7 , g6 );
buf ( n8 , g7 );
buf ( n9 , g8 );
buf ( n10 , g9 );
buf ( n11 , g10 );
buf ( n12 , g11 );
buf ( n13 , g12 );
buf ( n14 , g13 );
buf ( n15 , g14 );
buf ( n16 , g15 );
buf ( n17 , g16 );
buf ( n18 , g17 );
buf ( n19 , g18 );
buf ( n20 , g19 );
buf ( n21 , g20 );
buf ( n22 , g21 );
buf ( n23 , g22 );
buf ( n24 , g23 );
buf ( n25 , g24 );
buf ( n26 , g25 );
buf ( n27 , g26 );
buf ( n28 , g27 );
buf ( n29 , g28 );
buf ( n30 , g29 );
buf ( n31 , g30 );
buf ( n32 , g31 );
buf ( n33 , g32 );
buf ( n34 , g33 );
buf ( n35 , g34 );
buf ( n36 , g35 );
buf ( n37 , g36 );
buf ( n38 , g37 );
buf ( n39 , g38 );
buf ( n40 , g39 );
buf ( n41 , g40 );
buf ( n42 , g41 );
buf ( n43 , g42 );
buf ( n44 , g43 );
buf ( n45 , g44 );
buf ( n46 , g45 );
buf ( n47 , g46 );
buf ( n48 , g47 );
buf ( n49 , g48 );
buf ( n50 , g49 );
buf ( n51 , g50 );
buf ( n52 , g51 );
buf ( n53 , g52 );
buf ( n54 , g53 );
buf ( n55 , g54 );
buf ( n56 , g55 );
buf ( n57 , g56 );
buf ( n58 , g57 );
buf ( n59 , g58 );
buf ( n60 , g59 );
buf ( n61 , g60 );
buf ( n62 , g61 );
buf ( n63 , g62 );
buf ( n64 , g63 );
buf ( n65 , g64 );
buf ( n66 , g65 );
buf ( n67 , g66 );
buf ( n68 , g67 );
buf ( n69 , g68 );
buf ( n70 , g69 );
buf ( n71 , g70 );
buf ( n72 , g71 );
buf ( n73 , g72 );
buf ( n74 , g73 );
buf ( n75 , g74 );
buf ( n76 , g75 );
buf ( n77 , g76 );
buf ( n78 , g77 );
buf ( n79 , g78 );
buf ( n80 , g79 );
buf ( n81 , g80 );
buf ( n82 , g81 );
buf ( n83 , g82 );
buf ( n84 , g83 );
buf ( n85 , g84 );
buf ( n86 , g85 );
buf ( n87 , g86 );
buf ( n88 , g87 );
buf ( n89 , g88 );
buf ( n90 , g89 );
buf ( n91 , g90 );
buf ( n92 , g91 );
buf ( n93 , g92 );
buf ( n94 , g93 );
buf ( n95 , g94 );
buf ( n96 , g95 );
buf ( n97 , g96 );
buf ( n98 , g97 );
buf ( n99 , g98 );
buf ( n100 , g99 );
buf ( n101 , g100 );
buf ( n102 , g101 );
buf ( n103 , g102 );
buf ( n104 , g103 );
buf ( n105 , g104 );
buf ( n106 , g105 );
buf ( n107 , g106 );
buf ( n108 , g107 );
buf ( n109 , g108 );
buf ( n110 , g109 );
buf ( n111 , g110 );
buf ( n112 , g111 );
buf ( n113 , g112 );
buf ( n114 , g113 );
buf ( n115 , g114 );
buf ( n116 , g115 );
buf ( n117 , g116 );
buf ( n118 , g117 );
buf ( n119 , g118 );
buf ( n120 , g119 );
buf ( n121 , g120 );
buf ( n122 , g121 );
buf ( n123 , g122 );
buf ( n124 , g123 );
buf ( n125 , g124 );
buf ( n126 , g125 );
buf ( n127 , g126 );
buf ( n128 , g127 );
buf ( n129 , g128 );
buf ( n130 , g129 );
buf ( n131 , g130 );
buf ( n132 , g131 );
buf ( n133 , g132 );
buf ( n134 , g133 );
buf ( n135 , g134 );
buf ( n136 , g135 );
buf ( g136 , n137 );
buf ( g137 , n138 );
buf ( g138 , n139 );
buf ( g139 , n140 );
buf ( g140 , n141 );
buf ( g141 , n142 );
buf ( g142 , n143 );
buf ( g143 , n144 );
buf ( g144 , n145 );
buf ( g145 , n146 );
buf ( g146 , n147 );
buf ( g147 , n148 );
buf ( g148 , n149 );
buf ( g149 , n150 );
buf ( g150 , n151 );
buf ( g151 , n152 );
buf ( g152 , n153 );
buf ( g153 , n154 );
buf ( g154 , n155 );
buf ( g155 , n156 );
buf ( g156 , n157 );
buf ( g157 , n158 );
buf ( g158 , n159 );
buf ( g159 , n160 );
buf ( g160 , n161 );
buf ( g161 , n162 );
buf ( g162 , n163 );
buf ( g163 , n164 );
buf ( g164 , n165 );
buf ( g165 , n166 );
buf ( g166 , n167 );
buf ( n137 , n771 );
buf ( n138 , n363 );
buf ( n139 , n413 );
buf ( n140 , n1532 );
buf ( n141 , n905 );
buf ( n142 , n910 );
buf ( n143 , n1537 );
buf ( n144 , n1678 );
buf ( n145 , n810 );
buf ( n146 , n368 );
buf ( n147 , n863 );
buf ( n148 , n1990 );
buf ( n149 , n1257 );
buf ( n150 , n1112 );
buf ( n151 , n1734 );
buf ( n152 , n900 );
buf ( n153 , n408 );
buf ( n154 , n947 );
buf ( n155 , n1770 );
buf ( n156 , n2023 );
buf ( n157 , n1420 );
buf ( n158 , n1928 );
buf ( n159 , n1959 );
buf ( n160 , n1474 );
buf ( n161 , n2019 );
buf ( n162 , n1812 );
buf ( n163 , n578 );
buf ( n164 , n1872 );
buf ( n165 , n1905 );
buf ( n166 , n1506 );
buf ( n167 , n1910 );
xor ( n170 , n27 , n28 );
xor ( n171 , n29 , n30 );
nor ( n172 , n170 , n171 );
xor ( n173 , n24 , n23 );
xor ( n174 , n25 , n26 );
nor ( n175 , n173 , n174 );
and ( n176 , n172 , n175 );
not ( n177 , n176 );
xor ( n178 , n26 , n25 );
and ( n179 , n24 , n23 );
not ( n180 , n24 );
not ( n181 , n23 );
and ( n182 , n180 , n181 );
nor ( n183 , n179 , n182 );
nand ( n184 , n178 , n183 );
not ( n185 , n184 );
nand ( n186 , n185 , n172 );
nand ( n187 , n177 , n186 );
not ( n188 , n187 );
and ( n189 , n34 , n33 );
not ( n190 , n34 );
not ( n191 , n33 );
and ( n192 , n190 , n191 );
nor ( n193 , n189 , n192 );
not ( n194 , n193 );
xor ( n195 , n32 , n31 );
not ( n196 , n195 );
nand ( n197 , n194 , n196 );
not ( n198 , n197 );
not ( n199 , n198 );
not ( n200 , n171 );
not ( n201 , n175 );
and ( n202 , n200 , n201 );
xnor ( n203 , n25 , n26 );
nand ( n204 , n203 , n173 );
not ( n205 , n171 );
not ( n206 , n205 );
and ( n207 , n204 , n206 );
nor ( n208 , n202 , n207 );
not ( n209 , n170 );
nand ( n210 , n208 , n209 );
not ( n211 , n210 );
or ( n212 , n199 , n211 );
nand ( n213 , n195 , n193 );
not ( n214 , n213 );
not ( n215 , n171 );
nand ( n216 , n215 , n170 );
not ( n217 , n216 );
nor ( n218 , n173 , n174 );
and ( n219 , n217 , n218 );
not ( n220 , n219 );
or ( n221 , n214 , n220 );
nand ( n222 , n221 , n197 );
nand ( n223 , n212 , n222 );
not ( n224 , n213 );
nand ( n225 , n176 , n224 );
nor ( n226 , n197 , n209 );
nand ( n227 , n208 , n226 );
not ( n228 , n171 );
nor ( n229 , n228 , n170 );
not ( n230 , n193 );
nor ( n231 , n230 , n195 );
nand ( n232 , n229 , n231 , n185 );
and ( n233 , n225 , n227 , n232 );
nand ( n234 , n223 , n233 );
not ( n235 , n231 );
nand ( n236 , n229 , n218 );
nand ( n237 , n171 , n170 );
not ( n238 , n237 );
not ( n239 , n183 );
nand ( n240 , n239 , n178 );
not ( n241 , n240 );
nand ( n242 , n238 , n241 );
and ( n243 , n236 , n242 );
not ( n244 , n173 );
xor ( n245 , n25 , n26 );
nor ( n246 , n244 , n245 );
nand ( n247 , n217 , n246 );
nand ( n248 , n243 , n247 );
not ( n249 , n248 );
or ( n250 , n235 , n249 );
nor ( n251 , n171 , n170 );
nand ( n252 , n241 , n251 );
nand ( n253 , n252 , n195 );
not ( n254 , n241 );
not ( n255 , n216 );
not ( n256 , n255 );
or ( n257 , n254 , n256 );
nand ( n258 , n257 , n196 );
nand ( n259 , n253 , n258 , n193 );
nand ( n260 , n250 , n259 );
nor ( n261 , n234 , n260 );
not ( n262 , n261 );
not ( n263 , n236 );
nand ( n264 , n194 , n195 );
not ( n265 , n264 );
nand ( n266 , n263 , n265 );
nor ( n267 , n205 , n184 );
nand ( n268 , n267 , n170 );
not ( n269 , n268 );
nand ( n270 , n251 , n246 );
not ( n271 , n270 );
or ( n272 , n269 , n271 );
nand ( n273 , n272 , n195 );
nand ( n274 , n229 , n241 );
not ( n275 , n274 );
nand ( n276 , n275 , n198 );
nand ( n277 , n266 , n273 , n276 );
not ( n278 , n247 );
not ( n279 , n186 );
or ( n280 , n278 , n279 );
nand ( n281 , n280 , n198 );
nand ( n282 , n238 , n218 );
not ( n283 , n282 );
nand ( n284 , n255 , n241 );
not ( n285 , n284 );
or ( n286 , n283 , n285 );
nand ( n287 , n286 , n224 );
nand ( n288 , n281 , n287 );
nor ( n289 , n277 , n288 );
not ( n290 , n274 );
not ( n291 , n210 );
or ( n292 , n290 , n291 );
nand ( n293 , n292 , n194 );
nand ( n294 , n238 , n246 );
not ( n295 , n294 );
nand ( n296 , n255 , n185 );
not ( n297 , n296 );
or ( n298 , n295 , n297 );
nand ( n299 , n298 , n224 );
not ( n300 , n252 );
not ( n301 , n296 );
or ( n302 , n300 , n301 );
nand ( n303 , n302 , n198 );
not ( n304 , n186 );
nand ( n305 , n304 , n197 , n213 );
and ( n306 , n293 , n299 , n303 , n305 );
nand ( n307 , n289 , n306 );
nor ( n308 , n262 , n307 );
not ( n309 , n308 );
or ( n310 , n188 , n309 );
not ( n311 , n294 );
nor ( n312 , n311 , n253 );
not ( n313 , n268 );
or ( n314 , n258 , n313 );
nand ( n315 , n314 , n194 );
nor ( n316 , n312 , n315 );
and ( n317 , n219 , n224 );
nor ( n318 , n316 , n317 );
not ( n319 , n233 );
not ( n320 , n224 );
nand ( n321 , n236 , n247 );
not ( n322 , n321 );
or ( n323 , n320 , n322 );
not ( n324 , n270 );
not ( n325 , n264 );
and ( n326 , n324 , n325 );
not ( n327 , n282 );
and ( n328 , n327 , n198 );
nor ( n329 , n326 , n328 );
nand ( n330 , n323 , n329 );
nor ( n331 , n319 , n330 );
nand ( n332 , n318 , n331 );
not ( n333 , n265 );
not ( n334 , n267 );
nand ( n335 , n236 , n242 , n334 );
not ( n336 , n335 );
or ( n337 , n333 , n336 );
not ( n338 , n288 );
nand ( n339 , n337 , n338 );
not ( n340 , n277 );
not ( n341 , n243 );
nand ( n342 , n246 , n206 );
and ( n343 , n296 , n274 , n342 );
not ( n344 , n343 );
or ( n345 , n341 , n344 );
nand ( n346 , n345 , n231 );
nand ( n347 , n340 , n346 );
nor ( n348 , n332 , n339 , n347 );
nand ( n349 , n310 , n348 );
not ( n350 , n349 );
not ( n351 , n22 );
and ( n352 , n350 , n351 );
and ( n353 , n349 , n22 );
nor ( n354 , n352 , n353 );
nand ( n355 , n3 , n18 , n17 , n19 );
not ( n356 , n355 );
nand ( n357 , n354 , n356 );
and ( n358 , n355 , n3 );
and ( n359 , n358 , n21 );
not ( n360 , n3 );
and ( n361 , n360 , n20 );
nor ( n362 , n359 , n361 );
nand ( n363 , n357 , n362 );
not ( n364 , n354 );
or ( n365 , n364 , n356 );
not ( n366 , n74 );
or ( n367 , n355 , n366 );
nand ( n368 , n365 , n367 );
and ( n369 , n204 , n240 , n194 );
nor ( n370 , n369 , n187 );
nor ( n371 , n370 , n277 );
and ( n372 , n371 , n306 , n346 , n318 );
not ( n373 , n338 );
nor ( n374 , n373 , n234 );
not ( n375 , n187 );
nand ( n376 , n375 , n339 );
nand ( n377 , n372 , n374 , n376 );
and ( n378 , n339 , n241 );
not ( n379 , n274 );
not ( n380 , n231 );
and ( n381 , n379 , n380 );
and ( n382 , n313 , n265 );
nor ( n383 , n381 , n382 );
nand ( n384 , n281 , n383 );
nor ( n385 , n330 , n384 );
and ( n386 , n270 , n186 );
or ( n387 , n238 , n251 );
nand ( n388 , n387 , n241 );
nand ( n389 , n386 , n294 , n296 , n388 );
nand ( n390 , n389 , n231 );
not ( n391 , n177 );
and ( n392 , n296 , n342 );
not ( n393 , n392 );
or ( n394 , n391 , n393 );
nand ( n395 , n394 , n224 );
nand ( n396 , n385 , n390 , n395 , n223 );
nor ( n397 , n378 , n396 );
nand ( n398 , n377 , n397 );
not ( n399 , n398 );
not ( n400 , n37 );
and ( n401 , n399 , n400 );
and ( n402 , n398 , n37 );
nor ( n403 , n401 , n402 );
not ( n404 , n403 );
or ( n405 , n404 , n356 );
not ( n406 , n110 );
or ( n407 , n355 , n406 );
nand ( n408 , n405 , n407 );
nand ( n409 , n403 , n356 );
and ( n410 , n358 , n36 );
and ( n411 , n360 , n35 );
nor ( n412 , n410 , n411 );
nand ( n413 , n409 , n412 );
xor ( n414 , n40 , n41 );
not ( n415 , n414 );
xor ( n416 , n44 , n45 );
nand ( n417 , n415 , n416 );
not ( n418 , n417 );
not ( n419 , n418 );
not ( n420 , n49 );
not ( n421 , n48 );
or ( n422 , n420 , n421 );
not ( n423 , n48 );
not ( n424 , n49 );
nand ( n425 , n423 , n424 );
nand ( n426 , n422 , n425 );
not ( n427 , n426 );
xor ( n428 , n50 , n51 );
nand ( n429 , n427 , n428 );
not ( n430 , n429 );
not ( n431 , n46 );
not ( n432 , n47 );
and ( n433 , n431 , n432 );
and ( n434 , n46 , n47 );
nor ( n435 , n433 , n434 );
xor ( n436 , n43 , n42 );
nand ( n437 , n435 , n436 );
not ( n438 , n437 );
nand ( n439 , n430 , n438 );
nand ( n440 , n426 , n428 );
not ( n441 , n440 );
not ( n442 , n435 );
nand ( n443 , n442 , n436 );
not ( n444 , n443 );
nand ( n445 , n441 , n444 );
nand ( n446 , n439 , n445 );
not ( n447 , n446 );
or ( n448 , n419 , n447 );
not ( n449 , n435 );
not ( n450 , n436 );
nand ( n451 , n449 , n450 );
and ( n452 , n451 , n437 );
not ( n453 , n452 );
not ( n454 , n428 );
nand ( n455 , n454 , n426 );
not ( n456 , n455 );
nor ( n457 , n415 , n416 );
and ( n458 , n456 , n457 );
nand ( n459 , n453 , n458 );
nand ( n460 , n448 , n459 );
not ( n461 , n460 );
buf ( n462 , n449 );
not ( n463 , n462 );
not ( n464 , n463 );
nor ( n465 , n461 , n464 );
nor ( n466 , n442 , n436 );
nand ( n467 , n456 , n466 );
not ( n468 , n467 );
nand ( n469 , n414 , n416 );
not ( n470 , n469 );
and ( n471 , n468 , n470 );
not ( n472 , n440 );
not ( n473 , n451 );
nand ( n474 , n472 , n473 );
not ( n475 , n474 );
and ( n476 , n475 , n418 );
nor ( n477 , n471 , n476 );
nand ( n478 , n455 , n429 );
nor ( n479 , n436 , n416 );
not ( n480 , n416 );
nor ( n481 , n450 , n480 );
or ( n482 , n479 , n481 );
nand ( n483 , n482 , n462 );
nor ( n484 , n483 , n414 );
and ( n485 , n478 , n484 );
not ( n486 , n478 );
nor ( n487 , n443 , n469 );
and ( n488 , n486 , n487 );
nor ( n489 , n485 , n488 );
not ( n490 , n457 );
not ( n491 , n490 );
not ( n492 , n427 );
not ( n493 , n479 );
or ( n494 , n492 , n493 );
not ( n495 , n428 );
not ( n496 , n414 );
and ( n497 , n495 , n496 );
and ( n498 , n428 , n414 );
nor ( n499 , n497 , n498 );
not ( n500 , n499 );
nand ( n501 , n494 , n500 );
not ( n502 , n501 );
or ( n503 , n491 , n502 );
not ( n504 , n466 );
not ( n505 , n428 );
nand ( n506 , n505 , n427 );
not ( n507 , n506 );
not ( n508 , n507 );
or ( n509 , n504 , n508 );
nand ( n510 , n509 , n439 );
nand ( n511 , n503 , n510 );
nand ( n512 , n477 , n489 , n511 );
nor ( n513 , n465 , n512 );
nand ( n514 , n507 , n438 );
not ( n515 , n514 );
and ( n516 , n515 , n480 );
and ( n517 , n457 , n444 , n428 );
nor ( n518 , n516 , n517 );
not ( n519 , n518 );
not ( n520 , n464 );
not ( n521 , n478 );
or ( n522 , n520 , n521 );
nand ( n523 , n522 , n414 );
nand ( n524 , n519 , n523 );
nand ( n525 , n456 , n444 );
not ( n526 , n525 );
nand ( n527 , n453 , n441 );
not ( n528 , n527 );
or ( n529 , n526 , n528 );
nand ( n530 , n529 , n457 );
nor ( n531 , n455 , n437 );
nand ( n532 , n531 , n418 );
not ( n533 , n532 );
nor ( n534 , n414 , n416 );
not ( n535 , n534 );
not ( n536 , n531 );
or ( n537 , n535 , n536 );
not ( n538 , n469 );
nand ( n539 , n430 , n538 , n473 );
nand ( n540 , n537 , n539 );
and ( n541 , n441 , n438 , n538 );
nor ( n542 , n533 , n540 , n541 );
not ( n543 , n525 );
and ( n544 , n543 , n538 );
nand ( n545 , n441 , n466 );
nor ( n546 , n545 , n417 );
nor ( n547 , n544 , n546 );
and ( n548 , n524 , n530 , n542 , n547 );
nand ( n549 , n473 , n507 );
not ( n550 , n549 );
not ( n551 , n514 );
nand ( n552 , n430 , n466 );
not ( n553 , n552 );
or ( n554 , n551 , n553 );
nand ( n555 , n554 , n418 );
not ( n556 , n555 );
or ( n557 , n550 , n556 );
nand ( n558 , n557 , n500 );
nand ( n559 , n545 , n549 );
not ( n560 , n559 );
not ( n561 , n457 );
or ( n562 , n560 , n561 );
not ( n563 , n527 );
not ( n564 , n534 );
not ( n565 , n564 );
nand ( n566 , n563 , n565 );
nand ( n567 , n562 , n566 );
not ( n568 , n567 );
nand ( n569 , n513 , n548 , n558 , n568 );
not ( n570 , n128 );
and ( n571 , n569 , n570 );
not ( n572 , n569 );
and ( n573 , n572 , n128 );
nor ( n574 , n571 , n573 );
or ( n575 , n574 , n356 );
not ( n576 , n129 );
or ( n577 , n355 , n576 );
nand ( n578 , n575 , n577 );
not ( n579 , n4 );
not ( n580 , n579 );
xor ( n581 , n14 , n13 );
not ( n582 , n581 );
xor ( n583 , n15 , n16 );
nor ( n584 , n582 , n583 );
buf ( n585 , n584 );
not ( n586 , n585 );
xor ( n587 , n11 , n12 );
buf ( n588 , n587 );
not ( n589 , n588 );
and ( n590 , n10 , n9 );
not ( n591 , n10 );
not ( n592 , n9 );
and ( n593 , n591 , n592 );
nor ( n594 , n590 , n593 );
not ( n595 , n594 );
xor ( n596 , n7 , n8 );
nand ( n597 , n595 , n596 );
not ( n598 , n597 );
xor ( n599 , n5 , n6 );
not ( n600 , n599 );
nand ( n601 , n598 , n600 );
not ( n602 , n601 );
or ( n603 , n589 , n602 );
not ( n604 , n599 );
not ( n605 , n594 );
not ( n606 , n605 );
xor ( n607 , n8 , n7 );
nand ( n608 , n604 , n606 , n607 );
xnor ( n609 , n12 , n11 );
nand ( n610 , n608 , n609 );
nand ( n611 , n603 , n610 );
nand ( n612 , n598 , n599 );
not ( n613 , n612 );
and ( n614 , n588 , n613 );
not ( n615 , n588 );
not ( n616 , n596 );
buf ( n617 , n594 );
nand ( n618 , n616 , n617 , n599 );
not ( n619 , n618 );
and ( n620 , n615 , n619 );
nor ( n621 , n614 , n620 );
nand ( n622 , n611 , n621 );
not ( n623 , n622 );
or ( n624 , n586 , n623 );
not ( n625 , n5 );
not ( n626 , n6 );
and ( n627 , n625 , n626 );
and ( n628 , n5 , n6 );
nor ( n629 , n627 , n628 );
not ( n630 , n629 );
not ( n631 , n596 );
and ( n632 , n605 , n630 , n631 );
not ( n633 , n632 );
nand ( n634 , n633 , n618 );
nand ( n635 , n634 , n585 );
not ( n636 , n635 );
not ( n637 , n583 );
not ( n638 , n629 );
or ( n639 , n637 , n638 );
or ( n640 , n629 , n583 );
nand ( n641 , n639 , n640 );
not ( n642 , n581 );
nor ( n643 , n642 , n587 );
nand ( n644 , n641 , n643 );
not ( n645 , n644 );
and ( n646 , n636 , n645 );
not ( n647 , n612 );
not ( n648 , n618 );
or ( n649 , n647 , n648 );
not ( n650 , n583 );
nor ( n651 , n650 , n581 );
and ( n652 , n651 , n587 );
nand ( n653 , n649 , n652 );
not ( n654 , n653 );
nor ( n655 , n646 , n654 );
nand ( n656 , n624 , n655 );
not ( n657 , n656 );
not ( n658 , n644 );
nand ( n659 , n606 , n607 , n599 );
not ( n660 , n659 );
and ( n661 , n658 , n660 );
not ( n662 , n629 );
nor ( n663 , n662 , n596 , n617 );
buf ( n664 , n663 );
nor ( n665 , n581 , n583 );
nand ( n666 , n665 , n587 );
not ( n667 , n666 );
and ( n668 , n664 , n667 );
nor ( n669 , n661 , n668 );
nand ( n670 , n609 , n665 );
nand ( n671 , n669 , n670 );
not ( n672 , n663 );
nor ( n673 , n629 , n596 );
nand ( n674 , n606 , n673 );
nand ( n675 , n672 , n674 );
not ( n676 , n659 );
nor ( n677 , n675 , n676 );
not ( n678 , n677 );
and ( n679 , n671 , n678 );
not ( n680 , n664 );
nand ( n681 , n581 , n583 );
or ( n682 , n681 , n609 );
nor ( n683 , n680 , n682 );
not ( n684 , n652 );
not ( n685 , n676 );
or ( n686 , n684 , n685 );
nand ( n687 , n673 , n651 );
not ( n688 , n687 );
not ( n689 , n583 );
nor ( n690 , n689 , n607 );
not ( n691 , n607 );
nand ( n692 , n691 , n599 );
or ( n693 , n690 , n692 );
nand ( n694 , n600 , n607 );
or ( n695 , n694 , n689 );
nand ( n696 , n693 , n695 );
not ( n697 , n581 );
not ( n698 , n697 );
nand ( n699 , n696 , n698 );
not ( n700 , n699 );
or ( n701 , n688 , n700 );
buf ( n702 , n606 );
nor ( n703 , n588 , n702 );
nand ( n704 , n701 , n703 );
nand ( n705 , n686 , n704 );
nor ( n706 , n679 , n683 , n705 );
nand ( n707 , n618 , n601 );
not ( n708 , n707 );
not ( n709 , n682 );
nand ( n710 , n677 , n708 , n709 );
not ( n711 , n609 );
not ( n712 , n711 );
nand ( n713 , n613 , n712 );
not ( n714 , n713 );
nand ( n715 , n714 , n665 );
not ( n716 , n608 );
not ( n717 , n666 );
and ( n718 , n716 , n717 );
nand ( n719 , n651 , n609 );
not ( n720 , n719 );
and ( n721 , n707 , n720 );
nor ( n722 , n718 , n721 );
nand ( n723 , n710 , n715 , n722 );
not ( n724 , n723 );
nand ( n725 , n657 , n706 , n724 );
not ( n726 , n643 );
nand ( n727 , n587 , n697 );
nand ( n728 , n726 , n727 , n600 );
nand ( n729 , n728 , n690 );
nor ( n730 , n622 , n729 );
not ( n731 , n632 );
not ( n732 , n731 );
nand ( n733 , n730 , n732 );
not ( n734 , n681 );
nand ( n735 , n613 , n734 );
not ( n736 , n608 );
nand ( n737 , n736 , n651 );
nand ( n738 , n735 , n737 , n712 );
nand ( n739 , n659 , n674 );
not ( n740 , n739 );
not ( n741 , n585 );
or ( n742 , n740 , n741 );
buf ( n743 , n588 );
nand ( n744 , n742 , n743 );
and ( n745 , n738 , n744 );
not ( n746 , n743 );
not ( n747 , n601 );
not ( n748 , n747 );
or ( n749 , n746 , n748 );
not ( n750 , n682 );
and ( n751 , n719 , n666 );
not ( n752 , n751 );
or ( n753 , n750 , n752 );
not ( n754 , n674 );
nand ( n755 , n753 , n754 );
nand ( n756 , n749 , n755 );
not ( n757 , n665 );
not ( n758 , n757 );
and ( n759 , n756 , n758 );
nor ( n760 , n745 , n759 );
nand ( n761 , n733 , n760 );
nor ( n762 , n725 , n761 );
not ( n763 , n762 );
or ( n764 , n580 , n763 );
or ( n765 , n579 , n762 );
nand ( n766 , n764 , n765 );
or ( n767 , n766 , n355 );
and ( n768 , n358 , n2 );
and ( n769 , n360 , n1 );
nor ( n770 , n768 , n769 );
nand ( n771 , n767 , n770 );
not ( n772 , n73 );
not ( n773 , n356 );
or ( n774 , n772 , n773 );
not ( n775 , n439 );
and ( n776 , n775 , n565 );
and ( n777 , n457 , n507 , n444 );
nor ( n778 , n776 , n777 );
not ( n779 , n426 );
not ( n780 , n481 );
or ( n781 , n779 , n780 );
nand ( n782 , n781 , n499 );
and ( n783 , n501 , n782 , n463 );
nor ( n784 , n474 , n564 );
nor ( n785 , n783 , n784 );
not ( n786 , n467 );
not ( n787 , n490 );
and ( n788 , n786 , n787 );
and ( n789 , n430 , n444 , n534 );
nor ( n790 , n788 , n789 );
not ( n791 , n549 );
not ( n792 , n445 );
or ( n793 , n791 , n792 );
nand ( n794 , n793 , n418 );
nand ( n795 , n778 , n785 , n790 , n794 );
nor ( n796 , n510 , n475 );
nor ( n797 , n796 , n469 );
nor ( n798 , n795 , n797 );
or ( n799 , n559 , n543 );
nand ( n800 , n799 , n534 );
nand ( n801 , n786 , n418 );
nand ( n802 , n800 , n801 );
nand ( n803 , n538 , n456 , n473 );
nand ( n804 , n555 , n803 );
nor ( n805 , n802 , n804 );
nand ( n806 , n798 , n548 , n805 );
not ( n807 , n53 );
xor ( n808 , n806 , n807 );
or ( n809 , n808 , n356 );
nand ( n810 , n774 , n809 );
and ( n811 , n663 , n584 , n587 );
nor ( n812 , n731 , n666 );
nor ( n813 , n811 , n812 );
not ( n814 , n813 );
nor ( n815 , n588 , n681 );
not ( n816 , n815 );
not ( n817 , n619 );
or ( n818 , n816 , n817 );
nor ( n819 , n731 , n670 );
not ( n820 , n819 );
nand ( n821 , n818 , n820 );
nor ( n822 , n814 , n821 );
and ( n823 , n822 , n715 , n653 );
not ( n824 , n713 );
not ( n825 , n585 );
not ( n826 , n825 );
and ( n827 , n824 , n826 );
not ( n828 , n709 );
not ( n829 , n675 );
or ( n830 , n828 , n829 );
or ( n831 , n608 , n670 );
nand ( n832 , n830 , n831 );
nor ( n833 , n827 , n832 );
not ( n834 , n833 );
or ( n835 , n699 , n728 );
nand ( n836 , n835 , n669 );
nor ( n837 , n834 , n836 );
not ( n838 , n702 );
not ( n839 , n838 );
not ( n840 , n751 );
or ( n841 , n839 , n840 );
nand ( n842 , n841 , n730 );
nand ( n843 , n747 , n698 );
not ( n844 , n843 );
not ( n845 , n727 );
nand ( n846 , n845 , n619 );
not ( n847 , n846 );
or ( n848 , n844 , n847 );
nand ( n849 , n848 , n689 );
not ( n850 , n751 );
nand ( n851 , n850 , n676 );
and ( n852 , n849 , n851 );
nand ( n853 , n823 , n837 , n842 , n852 );
nor ( n854 , n853 , n761 );
and ( n855 , n854 , n75 );
not ( n856 , n854 );
not ( n857 , n75 );
and ( n858 , n856 , n857 );
nor ( n859 , n855 , n858 );
or ( n860 , n859 , n356 );
not ( n861 , n76 );
or ( n862 , n355 , n861 );
nand ( n863 , n860 , n862 );
not ( n864 , n635 );
not ( n865 , n737 );
or ( n866 , n864 , n865 );
nand ( n867 , n866 , n743 );
not ( n868 , n611 );
and ( n869 , n868 , n734 );
nand ( n870 , n719 , n757 );
and ( n871 , n739 , n870 );
nor ( n872 , n869 , n871 );
and ( n873 , n720 , n598 );
nor ( n874 , n873 , n819 );
and ( n875 , n867 , n833 , n872 , n874 );
not ( n876 , n734 );
not ( n877 , n712 );
not ( n878 , n618 );
or ( n879 , n877 , n878 );
nand ( n880 , n659 , n588 );
nand ( n881 , n879 , n880 );
nand ( n882 , n881 , n713 );
not ( n883 , n882 );
or ( n884 , n876 , n883 );
not ( n885 , n652 );
nand ( n886 , n885 , n670 );
nand ( n887 , n886 , n664 );
nand ( n888 , n884 , n887 );
not ( n889 , n888 );
nand ( n890 , n875 , n733 , n657 , n889 );
not ( n891 , n890 );
not ( n892 , n55 );
and ( n893 , n891 , n892 );
and ( n894 , n890 , n55 );
nor ( n895 , n893 , n894 );
not ( n896 , n895 );
or ( n897 , n896 , n356 );
not ( n898 , n109 );
or ( n899 , n355 , n898 );
nand ( n900 , n897 , n899 );
or ( n901 , n808 , n355 );
and ( n902 , n358 , n20 );
and ( n903 , n360 , n52 );
nor ( n904 , n902 , n903 );
nand ( n905 , n901 , n904 );
nand ( n906 , n895 , n356 );
and ( n907 , n358 , n35 );
and ( n908 , n360 , n54 );
nor ( n909 , n907 , n908 );
nand ( n910 , n906 , n909 );
not ( n911 , n540 );
not ( n912 , n483 );
and ( n913 , n912 , n414 , n430 );
nor ( n914 , n913 , n517 );
nand ( n915 , n911 , n477 , n778 , n914 );
not ( n916 , n915 );
not ( n917 , n538 );
not ( n918 , n552 );
not ( n919 , n918 );
or ( n920 , n917 , n919 );
not ( n921 , n541 );
nand ( n922 , n920 , n921 );
nor ( n923 , n922 , n460 );
not ( n924 , n514 );
not ( n925 , n525 );
or ( n926 , n924 , n925 );
nand ( n927 , n926 , n538 );
nand ( n928 , n441 , n438 );
not ( n929 , n928 );
not ( n930 , n467 );
or ( n931 , n929 , n930 );
nand ( n932 , n931 , n565 );
not ( n933 , n453 );
nand ( n934 , n933 , n507 , n418 );
nand ( n935 , n927 , n932 , n934 );
nor ( n936 , n796 , n490 );
nor ( n937 , n935 , n936 );
nand ( n938 , n916 , n923 , n937 , n805 );
not ( n939 , n111 );
and ( n940 , n938 , n939 );
not ( n941 , n938 );
and ( n942 , n941 , n111 );
nor ( n943 , n940 , n942 );
or ( n944 , n943 , n356 );
not ( n945 , n112 );
or ( n946 , n355 , n945 );
nand ( n947 , n944 , n946 );
and ( n948 , n64 , n104 );
not ( n949 , n64 );
not ( n950 , n104 );
and ( n951 , n949 , n950 );
nor ( n952 , n948 , n951 );
not ( n953 , n952 );
xor ( n954 , n62 , n103 );
nor ( n955 , n953 , n954 );
not ( n956 , n955 );
xor ( n957 , n101 , n102 );
not ( n958 , n957 );
not ( n959 , n98 );
not ( n960 , n99 );
and ( n961 , n959 , n960 );
and ( n962 , n98 , n99 );
nor ( n963 , n961 , n962 );
nor ( n964 , n958 , n963 );
not ( n965 , n964 );
nor ( n966 , n956 , n965 );
not ( n967 , n966 );
nor ( n968 , n963 , n957 );
nor ( n969 , n952 , n954 );
nand ( n970 , n968 , n969 );
nand ( n971 , n967 , n970 );
not ( n972 , n8 );
not ( n973 , n100 );
and ( n974 , n972 , n973 );
and ( n975 , n8 , n100 );
nor ( n976 , n974 , n975 );
xor ( n977 , n6 , n105 );
nand ( n978 , n976 , n977 );
not ( n979 , n978 );
and ( n980 , n971 , n979 );
and ( n981 , n964 , n969 );
not ( n982 , n981 );
not ( n983 , n976 );
not ( n984 , n983 );
not ( n985 , n977 );
nand ( n986 , n984 , n985 );
nor ( n987 , n982 , n986 );
nor ( n988 , n980 , n987 );
buf ( n989 , n957 );
not ( n990 , n989 );
not ( n991 , n990 );
not ( n992 , n963 );
not ( n993 , n992 );
and ( n994 , n969 , n993 );
not ( n995 , n994 );
or ( n996 , n991 , n995 );
nand ( n997 , n968 , n955 );
nand ( n998 , n996 , n997 );
nor ( n999 , n976 , n977 );
buf ( n1000 , n999 );
nand ( n1001 , n998 , n1000 );
nand ( n1002 , n988 , n1001 );
not ( n1003 , n986 );
not ( n1004 , n1003 );
not ( n1005 , n966 );
or ( n1006 , n1004 , n1005 );
and ( n1007 , n952 , n954 );
not ( n1008 , n963 );
nor ( n1009 , n1008 , n957 );
nand ( n1010 , n1007 , n1009 );
not ( n1011 , n1010 );
nand ( n1012 , n1011 , n979 );
nand ( n1013 , n1006 , n1012 );
not ( n1014 , n1000 );
nand ( n1015 , n955 , n1009 );
not ( n1016 , n1015 );
not ( n1017 , n1016 );
or ( n1018 , n1014 , n1017 );
nand ( n1019 , n955 , n993 );
not ( n1020 , n1019 );
not ( n1021 , n976 );
nand ( n1022 , n1021 , n977 );
not ( n1023 , n1022 );
nand ( n1024 , n1020 , n1023 , n989 );
nand ( n1025 , n1018 , n1024 );
nor ( n1026 , n1013 , n1025 );
nor ( n1027 , n957 , n977 );
nand ( n1028 , n969 , n1027 );
not ( n1029 , n1028 );
not ( n1030 , n978 );
nor ( n1031 , n1030 , n999 );
nor ( n1032 , n997 , n1031 );
not ( n1033 , n1032 );
not ( n1034 , n1033 );
or ( n1035 , n1029 , n1034 );
not ( n1036 , n983 );
buf ( n1037 , n1036 );
nand ( n1038 , n1035 , n1037 );
nand ( n1039 , n1026 , n1038 );
nor ( n1040 , n1002 , n1039 );
nand ( n1041 , n981 , n1023 );
nand ( n1042 , n994 , n999 , n989 );
and ( n1043 , n1041 , n1042 );
not ( n1044 , n952 );
not ( n1045 , n957 );
nand ( n1046 , n1044 , n1045 , n1036 );
nand ( n1047 , n1046 , n986 );
and ( n1048 , n957 , n954 );
nand ( n1049 , n1047 , n1048 );
not ( n1050 , n1049 );
not ( n1051 , n1044 );
not ( n1052 , n1051 );
nand ( n1053 , n1050 , n1052 );
nand ( n1054 , n1043 , n1053 );
and ( n1055 , n968 , n1007 );
not ( n1056 , n1055 );
not ( n1057 , n1056 );
not ( n1058 , n1009 );
nand ( n1059 , n1058 , n1044 , n954 , n965 );
not ( n1060 , n1059 );
or ( n1061 , n1057 , n1060 );
nand ( n1062 , n1061 , n1000 );
nand ( n1063 , n1048 , n1023 );
nand ( n1064 , n1062 , n1063 );
nor ( n1065 , n1054 , n1064 );
not ( n1066 , n989 );
not ( n1067 , n1020 );
or ( n1068 , n1066 , n1067 );
nand ( n1069 , n1068 , n1056 );
buf ( n1070 , n1003 );
nand ( n1071 , n1069 , n1070 );
nand ( n1072 , n1007 , n964 );
not ( n1073 , n1072 );
and ( n1074 , n1073 , n1000 );
nor ( n1075 , n1010 , n1022 );
nor ( n1076 , n1074 , n1075 );
not ( n1077 , n1044 );
not ( n1078 , n1077 );
not ( n1079 , n1045 );
and ( n1080 , n1078 , n1079 );
and ( n1081 , n1051 , n1045 );
nor ( n1082 , n1080 , n1081 );
not ( n1083 , n992 );
and ( n1084 , n1083 , n954 );
nand ( n1085 , n1082 , n1084 );
not ( n1086 , n1085 );
nand ( n1087 , n1086 , n979 );
nand ( n1088 , n1071 , n1076 , n1087 );
not ( n1089 , n1088 );
not ( n1090 , n954 );
nor ( n1091 , n1090 , n985 );
not ( n1092 , n1091 );
not ( n1093 , n1047 );
or ( n1094 , n1092 , n1093 );
nand ( n1095 , n1094 , n1049 );
and ( n1096 , n989 , n979 );
not ( n1097 , n989 );
and ( n1098 , n1097 , n1023 );
or ( n1099 , n1096 , n1098 );
and ( n1100 , n1099 , n969 );
or ( n1101 , n1095 , n1100 );
nand ( n1102 , n1101 , n1083 );
nand ( n1103 , n1040 , n1065 , n1089 , n1102 );
not ( n1104 , n97 );
and ( n1105 , n1103 , n1104 );
not ( n1106 , n1103 );
and ( n1107 , n1106 , n97 );
nor ( n1108 , n1105 , n1107 );
or ( n1109 , n1108 , n356 );
not ( n1110 , n106 );
or ( n1111 , n355 , n1110 );
nand ( n1112 , n1109 , n1111 );
xor ( n1113 , n90 , n91 );
not ( n1114 , n1113 );
xor ( n1115 , n88 , n89 );
nand ( n1116 , n1114 , n1115 );
not ( n1117 , n1116 );
not ( n1118 , n1117 );
and ( n1119 , n14 , n94 );
not ( n1120 , n14 );
not ( n1121 , n94 );
and ( n1122 , n1120 , n1121 );
nor ( n1123 , n1119 , n1122 );
not ( n1124 , n1123 );
xor ( n1125 , n16 , n95 );
nand ( n1126 , n1124 , n1125 );
not ( n1127 , n1126 );
xor ( n1128 , n26 , n93 );
not ( n1129 , n1128 );
nand ( n1130 , n1127 , n1129 );
not ( n1131 , n1130 );
not ( n1132 , n1131 );
or ( n1133 , n1118 , n1132 );
nand ( n1134 , n1128 , n1115 );
not ( n1135 , n1134 );
not ( n1136 , n1123 );
nor ( n1137 , n1136 , n1125 );
or ( n1138 , n1135 , n1137 );
nand ( n1139 , n1135 , n1126 );
not ( n1140 , n1128 );
not ( n1141 , n1115 );
and ( n1142 , n1140 , n1141 );
nor ( n1143 , n1142 , n1114 );
nand ( n1144 , n1138 , n1139 , n1143 );
nand ( n1145 , n1133 , n1144 );
not ( n1146 , n92 );
not ( n1147 , n24 );
or ( n1148 , n1146 , n1147 );
or ( n1149 , n24 , n92 );
nand ( n1150 , n1148 , n1149 );
buf ( n1151 , n1150 );
buf ( n1152 , n1151 );
and ( n1153 , n1145 , n1152 );
and ( n1154 , n1137 , n1129 );
not ( n1155 , n1154 );
not ( n1156 , n1113 );
nor ( n1157 , n1156 , n1115 );
nand ( n1158 , n1157 , n1150 );
not ( n1159 , n1158 );
not ( n1160 , n1159 );
or ( n1161 , n1155 , n1160 );
and ( n1162 , n1150 , n1114 , n1128 );
nand ( n1163 , n1162 , n1137 );
nand ( n1164 , n1161 , n1163 );
nor ( n1165 , n1113 , n1115 );
and ( n1166 , n1165 , n1150 );
and ( n1167 , n1164 , n1166 );
nor ( n1168 , n1153 , n1167 );
xor ( n1169 , n24 , n92 );
buf ( n1170 , n1169 );
not ( n1171 , n1170 );
nor ( n1172 , n1130 , n1115 );
not ( n1173 , n1172 );
or ( n1174 , n1171 , n1173 );
nor ( n1175 , n1128 , n1123 );
nand ( n1176 , n1159 , n1175 );
nand ( n1177 , n1174 , n1176 );
and ( n1178 , n1170 , n1114 );
nand ( n1179 , n1150 , n1115 );
nor ( n1180 , n1114 , n1179 );
nor ( n1181 , n1178 , n1180 );
not ( n1182 , n1123 );
nand ( n1183 , n1182 , n1128 );
not ( n1184 , n1183 );
not ( n1185 , n1125 );
nand ( n1186 , n1184 , n1185 );
nor ( n1187 , n1181 , n1186 );
nor ( n1188 , n1177 , n1187 );
nand ( n1189 , n1123 , n1125 );
not ( n1190 , n1189 );
nand ( n1191 , n1190 , n1128 );
and ( n1192 , n1191 , n1170 );
not ( n1193 , n1151 );
nand ( n1194 , n1129 , n1185 , n1182 );
not ( n1195 , n1194 );
or ( n1196 , n1193 , n1195 );
buf ( n1197 , n1165 );
nand ( n1198 , n1196 , n1197 );
nor ( n1199 , n1192 , n1198 );
nand ( n1200 , n1115 , n1169 );
nor ( n1201 , n1129 , n1200 );
not ( n1202 , n1201 );
not ( n1203 , n1137 );
nand ( n1204 , n1203 , n1113 );
not ( n1205 , n1204 );
or ( n1206 , n1202 , n1205 );
not ( n1207 , n1157 );
nor ( n1208 , n1191 , n1207 );
not ( n1209 , n1208 );
nand ( n1210 , n1206 , n1209 );
nor ( n1211 , n1137 , n1127 );
nor ( n1212 , n1200 , n1114 );
and ( n1213 , n1211 , n1212 , n1129 );
nor ( n1214 , n1199 , n1210 , n1213 );
not ( n1215 , n1154 );
and ( n1216 , n1151 , n1116 );
not ( n1217 , n1151 );
not ( n1218 , n1165 );
and ( n1219 , n1217 , n1218 );
nor ( n1220 , n1216 , n1219 );
not ( n1221 , n1220 );
or ( n1222 , n1215 , n1221 );
nor ( n1223 , n1186 , n1113 );
nand ( n1224 , n1190 , n1129 );
not ( n1225 , n1224 );
or ( n1226 , n1223 , n1225 );
not ( n1227 , n1179 );
nand ( n1228 , n1226 , n1227 );
nand ( n1229 , n1222 , n1228 );
not ( n1230 , n1229 );
nand ( n1231 , n1168 , n1188 , n1214 , n1230 );
nand ( n1232 , n1154 , n1117 );
not ( n1233 , n1157 );
not ( n1234 , n1233 );
not ( n1235 , n1194 );
nand ( n1236 , n1234 , n1235 );
nand ( n1237 , n1232 , n1236 );
nor ( n1238 , n1144 , n1185 );
or ( n1239 , n1237 , n1238 );
nand ( n1240 , n1239 , n1170 );
nor ( n1241 , n1183 , n1185 );
not ( n1242 , n1241 );
nand ( n1243 , n1242 , n1224 );
and ( n1244 , n1243 , n1166 );
and ( n1245 , n1208 , n1152 );
nor ( n1246 , n1244 , n1245 );
nand ( n1247 , n1240 , n1246 );
nor ( n1248 , n1231 , n1247 );
not ( n1249 , n1248 );
not ( n1250 , n87 );
and ( n1251 , n1249 , n1250 );
and ( n1252 , n1248 , n87 );
nor ( n1253 , n1251 , n1252 );
or ( n1254 , n1253 , n356 );
not ( n1255 , n96 );
or ( n1256 , n355 , n1255 );
nand ( n1257 , n1254 , n1256 );
and ( n1258 , n41 , n78 );
not ( n1259 , n41 );
not ( n1260 , n78 );
and ( n1261 , n1259 , n1260 );
nor ( n1262 , n1258 , n1261 );
xor ( n1263 , n80 , n81 );
nand ( n1264 , n1262 , n1263 );
xor ( n1265 , n45 , n79 );
not ( n1266 , n1265 );
xor ( n1267 , n70 , n85 );
nand ( n1268 , n1266 , n1267 );
nor ( n1269 , n1264 , n1268 );
not ( n1270 , n1269 );
nor ( n1271 , n1263 , n1262 );
not ( n1272 , n1271 );
and ( n1273 , n83 , n82 );
not ( n1274 , n83 );
not ( n1275 , n82 );
and ( n1276 , n1274 , n1275 );
nor ( n1277 , n1273 , n1276 );
not ( n1278 , n1277 );
not ( n1279 , n1278 );
and ( n1280 , n1272 , n1279 );
buf ( n1281 , n1278 );
and ( n1282 , n1264 , n1281 );
nor ( n1283 , n1280 , n1282 );
not ( n1284 , n84 );
not ( n1285 , n66 );
or ( n1286 , n1284 , n1285 );
or ( n1287 , n66 , n84 );
nand ( n1288 , n1286 , n1287 );
and ( n1289 , n1266 , n1288 );
not ( n1290 , n1266 );
xor ( n1291 , n66 , n84 );
and ( n1292 , n1290 , n1291 );
nor ( n1293 , n1289 , n1292 );
nand ( n1294 , n1283 , n1293 );
not ( n1295 , n1265 );
nand ( n1296 , n1295 , n1277 );
not ( n1297 , n1296 );
not ( n1298 , n1264 );
and ( n1299 , n1297 , n1298 );
not ( n1300 , n1299 );
not ( n1301 , n1262 );
nor ( n1302 , n1301 , n1263 );
nand ( n1303 , n1265 , n1277 );
not ( n1304 , n1303 );
nand ( n1305 , n1302 , n1304 );
not ( n1306 , n1262 );
nand ( n1307 , n1306 , n1263 );
not ( n1308 , n1307 );
nor ( n1309 , n1265 , n1277 );
nand ( n1310 , n1308 , n1309 );
nand ( n1311 , n1294 , n1300 , n1305 , n1310 );
not ( n1312 , n1311 );
not ( n1313 , n1312 );
or ( n1314 , n1270 , n1313 );
and ( n1315 , n1278 , n1265 );
nand ( n1316 , n1315 , n1302 );
not ( n1317 , n1316 );
nor ( n1318 , n1267 , n1291 );
not ( n1319 , n1318 );
not ( n1320 , n1319 );
nand ( n1321 , n1317 , n1320 );
buf ( n1322 , n1267 );
buf ( n1323 , n1288 );
nand ( n1324 , n1271 , n1297 , n1322 , n1323 );
not ( n1325 , n1310 );
nand ( n1326 , n1271 , n1315 );
not ( n1327 , n1326 );
or ( n1328 , n1325 , n1327 );
not ( n1329 , n1267 );
and ( n1330 , n1329 , n1291 );
nand ( n1331 , n1328 , n1330 );
nand ( n1332 , n1321 , n1324 , n1331 );
not ( n1333 , n1307 );
nand ( n1334 , n1333 , n1315 );
not ( n1335 , n1334 );
nand ( n1336 , n1309 , n1271 );
not ( n1337 , n1336 );
or ( n1338 , n1335 , n1337 );
nand ( n1339 , n1338 , n1320 );
not ( n1340 , n1326 );
and ( n1341 , n1288 , n1267 );
nand ( n1342 , n1340 , n1341 );
nand ( n1343 , n1339 , n1342 );
nor ( n1344 , n1332 , n1343 );
nand ( n1345 , n1314 , n1344 );
not ( n1346 , n1345 );
not ( n1347 , n1267 );
not ( n1348 , n1262 );
not ( n1349 , n1348 );
or ( n1350 , n1347 , n1349 );
or ( n1351 , n1348 , n1267 );
nand ( n1352 , n1350 , n1351 );
not ( n1353 , n1352 );
and ( n1354 , n1288 , n1265 , n1263 );
and ( n1355 , n1353 , n1354 );
and ( n1356 , n1269 , n1291 );
nor ( n1357 , n1355 , n1356 );
not ( n1358 , n1357 );
not ( n1359 , n1281 );
and ( n1360 , n1358 , n1359 );
not ( n1361 , n1322 );
not ( n1362 , n1361 );
and ( n1363 , n1271 , n1297 , n1288 );
not ( n1364 , n1363 );
or ( n1365 , n1362 , n1364 );
not ( n1366 , n1271 );
nand ( n1367 , n1366 , n1264 );
not ( n1368 , n1291 );
not ( n1369 , n1368 );
nand ( n1370 , n1367 , n1304 , n1369 );
nand ( n1371 , n1365 , n1370 );
nor ( n1372 , n1360 , n1371 );
nand ( n1373 , n1271 , n1304 );
not ( n1374 , n1373 );
not ( n1375 , n1316 );
or ( n1376 , n1374 , n1375 );
nand ( n1377 , n1291 , n1267 );
not ( n1378 , n1377 );
nand ( n1379 , n1376 , n1378 );
nand ( n1380 , n1299 , n1320 );
and ( n1381 , n1379 , n1380 );
not ( n1382 , n1322 );
not ( n1383 , n1315 );
nor ( n1384 , n1383 , n1264 );
not ( n1385 , n1384 );
or ( n1386 , n1382 , n1385 );
nand ( n1387 , n1386 , n1305 );
nand ( n1388 , n1387 , n1323 );
not ( n1389 , n1384 );
not ( n1390 , n1307 );
nand ( n1391 , n1390 , n1297 );
nand ( n1392 , n1389 , n1391 );
nand ( n1393 , n1297 , n1302 );
nand ( n1394 , n1336 , n1393 );
or ( n1395 , n1392 , n1394 );
nand ( n1396 , n1395 , n1330 );
nand ( n1397 , n1372 , n1381 , n1388 , n1396 );
nand ( n1398 , n1334 , n1391 );
nand ( n1399 , n1398 , n1378 );
and ( n1400 , n1309 , n1302 );
nor ( n1401 , n1341 , n1330 );
and ( n1402 , n1400 , n1401 );
nor ( n1403 , n1307 , n1303 );
and ( n1404 , n1403 , n1341 );
nor ( n1405 , n1402 , n1404 );
nand ( n1406 , n1299 , n1330 );
not ( n1407 , n1310 );
nand ( n1408 , n1407 , n1320 );
nand ( n1409 , n1399 , n1405 , n1406 , n1408 );
nor ( n1410 , n1397 , n1409 );
nand ( n1411 , n1346 , n1410 );
not ( n1412 , n116 );
and ( n1413 , n1411 , n1412 );
not ( n1414 , n1411 );
and ( n1415 , n1414 , n116 );
nor ( n1416 , n1413 , n1415 );
or ( n1417 , n1416 , n356 );
not ( n1418 , n117 );
or ( n1419 , n355 , n1418 );
nand ( n1420 , n1417 , n1419 );
not ( n1421 , n1023 );
not ( n1422 , n1055 );
or ( n1423 , n1421 , n1422 );
not ( n1424 , n986 );
nand ( n1425 , n1424 , n994 , n989 );
nand ( n1426 , n1423 , n1425 );
not ( n1427 , n1426 );
nor ( n1428 , n1085 , n1037 );
not ( n1429 , n1428 );
not ( n1430 , n1051 );
and ( n1431 , n1430 , n968 , n999 );
nor ( n1432 , n1032 , n1431 );
nand ( n1433 , n1072 , n1015 );
nand ( n1434 , n1433 , n1000 );
nand ( n1435 , n1427 , n1429 , n1432 , n1434 );
nor ( n1436 , n1435 , n1054 );
not ( n1437 , n1000 );
not ( n1438 , n1011 );
or ( n1439 , n1437 , n1438 );
or ( n1440 , n1433 , n981 );
nand ( n1441 , n1440 , n979 );
nand ( n1442 , n1439 , n1441 );
not ( n1443 , n1442 );
nand ( n1444 , n1436 , n1443 );
not ( n1445 , n1082 );
nand ( n1446 , n1023 , n1090 );
nor ( n1447 , n1445 , n1446 );
or ( n1448 , n1095 , n1447 );
not ( n1449 , n1083 );
nand ( n1450 , n1448 , n1449 );
not ( n1451 , n1059 );
nor ( n1452 , n990 , n1037 );
nand ( n1453 , n1451 , n1452 );
not ( n1454 , n1453 );
nand ( n1455 , n1010 , n970 );
nand ( n1456 , n1455 , n1037 );
not ( n1457 , n1456 );
or ( n1458 , n1454 , n1457 );
nand ( n1459 , n1458 , n977 );
or ( n1460 , n1069 , n994 );
nand ( n1461 , n1460 , n1070 );
and ( n1462 , n1047 , n1028 );
nand ( n1463 , n998 , n1462 );
nand ( n1464 , n1450 , n1459 , n1461 , n1463 );
nor ( n1465 , n1444 , n1464 );
not ( n1466 , n1465 );
not ( n1467 , n122 );
and ( n1468 , n1466 , n1467 );
and ( n1469 , n1465 , n122 );
nor ( n1470 , n1468 , n1469 );
or ( n1471 , n1470 , n356 );
not ( n1472 , n123 );
or ( n1473 , n355 , n1472 );
nand ( n1474 , n1471 , n1473 );
not ( n1475 , n645 );
not ( n1476 , n636 );
not ( n1477 , n675 );
nand ( n1478 , n1476 , n1477 );
not ( n1479 , n1478 );
or ( n1480 , n1475 , n1479 );
not ( n1481 , n584 );
nand ( n1482 , n1481 , n609 );
nor ( n1483 , n1482 , n608 );
not ( n1484 , n641 );
nand ( n1485 , n1484 , n598 );
nor ( n1486 , n1485 , n727 );
nor ( n1487 , n1483 , n1486 );
nand ( n1488 , n720 , n676 );
and ( n1489 , n813 , n1487 , n846 , n1488 );
nand ( n1490 , n1480 , n1489 );
nor ( n1491 , n1490 , n723 );
not ( n1492 , n881 );
nand ( n1493 , n1492 , n585 );
nand ( n1494 , n1493 , n755 , n849 );
nor ( n1495 , n1494 , n888 );
nand ( n1496 , n1491 , n1495 );
and ( n1497 , n1496 , n58 );
not ( n1498 , n1496 );
not ( n1499 , n58 );
and ( n1500 , n1498 , n1499 );
nor ( n1501 , n1497 , n1500 );
not ( n1502 , n1501 );
or ( n1503 , n1502 , n356 );
not ( n1504 , n134 );
or ( n1505 , n355 , n1504 );
nand ( n1506 , n1503 , n1505 );
nand ( n1507 , n430 , n479 , n415 , n463 );
nor ( n1508 , n506 , n480 );
nand ( n1509 , n452 , n1508 );
and ( n1510 , n1507 , n1509 , n532 );
nand ( n1511 , n1510 , n547 );
nor ( n1512 , n1511 , n567 );
nand ( n1513 , n441 , n538 );
not ( n1514 , n1513 );
nor ( n1515 , n417 , n436 );
nand ( n1516 , n478 , n1515 );
not ( n1517 , n1516 );
or ( n1518 , n1514 , n1517 );
nand ( n1519 , n1518 , n464 );
and ( n1520 , n1519 , n790 , n518 );
not ( n1521 , n802 );
nand ( n1522 , n1512 , n1520 , n923 , n1521 );
and ( n1523 , n1522 , n39 );
not ( n1524 , n1522 );
not ( n1525 , n39 );
and ( n1526 , n1524 , n1525 );
nor ( n1527 , n1523 , n1526 );
nand ( n1528 , n1527 , n356 );
and ( n1529 , n358 , n1 );
and ( n1530 , n360 , n38 );
nor ( n1531 , n1529 , n1530 );
nand ( n1532 , n1528 , n1531 );
nand ( n1533 , n1501 , n356 );
and ( n1534 , n358 , n57 );
and ( n1535 , n360 , n56 );
nor ( n1536 , n1534 , n1535 );
nand ( n1537 , n1533 , n1536 );
not ( n1538 , n61 );
not ( n1539 , n62 );
and ( n1540 , n1538 , n1539 );
and ( n1541 , n61 , n62 );
nor ( n1542 , n1540 , n1541 );
not ( n1543 , n1542 );
xor ( n1544 , n64 , n63 );
nor ( n1545 , n1543 , n1544 );
buf ( n1546 , n1545 );
not ( n1547 , n1546 );
xor ( n1548 , n66 , n65 );
not ( n1549 , n1548 );
xor ( n1550 , n69 , n70 );
nand ( n1551 , n1549 , n1550 );
not ( n1552 , n1551 );
xor ( n1553 , n72 , n71 );
xor ( n1554 , n67 , n68 );
nor ( n1555 , n1553 , n1554 );
nand ( n1556 , n1552 , n1555 );
not ( n1557 , n1550 );
nand ( n1558 , n1557 , n1548 );
not ( n1559 , n1558 );
not ( n1560 , n1553 );
nand ( n1561 , n1560 , n1554 );
not ( n1562 , n1561 );
nand ( n1563 , n1559 , n1562 );
nand ( n1564 , n1556 , n1563 );
not ( n1565 , n1550 );
not ( n1566 , n1554 );
or ( n1567 , n1565 , n1566 );
or ( n1568 , n1554 , n1550 );
nand ( n1569 , n1567 , n1568 );
buf ( n1570 , n1548 );
and ( n1571 , n1569 , n1553 , n1570 );
nor ( n1572 , n1564 , n1571 );
or ( n1573 , n1547 , n1572 );
nand ( n1574 , n1555 , n1559 );
not ( n1575 , n1574 );
and ( n1576 , n1550 , n1548 );
nand ( n1577 , n1562 , n1576 );
not ( n1578 , n1577 );
or ( n1579 , n1575 , n1578 );
not ( n1580 , n1544 );
nor ( n1581 , n1543 , n1580 );
nand ( n1582 , n1579 , n1581 );
nand ( n1583 , n1573 , n1582 );
or ( n1584 , n1542 , n1544 );
not ( n1585 , n1584 );
not ( n1586 , n1585 );
nand ( n1587 , n1555 , n1576 );
not ( n1588 , n1587 );
not ( n1589 , n1588 );
or ( n1590 , n1586 , n1589 );
and ( n1591 , n1553 , n1554 );
nand ( n1592 , n1552 , n1591 );
not ( n1593 , n1592 );
and ( n1594 , n1593 , n1585 );
nand ( n1595 , n1543 , n1544 );
not ( n1596 , n1595 );
nor ( n1597 , n1551 , n1561 );
and ( n1598 , n1596 , n1597 );
nor ( n1599 , n1594 , n1598 );
nand ( n1600 , n1590 , n1599 );
nor ( n1601 , n1583 , n1600 );
not ( n1602 , n1543 );
nand ( n1603 , n1551 , n1558 );
not ( n1604 , n1603 );
or ( n1605 , n1602 , n1604 );
nor ( n1606 , n1548 , n1550 );
nand ( n1607 , n1606 , n1542 );
nand ( n1608 , n1605 , n1607 );
buf ( n1609 , n1544 );
nor ( n1610 , n1542 , n1548 );
nor ( n1611 , n1609 , n1610 );
not ( n1612 , n1553 );
nor ( n1613 , n1612 , n1554 );
nand ( n1614 , n1608 , n1611 , n1613 );
not ( n1615 , n1563 );
not ( n1616 , n1595 );
and ( n1617 , n1615 , n1616 );
and ( n1618 , n1581 , n1606 , n1555 );
nor ( n1619 , n1617 , n1618 );
nand ( n1620 , n1614 , n1619 );
nand ( n1621 , n1606 , n1591 );
nand ( n1622 , n1621 , n1577 );
nand ( n1623 , n1622 , n1543 );
not ( n1624 , n1556 );
not ( n1625 , n1584 );
and ( n1626 , n1624 , n1625 );
and ( n1627 , n1610 , n1569 , n1609 );
nor ( n1628 , n1626 , n1627 );
nand ( n1629 , n1559 , n1591 );
nand ( n1630 , n1587 , n1629 );
nand ( n1631 , n1630 , n1545 );
nand ( n1632 , n1623 , n1628 , n1631 );
nor ( n1633 , n1620 , n1632 );
not ( n1634 , n1629 );
not ( n1635 , n1581 );
not ( n1636 , n1635 );
and ( n1637 , n1634 , n1636 );
nand ( n1638 , n1613 , n1576 );
not ( n1639 , n1638 );
and ( n1640 , n1639 , n1545 );
nor ( n1641 , n1637 , n1640 );
and ( n1642 , n1597 , n1545 );
nand ( n1643 , n1606 , n1562 );
not ( n1644 , n1643 );
and ( n1645 , n1644 , n1581 );
nor ( n1646 , n1642 , n1645 );
nand ( n1647 , n1641 , n1646 );
nand ( n1648 , n1552 , n1613 );
not ( n1649 , n1648 );
not ( n1650 , n1587 );
or ( n1651 , n1649 , n1650 );
nand ( n1652 , n1651 , n1581 );
not ( n1653 , n1574 );
not ( n1654 , n1584 );
and ( n1655 , n1653 , n1654 );
nand ( n1656 , n1606 , n1613 );
not ( n1657 , n1656 );
and ( n1658 , n1657 , n1596 );
nor ( n1659 , n1655 , n1658 );
nand ( n1660 , n1652 , n1659 );
nor ( n1661 , n1647 , n1660 );
not ( n1662 , n1610 );
not ( n1663 , n1596 );
and ( n1664 , n1662 , n1663 );
and ( n1665 , n1629 , n1638 , n1656 );
nor ( n1666 , n1664 , n1665 );
nand ( n1667 , n1570 , n1666 );
nand ( n1668 , n1601 , n1633 , n1661 , n1667 );
and ( n1669 , n1668 , n60 );
not ( n1670 , n1668 );
not ( n1671 , n60 );
and ( n1672 , n1670 , n1671 );
nor ( n1673 , n1669 , n1672 );
nand ( n1674 , n1673 , n356 );
and ( n1675 , n358 , n38 );
and ( n1676 , n360 , n59 );
nor ( n1677 , n1675 , n1676 );
nand ( n1678 , n1674 , n1677 );
not ( n1679 , n1609 );
and ( n1680 , n1610 , n1569 , n1679 );
or ( n1681 , n1600 , n1680 );
not ( n1682 , n1553 );
nand ( n1683 , n1681 , n1682 );
not ( n1684 , n1621 );
nand ( n1685 , n1684 , n1596 );
not ( n1686 , n1556 );
nor ( n1687 , n1596 , n1545 );
nand ( n1688 , n1686 , n1687 );
and ( n1689 , n1550 , n1682 );
not ( n1690 , n1550 );
and ( n1691 , n1690 , n1553 );
nor ( n1692 , n1689 , n1691 );
nand ( n1693 , n1692 , n1576 , n1609 );
not ( n1694 , n1693 );
nand ( n1695 , n1543 , n1554 );
not ( n1696 , n1695 );
nand ( n1697 , n1694 , n1696 );
and ( n1698 , n1685 , n1688 , n1697 );
not ( n1699 , n1665 );
nand ( n1700 , n1699 , n1585 );
nand ( n1701 , n1657 , n1581 );
and ( n1702 , n1698 , n1700 , n1701 );
nand ( n1703 , n1622 , n1546 );
not ( n1704 , n1621 );
not ( n1705 , n1584 );
and ( n1706 , n1704 , n1705 );
and ( n1707 , n1571 , n1581 );
nor ( n1708 , n1706 , n1707 );
nand ( n1709 , n1643 , n1648 );
nand ( n1710 , n1709 , n1596 );
nand ( n1711 , n1703 , n1708 , n1710 );
not ( n1712 , n1574 );
not ( n1713 , n1592 );
or ( n1714 , n1712 , n1713 );
nand ( n1715 , n1714 , n1546 );
not ( n1716 , n1577 );
nand ( n1717 , n1716 , n1596 );
nand ( n1718 , n1641 , n1715 , n1717 );
nor ( n1719 , n1711 , n1718 );
not ( n1720 , n1546 );
not ( n1721 , n1564 );
or ( n1722 , n1720 , n1721 );
nand ( n1723 , n1722 , n1652 );
nor ( n1724 , n1723 , n1620 );
nand ( n1725 , n1683 , n1702 , n1719 , n1724 );
not ( n1726 , n107 );
and ( n1727 , n1725 , n1726 );
not ( n1728 , n1725 );
and ( n1729 , n1728 , n107 );
nor ( n1730 , n1727 , n1729 );
or ( n1731 , n1730 , n356 );
not ( n1732 , n108 );
or ( n1733 , n355 , n1732 );
nand ( n1734 , n1731 , n1733 );
nor ( n1735 , n1002 , n1088 );
and ( n1736 , n966 , n1000 );
nor ( n1737 , n1426 , n1736 );
not ( n1738 , n1737 );
nor ( n1739 , n1738 , n1442 );
not ( n1740 , n1099 );
not ( n1741 , n1428 );
or ( n1742 , n1740 , n1741 );
not ( n1743 , n1011 );
nand ( n1744 , n1743 , n1059 );
nand ( n1745 , n1070 , n1744 );
nand ( n1746 , n1742 , n1745 );
nor ( n1747 , n978 , n1090 );
not ( n1748 , n1747 );
nand ( n1749 , n1748 , n1446 );
not ( n1750 , n1009 );
nand ( n1751 , n1749 , n1445 , n965 , n1750 );
not ( n1752 , n1063 );
not ( n1753 , n1051 );
and ( n1754 , n1752 , n1753 );
nor ( n1755 , n1754 , n1431 );
nand ( n1756 , n1044 , n992 , n954 );
not ( n1757 , n1756 );
nand ( n1758 , n1757 , n1000 , n989 );
nand ( n1759 , n1751 , n1755 , n1024 , n1758 );
nor ( n1760 , n1746 , n1759 );
nand ( n1761 , n1735 , n1739 , n1760 );
not ( n1762 , n113 );
and ( n1763 , n1761 , n1762 );
not ( n1764 , n1761 );
and ( n1765 , n1764 , n113 );
nor ( n1766 , n1763 , n1765 );
or ( n1767 , n1766 , n356 );
not ( n1768 , n114 );
or ( n1769 , n355 , n1768 );
nand ( n1770 , n1767 , n1769 );
not ( n1771 , n1332 );
or ( n1772 , n1394 , n1403 );
nand ( n1773 , n1772 , n1378 );
not ( n1774 , n1393 );
and ( n1775 , n1774 , n1320 );
and ( n1776 , n1400 , n1341 );
nor ( n1777 , n1775 , n1776 );
and ( n1778 , n1773 , n1777 );
not ( n1779 , n1294 );
not ( n1780 , n1322 );
and ( n1781 , n1779 , n1780 );
not ( n1782 , n1330 );
not ( n1783 , n1263 );
or ( n1784 , n1303 , n1783 );
nand ( n1785 , n1784 , n1316 );
not ( n1786 , n1785 );
or ( n1787 , n1782 , n1786 );
nand ( n1788 , n1398 , n1320 );
nand ( n1789 , n1787 , n1788 );
nor ( n1790 , n1781 , n1789 );
not ( n1791 , n1369 );
not ( n1792 , n1384 );
or ( n1793 , n1791 , n1792 );
nand ( n1794 , n1793 , n1379 );
nor ( n1795 , n1361 , n1348 );
nand ( n1796 , n1794 , n1795 );
nand ( n1797 , n1771 , n1778 , n1790 , n1796 );
not ( n1798 , n1341 );
not ( n1799 , n1311 );
or ( n1800 , n1798 , n1799 );
not ( n1801 , n1409 );
nand ( n1802 , n1800 , n1801 );
nor ( n1803 , n1797 , n1802 );
not ( n1804 , n1803 );
not ( n1805 , n126 );
and ( n1806 , n1804 , n1805 );
and ( n1807 , n1803 , n126 );
nor ( n1808 , n1806 , n1807 );
or ( n1809 , n1808 , n356 );
not ( n1810 , n127 );
or ( n1811 , n355 , n1810 );
nand ( n1812 , n1809 , n1811 );
not ( n1813 , n1188 );
not ( n1814 , n1115 );
not ( n1815 , n1814 );
nand ( n1816 , n1813 , n1815 );
not ( n1817 , n1247 );
not ( n1818 , n1227 );
not ( n1819 , n1235 );
or ( n1820 , n1818 , n1819 );
and ( n1821 , n1125 , n1169 );
not ( n1822 , n1125 );
and ( n1823 , n1822 , n1150 );
nor ( n1824 , n1821 , n1823 );
and ( n1825 , n1128 , n1814 , n1123 );
nand ( n1826 , n1824 , n1825 );
nand ( n1827 , n1820 , n1826 );
and ( n1828 , n1827 , n1114 );
not ( n1829 , n1129 );
not ( n1830 , n1180 );
or ( n1831 , n1829 , n1830 );
not ( n1832 , n1201 );
nand ( n1833 , n1831 , n1832 );
and ( n1834 , n1833 , n1190 );
nor ( n1835 , n1828 , n1834 );
nand ( n1836 , n1197 , n1170 );
not ( n1837 , n1836 );
not ( n1838 , n1180 );
and ( n1839 , n1158 , n1838 );
not ( n1840 , n1839 );
or ( n1841 , n1837 , n1840 );
nand ( n1842 , n1841 , n1131 );
nand ( n1843 , n1835 , n1842 );
not ( n1844 , n1152 );
not ( n1845 , n1232 );
not ( n1846 , n1845 );
or ( n1847 , n1844 , n1846 );
nand ( n1848 , n1235 , n1197 );
nand ( n1849 , n1847 , n1848 );
nor ( n1850 , n1224 , n1151 );
not ( n1851 , n1850 );
and ( n1852 , n1851 , n1186 );
nor ( n1853 , n1852 , n1207 );
nor ( n1854 , n1843 , n1849 , n1853 );
not ( n1855 , n1164 );
not ( n1856 , n1203 );
not ( n1857 , n1130 );
or ( n1858 , n1856 , n1857 );
nand ( n1859 , n1858 , n1212 );
nand ( n1860 , n1850 , n1117 );
nand ( n1861 , n1220 , n1241 );
and ( n1862 , n1855 , n1859 , n1860 , n1861 );
nand ( n1863 , n1816 , n1817 , n1854 , n1862 );
not ( n1864 , n130 );
and ( n1865 , n1863 , n1864 );
not ( n1866 , n1863 );
and ( n1867 , n1866 , n130 );
nor ( n1868 , n1865 , n1867 );
or ( n1869 , n1868 , n356 );
not ( n1870 , n131 );
or ( n1871 , n355 , n1870 );
nand ( n1872 , n1869 , n1871 );
not ( n1873 , n1611 );
not ( n1874 , n1622 );
or ( n1875 , n1873 , n1874 );
nand ( n1876 , n1875 , n1659 );
nor ( n1877 , n1647 , n1876 );
nand ( n1878 , n1592 , n1587 );
not ( n1879 , n1878 );
not ( n1880 , n1542 );
or ( n1881 , n1879 , n1880 );
nand ( n1882 , n1881 , n1563 );
and ( n1883 , n1608 , n1555 );
or ( n1884 , n1882 , n1883 );
not ( n1885 , n1679 );
nand ( n1886 , n1884 , n1885 );
nand ( n1887 , n1709 , n1585 );
not ( n1888 , n1682 );
not ( n1889 , n1606 );
or ( n1890 , n1888 , n1889 );
nand ( n1891 , n1890 , n1693 );
nor ( n1892 , n1543 , n1554 );
nand ( n1893 , n1891 , n1892 );
nand ( n1894 , n1571 , n1545 );
and ( n1895 , n1599 , n1887 , n1893 , n1894 );
nand ( n1896 , n1702 , n1877 , n1886 , n1895 );
not ( n1897 , n132 );
and ( n1898 , n1896 , n1897 );
not ( n1899 , n1896 );
and ( n1900 , n1899 , n132 );
nor ( n1901 , n1898 , n1900 );
or ( n1902 , n1901 , n356 );
not ( n1903 , n133 );
or ( n1904 , n355 , n1903 );
nand ( n1905 , n1902 , n1904 );
xor ( n1906 , n135 , n308 );
or ( n1907 , n1906 , n356 );
not ( n1908 , n136 );
or ( n1909 , n355 , n1908 );
nand ( n1910 , n1907 , n1909 );
not ( n1911 , n1666 );
or ( n1912 , n1569 , n1570 );
nand ( n1913 , n1912 , n1695 );
and ( n1914 , n1611 , n1913 , n1692 );
and ( n1915 , n1585 , n1639 );
nor ( n1916 , n1914 , n1915 );
nand ( n1917 , n1911 , n1916 );
nor ( n1918 , n1917 , n1711 );
nand ( n1919 , n1918 , n1601 , n1886 );
not ( n1920 , n118 );
and ( n1921 , n1919 , n1920 );
not ( n1922 , n1919 );
and ( n1923 , n1922 , n118 );
nor ( n1924 , n1921 , n1923 );
or ( n1925 , n1924 , n356 );
not ( n1926 , n119 );
or ( n1927 , n355 , n1926 );
nand ( n1928 , n1925 , n1927 );
not ( n1929 , n1172 );
or ( n1930 , n1186 , n1200 );
nand ( n1931 , n1190 , n1152 );
nand ( n1932 , n1929 , n1930 , n1931 );
and ( n1933 , n1932 , n1113 );
not ( n1934 , n1200 );
nand ( n1935 , n1934 , n1114 );
nand ( n1936 , n1839 , n1935 );
and ( n1937 , n1936 , n1235 );
nor ( n1938 , n1933 , n1937 );
not ( n1939 , n1826 );
not ( n1940 , n1114 );
and ( n1941 , n1939 , n1940 );
and ( n1942 , n1131 , n1166 );
nor ( n1943 , n1941 , n1942 );
not ( n1944 , n1211 );
and ( n1945 , n1944 , n1201 );
and ( n1946 , n1159 , n1184 );
nor ( n1947 , n1945 , n1946 );
nand ( n1948 , n1943 , n1947 );
nor ( n1949 , n1948 , n1199 );
nand ( n1950 , n1938 , n1862 , n1230 , n1949 );
not ( n1951 , n120 );
and ( n1952 , n1950 , n1951 );
not ( n1953 , n1950 );
and ( n1954 , n1953 , n120 );
nor ( n1955 , n1952 , n1954 );
or ( n1956 , n1955 , n356 );
not ( n1957 , n121 );
or ( n1958 , n355 , n1957 );
nand ( n1959 , n1956 , n1958 );
or ( n1960 , n1305 , n1322 );
or ( n1961 , n1369 , n1391 );
not ( n1962 , n1318 );
nand ( n1963 , n1962 , n1377 );
nand ( n1964 , n1963 , n1304 , n1298 );
nand ( n1965 , n1960 , n1961 , n1964 );
not ( n1966 , n1341 );
nor ( n1967 , n1966 , n1294 );
nor ( n1968 , n1965 , n1967 );
not ( n1969 , n1309 );
or ( n1970 , n1319 , n1969 , n1264 );
and ( n1971 , n1354 , n1281 );
and ( n1972 , n1309 , n1291 );
nor ( n1973 , n1971 , n1972 );
nand ( n1974 , n1352 , n1264 );
or ( n1975 , n1973 , n1974 );
nand ( n1976 , n1970 , n1975 );
nor ( n1977 , n1794 , n1976 );
or ( n1978 , n1398 , n1299 );
nand ( n1979 , n1978 , n1330 );
nand ( n1980 , n1778 , n1968 , n1977 , n1979 );
nor ( n1981 , n1345 , n1980 );
not ( n1982 , n1981 );
not ( n1983 , n77 );
and ( n1984 , n1982 , n1983 );
and ( n1985 , n1981 , n77 );
nor ( n1986 , n1984 , n1985 );
or ( n1987 , n1986 , n356 );
not ( n1988 , n86 );
or ( n1989 , n355 , n1988 );
nand ( n1990 , n1987 , n1989 );
nor ( n1991 , n1085 , n1023 );
nand ( n1992 , n1028 , n1072 );
or ( n1993 , n1991 , n1992 );
not ( n1994 , n1070 );
nand ( n1995 , n1993 , n1994 );
nand ( n1996 , n1737 , n1026 , n1463 , n1995 );
not ( n1997 , n1756 );
not ( n1998 , n1019 );
or ( n1999 , n1997 , n1998 );
nand ( n2000 , n1999 , n1099 );
and ( n2001 , n1453 , n2000 , n1041 , n1758 );
not ( n2002 , n1756 );
not ( n2003 , n1056 );
or ( n2004 , n2002 , n2003 );
nand ( n2005 , n2004 , n1070 );
not ( n2006 , n1455 );
nand ( n2007 , n2005 , n2006 );
nand ( n2008 , n1047 , n2007 );
nand ( n2009 , n2001 , n2008 );
nor ( n2010 , n1996 , n2009 );
not ( n2011 , n2010 );
not ( n2012 , n124 );
and ( n2013 , n2011 , n2012 );
and ( n2014 , n2010 , n124 );
nor ( n2015 , n2013 , n2014 );
or ( n2016 , n2015 , n356 );
not ( n2017 , n125 );
or ( n2018 , n355 , n2017 );
nand ( n2019 , n2016 , n2018 );
or ( n2020 , n766 , n356 );
not ( n2021 , n355 );
nand ( n2022 , n2021 , n115 );
nand ( n2023 , n2020 , n2022 );
endmodule
