//NOTE: no-implementation module stub

module REG2D8L (
    input wire DSPCLK,
    input wire CLKmr2renb,
    input wire MR2r_we,
    input wire [7:0] MR2rin,
    input wire [7:0] MACin,
    output reg [7:0] MR2r
);

endmodule
