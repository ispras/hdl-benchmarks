module mcst50 

















































( 

C, S, 

A0, A1, A2, A3, A4, A5 
); 

input [49:0] A0; 
input [49:0] A1; 
input [49:0] A2; 
input [49:0] A3; 
input [49:0] A4; 
input [49:0] A5; 

output [49:0] C; 
output [49:0] S; 

wire [48:0] C0; 
wire [48:0] C1; 
wire [48:0] C2; 


wire [2:0] DUMMY; 



























mcsa6 mcsa00 ( 
.S (S [00]), 
.C (C [00]), 
.COUT ({C2[00], 
C1[00], 
C0[00]}), 
.A ({A5[00], 
A4[00], 
A3[00], 
A2[00], 
A1[00], 
A0[00]}), 
.CIN ({1'B0, 
1'B0, 
1'B0 }) 
); 

mcsa6 mcsa01 ( 
.S ( S [01]), 
.C ( C [01]), 
.COUT ({C2[01], 
C1[01], 
C0[01]}), 
.A ({A5[01], 
A4[01], 
A3[01], 
A2[01], 
A1[01], 
A0[01]}), 
.CIN ({C2[00], 
C1[00], 
C0[00]}) 
); 

mcsa6 mcsa02 ( 
.S ( S [02]), 
.C ( C [02]), 
.COUT ({C2[02], 
C1[02], 
C0[02]}), 
.A ({A5[02], 
A4[02], 
A3[02], 
A2[02], 
A1[02], 
A0[02]}), 
.CIN ({C2[01], 
C1[01], 
C0[01]}) 
); 

mcsa6 mcsa03 ( 
.S ( S [03]), 
.C ( C [03]), 
.COUT ({C2[03], 
C1[03], 
C0[03]}), 
.A ({A5[03], 
A4[03], 
A3[03], 
A2[03], 
A1[03], 
A0[03]}), 
.CIN ({C2[02], 
C1[02], 
C0[02]}) 
); 

mcsa6 mcsa04 ( 
.S ( S [04]), 
.C ( C [04]), 
.COUT ({C2[04], 
C1[04], 
C0[04]}), 
.A ({A5[04], 
A4[04], 
A3[04], 
A2[04], 
A1[04], 
A0[04]}), 
.CIN ({C2[03], 
C1[03], 
C0[03]}) 
); 

mcsa6 mcsa05 ( 
.S ( S [05]), 
.C ( C [05]), 
.COUT ({C2[05], 
C1[05], 
C0[05]}), 
.A ({A5[05], 
A4[05], 
A3[05], 
A2[05], 
A1[05], 
A0[05]}), 
.CIN ({C2[04], 
C1[04], 
C0[04]}) 
); 

mcsa6 mcsa06 ( 
.S ( S [06]), 
.C ( C [06]), 
.COUT ({C2[06], 
C1[06], 
C0[06]}), 
.A ({A5[06], 
A4[06], 
A3[06], 
A2[06], 
A1[06], 
A0[06]}), 
.CIN ({C2[05], 
C1[05], 
C0[05]}) 
); 

mcsa6 mcsa07 ( 
.S ( S [07]), 
.C ( C [07]), 
.COUT ({C2[07], 
C1[07], 
C0[07]}), 
.A ({A5[07], 
A4[07], 
A3[07], 
A2[07], 
A1[07], 
A0[07]}), 
.CIN ({C2[06], 
C1[06], 
C0[06]}) 
); 

mcsa6 mcsa08 ( 
.S ( S [08]), 
.C ( C [08]), 
.COUT ({C2[08], 
C1[08], 
C0[08]}), 
.A ({A5[08], 
A4[08], 
A3[08], 
A2[08], 
A1[08], 
A0[08]}), 
.CIN ({C2[07], 
C1[07], 
C0[07]}) 
); 

mcsa6 mcsa09 ( 
.S ( S [09]), 
.C ( C [09]), 
.COUT ({C2[09], 
C1[09], 
C0[09]}), 
.A ({A5[09], 
A4[09], 
A3[09], 
A2[09], 
A1[09], 
A0[09]}), 
.CIN ({C2[08], 
C1[08], 
C0[08]}) 
); 

mcsa6 mcsa10 ( 
.S ( S [10]), 
.C ( C [10]), 
.COUT ({C2[10], 
C1[10], 
C0[10]}), 
.A ({A5[10], 
A4[10], 
A3[10], 
A2[10], 
A1[10], 
A0[10]}), 
.CIN ({C2[09], 
C1[09], 
C0[09]}) 
); 

mcsa6 mcsa11 ( 
.S ( S [11]), 
.C ( C [11]), 
.COUT ({C2[11], 
C1[11], 
C0[11]}), 
.A ({A5[11], 
A4[11], 
A3[11], 
A2[11], 
A1[11], 
A0[11]}), 
.CIN ({C2[10], 
C1[10], 
C0[10]}) 
); 

mcsa6 mcsa12 ( 
.S ( S [12]), 
.C ( C [12]), 
.COUT ({C2[12], 
C1[12], 
C0[12]}), 
.A ({A5[12], 
A4[12], 
A3[12], 
A2[12], 
A1[12], 
A0[12]}), 
.CIN ({C2[11], 
C1[11], 
C0[11]}) 
); 

mcsa6 mcsa13 ( 
.S ( S [13]), 
.C ( C [13]), 
.COUT ({C2[13], 
C1[13], 
C0[13]}), 
.A ({A5[13], 
A4[13], 
A3[13], 
A2[13], 
A1[13], 
A0[13]}), 
.CIN ({C2[12], 
C1[12], 
C0[12]}) 
); 

mcsa6 mcsa14 ( 
.S ( S [14]), 
.C ( C [14]), 
.COUT ({C2[14], 
C1[14], 
C0[14]}), 
.A ({A5[14], 
A4[14], 
A3[14], 
A2[14], 
A1[14], 
A0[14]}), 
.CIN ({C2[13], 
C1[13], 
C0[13]}) 
); 

mcsa6 mcsa15 ( 
.S ( S [15]), 
.C ( C [15]), 
.COUT ({C2[15], 
C1[15], 
C0[15]}), 
.A ({A5[15], 
A4[15], 
A3[15], 
A2[15], 
A1[15], 
A0[15]}), 
.CIN ({C2[14], 
C1[14], 
C0[14]}) 
); 

mcsa6 mcsa16 ( 
.S ( S [16]), 
.C ( C [16]), 
.COUT ({C2[16], 
C1[16], 
C0[16]}), 
.A ({A5[16], 
A4[16], 
A3[16], 
A2[16], 
A1[16], 
A0[16]}), 
.CIN ({C2[15], 
C1[15], 
C0[15]}) 
); 

mcsa6 mcsa17 ( 
.S ( S [17]), 
.C ( C [17]), 
.COUT ({C2[17], 
C1[17], 
C0[17]}), 
.A ({A5[17], 
A4[17], 
A3[17], 
A2[17], 
A1[17], 
A0[17]}), 
.CIN ({C2[16], 
C1[16], 
C0[16]}) 
); 

mcsa6 mcsa18 ( 
.S ( S [18]), 
.C ( C [18]), 
.COUT ({C2[18], 
C1[18], 
C0[18]}), 
.A ({A5[18], 
A4[18], 
A3[18], 
A2[18], 
A1[18], 
A0[18]}), 
.CIN ({C2[17], 
C1[17], 
C0[17]}) 
); 

mcsa6 mcsa19 ( 
.S ( S [19]), 
.C ( C [19]), 
.COUT ({C2[19], 
C1[19], 
C0[19]}), 
.A ({A5[19], 
A4[19], 
A3[19], 
A2[19], 
A1[19], 
A0[19]}), 
.CIN ({C2[18], 
C1[18], 
C0[18]}) 
); 

mcsa6 mcsa20 ( 
.S ( S [20]), 
.C ( C [20]), 
.COUT ({C2[20], 
C1[20], 
C0[20]}), 
.A ({A5[20], 
A4[20], 
A3[20], 
A2[20], 
A1[20], 
A0[20]}), 
.CIN ({C2[19], 
C1[19], 
C0[19]}) 
); 

mcsa6 mcsa21 ( 
.S ( S [21]), 
.C ( C [21]), 
.COUT ({C2[21], 
C1[21], 
C0[21]}), 
.A ({A5[21], 
A4[21], 
A3[21], 
A2[21], 
A1[21], 
A0[21]}), 
.CIN ({C2[20], 
C1[20], 
C0[20]}) 
); 

mcsa6 mcsa22 ( 
.S ( S [22]), 
.C ( C [22]), 
.COUT ({C2[22], 
C1[22], 
C0[22]}), 
.A ({A5[22], 
A4[22], 
A3[22], 
A2[22], 
A1[22], 
A0[22]}), 
.CIN ({C2[21], 
C1[21], 
C0[21]}) 
); 

mcsa6 mcsa23 ( 
.S ( S [23]), 
.C ( C [23]), 
.COUT ({C2[23], 
C1[23], 
C0[23]}), 
.A ({A5[23], 
A4[23], 
A3[23], 
A2[23], 
A1[23], 
A0[23]}), 
.CIN ({C2[22], 
C1[22], 
C0[22]}) 
); 

mcsa6 mcsa24 ( 
.S ( S [24]), 
.C ( C [24]), 
.COUT ({C2[24], 
C1[24], 
C0[24]}), 
.A ({A5[24], 
A4[24], 
A3[24], 
A2[24], 
A1[24], 
A0[24]}), 
.CIN ({C2[23], 
C1[23], 
C0[23]}) 
); 

mcsa6 mcsa25 ( 
.S ( S [25]), 
.C ( C [25]), 
.COUT ({C2[25], 
C1[25], 
C0[25]}), 
.A ({A5[25], 
A4[25], 
A3[25], 
A2[25], 
A1[25], 
A0[25]}), 
.CIN ({C2[24], 
C1[24], 
C0[24]}) 
); 

mcsa6 mcsa26 ( 
.S ( S [26]), 
.C ( C [26]), 
.COUT ({C2[26], 
C1[26], 
C0[26]}), 
.A ({A5[26], 
A4[26], 
A3[26], 
A2[26], 
A1[26], 
A0[26]}), 
.CIN ({C2[25], 
C1[25], 
C0[25]}) 
); 

mcsa6 mcsa27 ( 
.S ( S [27]), 
.C ( C [27]), 
.COUT ({C2[27], 
C1[27], 
C0[27]}), 
.A ({A5[27], 
A4[27], 
A3[27], 
A2[27], 
A1[27], 
A0[27]}), 
.CIN ({C2[26], 
C1[26], 
C0[26]}) 
); 

mcsa6 mcsa28 ( 
.S ( S [28]), 
.C ( C [28]), 
.COUT ({C2[28], 
C1[28], 
C0[28]}), 
.A ({A5[28], 
A4[28], 
A3[28], 
A2[28], 
A1[28], 
A0[28]}), 
.CIN ({C2[27], 
C1[27], 
C0[27]}) 
); 

mcsa6 mcsa29 ( 
.S ( S [29]), 
.C ( C [29]), 
.COUT ({C2[29], 
C1[29], 
C0[29]}), 
.A ({A5[29], 
A4[29], 
A3[29], 
A2[29], 
A1[29], 
A0[29]}), 
.CIN ({C2[28], 
C1[28], 
C0[28]}) 
); 

mcsa6 mcsa30 ( 
.S ( S [30]), 
.C ( C [30]), 
.COUT ({C2[30], 
C1[30], 
C0[30]}), 
.A ({A5[30], 
A4[30], 
A3[30], 
A2[30], 
A1[30], 
A0[30]}), 
.CIN ({C2[29], 
C1[29], 
C0[29]}) 
); 

mcsa6 mcsa31 ( 
.S ( S [31]), 
.C ( C [31]), 
.COUT ({C2[31], 
C1[31], 
C0[31]}), 
.A ({A5[31], 
A4[31], 
A3[31], 
A2[31], 
A1[31], 
A0[31]}), 
.CIN ({C2[30], 
C1[30], 
C0[30]}) 
); 

mcsa6 mcsa32 ( 
.S ( S [32]), 
.C ( C [32]), 
.COUT ({C2[32], 
C1[32], 
C0[32]}), 
.A ({A5[32], 
A4[32], 
A3[32], 
A2[32], 
A1[32], 
A0[32]}), 
.CIN ({C2[31], 
C1[31], 
C0[31]}) 
); 

mcsa6 mcsa33 ( 
.S ( S [33]), 
.C ( C [33]), 
.COUT ({C2[33], 
C1[33], 
C0[33]}), 
.A ({A5[33], 
A4[33], 
A3[33], 
A2[33], 
A1[33], 
A0[33]}), 
.CIN ({C2[32], 
C1[32], 
C0[32]}) 
); 

mcsa6 mcsa34 ( 
.S ( S [34]), 
.C ( C [34]), 
.COUT ({C2[34], 
C1[34], 
C0[34]}), 
.A ({A5[34], 
A4[34], 
A3[34], 
A2[34], 
A1[34], 
A0[34]}), 
.CIN ({C2[33], 
C1[33], 
C0[33]}) 
); 

mcsa6 mcsa35 ( 
.S ( S [35]), 
.C ( C [35]), 
.COUT ({C2[35], 
C1[35], 
C0[35]}), 
.A ({A5[35], 
A4[35], 
A3[35], 
A2[35], 
A1[35], 
A0[35]}), 
.CIN ({C2[34], 
C1[34], 
C0[34]}) 
); 

mcsa6 mcsa36 ( 
.S ( S [36]), 
.C ( C [36]), 
.COUT ({C2[36], 
C1[36], 
C0[36]}), 
.A ({A5[36], 
A4[36], 
A3[36], 
A2[36], 
A1[36], 
A0[36]}), 
.CIN ({C2[35], 
C1[35], 
C0[35]}) 
); 

mcsa6 mcsa37 ( 
.S ( S [37]), 
.C ( C [37]), 
.COUT ({C2[37], 
C1[37], 
C0[37]}), 
.A ({A5[37], 
A4[37], 
A3[37], 
A2[37], 
A1[37], 
A0[37]}), 
.CIN ({C2[36], 
C1[36], 
C0[36]}) 
); 

mcsa6 mcsa38 ( 
.S ( S [38]), 
.C ( C [38]), 
.COUT ({C2[38], 
C1[38], 
C0[38]}), 
.A ({A5[38], 
A4[38], 
A3[38], 
A2[38], 
A1[38], 
A0[38]}), 
.CIN ({C2[37], 
C1[37], 
C0[37]}) 
); 

mcsa6 mcsa39 ( 
.S ( S [39]), 
.C ( C [39]), 
.COUT ({C2[39], 
C1[39], 
C0[39]}), 
.A ({A5[39], 
A4[39], 
A3[39], 
A2[39], 
A1[39], 
A0[39]}), 
.CIN ({C2[38], 
C1[38], 
C0[38]}) 
); 

mcsa6 mcsa40 ( 
.S ( S [40]), 
.C ( C [40]), 
.COUT ({C2[40], 
C1[40], 
C0[40]}), 
.A ({A5[40], 
A4[40], 
A3[40], 
A2[40], 
A1[40], 
A0[40]}), 
.CIN ({C2[39], 
C1[39], 
C0[39]}) 
); 

mcsa6 mcsa41 ( 
.S ( S [41]), 
.C ( C [41]), 
.COUT ({C2[41], 
C1[41], 
C0[41]}), 
.A ({A5[41], 
A4[41], 
A3[41], 
A2[41], 
A1[41], 
A0[41]}), 
.CIN ({C2[40], 
C1[40], 
C0[40]}) 
); 

mcsa6 mcsa42 ( 
.S ( S [42]), 
.C ( C [42]), 
.COUT ({C2[42], 
C1[42], 
C0[42]}), 
.A ({A5[42], 
A4[42], 
A3[42], 
A2[42], 
A1[42], 
A0[42]}), 
.CIN ({C2[41], 
C1[41], 
C0[41]}) 
); 

mcsa6 mcsa43 ( 
.S ( S [43]), 
.C ( C [43]), 
.COUT ({C2[43], 
C1[43], 
C0[43]}), 
.A ({A5[43], 
A4[43], 
A3[43], 
A2[43], 
A1[43], 
A0[43]}), 
.CIN ({C2[42], 
C1[42], 
C0[42]}) 
); 

mcsa6 mcsa44 ( 
.S ( S [44]), 
.C ( C [44]), 
.COUT ({C2[44], 
C1[44], 
C0[44]}), 
.A ({A5[44], 
A4[44], 
A3[44], 
A2[44], 
A1[44], 
A0[44]}), 
.CIN ({C2[43], 
C1[43], 
C0[43]}) 
); 

mcsa6 mcsa45 ( 
.S ( S [45]), 
.C ( C [45]), 
.COUT ({C2[45], 
C1[45], 
C0[45]}), 
.A ({A5[45], 
A4[45], 
A3[45], 
A2[45], 
A1[45], 
A0[45]}), 
.CIN ({C2[44], 
C1[44], 
C0[44]}) 
); 

mcsa6 mcsa46 ( 
.S ( S [46]), 
.C ( C [46]), 
.COUT ({C2[46], 
C1[46], 
C0[46]}), 
.A ({A5[46], 
A4[46], 
A3[46], 
A2[46], 
A1[46], 
A0[46]}), 
.CIN ({C2[45], 
C1[45], 
C0[45]}) 
); 

mcsa6 mcsa47 ( 
.S ( S [47]), 
.C ( C [47]), 
.COUT ({C2[47], 
C1[47], 
C0[47]}), 
.A ({A5[47], 
A4[47], 
A3[47], 
A2[47], 
A1[47], 
A0[47]}), 
.CIN ({C2[46], 
C1[46], 
C0[46]}) 
); 

mcsa6 mcsa48 ( 
.S ( S [48]), 
.C ( C [48]), 
.COUT ({C2[48], 
C1[48], 
C0[48]}), 
.A ({A5[48], 
A4[48], 
A3[48], 
A2[48], 
A1[48], 
A0[48]}), 
.CIN ({C2[47], 
C1[47], 
C0[47]}) 
); 

mcsa6 mcsa49 ( 
.S ( S [49]), 
.C ( C [49]), 
.COUT ({DUMMY[2] , 
DUMMY[1] , 
DUMMY[0] }), 
.A ({A5[49], 
A4[49], 
A3[49], 
A2[49], 
A1[49], 
A0[49]}), 
.CIN ({C2[48], 
C1[48], 
C0[48]}) 
); 

endmodule 
