// IWLS benchmark module "MultiplierB_16" printed on Wed May 29 22:12:32 2002
module MultiplierB_16(\1 , \3 , \4 , \5 , \6 , \7 , \8 , \9 , \10 , \11 , \12 , \13 , \14 , \15 , \16 , \17 , \18 , \50 );
input
  \1 ,
  \3 ,
  \4 ,
  \5 ,
  \6 ,
  \7 ,
  \8 ,
  \9 ,
  \10 ,
  \11 ,
  \12 ,
  \13 ,
  \14 ,
  \15 ,
  \16 ,
  \17 ,
  \18 ;
output
  \50 ;
reg
  \2 ,
  \20 ,
  \21 ,
  \22 ,
  \23 ,
  \24 ,
  \25 ,
  \26 ,
  \27 ,
  \28 ,
  \29 ,
  \30 ,
  \31 ,
  \32 ,
  \33 ,
  \34 ,
  \35 ,
  \36 ,
  \37 ,
  \38 ,
  \39 ,
  \40 ,
  \41 ,
  \42 ,
  \43 ,
  \44 ,
  \45 ,
  \46 ,
  \47 ,
  \48 ;
wire
  \[59] ,
  \[60] ,
  \100 ,
  \101 ,
  \102 ,
  \103 ,
  \104 ,
  \105 ,
  \106 ,
  \107 ,
  \108 ,
  \109 ,
  \110 ,
  \111 ,
  \112 ,
  \113 ,
  \114 ,
  \115 ,
  \116 ,
  \117 ,
  \118 ,
  \119 ,
  \120 ,
  \121 ,
  \122 ,
  \123 ,
  \124 ,
  \125 ,
  \126 ,
  \127 ,
  \128 ,
  \129 ,
  \130 ,
  \131 ,
  \132 ,
  \133 ,
  \134 ,
  \135 ,
  \136 ,
  \137 ,
  \138 ,
  \139 ,
  \140 ,
  \141 ,
  \142 ,
  \143 ,
  \144 ,
  \145 ,
  \146 ,
  \147 ,
  \148 ,
  \149 ,
  \150 ,
  \151 ,
  \152 ,
  \153 ,
  \154 ,
  \155 ,
  \156 ,
  \157 ,
  \158 ,
  \159 ,
  \160 ,
  \161 ,
  \162 ,
  \163 ,
  \164 ,
  \165 ,
  \166 ,
  \167 ,
  \168 ,
  \169 ,
  \170 ,
  \171 ,
  \172 ,
  \173 ,
  \174 ,
  \175 ,
  \176 ,
  \177 ,
  \178 ,
  \179 ,
  \180 ,
  \181 ,
  \182 ,
  \183 ,
  \184 ,
  \185 ,
  \186 ,
  \187 ,
  \188 ,
  \189 ,
  \190 ,
  \191 ,
  \192 ,
  \193 ,
  \194 ,
  \195 ,
  \196 ,
  \197 ,
  \198 ,
  \199 ,
  \[31] ,
  \[32] ,
  \[33] ,
  \[34] ,
  \[35] ,
  \200 ,
  \201 ,
  \202 ,
  \203 ,
  \204 ,
  \205 ,
  \206 ,
  \207 ,
  \208 ,
  \209 ,
  \[36] ,
  \210 ,
  \211 ,
  \212 ,
  \213 ,
  \214 ,
  \215 ,
  \216 ,
  \217 ,
  \218 ,
  \219 ,
  \[37] ,
  \220 ,
  \221 ,
  \222 ,
  \223 ,
  \224 ,
  \225 ,
  \226 ,
  \227 ,
  \228 ,
  \229 ,
  \[38] ,
  \230 ,
  \231 ,
  \232 ,
  \233 ,
  \234 ,
  \235 ,
  \236 ,
  \237 ,
  \238 ,
  \239 ,
  \[39] ,
  \240 ,
  \241 ,
  \242 ,
  \243 ,
  \244 ,
  \245 ,
  \246 ,
  \247 ,
  \248 ,
  \249 ,
  \250 ,
  \251 ,
  \252 ,
  \253 ,
  \254 ,
  \255 ,
  \256 ,
  \257 ,
  \258 ,
  \259 ,
  \260 ,
  \261 ,
  \262 ,
  \263 ,
  \264 ,
  \265 ,
  \266 ,
  \[40] ,
  \[41] ,
  \[42] ,
  \[43] ,
  \[44] ,
  \[45] ,
  \[46] ,
  \[47] ,
  \[48] ,
  \[49] ,
  \49 ,
  \80 ,
  \81 ,
  \82 ,
  \83 ,
  \84 ,
  \85 ,
  \86 ,
  \87 ,
  \[50] ,
  \88 ,
  \89 ,
  \90 ,
  \91 ,
  \92 ,
  \93 ,
  \94 ,
  \95 ,
  \96 ,
  \97 ,
  \[51] ,
  \98 ,
  \99 ,
  \[52] ,
  \[53] ,
  \[54] ,
  \[55] ,
  \[56] ,
  \[57] ,
  \[58] ;
assign
  \[59]  = \183 ,
  \[60]  = \188 ,
  \100  = 0,
  \101  = 0,
  \102  = 0,
  \103  = 0,
  \104  = 0,
  \105  = 0,
  \106  = 0,
  \107  = 0,
  \108  = 0,
  \109  = 0,
  \110  = 0,
  \111  = 0,
  \112  = \18 ,
  \113  = 0,
  \114  = (~\191  & \190 ) | (\191  & ~\190 ),
  \115  = \190  & \20 ,
  \116  = \190  & \34 ,
  \117  = \20  & \34 ,
  \118  = \192  | \117 ,
  \119  = (~\194  & \193 ) | (\194  & ~\193 ),
  \120  = \193  & \21 ,
  \121  = \193  & \35 ,
  \122  = \21  & \35 ,
  \123  = \195  | \122 ,
  \124  = (~\197  & \196 ) | (\197  & ~\196 ),
  \125  = \196  & \22 ,
  \126  = \196  & \36 ,
  \127  = \22  & \36 ,
  \128  = \198  | \127 ,
  \129  = (~\200  & \199 ) | (\200  & ~\199 ),
  \130  = \199  & \23 ,
  \131  = \199  & \37 ,
  \132  = \23  & \37 ,
  \133  = \201  | \132 ,
  \134  = (~\203  & \202 ) | (\203  & ~\202 ),
  \135  = \202  & \24 ,
  \136  = \202  & \38 ,
  \137  = \24  & \38 ,
  \138  = \204  | \137 ,
  \139  = (~\206  & \205 ) | (\206  & ~\205 ),
  \140  = \205  & \25 ,
  \141  = \205  & \39 ,
  \142  = \25  & \39 ,
  \143  = \207  | \142 ,
  \144  = (~\209  & \208 ) | (\209  & ~\208 ),
  \145  = \208  & \26 ,
  \146  = \208  & \40 ,
  \147  = \26  & \40 ,
  \148  = \210  | \147 ,
  \149  = (~\212  & \211 ) | (\212  & ~\211 ),
  \150  = \211  & \27 ,
  \151  = \211  & \41 ,
  \152  = \27  & \41 ,
  \153  = \213  | \152 ,
  \154  = (~\215  & \214 ) | (\215  & ~\214 ),
  \155  = \214  & \28 ,
  \156  = \214  & \42 ,
  \157  = \28  & \42 ,
  \158  = \216  | \157 ,
  \159  = (~\218  & \217 ) | (\218  & ~\217 ),
  \160  = \217  & \29 ,
  \161  = \217  & \43 ,
  \162  = \29  & \43 ,
  \163  = \219  | \162 ,
  \164  = (~\221  & \220 ) | (\221  & ~\220 ),
  \165  = \220  & \30 ,
  \166  = \220  & \44 ,
  \167  = \30  & \44 ,
  \168  = \222  | \167 ,
  \169  = (~\224  & \223 ) | (\224  & ~\223 ),
  \170  = \223  & \31 ,
  \171  = \223  & \45 ,
  \172  = \31  & \45 ,
  \173  = \225  | \172 ,
  \174  = (~\227  & \226 ) | (\227  & ~\226 ),
  \175  = \226  & \32 ,
  \176  = \226  & \46 ,
  \177  = \32  & \46 ,
  \178  = \228  | \177 ,
  \179  = (~\230  & \229 ) | (\230  & ~\229 ),
  \180  = \229  & \33 ,
  \181  = \229  & \47 ,
  \182  = \33  & \47 ,
  \183  = \231  | \182 ,
  \184  = (~\233  & \232 ) | (\233  & ~\232 ),
  \185  = \232  & \2 ,
  \186  = \232  & \48 ,
  \187  = \2  & \48 ,
  \188  = \234  | \187 ,
  \189  = 0,
  \190  = \266  | \265 ,
  \191  = (~\20  & \34 ) | (\20  & ~\34 ),
  \192  = \116  | \115 ,
  \193  = \264  | \263 ,
  \194  = (~\21  & \35 ) | (\21  & ~\35 ),
  \195  = \121  | \120 ,
  \196  = \262  | \261 ,
  \197  = (~\22  & \36 ) | (\22  & ~\36 ),
  \198  = \126  | \125 ,
  \199  = \260  | \259 ,
  \[31]  = \49 ,
  \[32]  = \119 ,
  \[33]  = \124 ,
  \[34]  = \129 ,
  \[35]  = \134 ,
  \200  = (~\23  & \37 ) | (\23  & ~\37 ),
  \201  = \131  | \130 ,
  \202  = \258  | \257 ,
  \203  = (~\24  & \38 ) | (\24  & ~\38 ),
  \204  = \136  | \135 ,
  \205  = \256  | \255 ,
  \206  = (~\25  & \39 ) | (\25  & ~\39 ),
  \207  = \141  | \140 ,
  \208  = \254  | \253 ,
  \209  = (~\26  & \40 ) | (\26  & ~\40 ),
  \[36]  = \139 ,
  \210  = \146  | \145 ,
  \211  = \252  | \251 ,
  \212  = (~\27  & \41 ) | (\27  & ~\41 ),
  \213  = \151  | \150 ,
  \214  = \250  | \249 ,
  \215  = (~\28  & \42 ) | (\28  & ~\42 ),
  \216  = \156  | \155 ,
  \217  = \248  | \247 ,
  \218  = (~\29  & \43 ) | (\29  & ~\43 ),
  \219  = \161  | \160 ,
  \[37]  = \144 ,
  \220  = \246  | \245 ,
  \221  = (~\30  & \44 ) | (\30  & ~\44 ),
  \222  = \166  | \165 ,
  \223  = \244  | \243 ,
  \224  = (~\31  & \45 ) | (\31  & ~\45 ),
  \225  = \171  | \170 ,
  \226  = \242  | \241 ,
  \227  = (~\32  & \46 ) | (\32  & ~\46 ),
  \228  = \176  | \175 ,
  \229  = \240  | \239 ,
  \[38]  = \149 ,
  \230  = (~\33  & \47 ) | (\33  & ~\47 ),
  \231  = \181  | \180 ,
  \232  = \238  | \237 ,
  \233  = (~\2  & \48 ) | (\2  & ~\48 ),
  \234  = \186  | \185 ,
  \235  = \112  & \80 ,
  \236  = \113  & \81 ,
  \237  = \96  & \80 ,
  \238  = \111  & \81 ,
  \239  = \95  & \80 ,
  \[39]  = \154 ,
  \240  = \110  & \81 ,
  \241  = \94  & \80 ,
  \242  = \109  & \81 ,
  \243  = \93  & \80 ,
  \244  = \108  & \81 ,
  \245  = \92  & \80 ,
  \246  = \107  & \81 ,
  \247  = \91  & \80 ,
  \248  = \106  & \81 ,
  \249  = \90  & \80 ,
  \250  = \105  & \81 ,
  \251  = \89  & \80 ,
  \252  = \104  & \81 ,
  \253  = \88  & \80 ,
  \254  = \103  & \81 ,
  \255  = \87  & \80 ,
  \256  = \102  & \81 ,
  \257  = \86  & \80 ,
  \258  = \101  & \81 ,
  \259  = \85  & \80 ,
  \260  = \100  & \81 ,
  \261  = \84  & \80 ,
  \262  = \99  & \81 ,
  \263  = \83  & \80 ,
  \264  = \98  & \81 ,
  \265  = \82  & \80 ,
  \266  = \97  & \81 ,
  \[40]  = \159 ,
  \[41]  = \164 ,
  \[42]  = \169 ,
  \[43]  = \174 ,
  \[44]  = \179 ,
  \[45]  = \184 ,
  \[46]  = \118 ,
  \[47]  = \123 ,
  \[48]  = \128 ,
  \[49]  = \133 ,
  \49  = \236  | \235 ,
  \50  = \114 ,
  \80  = ~\81 ,
  \81  = (~\189  & ~\1 ) | (\189  & \1 ),
  \82  = \3 ,
  \83  = \4 ,
  \84  = \5 ,
  \85  = \6 ,
  \86  = \7 ,
  \87  = \8 ,
  \[50]  = \138 ,
  \88  = \9 ,
  \89  = \10 ,
  \90  = \11 ,
  \91  = \12 ,
  \92  = \13 ,
  \93  = \14 ,
  \94  = \15 ,
  \95  = \16 ,
  \96  = \17 ,
  \97  = 0,
  \[51]  = \143 ,
  \98  = 0,
  \99  = 0,
  \[52]  = \148 ,
  \[53]  = \153 ,
  \[54]  = \158 ,
  \[55]  = \163 ,
  \[56]  = \168 ,
  \[57]  = \173 ,
  \[58]  = \178 ;
always begin
  \2  = \[31] ;
  \20  = \[32] ;
  \21  = \[33] ;
  \22  = \[34] ;
  \23  = \[35] ;
  \24  = \[36] ;
  \25  = \[37] ;
  \26  = \[38] ;
  \27  = \[39] ;
  \28  = \[40] ;
  \29  = \[41] ;
  \30  = \[42] ;
  \31  = \[43] ;
  \32  = \[44] ;
  \33  = \[45] ;
  \34  = \[46] ;
  \35  = \[47] ;
  \36  = \[48] ;
  \37  = \[49] ;
  \38  = \[50] ;
  \39  = \[51] ;
  \40  = \[52] ;
  \41  = \[53] ;
  \42  = \[54] ;
  \43  = \[55] ;
  \44  = \[56] ;
  \45  = \[57] ;
  \46  = \[58] ;
  \47  = \[59] ;
  \48  = \[60] ;
end
initial begin
  \2  = 0;
  \20  = 0;
  \21  = 0;
  \22  = 0;
  \23  = 0;
  \24  = 0;
  \25  = 0;
  \26  = 0;
  \27  = 0;
  \28  = 0;
  \29  = 0;
  \30  = 0;
  \31  = 0;
  \32  = 0;
  \33  = 0;
  \34  = 0;
  \35  = 0;
  \36  = 0;
  \37  = 0;
  \38  = 0;
  \39  = 0;
  \40  = 0;
  \41  = 0;
  \42  = 0;
  \43  = 0;
  \44  = 0;
  \45  = 0;
  \46  = 0;
  \47  = 0;
  \48  = 0;
end
endmodule

