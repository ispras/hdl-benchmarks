//NOTE: no-implementation module stub

module UROSCAHB (
    inout wire IO,
    input wire I,
    input wire E,
    output wire O,
    input wire FEB,
    input wire EB,
    input wire S0,
    input wire S1
);
endmodule

module XFAB (
    output wire O,
    input wire I,
    input wire PU,
    input wire PD,
    input wire SMT
);
endmodule

module INV1 (
    output wire O,
    input wire I
);
endmodule

module AN2P (
    output wire O,
    input wire I1,
    input wire I2
);
endmodule

module BUF4 (
    output wire O,
    input wire I
);
endmodule

module YFA2GSB (
    output wire O,
    input wire I,
    input wire E,
    input wire E2,
    input wire E4,
    input wire E8,
    input wire SR
);
endmodule

module OR2P (
    output wire O,
    input wire I1,
    input wire I2
);
endmodule

module AO12P (
    output wire O,
    input wire A1,
    input wire B1,
    input wire B2
);
endmodule

module ZFA2GSB (
    inout wire IO,
    output wire O,
    input wire I,
    input wire E,
    input wire E8,
    input wire E4,
    input wire E2,
    input wire SMT,
    input wire PU,
    input wire PD,
    input wire SR
);
endmodule

module INV2 (
    output wire O,
    input wire I
);
endmodule
