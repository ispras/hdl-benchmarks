module RAMB4_S4_S4 (CLKA, CLKB, RSTB, RSTA, DOA, ADDRA, DIA, ENA, WEA, DOB, ADDRB, DIB, ENB, WEB);
  input CLKA;
  input CLKB;
  input RSTB;
  input RSTA;
  output [3:0] DOA;
  output [9:0] ADDRA;
  input DIA;
  output ENA;
  input WEA;
  output [3:0] DOB;
  output [9:0] ADDRB;
  output [3:0] DIB;
  output ENB;
  output WEB;
endmodule
